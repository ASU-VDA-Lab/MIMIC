module real_aes_6997_n_270 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_270);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_270;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_852;
wire n_857;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_372;
wire n_528;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_352;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_755;
wire n_284;
wire n_316;
wire n_656;
wire n_532;
wire n_746;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_278;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_713;
wire n_404;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_692;
wire n_789;
wire n_544;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_472;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_753;
wire n_283;
wire n_314;
wire n_741;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_554;
wire n_475;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_SL g557 ( .A1(n_0), .A2(n_239), .B1(n_558), .B2(n_559), .Y(n_557) );
AOI22xp33_ASAP7_75t_SL g560 ( .A1(n_1), .A2(n_109), .B1(n_366), .B2(n_561), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_2), .A2(n_249), .B1(n_355), .B2(n_640), .Y(n_639) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_3), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_4), .B(n_334), .Y(n_385) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_5), .Y(n_499) );
AOI22xp33_ASAP7_75t_SL g583 ( .A1(n_6), .A2(n_98), .B1(n_343), .B2(n_464), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_7), .A2(n_158), .B1(n_351), .B2(n_726), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_8), .B(n_325), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_9), .A2(n_75), .B1(n_355), .B2(n_501), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_10), .A2(n_266), .B1(n_325), .B2(n_332), .Y(n_324) );
XOR2x2_ASAP7_75t_L g459 ( .A(n_11), .B(n_460), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_12), .Y(n_813) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_13), .A2(n_172), .B1(n_463), .B2(n_464), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g605 ( .A(n_14), .Y(n_605) );
AOI22xp33_ASAP7_75t_SL g396 ( .A1(n_15), .A2(n_116), .B1(n_351), .B2(n_397), .Y(n_396) );
CKINVDCx20_ASAP7_75t_R g377 ( .A(n_16), .Y(n_377) );
AOI22xp33_ASAP7_75t_SL g564 ( .A1(n_17), .A2(n_214), .B1(n_393), .B2(n_565), .Y(n_564) );
AOI22xp33_ASAP7_75t_SL g687 ( .A1(n_18), .A2(n_133), .B1(n_339), .B2(n_400), .Y(n_687) );
AOI22xp33_ASAP7_75t_SL g390 ( .A1(n_19), .A2(n_181), .B1(n_339), .B2(n_391), .Y(n_390) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_20), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_21), .A2(n_31), .B1(n_380), .B2(n_669), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_22), .A2(n_493), .B1(n_530), .B2(n_531), .Y(n_492) );
INVx1_ASAP7_75t_L g531 ( .A(n_22), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_23), .A2(n_260), .B1(n_550), .B2(n_669), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_24), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_25), .A2(n_33), .B1(n_472), .B2(n_618), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_26), .A2(n_123), .B1(n_339), .B2(n_590), .Y(n_855) );
AO22x2_ASAP7_75t_L g291 ( .A1(n_27), .A2(n_85), .B1(n_292), .B2(n_293), .Y(n_291) );
INVx1_ASAP7_75t_L g802 ( .A(n_27), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_28), .A2(n_46), .B1(n_585), .B2(n_587), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g379 ( .A1(n_29), .A2(n_36), .B1(n_380), .B2(n_381), .Y(n_379) );
AOI22xp33_ASAP7_75t_SL g616 ( .A1(n_30), .A2(n_48), .B1(n_450), .B2(n_466), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_32), .B(n_661), .Y(n_660) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_34), .Y(n_778) );
CKINVDCx20_ASAP7_75t_R g842 ( .A(n_35), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_37), .A2(n_79), .B1(n_507), .B2(n_509), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_38), .A2(n_185), .B1(n_443), .B2(n_445), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_39), .A2(n_160), .B1(n_311), .B2(n_574), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_40), .A2(n_257), .B1(n_348), .B2(n_351), .Y(n_347) );
AO22x1_ASAP7_75t_L g405 ( .A1(n_41), .A2(n_406), .B1(n_457), .B2(n_458), .Y(n_405) );
INVx1_ASAP7_75t_L g457 ( .A(n_41), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g409 ( .A(n_42), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_43), .A2(n_218), .B1(n_449), .B2(n_450), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_44), .A2(n_262), .B1(n_318), .B2(n_518), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_45), .A2(n_235), .B1(n_473), .B2(n_614), .Y(n_613) );
AO22x2_ASAP7_75t_L g295 ( .A1(n_47), .A2(n_88), .B1(n_292), .B2(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g803 ( .A(n_47), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_49), .A2(n_58), .B1(n_765), .B2(n_766), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_50), .A2(n_182), .B1(n_359), .B2(n_724), .Y(n_723) );
AOI22xp33_ASAP7_75t_SL g315 ( .A1(n_51), .A2(n_195), .B1(n_316), .B2(n_321), .Y(n_315) );
AOI22xp33_ASAP7_75t_SL g721 ( .A1(n_52), .A2(n_99), .B1(n_443), .B2(n_509), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_53), .Y(n_763) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_54), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_55), .A2(n_269), .B1(n_360), .B2(n_473), .Y(n_688) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_56), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_57), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_59), .A2(n_252), .B1(n_439), .B2(n_440), .Y(n_438) );
XNOR2x1_ASAP7_75t_L g598 ( .A(n_60), .B(n_599), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_61), .A2(n_106), .B1(n_463), .B2(n_822), .Y(n_821) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_62), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g603 ( .A(n_63), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_64), .A2(n_240), .B1(n_348), .B2(n_470), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_65), .A2(n_113), .B1(n_387), .B2(n_849), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_66), .A2(n_120), .B1(n_350), .B2(n_675), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_67), .A2(n_184), .B1(n_357), .B2(n_391), .Y(n_749) );
AOI22xp33_ASAP7_75t_SL g663 ( .A1(n_68), .A2(n_142), .B1(n_580), .B2(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_69), .B(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g483 ( .A(n_70), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_71), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_72), .A2(n_196), .B1(n_467), .B2(n_561), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_73), .A2(n_125), .B1(n_339), .B2(n_343), .Y(n_338) );
CKINVDCx20_ASAP7_75t_R g626 ( .A(n_74), .Y(n_626) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_76), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_77), .A2(n_151), .B1(n_399), .B2(n_400), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_78), .A2(n_253), .B1(n_312), .B2(n_387), .Y(n_484) );
AOI22xp33_ASAP7_75t_SL g642 ( .A1(n_80), .A2(n_238), .B1(n_507), .B2(n_643), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_81), .A2(n_207), .B1(n_355), .B2(n_359), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_82), .A2(n_203), .B1(n_321), .B2(n_479), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_83), .A2(n_121), .B1(n_472), .B2(n_473), .Y(n_471) );
AOI22xp33_ASAP7_75t_SL g589 ( .A1(n_84), .A2(n_138), .B1(n_363), .B2(n_590), .Y(n_589) );
CKINVDCx20_ASAP7_75t_R g852 ( .A(n_86), .Y(n_852) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_87), .Y(n_701) );
CKINVDCx20_ASAP7_75t_R g667 ( .A(n_89), .Y(n_667) );
AOI22xp33_ASAP7_75t_SL g720 ( .A1(n_90), .A2(n_171), .B1(n_343), .B2(n_355), .Y(n_720) );
INVx1_ASAP7_75t_L g278 ( .A(n_91), .Y(n_278) );
AOI22xp33_ASAP7_75t_SL g672 ( .A1(n_92), .A2(n_149), .B1(n_587), .B2(n_673), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_93), .A2(n_189), .B1(n_380), .B2(n_664), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_94), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_95), .A2(n_179), .B1(n_399), .B2(n_400), .Y(n_737) );
INVx1_ASAP7_75t_L g276 ( .A(n_96), .Y(n_276) );
AOI22xp33_ASAP7_75t_SL g579 ( .A1(n_97), .A2(n_223), .B1(n_387), .B2(n_580), .Y(n_579) );
AOI22xp33_ASAP7_75t_SL g825 ( .A1(n_100), .A2(n_231), .B1(n_363), .B2(n_467), .Y(n_825) );
AOI22xp33_ASAP7_75t_SL g681 ( .A1(n_101), .A2(n_111), .B1(n_467), .B2(n_472), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_102), .A2(n_226), .B1(n_464), .B2(n_587), .Y(n_612) );
CKINVDCx20_ASAP7_75t_R g420 ( .A(n_103), .Y(n_420) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_104), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_105), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_107), .A2(n_119), .B1(n_453), .B2(n_456), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_108), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g624 ( .A(n_110), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_112), .A2(n_128), .B1(n_318), .B2(n_387), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_114), .A2(n_208), .B1(n_449), .B2(n_585), .Y(n_773) );
AOI22xp33_ASAP7_75t_SL g824 ( .A1(n_115), .A2(n_229), .B1(n_399), .B2(n_470), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_117), .B(n_578), .Y(n_577) );
AOI22xp33_ASAP7_75t_SL g736 ( .A1(n_118), .A2(n_213), .B1(n_352), .B2(n_444), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_122), .A2(n_256), .B1(n_312), .B2(n_381), .Y(n_606) );
AOI22xp33_ASAP7_75t_SL g820 ( .A1(n_124), .A2(n_153), .B1(n_565), .B2(n_726), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_126), .A2(n_198), .B1(n_549), .B2(n_631), .Y(n_630) );
XOR2x2_ASAP7_75t_L g702 ( .A(n_127), .B(n_703), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_129), .A2(n_211), .B1(n_359), .B2(n_453), .Y(n_566) );
CKINVDCx20_ASAP7_75t_R g553 ( .A(n_130), .Y(n_553) );
AOI22xp33_ASAP7_75t_SL g678 ( .A1(n_131), .A2(n_150), .B1(n_679), .B2(n_680), .Y(n_678) );
CKINVDCx20_ASAP7_75t_R g847 ( .A(n_132), .Y(n_847) );
INVx2_ASAP7_75t_L g279 ( .A(n_134), .Y(n_279) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_135), .Y(n_430) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_136), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_137), .A2(n_143), .B1(n_467), .B2(n_592), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_139), .A2(n_227), .B1(n_348), .B2(n_559), .Y(n_647) );
OA22x2_ASAP7_75t_L g655 ( .A1(n_140), .A2(n_656), .B1(n_657), .B2(n_682), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_140), .Y(n_656) );
INVx1_ASAP7_75t_L g402 ( .A(n_141), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_144), .B(n_334), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_145), .B(n_476), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_146), .A2(n_263), .B1(n_443), .B2(n_618), .Y(n_774) );
AND2x6_ASAP7_75t_L g275 ( .A(n_147), .B(n_276), .Y(n_275) );
HB1xp67_ASAP7_75t_L g796 ( .A(n_147), .Y(n_796) );
AO22x2_ASAP7_75t_L g299 ( .A1(n_148), .A2(n_222), .B1(n_292), .B2(n_296), .Y(n_299) );
CKINVDCx20_ASAP7_75t_R g707 ( .A(n_152), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_154), .A2(n_250), .B1(n_550), .B2(n_669), .Y(n_692) );
CKINVDCx20_ASAP7_75t_R g302 ( .A(n_155), .Y(n_302) );
CKINVDCx20_ASAP7_75t_R g633 ( .A(n_156), .Y(n_633) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_157), .Y(n_545) );
AOI211xp5_ASAP7_75t_L g270 ( .A1(n_159), .A2(n_271), .B(n_280), .C(n_804), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_161), .A2(n_206), .B1(n_305), .B2(n_318), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g809 ( .A(n_162), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g423 ( .A(n_163), .Y(n_423) );
CKINVDCx20_ASAP7_75t_R g572 ( .A(n_164), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_165), .B(n_384), .Y(n_383) );
CKINVDCx20_ASAP7_75t_R g629 ( .A(n_166), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g805 ( .A1(n_167), .A2(n_806), .B1(n_826), .B2(n_827), .Y(n_805) );
CKINVDCx20_ASAP7_75t_R g826 ( .A(n_167), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_168), .A2(n_268), .B1(n_476), .B2(n_477), .Y(n_475) );
XNOR2x1_ASAP7_75t_L g567 ( .A(n_169), .B(n_568), .Y(n_567) );
AO22x2_ASAP7_75t_L g301 ( .A1(n_170), .A2(n_241), .B1(n_292), .B2(n_293), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_173), .A2(n_265), .B1(n_357), .B2(n_363), .Y(n_700) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_174), .Y(n_810) );
CKINVDCx20_ASAP7_75t_R g414 ( .A(n_175), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_176), .A2(n_219), .B1(n_357), .B2(n_393), .Y(n_392) );
AOI22xp5_ASAP7_75t_L g465 ( .A1(n_177), .A2(n_251), .B1(n_466), .B2(n_467), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g602 ( .A(n_178), .Y(n_602) );
AOI22xp33_ASAP7_75t_SL g303 ( .A1(n_180), .A2(n_197), .B1(n_304), .B2(n_310), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_183), .A2(n_209), .B1(n_675), .B2(n_676), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_186), .Y(n_523) );
XNOR2x1_ASAP7_75t_L g620 ( .A(n_187), .B(n_621), .Y(n_620) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_188), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g817 ( .A(n_190), .Y(n_817) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_191), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_192), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_193), .A2(n_258), .B1(n_363), .B2(n_366), .Y(n_362) );
CKINVDCx20_ASAP7_75t_R g853 ( .A(n_194), .Y(n_853) );
CKINVDCx20_ASAP7_75t_R g635 ( .A(n_199), .Y(n_635) );
AOI22xp33_ASAP7_75t_SL g698 ( .A1(n_200), .A2(n_264), .B1(n_351), .B2(n_699), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g857 ( .A1(n_201), .A2(n_245), .B1(n_640), .B2(n_858), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_202), .B(n_384), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g609 ( .A(n_204), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_205), .B(n_334), .Y(n_695) );
OA22x2_ASAP7_75t_L g283 ( .A1(n_210), .A2(n_284), .B1(n_285), .B2(n_368), .Y(n_283) );
CKINVDCx20_ASAP7_75t_R g284 ( .A(n_210), .Y(n_284) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_212), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_215), .Y(n_785) );
CKINVDCx20_ASAP7_75t_R g836 ( .A(n_216), .Y(n_836) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_217), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_220), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_221), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g800 ( .A(n_222), .B(n_801), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_224), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_225), .Y(n_706) );
CKINVDCx20_ASAP7_75t_R g691 ( .A(n_228), .Y(n_691) );
AOI22xp33_ASAP7_75t_SL g645 ( .A1(n_230), .A2(n_236), .B1(n_339), .B2(n_646), .Y(n_645) );
CKINVDCx20_ASAP7_75t_R g425 ( .A(n_232), .Y(n_425) );
AOI22xp33_ASAP7_75t_SL g748 ( .A1(n_233), .A2(n_267), .B1(n_350), .B2(n_455), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g843 ( .A(n_234), .Y(n_843) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_237), .Y(n_514) );
INVx1_ASAP7_75t_L g799 ( .A(n_241), .Y(n_799) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_242), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_243), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_244), .B(n_631), .Y(n_713) );
OA22x2_ASAP7_75t_L g752 ( .A1(n_246), .A2(n_753), .B1(n_754), .B2(n_755), .Y(n_752) );
CKINVDCx16_ASAP7_75t_R g753 ( .A(n_246), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g776 ( .A(n_247), .Y(n_776) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_248), .Y(n_540) );
INVx1_ASAP7_75t_L g292 ( .A(n_254), .Y(n_292) );
INVx1_ASAP7_75t_L g294 ( .A(n_254), .Y(n_294) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_255), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g608 ( .A(n_259), .Y(n_608) );
CKINVDCx20_ASAP7_75t_R g427 ( .A(n_261), .Y(n_427) );
CKINVDCx20_ASAP7_75t_R g271 ( .A(n_272), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_273), .Y(n_272) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
HB1xp67_ASAP7_75t_L g795 ( .A(n_276), .Y(n_795) );
OAI21xp5_ASAP7_75t_L g834 ( .A1(n_277), .A2(n_794), .B(n_835), .Y(n_834) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
AOI221xp5_ASAP7_75t_SL g280 ( .A1(n_281), .A2(n_595), .B1(n_789), .B2(n_790), .C(n_791), .Y(n_280) );
INVx1_ASAP7_75t_L g789 ( .A(n_281), .Y(n_789) );
XOR2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_488), .Y(n_281) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_369), .B1(n_486), .B2(n_487), .Y(n_282) );
INVx1_ASAP7_75t_L g486 ( .A(n_283), .Y(n_486) );
INVx2_ASAP7_75t_L g368 ( .A(n_285), .Y(n_368) );
NAND2x1_ASAP7_75t_L g285 ( .A(n_286), .B(n_336), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_287), .B(n_314), .Y(n_286) );
OAI21xp5_ASAP7_75t_SL g287 ( .A1(n_288), .A2(n_302), .B(n_303), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g378 ( .A(n_289), .Y(n_378) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_289), .Y(n_422) );
BUFx3_ASAP7_75t_L g482 ( .A(n_289), .Y(n_482) );
INVx2_ASAP7_75t_SL g546 ( .A(n_289), .Y(n_546) );
INVx4_ASAP7_75t_L g571 ( .A(n_289), .Y(n_571) );
AND2x6_ASAP7_75t_L g289 ( .A(n_290), .B(n_297), .Y(n_289) );
AND2x4_ASAP7_75t_L g321 ( .A(n_290), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g434 ( .A(n_290), .Y(n_434) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_295), .Y(n_290) );
AND2x2_ASAP7_75t_L g309 ( .A(n_291), .B(n_299), .Y(n_309) );
INVx2_ASAP7_75t_L g331 ( .A(n_291), .Y(n_331) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g296 ( .A(n_294), .Y(n_296) );
INVx2_ASAP7_75t_L g308 ( .A(n_295), .Y(n_308) );
INVx1_ASAP7_75t_L g320 ( .A(n_295), .Y(n_320) );
OR2x2_ASAP7_75t_L g330 ( .A(n_295), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g335 ( .A(n_295), .B(n_331), .Y(n_335) );
AND2x6_ASAP7_75t_L g350 ( .A(n_297), .B(n_329), .Y(n_350) );
AND2x4_ASAP7_75t_L g352 ( .A(n_297), .B(n_335), .Y(n_352) );
AND2x2_ASAP7_75t_L g358 ( .A(n_297), .B(n_342), .Y(n_358) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_300), .Y(n_297) );
AND2x2_ASAP7_75t_L g328 ( .A(n_298), .B(n_301), .Y(n_328) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g341 ( .A(n_299), .B(n_323), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_299), .B(n_301), .Y(n_346) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g307 ( .A(n_301), .Y(n_307) );
INVx1_ASAP7_75t_L g323 ( .A(n_301), .Y(n_323) );
INVx1_ASAP7_75t_L g419 ( .A(n_304), .Y(n_419) );
BUFx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_305), .Y(n_387) );
BUFx4f_ASAP7_75t_SL g518 ( .A(n_305), .Y(n_518) );
BUFx6f_ASAP7_75t_L g631 ( .A(n_305), .Y(n_631) );
BUFx6f_ASAP7_75t_L g664 ( .A(n_305), .Y(n_664) );
AND2x4_ASAP7_75t_L g305 ( .A(n_306), .B(n_309), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx1_ASAP7_75t_L g313 ( .A(n_307), .Y(n_313) );
AND2x2_ASAP7_75t_L g342 ( .A(n_308), .B(n_331), .Y(n_342) );
INVx1_ASAP7_75t_L g401 ( .A(n_308), .Y(n_401) );
AND2x4_ASAP7_75t_L g312 ( .A(n_309), .B(n_313), .Y(n_312) );
AND2x4_ASAP7_75t_L g318 ( .A(n_309), .B(n_319), .Y(n_318) );
NAND2x1p5_ASAP7_75t_L g429 ( .A(n_309), .B(n_401), .Y(n_429) );
INVx2_ASAP7_75t_L g424 ( .A(n_310), .Y(n_424) );
BUFx3_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g851 ( .A(n_311), .Y(n_851) );
BUFx6f_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
BUFx12f_ASAP7_75t_L g380 ( .A(n_312), .Y(n_380) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_312), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_324), .Y(n_314) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
BUFx3_ASAP7_75t_L g479 ( .A(n_318), .Y(n_479) );
BUFx2_ASAP7_75t_L g580 ( .A(n_318), .Y(n_580) );
BUFx2_ASAP7_75t_L g849 ( .A(n_318), .Y(n_849) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
OR2x6_ASAP7_75t_L g367 ( .A(n_320), .B(n_346), .Y(n_367) );
BUFx3_ASAP7_75t_L g381 ( .A(n_321), .Y(n_381) );
BUFx2_ASAP7_75t_SL g574 ( .A(n_321), .Y(n_574) );
BUFx6f_ASAP7_75t_L g669 ( .A(n_321), .Y(n_669) );
INVx1_ASAP7_75t_L g435 ( .A(n_322), .Y(n_435) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g384 ( .A(n_326), .Y(n_384) );
INVx2_ASAP7_75t_L g476 ( .A(n_326), .Y(n_476) );
INVx5_ASAP7_75t_L g744 ( .A(n_326), .Y(n_744) );
INVx4_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
AND2x6_ASAP7_75t_L g334 ( .A(n_328), .B(n_335), .Y(n_334) );
AND2x4_ASAP7_75t_L g361 ( .A(n_328), .B(n_342), .Y(n_361) );
INVx1_ASAP7_75t_L g413 ( .A(n_328), .Y(n_413) );
NAND2x1p5_ASAP7_75t_L g417 ( .A(n_328), .B(n_335), .Y(n_417) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g412 ( .A(n_330), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_SL g661 ( .A(n_333), .Y(n_661) );
INVx1_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
BUFx4f_ASAP7_75t_L g477 ( .A(n_334), .Y(n_477) );
BUFx2_ASAP7_75t_L g578 ( .A(n_334), .Y(n_578) );
AND2x2_ASAP7_75t_L g365 ( .A(n_335), .B(n_341), .Y(n_365) );
NOR2x1_ASAP7_75t_L g336 ( .A(n_337), .B(n_353), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_338), .B(n_347), .Y(n_337) );
BUFx3_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
BUFx3_ASAP7_75t_L g455 ( .A(n_340), .Y(n_455) );
BUFx3_ASAP7_75t_L g464 ( .A(n_340), .Y(n_464) );
BUFx3_ASAP7_75t_L g673 ( .A(n_340), .Y(n_673) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_341), .B(n_342), .Y(n_781) );
AND2x4_ASAP7_75t_L g344 ( .A(n_342), .B(n_345), .Y(n_344) );
BUFx2_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
BUFx3_ASAP7_75t_L g391 ( .A(n_344), .Y(n_391) );
BUFx3_ASAP7_75t_L g456 ( .A(n_344), .Y(n_456) );
BUFx3_ASAP7_75t_L g473 ( .A(n_344), .Y(n_473) );
INVx1_ASAP7_75t_L g504 ( .A(n_344), .Y(n_504) );
BUFx2_ASAP7_75t_SL g565 ( .A(n_344), .Y(n_565) );
BUFx2_ASAP7_75t_L g676 ( .A(n_344), .Y(n_676) );
AND2x2_ASAP7_75t_L g400 ( .A(n_345), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx4_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_SL g724 ( .A(n_349), .Y(n_724) );
INVx3_ASAP7_75t_L g822 ( .A(n_349), .Y(n_822) );
INVx11_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx11_ASAP7_75t_L g394 ( .A(n_350), .Y(n_394) );
INVx3_ASAP7_75t_L g498 ( .A(n_351), .Y(n_498) );
BUFx3_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx6_ASAP7_75t_L g451 ( .A(n_352), .Y(n_451) );
BUFx3_ASAP7_75t_L g559 ( .A(n_352), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_362), .Y(n_353) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx3_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx3_ASAP7_75t_L g439 ( .A(n_357), .Y(n_439) );
BUFx3_ASAP7_75t_L g558 ( .A(n_357), .Y(n_558) );
BUFx6f_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
BUFx2_ASAP7_75t_SL g470 ( .A(n_358), .Y(n_470) );
INVx2_ASAP7_75t_L g586 ( .A(n_358), .Y(n_586) );
BUFx2_ASAP7_75t_SL g675 ( .A(n_358), .Y(n_675) );
BUFx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
BUFx3_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_361), .Y(n_399) );
INVx2_ASAP7_75t_L g441 ( .A(n_361), .Y(n_441) );
BUFx3_ASAP7_75t_L g472 ( .A(n_361), .Y(n_472) );
BUFx3_ASAP7_75t_L g592 ( .A(n_361), .Y(n_592) );
INVx3_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx5_ASAP7_75t_L g397 ( .A(n_364), .Y(n_397) );
INVx4_ASAP7_75t_L g444 ( .A(n_364), .Y(n_444) );
INVx2_ASAP7_75t_L g466 ( .A(n_364), .Y(n_466) );
BUFx3_ASAP7_75t_L g508 ( .A(n_364), .Y(n_508) );
INVx1_ASAP7_75t_L g680 ( .A(n_364), .Y(n_680) );
INVx8_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
INVx6_ASAP7_75t_SL g446 ( .A(n_367), .Y(n_446) );
INVx1_ASAP7_75t_L g509 ( .A(n_367), .Y(n_509) );
INVx1_ASAP7_75t_SL g643 ( .A(n_367), .Y(n_643) );
INVx1_ASAP7_75t_L g487 ( .A(n_369), .Y(n_487) );
XOR2xp5_ASAP7_75t_L g369 ( .A(n_370), .B(n_403), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx3_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
XOR2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_402), .Y(n_373) );
NAND2x1p5_ASAP7_75t_L g374 ( .A(n_375), .B(n_388), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_376), .B(n_382), .Y(n_375) );
OAI21xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_378), .B(n_379), .Y(n_376) );
OAI222xp33_ASAP7_75t_L g516 ( .A1(n_378), .A2(n_517), .B1(n_519), .B2(n_520), .C1(n_521), .C2(n_523), .Y(n_516) );
OAI21xp33_ASAP7_75t_SL g628 ( .A1(n_378), .A2(n_629), .B(n_630), .Y(n_628) );
OAI221xp5_ASAP7_75t_L g710 ( .A1(n_378), .A2(n_424), .B1(n_711), .B2(n_712), .C(n_713), .Y(n_710) );
BUFx4f_ASAP7_75t_SL g527 ( .A(n_380), .Y(n_527) );
INVx2_ASAP7_75t_L g767 ( .A(n_380), .Y(n_767) );
NAND3xp33_ASAP7_75t_L g382 ( .A(n_383), .B(n_385), .C(n_386), .Y(n_382) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_387), .Y(n_544) );
NOR2x1_ASAP7_75t_L g388 ( .A(n_389), .B(n_395), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
INVx2_ASAP7_75t_L g859 ( .A(n_391), .Y(n_859) );
INVx5_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g449 ( .A(n_394), .Y(n_449) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_394), .Y(n_496) );
INVx4_ASAP7_75t_L g587 ( .A(n_394), .Y(n_587) );
INVx2_ASAP7_75t_SL g699 ( .A(n_394), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_396), .B(n_398), .Y(n_395) );
INVx4_ASAP7_75t_L g641 ( .A(n_399), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_405), .B1(n_459), .B2(n_485), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_SL g458 ( .A(n_406), .Y(n_458) );
AND2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_436), .Y(n_406) );
NOR3xp33_ASAP7_75t_L g407 ( .A(n_408), .B(n_418), .C(n_426), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B1(n_414), .B2(n_415), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g705 ( .A1(n_410), .A2(n_706), .B1(n_707), .B2(n_708), .Y(n_705) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_SL g513 ( .A(n_411), .Y(n_513) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_412), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_412), .A2(n_415), .B1(n_602), .B2(n_603), .Y(n_601) );
BUFx3_ASAP7_75t_L g625 ( .A(n_412), .Y(n_625) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g811 ( .A(n_416), .Y(n_811) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx3_ASAP7_75t_L g515 ( .A(n_417), .Y(n_515) );
OAI222xp33_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_420), .B1(n_421), .B2(n_423), .C1(n_424), .C2(n_425), .Y(n_418) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_419), .A2(n_521), .B1(n_608), .B2(n_609), .Y(n_607) );
INVx2_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_428), .B1(n_430), .B2(n_431), .Y(n_426) );
OAI22xp5_ASAP7_75t_SL g552 ( .A1(n_428), .A2(n_431), .B1(n_553), .B2(n_554), .Y(n_552) );
BUFx3_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx4_ASAP7_75t_L g522 ( .A(n_429), .Y(n_522) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_429), .Y(n_716) );
OAI22xp33_ASAP7_75t_SL g768 ( .A1(n_429), .A2(n_431), .B1(n_769), .B2(n_770), .Y(n_768) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_431), .A2(n_715), .B1(n_716), .B2(n_717), .Y(n_714) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g636 ( .A(n_432), .Y(n_636) );
CKINVDCx16_ASAP7_75t_R g432 ( .A(n_433), .Y(n_432) );
BUFx2_ASAP7_75t_L g529 ( .A(n_433), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_433), .A2(n_634), .B1(n_816), .B2(n_817), .Y(n_815) );
OR2x6_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_437), .B(n_447), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_442), .Y(n_437) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OAI221xp5_ASAP7_75t_SL g502 ( .A1(n_441), .A2(n_503), .B1(n_504), .B2(n_505), .C(n_506), .Y(n_502) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g562 ( .A(n_444), .Y(n_562) );
BUFx4f_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
BUFx2_ASAP7_75t_L g467 ( .A(n_446), .Y(n_467) );
BUFx2_ASAP7_75t_L g618 ( .A(n_446), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g447 ( .A(n_448), .B(n_452), .Y(n_447) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g463 ( .A(n_451), .Y(n_463) );
INVx3_ASAP7_75t_L g590 ( .A(n_451), .Y(n_590) );
INVx2_ASAP7_75t_L g679 ( .A(n_451), .Y(n_679) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx4f_ASAP7_75t_SL g726 ( .A(n_455), .Y(n_726) );
INVx1_ASAP7_75t_SL g485 ( .A(n_459), .Y(n_485) );
NOR4xp75_ASAP7_75t_L g460 ( .A(n_461), .B(n_468), .C(n_474), .D(n_480), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_462), .B(n_465), .Y(n_461) );
INVx2_ASAP7_75t_L g777 ( .A(n_463), .Y(n_777) );
BUFx3_ASAP7_75t_L g501 ( .A(n_464), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_469), .B(n_471), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_475), .B(n_478), .Y(n_474) );
OAI21xp5_ASAP7_75t_SL g480 ( .A1(n_481), .A2(n_483), .B(n_484), .Y(n_480) );
OAI21xp33_ASAP7_75t_L g604 ( .A1(n_481), .A2(n_605), .B(n_606), .Y(n_604) );
OAI21xp33_ASAP7_75t_SL g762 ( .A1(n_481), .A2(n_763), .B(n_764), .Y(n_762) );
INVx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_492), .B1(n_532), .B2(n_533), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g530 ( .A(n_493), .Y(n_530) );
AND2x2_ASAP7_75t_SL g493 ( .A(n_494), .B(n_510), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_495), .B(n_502), .Y(n_494) );
OAI221xp5_ASAP7_75t_SL g495 ( .A1(n_496), .A2(n_497), .B1(n_498), .B2(n_499), .C(n_500), .Y(n_495) );
INVx1_ASAP7_75t_L g646 ( .A(n_504), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g782 ( .A1(n_504), .A2(n_783), .B1(n_784), .B2(n_785), .Y(n_782) );
INVx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NOR3xp33_ASAP7_75t_L g510 ( .A(n_511), .B(n_516), .C(n_524), .Y(n_510) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_513), .B1(n_514), .B2(n_515), .Y(n_511) );
OAI22xp5_ASAP7_75t_SL g538 ( .A1(n_515), .A2(n_539), .B1(n_540), .B2(n_541), .Y(n_538) );
BUFx3_ASAP7_75t_L g627 ( .A(n_515), .Y(n_627) );
INVx2_ASAP7_75t_L g709 ( .A(n_515), .Y(n_709) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx3_ASAP7_75t_SL g634 ( .A(n_522), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_526), .B1(n_528), .B2(n_529), .Y(n_524) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
OAI22xp5_ASAP7_75t_SL g850 ( .A1(n_529), .A2(n_851), .B1(n_852), .B2(n_853), .Y(n_850) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
OAI22xp5_ASAP7_75t_SL g533 ( .A1(n_534), .A2(n_567), .B1(n_593), .B2(n_594), .Y(n_533) );
INVx2_ASAP7_75t_L g593 ( .A(n_534), .Y(n_593) );
XNOR2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_555), .Y(n_536) );
NOR3xp33_ASAP7_75t_L g537 ( .A(n_538), .B(n_542), .C(n_552), .Y(n_537) );
INVx1_ASAP7_75t_L g759 ( .A(n_539), .Y(n_759) );
OAI22xp5_ASAP7_75t_L g808 ( .A1(n_539), .A2(n_809), .B1(n_810), .B2(n_811), .Y(n_808) );
OAI222xp33_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_545), .B1(n_546), .B2(n_547), .C1(n_548), .C2(n_551), .Y(n_542) );
INVx2_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
OAI21xp5_ASAP7_75t_SL g812 ( .A1(n_546), .A2(n_813), .B(n_814), .Y(n_812) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
BUFx4f_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_556), .B(n_563), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_560), .Y(n_556) );
INVx3_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_566), .Y(n_563) );
INVx2_ASAP7_75t_L g594 ( .A(n_567), .Y(n_594) );
AND2x4_ASAP7_75t_L g568 ( .A(n_569), .B(n_581), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_570), .B(n_575), .Y(n_569) );
OAI21xp5_ASAP7_75t_SL g570 ( .A1(n_571), .A2(n_572), .B(n_573), .Y(n_570) );
BUFx2_ASAP7_75t_L g666 ( .A(n_571), .Y(n_666) );
OAI21xp5_ASAP7_75t_L g690 ( .A1(n_571), .A2(n_691), .B(n_692), .Y(n_690) );
OAI21xp5_ASAP7_75t_L g739 ( .A1(n_571), .A2(n_740), .B(n_741), .Y(n_739) );
INVx4_ASAP7_75t_L g846 ( .A(n_571), .Y(n_846) );
NAND3xp33_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .C(n_579), .Y(n_575) );
NOR2x1_ASAP7_75t_L g581 ( .A(n_582), .B(n_588), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
INVx3_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx3_ASAP7_75t_L g614 ( .A(n_586), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_591), .Y(n_588) );
INVx1_ASAP7_75t_L g784 ( .A(n_592), .Y(n_784) );
INVx1_ASAP7_75t_L g790 ( .A(n_595), .Y(n_790) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_648), .B1(n_787), .B2(n_788), .Y(n_595) );
CKINVDCx20_ASAP7_75t_R g787 ( .A(n_596), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B1(n_619), .B2(n_620), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_610), .Y(n_599) );
NOR3xp33_ASAP7_75t_L g600 ( .A(n_601), .B(n_604), .C(n_607), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_611), .B(n_615), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_637), .Y(n_621) );
NOR3xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_628), .C(n_632), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_625), .B1(n_626), .B2(n_627), .Y(n_623) );
OAI22xp5_ASAP7_75t_SL g757 ( .A1(n_627), .A2(n_758), .B1(n_760), .B2(n_761), .Y(n_757) );
BUFx2_ASAP7_75t_L g765 ( .A(n_631), .Y(n_765) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_634), .B1(n_635), .B2(n_636), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_638), .B(n_644), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_639), .B(n_642), .Y(n_638) );
INVx4_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_647), .Y(n_644) );
INVx1_ASAP7_75t_L g788 ( .A(n_648), .Y(n_788) );
XOR2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_728), .Y(n_648) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_653), .B1(n_702), .B2(n_727), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OAI22xp5_ASAP7_75t_SL g653 ( .A1(n_654), .A2(n_655), .B1(n_683), .B2(n_684), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx2_ASAP7_75t_SL g682 ( .A(n_657), .Y(n_682) );
NAND2x1p5_ASAP7_75t_L g657 ( .A(n_658), .B(n_670), .Y(n_657) );
NOR2xp67_ASAP7_75t_SL g658 ( .A(n_659), .B(n_665), .Y(n_658) );
NAND3xp33_ASAP7_75t_L g659 ( .A(n_660), .B(n_662), .C(n_663), .Y(n_659) );
OAI21xp5_ASAP7_75t_SL g665 ( .A1(n_666), .A2(n_667), .B(n_668), .Y(n_665) );
NOR2x1_ASAP7_75t_L g670 ( .A(n_671), .B(n_677), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_672), .B(n_674), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_681), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_683), .A2(n_729), .B1(n_730), .B2(n_731), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_683), .Y(n_729) );
INVx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
XOR2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_701), .Y(n_684) );
NAND3x1_ASAP7_75t_L g685 ( .A(n_686), .B(n_689), .C(n_697), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
NOR2x1_ASAP7_75t_L g689 ( .A(n_690), .B(n_693), .Y(n_689) );
NAND3xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .C(n_696), .Y(n_693) );
AND2x2_ASAP7_75t_L g697 ( .A(n_698), .B(n_700), .Y(n_697) );
INVx2_ASAP7_75t_L g727 ( .A(n_702), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_704), .B(n_718), .Y(n_703) );
NOR3xp33_ASAP7_75t_L g704 ( .A(n_705), .B(n_710), .C(n_714), .Y(n_704) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_719), .B(n_722), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_723), .B(n_725), .Y(n_722) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_751), .B1(n_752), .B2(n_786), .Y(n_732) );
INVx3_ASAP7_75t_L g786 ( .A(n_733), .Y(n_786) );
XOR2x2_ASAP7_75t_L g733 ( .A(n_734), .B(n_750), .Y(n_733) );
NAND3x1_ASAP7_75t_SL g734 ( .A(n_735), .B(n_738), .C(n_747), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
NOR2x1_ASAP7_75t_L g738 ( .A(n_739), .B(n_742), .Y(n_738) );
NAND3xp33_ASAP7_75t_L g742 ( .A(n_743), .B(n_745), .C(n_746), .Y(n_742) );
AND2x2_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .Y(n_747) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
AND2x2_ASAP7_75t_L g755 ( .A(n_756), .B(n_771), .Y(n_755) );
NOR3xp33_ASAP7_75t_L g756 ( .A(n_757), .B(n_762), .C(n_768), .Y(n_756) );
OAI22xp5_ASAP7_75t_L g841 ( .A1(n_758), .A2(n_811), .B1(n_842), .B2(n_843), .Y(n_841) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx3_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
NOR3xp33_ASAP7_75t_L g771 ( .A(n_772), .B(n_775), .C(n_782), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_773), .B(n_774), .Y(n_772) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_777), .B1(n_778), .B2(n_779), .Y(n_775) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_SL g791 ( .A(n_792), .Y(n_791) );
NOR2x1_ASAP7_75t_L g792 ( .A(n_793), .B(n_797), .Y(n_792) );
OR2x2_ASAP7_75t_SL g863 ( .A(n_793), .B(n_798), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_794), .B(n_796), .Y(n_793) );
CKINVDCx20_ASAP7_75t_R g829 ( .A(n_794), .Y(n_829) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_795), .B(n_832), .Y(n_835) );
CKINVDCx16_ASAP7_75t_R g832 ( .A(n_796), .Y(n_832) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_798), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_802), .B(n_803), .Y(n_801) );
OAI322xp33_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_828), .A3(n_830), .B1(n_833), .B2(n_836), .C1(n_837), .C2(n_861), .Y(n_804) );
INVx2_ASAP7_75t_L g827 ( .A(n_806), .Y(n_827) );
AND2x2_ASAP7_75t_L g806 ( .A(n_807), .B(n_818), .Y(n_806) );
NOR3xp33_ASAP7_75t_L g807 ( .A(n_808), .B(n_812), .C(n_815), .Y(n_807) );
NOR2xp33_ASAP7_75t_L g818 ( .A(n_819), .B(n_823), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_820), .B(n_821), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_824), .B(n_825), .Y(n_823) );
HB1xp67_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
HB1xp67_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
CKINVDCx20_ASAP7_75t_R g833 ( .A(n_834), .Y(n_833) );
XNOR2x1_ASAP7_75t_L g838 ( .A(n_836), .B(n_839), .Y(n_838) );
HB1xp67_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
AND2x2_ASAP7_75t_L g839 ( .A(n_840), .B(n_854), .Y(n_839) );
NOR3xp33_ASAP7_75t_L g840 ( .A(n_841), .B(n_844), .C(n_850), .Y(n_840) );
OAI21xp33_ASAP7_75t_SL g844 ( .A1(n_845), .A2(n_847), .B(n_848), .Y(n_844) );
INVx2_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
AND4x1_ASAP7_75t_L g854 ( .A(n_855), .B(n_856), .C(n_857), .D(n_860), .Y(n_854) );
INVx2_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
CKINVDCx20_ASAP7_75t_R g861 ( .A(n_862), .Y(n_861) );
CKINVDCx20_ASAP7_75t_R g862 ( .A(n_863), .Y(n_862) );
endmodule