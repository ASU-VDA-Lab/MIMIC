module fake_jpeg_20287_n_129 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_129);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_5),
.B(n_8),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_19),
.Y(n_39)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_27),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_35),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_37),
.B(n_21),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_39),
.A2(n_50),
.B1(n_16),
.B2(n_32),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_35),
.A2(n_17),
.B1(n_20),
.B2(n_22),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_42),
.A2(n_35),
.B1(n_32),
.B2(n_28),
.Y(n_73)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_29),
.A2(n_20),
.B1(n_17),
.B2(n_26),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_31),
.B(n_19),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_48),
.B(n_23),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_29),
.A2(n_20),
.B1(n_26),
.B2(n_16),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_60),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_34),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_54),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_45),
.B(n_37),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_33),
.B(n_21),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_34),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_62),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_40),
.B(n_25),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_30),
.B1(n_32),
.B2(n_28),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_65),
.B1(n_22),
.B2(n_18),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_49),
.B(n_37),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_30),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_68),
.C(n_21),
.Y(n_83)
);

FAx1_ASAP7_75t_SL g64 ( 
.A(n_38),
.B(n_33),
.CI(n_37),
.CON(n_64),
.SN(n_64)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_66),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_38),
.B(n_25),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_47),
.B(n_15),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_69),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_41),
.A2(n_13),
.B(n_14),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_39),
.B(n_36),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_15),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_73),
.B1(n_55),
.B2(n_58),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_22),
.B1(n_36),
.B2(n_14),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_75),
.A2(n_76),
.B1(n_88),
.B2(n_54),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_80),
.B(n_83),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_56),
.A2(n_36),
.B1(n_23),
.B2(n_18),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_93),
.B1(n_98),
.B2(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_87),
.B(n_72),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_91),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_59),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_53),
.B1(n_69),
.B2(n_65),
.Y(n_93)
);

OAI21xp33_ASAP7_75t_L g94 ( 
.A1(n_78),
.A2(n_59),
.B(n_63),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_99),
.C(n_86),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_74),
.A2(n_68),
.B(n_71),
.Y(n_95)
);

OAI22x1_ASAP7_75t_L g103 ( 
.A1(n_95),
.A2(n_64),
.B1(n_76),
.B2(n_61),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_62),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_64),
.C(n_81),
.Y(n_104)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_97),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_82),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_78),
.A2(n_83),
.B(n_77),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_99),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_102),
.A2(n_52),
.B1(n_57),
.B2(n_84),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_103),
.A2(n_89),
.B1(n_93),
.B2(n_51),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_105),
.C(n_24),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_79),
.C(n_81),
.Y(n_105)
);

AOI321xp33_ASAP7_75t_L g115 ( 
.A1(n_108),
.A2(n_111),
.A3(n_107),
.B1(n_21),
.B2(n_12),
.C(n_11),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_96),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_110),
.Y(n_119)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

OAI322xp33_ASAP7_75t_L g111 ( 
.A1(n_106),
.A2(n_104),
.A3(n_107),
.B1(n_91),
.B2(n_79),
.C1(n_95),
.C2(n_97),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_113),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_114),
.B(n_36),
.Y(n_118)
);

AOI31xp67_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_116),
.A3(n_2),
.B(n_4),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_110),
.A2(n_10),
.B(n_1),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_114),
.C(n_108),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_121),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_119),
.B(n_109),
.Y(n_121)
);

AOI322xp5_ASAP7_75t_L g122 ( 
.A1(n_117),
.A2(n_112),
.A3(n_113),
.B1(n_84),
.B2(n_5),
.C1(n_6),
.C2(n_0),
.Y(n_122)
);

AOI31xp33_ASAP7_75t_L g125 ( 
.A1(n_122),
.A2(n_123),
.A3(n_4),
.B(n_6),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_4),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_7),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_124),
.C(n_21),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_125),
.Y(n_129)
);


endmodule