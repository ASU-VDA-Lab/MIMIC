module fake_ariane_1027_n_2394 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_332, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_528, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_550, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_511, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_53, n_260, n_362, n_543, n_310, n_236, n_565, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_546, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_448, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_560, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_555, n_234, n_492, n_280, n_215, n_252, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_540, n_216, n_544, n_5, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_506, n_558, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_127, n_531, n_2394);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_332;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_528;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_511;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_565;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_546;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_555;
input n_234;
input n_492;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_506;
input n_558;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_127;
input n_531;

output n_2394;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_2334;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_690;
wire n_1109;
wire n_1430;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_2376;
wire n_2367;
wire n_1706;
wire n_2207;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_1682;
wire n_1836;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_2248;
wire n_813;
wire n_1985;
wire n_2288;
wire n_995;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_2322;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_2233;
wire n_2370;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_770;
wire n_1514;
wire n_1528;
wire n_901;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_1703;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_661;
wire n_2098;
wire n_1751;
wire n_1917;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_1112;
wire n_1159;
wire n_700;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_652;
wire n_1819;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_696;
wire n_1442;
wire n_798;
wire n_577;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_2185;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_1240;
wire n_1087;
wire n_632;
wire n_650;
wire n_2388;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2294;
wire n_2274;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_2328;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2144;
wire n_1029;
wire n_1247;
wire n_760;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_2262;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_706;
wire n_2120;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2168;
wire n_2312;
wire n_670;
wire n_1826;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_2122;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_600;
wire n_1609;
wire n_1053;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_2195;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_604;
wire n_677;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_727;
wire n_590;
wire n_699;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_1156;
wire n_2184;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_957;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_1005;
wire n_2379;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_2300;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2266;
wire n_890;
wire n_842;
wire n_1898;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_2366;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2211;
wire n_2292;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_2348;
wire n_1281;
wire n_2364;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_726;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_2383;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_2386;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2320;
wire n_979;
wire n_2329;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_802;
wire n_1151;
wire n_960;
wire n_2352;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2314;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2203;
wire n_2133;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_2158;
wire n_2285;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_2173;
wire n_1035;
wire n_1143;
wire n_2070;
wire n_2136;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_1103;
wire n_825;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_2020;
wire n_748;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_1165;
wire n_1641;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2331;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_601;
wire n_683;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2303;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_1814;
wire n_2154;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_692;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1910;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_1785;
wire n_792;
wire n_1262;
wire n_2180;
wire n_1942;
wire n_580;
wire n_1579;
wire n_2181;
wire n_2014;
wire n_975;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2270;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_2251;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2321;
wire n_1077;
wire n_607;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_917;
wire n_1271;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2252;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_1136;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_2097;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_574;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_1967;
wire n_2384;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_1063;
wire n_991;
wire n_2205;
wire n_2183;
wire n_2275;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_2209;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_937;
wire n_1474;
wire n_2081;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_1102;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_1010;
wire n_882;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2336;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_573;
wire n_796;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g570 ( 
.A(n_539),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_194),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_327),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_508),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_119),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_439),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_68),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_514),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_148),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_285),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_425),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_486),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_37),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_214),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_362),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_503),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_207),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_241),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_371),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_465),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_350),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_459),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_129),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_19),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_271),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_104),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_210),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_406),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_448),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_205),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_541),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_281),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_226),
.Y(n_602)
);

INVx1_ASAP7_75t_SL g603 ( 
.A(n_261),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_79),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_229),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_240),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_53),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_197),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_512),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_427),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_446),
.Y(n_611)
);

INVx1_ASAP7_75t_SL g612 ( 
.A(n_82),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_395),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_89),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_369),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_532),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_238),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_401),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_340),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_306),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_550),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_19),
.Y(n_622)
);

CKINVDCx16_ASAP7_75t_R g623 ( 
.A(n_366),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_213),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_231),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_513),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_557),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_566),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_150),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_454),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_561),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_172),
.Y(n_632)
);

BUFx8_ASAP7_75t_SL g633 ( 
.A(n_526),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_126),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_257),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_27),
.Y(n_636)
);

BUFx10_ASAP7_75t_L g637 ( 
.A(n_99),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_417),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_295),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_288),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_182),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_193),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_49),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_156),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_299),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_521),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_154),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_37),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_196),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_83),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_175),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_142),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_564),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_384),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_170),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_286),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_298),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_480),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_543),
.Y(n_659)
);

CKINVDCx16_ASAP7_75t_R g660 ( 
.A(n_98),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_125),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_407),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_298),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_397),
.Y(n_664)
);

BUFx2_ASAP7_75t_L g665 ( 
.A(n_162),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_545),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_510),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_385),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_547),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_429),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_8),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_146),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_116),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_485),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_283),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_221),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_100),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_375),
.Y(n_678)
);

CKINVDCx20_ASAP7_75t_R g679 ( 
.A(n_409),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_260),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_559),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_400),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_499),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_206),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_315),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_445),
.Y(n_686)
);

CKINVDCx20_ASAP7_75t_R g687 ( 
.A(n_299),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_29),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_327),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_173),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_342),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_555),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_92),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_391),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_233),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_31),
.Y(n_696)
);

HB1xp67_ASAP7_75t_L g697 ( 
.A(n_435),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_56),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_419),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_124),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_54),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_471),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_131),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_221),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_383),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_32),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_318),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_519),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_390),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_2),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_490),
.Y(n_711)
);

BUFx10_ASAP7_75t_L g712 ( 
.A(n_540),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_333),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_497),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_536),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_529),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_418),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_405),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_236),
.Y(n_719)
);

BUFx10_ASAP7_75t_L g720 ( 
.A(n_292),
.Y(n_720)
);

BUFx2_ASAP7_75t_L g721 ( 
.A(n_38),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_356),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_48),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_267),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_352),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_171),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_213),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_556),
.Y(n_728)
);

INVx1_ASAP7_75t_SL g729 ( 
.A(n_248),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_132),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_10),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_306),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_472),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_354),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_433),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_8),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_533),
.Y(n_737)
);

HB1xp67_ASAP7_75t_L g738 ( 
.A(n_387),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_247),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_300),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_20),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_204),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_225),
.Y(n_743)
);

CKINVDCx20_ASAP7_75t_R g744 ( 
.A(n_452),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_76),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_41),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_5),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_468),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_25),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_558),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_334),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_127),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_370),
.Y(n_753)
);

CKINVDCx14_ASAP7_75t_R g754 ( 
.A(n_361),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_202),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_246),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_220),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_31),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_143),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_531),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_542),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_202),
.Y(n_762)
);

CKINVDCx20_ASAP7_75t_R g763 ( 
.A(n_462),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_426),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_262),
.Y(n_765)
);

BUFx2_ASAP7_75t_L g766 ( 
.A(n_276),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_235),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_100),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_159),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_365),
.Y(n_770)
);

BUFx8_ASAP7_75t_SL g771 ( 
.A(n_175),
.Y(n_771)
);

INVx1_ASAP7_75t_SL g772 ( 
.A(n_222),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_61),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_272),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_422),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_256),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_211),
.Y(n_777)
);

BUFx10_ASAP7_75t_L g778 ( 
.A(n_368),
.Y(n_778)
);

CKINVDCx14_ASAP7_75t_R g779 ( 
.A(n_378),
.Y(n_779)
);

CKINVDCx20_ASAP7_75t_R g780 ( 
.A(n_88),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_552),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_197),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_82),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_515),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_174),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_267),
.Y(n_786)
);

CKINVDCx16_ASAP7_75t_R g787 ( 
.A(n_377),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_191),
.Y(n_788)
);

CKINVDCx20_ASAP7_75t_R g789 ( 
.A(n_436),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_269),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_582),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_582),
.Y(n_792)
);

INVxp67_ASAP7_75t_SL g793 ( 
.A(n_690),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_690),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_727),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_771),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_632),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_727),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_610),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_771),
.Y(n_800)
);

CKINVDCx20_ASAP7_75t_R g801 ( 
.A(n_576),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_572),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_578),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_579),
.Y(n_804)
);

CKINVDCx20_ASAP7_75t_R g805 ( 
.A(n_576),
.Y(n_805)
);

INVxp33_ASAP7_75t_SL g806 ( 
.A(n_710),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_587),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_666),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_596),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_592),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_623),
.Y(n_811)
);

INVxp67_ASAP7_75t_L g812 ( 
.A(n_665),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_787),
.Y(n_813)
);

INVxp67_ASAP7_75t_SL g814 ( 
.A(n_632),
.Y(n_814)
);

BUFx2_ASAP7_75t_L g815 ( 
.A(n_721),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_632),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_593),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_633),
.Y(n_818)
);

BUFx3_ASAP7_75t_L g819 ( 
.A(n_666),
.Y(n_819)
);

INVxp33_ASAP7_75t_SL g820 ( 
.A(n_697),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_595),
.Y(n_821)
);

INVx4_ASAP7_75t_R g822 ( 
.A(n_692),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_605),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_632),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_619),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_634),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_639),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_640),
.Y(n_828)
);

INVx1_ASAP7_75t_SL g829 ( 
.A(n_596),
.Y(n_829)
);

INVxp33_ASAP7_75t_L g830 ( 
.A(n_766),
.Y(n_830)
);

CKINVDCx20_ASAP7_75t_R g831 ( 
.A(n_601),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_641),
.Y(n_832)
);

CKINVDCx16_ASAP7_75t_R g833 ( 
.A(n_660),
.Y(n_833)
);

INVxp33_ASAP7_75t_SL g834 ( 
.A(n_738),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_642),
.Y(n_835)
);

NOR2xp67_ASAP7_75t_L g836 ( 
.A(n_602),
.B(n_0),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_692),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_633),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_672),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_573),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_601),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_608),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_573),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_673),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_597),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_597),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_684),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_688),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_698),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_701),
.Y(n_850)
);

CKINVDCx20_ASAP7_75t_R g851 ( 
.A(n_608),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_703),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_704),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_719),
.Y(n_854)
);

INVxp33_ASAP7_75t_L g855 ( 
.A(n_723),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_732),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_740),
.Y(n_857)
);

OR2x2_ASAP7_75t_L g858 ( 
.A(n_583),
.B(n_0),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_741),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_610),
.Y(n_860)
);

CKINVDCx16_ASAP7_75t_R g861 ( 
.A(n_637),
.Y(n_861)
);

INVxp33_ASAP7_75t_L g862 ( 
.A(n_742),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_743),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_602),
.B(n_1),
.Y(n_864)
);

INVxp67_ASAP7_75t_SL g865 ( 
.A(n_583),
.Y(n_865)
);

CKINVDCx14_ASAP7_75t_R g866 ( 
.A(n_754),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_746),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_747),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_735),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_757),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_765),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_774),
.Y(n_872)
);

INVxp67_ASAP7_75t_SL g873 ( 
.A(n_614),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_735),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_570),
.Y(n_875)
);

INVxp67_ASAP7_75t_SL g876 ( 
.A(n_614),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_783),
.Y(n_877)
);

INVxp33_ASAP7_75t_SL g878 ( 
.A(n_574),
.Y(n_878)
);

INVxp33_ASAP7_75t_SL g879 ( 
.A(n_574),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_786),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_788),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_575),
.Y(n_882)
);

CKINVDCx14_ASAP7_75t_R g883 ( 
.A(n_779),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_659),
.Y(n_884)
);

INVxp67_ASAP7_75t_SL g885 ( 
.A(n_649),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_649),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_661),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_661),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_663),
.Y(n_889)
);

OAI22xp5_ASAP7_75t_R g890 ( 
.A1(n_840),
.A2(n_687),
.B1(n_780),
.B2(n_617),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_829),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_816),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_797),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_799),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_799),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_796),
.Y(n_896)
);

CKINVDCx6p67_ASAP7_75t_R g897 ( 
.A(n_833),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_816),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_811),
.B(n_712),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_797),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_799),
.Y(n_901)
);

OR2x2_ASAP7_75t_L g902 ( 
.A(n_815),
.B(n_571),
.Y(n_902)
);

BUFx12f_ASAP7_75t_L g903 ( 
.A(n_818),
.Y(n_903)
);

HB1xp67_ASAP7_75t_L g904 ( 
.A(n_796),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_793),
.B(n_590),
.Y(n_905)
);

BUFx8_ASAP7_75t_SL g906 ( 
.A(n_801),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_824),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_824),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_820),
.A2(n_687),
.B1(n_780),
.B2(n_617),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_799),
.Y(n_910)
);

BUFx8_ASAP7_75t_SL g911 ( 
.A(n_801),
.Y(n_911)
);

BUFx8_ASAP7_75t_L g912 ( 
.A(n_837),
.Y(n_912)
);

BUFx2_ASAP7_75t_L g913 ( 
.A(n_818),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_797),
.Y(n_914)
);

AOI22x1_ASAP7_75t_SL g915 ( 
.A1(n_805),
.A2(n_594),
.B1(n_604),
.B2(n_599),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_865),
.B(n_637),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_814),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_808),
.B(n_675),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_L g919 ( 
.A1(n_820),
.A2(n_834),
.B1(n_806),
.B2(n_812),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_875),
.Y(n_920)
);

INVx4_ASAP7_75t_L g921 ( 
.A(n_799),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_875),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_860),
.Y(n_923)
);

BUFx6f_ASAP7_75t_L g924 ( 
.A(n_860),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_808),
.B(n_675),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_860),
.Y(n_926)
);

BUFx3_ASAP7_75t_L g927 ( 
.A(n_819),
.Y(n_927)
);

OAI22xp5_ASAP7_75t_L g928 ( 
.A1(n_834),
.A2(n_612),
.B1(n_729),
.B2(n_603),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_860),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_882),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_860),
.Y(n_931)
);

AOI22xp5_ASAP7_75t_L g932 ( 
.A1(n_806),
.A2(n_879),
.B1(n_878),
.B2(n_679),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_882),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_878),
.A2(n_679),
.B1(n_744),
.B2(n_659),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_837),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_869),
.Y(n_936)
);

BUFx6f_ASAP7_75t_L g937 ( 
.A(n_869),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_819),
.B(n_696),
.Y(n_938)
);

INVx5_ASAP7_75t_L g939 ( 
.A(n_874),
.Y(n_939)
);

OAI21x1_ASAP7_75t_L g940 ( 
.A1(n_791),
.A2(n_598),
.B(n_591),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_886),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_887),
.Y(n_942)
);

BUFx3_ASAP7_75t_L g943 ( 
.A(n_874),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_888),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_889),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_802),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_803),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_866),
.Y(n_948)
);

HB1xp67_ASAP7_75t_L g949 ( 
.A(n_800),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_804),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_883),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_800),
.Y(n_952)
);

INVxp67_ASAP7_75t_L g953 ( 
.A(n_838),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_792),
.B(n_600),
.Y(n_954)
);

AND2x4_ASAP7_75t_L g955 ( 
.A(n_927),
.B(n_873),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_947),
.Y(n_956)
);

CKINVDCx20_ASAP7_75t_R g957 ( 
.A(n_906),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_R g958 ( 
.A(n_948),
.B(n_838),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_947),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_927),
.B(n_876),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_917),
.B(n_811),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_914),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_903),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_917),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_916),
.B(n_813),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_946),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_903),
.Y(n_967)
);

NOR2x1_ASAP7_75t_L g968 ( 
.A(n_943),
.B(n_744),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_946),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_950),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_916),
.B(n_943),
.Y(n_971)
);

CKINVDCx20_ASAP7_75t_R g972 ( 
.A(n_911),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_948),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_891),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_914),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_936),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_950),
.Y(n_977)
);

HB1xp67_ASAP7_75t_L g978 ( 
.A(n_902),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_951),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_921),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_935),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_936),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_935),
.B(n_813),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_941),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_951),
.Y(n_985)
);

INVxp67_ASAP7_75t_L g986 ( 
.A(n_902),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_897),
.Y(n_987)
);

CKINVDCx20_ASAP7_75t_R g988 ( 
.A(n_934),
.Y(n_988)
);

HB1xp67_ASAP7_75t_L g989 ( 
.A(n_909),
.Y(n_989)
);

CKINVDCx20_ASAP7_75t_R g990 ( 
.A(n_934),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_941),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_893),
.B(n_864),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_918),
.B(n_879),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_918),
.B(n_861),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_944),
.Y(n_995)
);

CKINVDCx16_ASAP7_75t_R g996 ( 
.A(n_932),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_918),
.B(n_925),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_897),
.Y(n_998)
);

BUFx3_ASAP7_75t_L g999 ( 
.A(n_936),
.Y(n_999)
);

CKINVDCx16_ASAP7_75t_R g1000 ( 
.A(n_932),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_R g1001 ( 
.A(n_913),
.B(n_840),
.Y(n_1001)
);

HB1xp67_ASAP7_75t_L g1002 ( 
.A(n_913),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_936),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_936),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_890),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_890),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_937),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_896),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_904),
.Y(n_1009)
);

AND2x4_ASAP7_75t_L g1010 ( 
.A(n_918),
.B(n_885),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_949),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_944),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_893),
.B(n_794),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_925),
.B(n_836),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_952),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_893),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_900),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_953),
.Y(n_1018)
);

CKINVDCx20_ASAP7_75t_R g1019 ( 
.A(n_919),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_925),
.B(n_830),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_937),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_900),
.B(n_795),
.Y(n_1022)
);

INVxp67_ASAP7_75t_L g1023 ( 
.A(n_925),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_938),
.B(n_588),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_921),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_915),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_921),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_938),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_900),
.B(n_912),
.Y(n_1029)
);

CKINVDCx20_ASAP7_75t_R g1030 ( 
.A(n_915),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_937),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_899),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_937),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_937),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_928),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_912),
.Y(n_1036)
);

OA21x2_ASAP7_75t_L g1037 ( 
.A1(n_940),
.A2(n_669),
.B(n_638),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_938),
.B(n_855),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_912),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_912),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_962),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_965),
.B(n_939),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_971),
.B(n_983),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_962),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_997),
.B(n_939),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_975),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_975),
.Y(n_1047)
);

AOI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_961),
.A2(n_789),
.B1(n_763),
.B2(n_748),
.Y(n_1048)
);

HB1xp67_ASAP7_75t_L g1049 ( 
.A(n_974),
.Y(n_1049)
);

INVxp67_ASAP7_75t_SL g1050 ( 
.A(n_980),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_980),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_964),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_981),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_997),
.B(n_939),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_1016),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_966),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_997),
.B(n_938),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1017),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_969),
.Y(n_1059)
);

OR2x6_ASAP7_75t_L g1060 ( 
.A(n_986),
.B(n_858),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_976),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_970),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_976),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_992),
.A2(n_940),
.B(n_905),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_982),
.Y(n_1065)
);

INVx4_ASAP7_75t_L g1066 ( 
.A(n_1036),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_977),
.Y(n_1067)
);

NAND3xp33_ASAP7_75t_L g1068 ( 
.A(n_1018),
.B(n_845),
.C(n_843),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_L g1069 ( 
.A1(n_989),
.A2(n_858),
.B1(n_930),
.B2(n_920),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_1010),
.B(n_922),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_SL g1071 ( 
.A(n_955),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_982),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1010),
.B(n_922),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_984),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_991),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_1004),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_1004),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_1021),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_995),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_993),
.B(n_748),
.Y(n_1080)
);

BUFx10_ASAP7_75t_L g1081 ( 
.A(n_979),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_1023),
.B(n_763),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_980),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1021),
.Y(n_1084)
);

INVx8_ASAP7_75t_L g1085 ( 
.A(n_987),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_956),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1012),
.Y(n_1087)
);

NAND3xp33_ASAP7_75t_L g1088 ( 
.A(n_1018),
.B(n_845),
.C(n_843),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_959),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1010),
.B(n_922),
.Y(n_1090)
);

AND3x2_ASAP7_75t_L g1091 ( 
.A(n_978),
.B(n_809),
.C(n_805),
.Y(n_1091)
);

INVx2_ASAP7_75t_SL g1092 ( 
.A(n_1038),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1013),
.Y(n_1093)
);

AO21x2_ASAP7_75t_L g1094 ( 
.A1(n_1033),
.A2(n_611),
.B(n_609),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1022),
.Y(n_1095)
);

INVxp67_ASAP7_75t_SL g1096 ( 
.A(n_1025),
.Y(n_1096)
);

BUFx2_ASAP7_75t_L g1097 ( 
.A(n_1001),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_1025),
.B(n_939),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_955),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_1028),
.B(n_789),
.Y(n_1100)
);

NOR3xp33_ASAP7_75t_L g1101 ( 
.A(n_996),
.B(n_884),
.C(n_846),
.Y(n_1101)
);

AND3x2_ASAP7_75t_L g1102 ( 
.A(n_1002),
.B(n_831),
.C(n_809),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_1025),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_1020),
.B(n_846),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1034),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_955),
.B(n_920),
.Y(n_1106)
);

AND2x6_ASAP7_75t_L g1107 ( 
.A(n_968),
.B(n_638),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_1027),
.B(n_939),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_1035),
.A2(n_930),
.B1(n_933),
.B2(n_862),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_960),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_1008),
.B(n_884),
.Y(n_1111)
);

INVx3_ASAP7_75t_L g1112 ( 
.A(n_1027),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_985),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1007),
.Y(n_1114)
);

AND2x6_ASAP7_75t_L g1115 ( 
.A(n_1029),
.B(n_669),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_1019),
.A2(n_933),
.B1(n_945),
.B2(n_942),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1007),
.Y(n_1117)
);

OR2x6_ASAP7_75t_L g1118 ( 
.A(n_994),
.B(n_954),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_960),
.Y(n_1119)
);

AOI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_1014),
.A2(n_715),
.B1(n_589),
.B2(n_588),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_1027),
.B(n_939),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1007),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_960),
.Y(n_1123)
);

NAND3xp33_ASAP7_75t_L g1124 ( 
.A(n_1008),
.B(n_599),
.C(n_594),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1007),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_999),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_999),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_1007),
.B(n_589),
.Y(n_1128)
);

INVx3_ASAP7_75t_L g1129 ( 
.A(n_1003),
.Y(n_1129)
);

BUFx3_ASAP7_75t_L g1130 ( 
.A(n_1003),
.Y(n_1130)
);

CKINVDCx20_ASAP7_75t_R g1131 ( 
.A(n_1000),
.Y(n_1131)
);

INVxp67_ASAP7_75t_SL g1132 ( 
.A(n_1031),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1031),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_1032),
.B(n_770),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1024),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_1036),
.B(n_770),
.Y(n_1136)
);

INVx2_ASAP7_75t_SL g1137 ( 
.A(n_1009),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1037),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1039),
.B(n_1040),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1037),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1037),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1039),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1040),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1009),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_987),
.Y(n_1145)
);

INVx4_ASAP7_75t_L g1146 ( 
.A(n_998),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1011),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1011),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1015),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_1015),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_973),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_973),
.B(n_958),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1019),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_988),
.B(n_942),
.Y(n_1154)
);

AND2x6_ASAP7_75t_L g1155 ( 
.A(n_963),
.B(n_683),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_963),
.B(n_942),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_967),
.B(n_942),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_988),
.A2(n_945),
.B1(n_942),
.B2(n_790),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_990),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_967),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_990),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1026),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1005),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1030),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_1006),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1006),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_957),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_L g1168 ( 
.A1(n_1030),
.A2(n_945),
.B1(n_790),
.B2(n_696),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_957),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_972),
.Y(n_1170)
);

NAND3xp33_ASAP7_75t_L g1171 ( 
.A(n_972),
.B(n_680),
.C(n_604),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_962),
.Y(n_1172)
);

INVx1_ASAP7_75t_SL g1173 ( 
.A(n_974),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_962),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_962),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_980),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_1148),
.B(n_775),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_1148),
.B(n_775),
.Y(n_1178)
);

BUFx8_ASAP7_75t_L g1179 ( 
.A(n_1097),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1043),
.B(n_945),
.Y(n_1180)
);

NAND2xp33_ASAP7_75t_L g1181 ( 
.A(n_1051),
.B(n_680),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1070),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_1100),
.B(n_831),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1043),
.B(n_945),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1070),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_1100),
.B(n_841),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1093),
.B(n_892),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_1048),
.B(n_841),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1095),
.B(n_892),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1052),
.B(n_898),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_1113),
.Y(n_1191)
);

INVx2_ASAP7_75t_SL g1192 ( 
.A(n_1173),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1056),
.B(n_1059),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1062),
.B(n_898),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1067),
.B(n_907),
.Y(n_1195)
);

AO221x1_ASAP7_75t_L g1196 ( 
.A1(n_1145),
.A2(n_663),
.B1(n_736),
.B2(n_691),
.C(n_676),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1074),
.B(n_907),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1070),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1099),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1075),
.B(n_908),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1110),
.B(n_772),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1119),
.B(n_1123),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_L g1203 ( 
.A(n_1080),
.B(n_842),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1069),
.B(n_773),
.Y(n_1204)
);

INVxp33_ASAP7_75t_L g1205 ( 
.A(n_1111),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_1080),
.B(n_842),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1060),
.B(n_851),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1082),
.B(n_851),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1073),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1069),
.B(n_773),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1082),
.B(n_776),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_1149),
.B(n_776),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1061),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1106),
.B(n_777),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1061),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_1149),
.B(n_777),
.Y(n_1216)
);

NAND3xp33_ASAP7_75t_L g1217 ( 
.A(n_1144),
.B(n_785),
.C(n_635),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1090),
.B(n_785),
.Y(n_1218)
);

OAI21xp33_ASAP7_75t_L g1219 ( 
.A1(n_1137),
.A2(n_636),
.B(n_624),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1079),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_1150),
.B(n_586),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1150),
.B(n_606),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1060),
.B(n_1104),
.Y(n_1223)
);

INVxp67_ASAP7_75t_L g1224 ( 
.A(n_1049),
.Y(n_1224)
);

XOR2xp5_ASAP7_75t_L g1225 ( 
.A(n_1113),
.B(n_798),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1087),
.B(n_908),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_SL g1227 ( 
.A(n_1057),
.B(n_1147),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_1130),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1063),
.Y(n_1229)
);

OR2x6_ASAP7_75t_L g1230 ( 
.A(n_1085),
.B(n_823),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1109),
.B(n_676),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1109),
.B(n_1057),
.Y(n_1232)
);

HB1xp67_ASAP7_75t_L g1233 ( 
.A(n_1071),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1063),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1060),
.B(n_1153),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_1151),
.B(n_607),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1041),
.Y(n_1237)
);

BUFx5_ASAP7_75t_L g1238 ( 
.A(n_1141),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_SL g1239 ( 
.A(n_1057),
.B(n_620),
.Y(n_1239)
);

NOR2xp67_ASAP7_75t_L g1240 ( 
.A(n_1146),
.B(n_807),
.Y(n_1240)
);

INVx2_ASAP7_75t_SL g1241 ( 
.A(n_1081),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1065),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1139),
.B(n_622),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1154),
.B(n_810),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1044),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1154),
.B(n_691),
.Y(n_1246)
);

OR2x6_ASAP7_75t_L g1247 ( 
.A(n_1085),
.B(n_872),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1086),
.B(n_1046),
.Y(n_1248)
);

NAND3xp33_ASAP7_75t_L g1249 ( 
.A(n_1068),
.B(n_657),
.C(n_648),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1065),
.Y(n_1250)
);

NOR2x1p5_ASAP7_75t_L g1251 ( 
.A(n_1146),
.B(n_1167),
.Y(n_1251)
);

NOR3xp33_ASAP7_75t_L g1252 ( 
.A(n_1088),
.B(n_1152),
.C(n_1171),
.Y(n_1252)
);

INVxp67_ASAP7_75t_L g1253 ( 
.A(n_1071),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1047),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_SL g1255 ( 
.A(n_1066),
.B(n_625),
.Y(n_1255)
);

OR2x2_ASAP7_75t_L g1256 ( 
.A(n_1159),
.B(n_817),
.Y(n_1256)
);

BUFx8_ASAP7_75t_L g1257 ( 
.A(n_1160),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1172),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1174),
.Y(n_1259)
);

HB1xp67_ASAP7_75t_L g1260 ( 
.A(n_1092),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_SL g1261 ( 
.A(n_1066),
.B(n_629),
.Y(n_1261)
);

NOR3xp33_ASAP7_75t_L g1262 ( 
.A(n_1152),
.B(n_1136),
.C(n_1124),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1086),
.B(n_1175),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1134),
.B(n_643),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1072),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1055),
.B(n_616),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_1134),
.B(n_644),
.Y(n_1267)
);

NOR3xp33_ASAP7_75t_L g1268 ( 
.A(n_1136),
.B(n_647),
.C(n_645),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1072),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_L g1270 ( 
.A(n_1130),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_SL g1271 ( 
.A(n_1160),
.B(n_650),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1053),
.Y(n_1272)
);

AO221x1_ASAP7_75t_L g1273 ( 
.A1(n_1145),
.A2(n_782),
.B1(n_736),
.B2(n_722),
.C(n_615),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1076),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1116),
.A2(n_712),
.B1(n_778),
.B2(n_720),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1159),
.B(n_821),
.Y(n_1276)
);

AOI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1118),
.A2(n_715),
.B1(n_631),
.B2(n_646),
.Y(n_1277)
);

INVx1_ASAP7_75t_SL g1278 ( 
.A(n_1161),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1053),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1089),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1129),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1116),
.B(n_782),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1076),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1155),
.B(n_651),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1077),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_1142),
.B(n_652),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1055),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1077),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1078),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_L g1290 ( 
.A(n_1142),
.B(n_655),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1078),
.Y(n_1291)
);

CKINVDCx20_ASAP7_75t_R g1292 ( 
.A(n_1085),
.Y(n_1292)
);

BUFx6f_ASAP7_75t_L g1293 ( 
.A(n_1129),
.Y(n_1293)
);

INVxp67_ASAP7_75t_L g1294 ( 
.A(n_1160),
.Y(n_1294)
);

INVxp67_ASAP7_75t_L g1295 ( 
.A(n_1160),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1058),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1133),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1155),
.B(n_656),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1155),
.B(n_671),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1084),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_SL g1301 ( 
.A(n_1145),
.B(n_677),
.Y(n_1301)
);

INVxp67_ASAP7_75t_L g1302 ( 
.A(n_1118),
.Y(n_1302)
);

NAND2xp33_ASAP7_75t_L g1303 ( 
.A(n_1051),
.B(n_685),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1058),
.B(n_618),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1064),
.B(n_653),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1083),
.B(n_654),
.Y(n_1306)
);

BUFx6f_ASAP7_75t_L g1307 ( 
.A(n_1133),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_SL g1308 ( 
.A(n_1145),
.B(n_689),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1105),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1105),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_1143),
.B(n_693),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1155),
.B(n_695),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1084),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1155),
.B(n_700),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1135),
.B(n_706),
.Y(n_1315)
);

A2O1A1Ixp33_ASAP7_75t_L g1316 ( 
.A1(n_1083),
.A2(n_668),
.B(n_670),
.C(n_662),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_SL g1317 ( 
.A(n_1081),
.B(n_707),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1126),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1114),
.Y(n_1319)
);

INVxp33_ASAP7_75t_SL g1320 ( 
.A(n_1170),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1050),
.B(n_713),
.Y(n_1321)
);

NOR2xp33_ASAP7_75t_L g1322 ( 
.A(n_1118),
.B(n_724),
.Y(n_1322)
);

INVx2_ASAP7_75t_SL g1323 ( 
.A(n_1081),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1127),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1114),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1103),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_SL g1327 ( 
.A(n_1156),
.B(n_726),
.Y(n_1327)
);

NAND3xp33_ASAP7_75t_L g1328 ( 
.A(n_1120),
.B(n_751),
.C(n_731),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1096),
.B(n_730),
.Y(n_1329)
);

AOI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1098),
.A2(n_1121),
.B(n_1108),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1117),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1158),
.B(n_1107),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1168),
.B(n_825),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_L g1334 ( 
.A(n_1157),
.B(n_739),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_1103),
.B(n_745),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_SL g1336 ( 
.A(n_1112),
.B(n_749),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1112),
.B(n_1176),
.Y(n_1337)
);

NAND3xp33_ASAP7_75t_L g1338 ( 
.A(n_1128),
.B(n_759),
.C(n_755),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1158),
.B(n_752),
.Y(n_1339)
);

BUFx3_ASAP7_75t_L g1340 ( 
.A(n_1131),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1176),
.B(n_686),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1107),
.B(n_709),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1117),
.Y(n_1343)
);

NAND3xp33_ASAP7_75t_L g1344 ( 
.A(n_1128),
.B(n_767),
.C(n_758),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_L g1345 ( 
.A(n_1170),
.B(n_756),
.Y(n_1345)
);

AO221x1_ASAP7_75t_L g1346 ( 
.A1(n_1165),
.A2(n_722),
.B1(n_615),
.B2(n_610),
.C(n_714),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1122),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_1102),
.B(n_762),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1122),
.Y(n_1349)
);

NOR2xp67_ASAP7_75t_L g1350 ( 
.A(n_1162),
.B(n_826),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1125),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1125),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1131),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1138),
.Y(n_1354)
);

AO221x1_ASAP7_75t_L g1355 ( 
.A1(n_1165),
.A2(n_1166),
.B1(n_1163),
.B2(n_1169),
.C(n_1168),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1107),
.B(n_711),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_SL g1357 ( 
.A(n_1132),
.B(n_1101),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1045),
.B(n_768),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1107),
.B(n_718),
.Y(n_1359)
);

NAND2xp33_ASAP7_75t_L g1360 ( 
.A(n_1115),
.B(n_769),
.Y(n_1360)
);

AND2x4_ASAP7_75t_L g1361 ( 
.A(n_1045),
.B(n_827),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1107),
.B(n_764),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1138),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_SL g1364 ( 
.A(n_1054),
.B(n_712),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1042),
.B(n_781),
.Y(n_1365)
);

NAND2xp33_ASAP7_75t_R g1366 ( 
.A(n_1091),
.B(n_822),
.Y(n_1366)
);

INVxp67_ASAP7_75t_L g1367 ( 
.A(n_1164),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1042),
.B(n_683),
.Y(n_1368)
);

INVx2_ASAP7_75t_SL g1369 ( 
.A(n_1164),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1140),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1054),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1140),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1094),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_SL g1374 ( 
.A(n_1098),
.B(n_778),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1094),
.Y(n_1375)
);

INVxp67_ASAP7_75t_L g1376 ( 
.A(n_1192),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_SL g1377 ( 
.A(n_1278),
.B(n_637),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1220),
.Y(n_1378)
);

INVx2_ASAP7_75t_SL g1379 ( 
.A(n_1257),
.Y(n_1379)
);

NAND2x1p5_ASAP7_75t_L g1380 ( 
.A(n_1228),
.B(n_1108),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_SL g1381 ( 
.A(n_1278),
.B(n_720),
.Y(n_1381)
);

AO22x2_ASAP7_75t_L g1382 ( 
.A1(n_1373),
.A2(n_832),
.B1(n_835),
.B2(n_828),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1193),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1244),
.B(n_1115),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1188),
.A2(n_1206),
.B1(n_1203),
.B2(n_1208),
.Y(n_1385)
);

AO22x2_ASAP7_75t_L g1386 ( 
.A1(n_1375),
.A2(n_844),
.B1(n_847),
.B2(n_839),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1211),
.B(n_1115),
.Y(n_1387)
);

BUFx6f_ASAP7_75t_SL g1388 ( 
.A(n_1340),
.Y(n_1388)
);

INVx4_ASAP7_75t_L g1389 ( 
.A(n_1191),
.Y(n_1389)
);

AO22x2_ASAP7_75t_L g1390 ( 
.A1(n_1207),
.A2(n_849),
.B1(n_850),
.B2(n_848),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1257),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1193),
.Y(n_1392)
);

AO22x2_ASAP7_75t_L g1393 ( 
.A1(n_1332),
.A2(n_853),
.B1(n_854),
.B2(n_852),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1213),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1215),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1229),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1232),
.B(n_1115),
.Y(n_1397)
);

AO22x2_ASAP7_75t_L g1398 ( 
.A1(n_1231),
.A2(n_857),
.B1(n_859),
.B2(n_856),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1234),
.Y(n_1399)
);

OAI221xp5_ASAP7_75t_L g1400 ( 
.A1(n_1183),
.A2(n_868),
.B1(n_870),
.B2(n_867),
.C(n_863),
.Y(n_1400)
);

AO22x2_ASAP7_75t_L g1401 ( 
.A1(n_1333),
.A2(n_877),
.B1(n_880),
.B2(n_871),
.Y(n_1401)
);

BUFx3_ASAP7_75t_L g1402 ( 
.A(n_1179),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1242),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1230),
.B(n_881),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1280),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1186),
.B(n_720),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1199),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1237),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1245),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1254),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1276),
.B(n_1115),
.Y(n_1411)
);

NOR2xp67_ASAP7_75t_L g1412 ( 
.A(n_1241),
.B(n_1121),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1258),
.Y(n_1413)
);

AO22x2_ASAP7_75t_L g1414 ( 
.A1(n_1235),
.A2(n_784),
.B1(n_734),
.B2(n_778),
.Y(n_1414)
);

NAND2x1p5_ASAP7_75t_L g1415 ( 
.A(n_1228),
.B(n_910),
.Y(n_1415)
);

AO22x2_ASAP7_75t_L g1416 ( 
.A1(n_1342),
.A2(n_784),
.B1(n_734),
.B2(n_3),
.Y(n_1416)
);

AO22x2_ASAP7_75t_L g1417 ( 
.A1(n_1342),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1250),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1259),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1272),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1209),
.B(n_4),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1279),
.Y(n_1422)
);

AO22x2_ASAP7_75t_L g1423 ( 
.A1(n_1356),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_1423)
);

AO22x2_ASAP7_75t_L g1424 ( 
.A1(n_1356),
.A2(n_1362),
.B1(n_1359),
.B2(n_1210),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1243),
.B(n_6),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1287),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1334),
.B(n_7),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1296),
.Y(n_1428)
);

AO22x2_ASAP7_75t_L g1429 ( 
.A1(n_1359),
.A2(n_10),
.B1(n_7),
.B2(n_9),
.Y(n_1429)
);

OAI221xp5_ASAP7_75t_L g1430 ( 
.A1(n_1322),
.A2(n_581),
.B1(n_584),
.B2(n_580),
.C(n_577),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1309),
.Y(n_1431)
);

AO22x2_ASAP7_75t_L g1432 ( 
.A1(n_1362),
.A2(n_12),
.B1(n_9),
.B2(n_11),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1310),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1361),
.B(n_11),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1202),
.Y(n_1435)
);

NAND2x1p5_ASAP7_75t_L g1436 ( 
.A(n_1228),
.B(n_910),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1223),
.B(n_1205),
.Y(n_1437)
);

AO22x2_ASAP7_75t_L g1438 ( 
.A1(n_1204),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1320),
.B(n_585),
.Y(n_1439)
);

AND2x6_ASAP7_75t_L g1440 ( 
.A(n_1182),
.B(n_610),
.Y(n_1440)
);

AOI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1264),
.A2(n_621),
.B1(n_626),
.B2(n_613),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1361),
.B(n_13),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1248),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1185),
.B(n_14),
.Y(n_1444)
);

A2O1A1Ixp33_ASAP7_75t_L g1445 ( 
.A1(n_1267),
.A2(n_926),
.B(n_929),
.C(n_923),
.Y(n_1445)
);

NAND2x1p5_ASAP7_75t_L g1446 ( 
.A(n_1270),
.B(n_923),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1224),
.B(n_1230),
.Y(n_1447)
);

AO22x2_ASAP7_75t_L g1448 ( 
.A1(n_1367),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_SL g1449 ( 
.A(n_1270),
.B(n_627),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_L g1450 ( 
.A(n_1302),
.B(n_628),
.Y(n_1450)
);

INVx3_ASAP7_75t_L g1451 ( 
.A(n_1179),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1248),
.Y(n_1452)
);

AOI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1262),
.A2(n_630),
.B1(n_664),
.B2(n_658),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_1292),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1230),
.B(n_15),
.Y(n_1455)
);

BUFx6f_ASAP7_75t_L g1456 ( 
.A(n_1270),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_1366),
.Y(n_1457)
);

NAND2xp33_ASAP7_75t_SL g1458 ( 
.A(n_1323),
.B(n_667),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1247),
.B(n_16),
.Y(n_1459)
);

AOI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1286),
.A2(n_674),
.B1(n_681),
.B2(n_678),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1263),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_1247),
.Y(n_1462)
);

INVxp67_ASAP7_75t_L g1463 ( 
.A(n_1260),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1263),
.Y(n_1464)
);

BUFx3_ASAP7_75t_L g1465 ( 
.A(n_1353),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1265),
.Y(n_1466)
);

AO22x2_ASAP7_75t_L g1467 ( 
.A1(n_1225),
.A2(n_20),
.B1(n_17),
.B2(n_18),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1269),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1190),
.Y(n_1469)
);

NAND2x1p5_ASAP7_75t_L g1470 ( 
.A(n_1198),
.B(n_926),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1214),
.B(n_18),
.Y(n_1471)
);

AO22x2_ASAP7_75t_L g1472 ( 
.A1(n_1369),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_1472)
);

AO22x2_ASAP7_75t_L g1473 ( 
.A1(n_1339),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_1473)
);

AO22x2_ASAP7_75t_L g1474 ( 
.A1(n_1282),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_1474)
);

AO22x2_ASAP7_75t_L g1475 ( 
.A1(n_1256),
.A2(n_27),
.B1(n_24),
.B2(n_26),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1190),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1221),
.B(n_28),
.Y(n_1477)
);

AO22x2_ASAP7_75t_L g1478 ( 
.A1(n_1305),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_1478)
);

NOR2xp67_ASAP7_75t_L g1479 ( 
.A(n_1294),
.B(n_682),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1222),
.B(n_30),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1212),
.B(n_32),
.Y(n_1481)
);

NAND2x1p5_ASAP7_75t_L g1482 ( 
.A(n_1251),
.B(n_929),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1194),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1274),
.Y(n_1484)
);

OR2x6_ASAP7_75t_L g1485 ( 
.A(n_1247),
.B(n_615),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_R g1486 ( 
.A(n_1303),
.B(n_694),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1283),
.Y(n_1487)
);

AOI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1290),
.A2(n_699),
.B1(n_705),
.B2(n_702),
.Y(n_1488)
);

OAI221xp5_ASAP7_75t_L g1489 ( 
.A1(n_1216),
.A2(n_716),
.B1(n_725),
.B2(n_717),
.C(n_708),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1246),
.B(n_33),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1194),
.Y(n_1491)
);

AO22x2_ASAP7_75t_L g1492 ( 
.A1(n_1305),
.A2(n_1324),
.B1(n_1318),
.B2(n_1371),
.Y(n_1492)
);

BUFx8_ASAP7_75t_L g1493 ( 
.A(n_1281),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1195),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1218),
.B(n_33),
.Y(n_1495)
);

AND2x2_ASAP7_75t_SL g1496 ( 
.A(n_1275),
.B(n_615),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1195),
.Y(n_1497)
);

OAI221xp5_ASAP7_75t_L g1498 ( 
.A1(n_1277),
.A2(n_733),
.B1(n_750),
.B2(n_737),
.C(n_728),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1285),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1197),
.Y(n_1500)
);

INVx2_ASAP7_75t_SL g1501 ( 
.A(n_1233),
.Y(n_1501)
);

BUFx2_ASAP7_75t_L g1502 ( 
.A(n_1253),
.Y(n_1502)
);

OAI221xp5_ASAP7_75t_L g1503 ( 
.A1(n_1236),
.A2(n_760),
.B1(n_761),
.B2(n_753),
.C(n_722),
.Y(n_1503)
);

NAND2x1p5_ASAP7_75t_L g1504 ( 
.A(n_1227),
.B(n_722),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1197),
.Y(n_1505)
);

OAI221xp5_ASAP7_75t_L g1506 ( 
.A1(n_1311),
.A2(n_1345),
.B1(n_1315),
.B2(n_1219),
.C(n_1252),
.Y(n_1506)
);

NAND2xp33_ASAP7_75t_L g1507 ( 
.A(n_1281),
.B(n_894),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1200),
.Y(n_1508)
);

AND2x4_ASAP7_75t_L g1509 ( 
.A(n_1295),
.B(n_34),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1288),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1180),
.B(n_34),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1200),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1226),
.Y(n_1513)
);

INVxp67_ASAP7_75t_L g1514 ( 
.A(n_1350),
.Y(n_1514)
);

AO22x2_ASAP7_75t_L g1515 ( 
.A1(n_1354),
.A2(n_38),
.B1(n_35),
.B2(n_36),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1226),
.Y(n_1516)
);

AOI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1355),
.A2(n_895),
.B1(n_901),
.B2(n_894),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1187),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1187),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1189),
.Y(n_1520)
);

AOI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1181),
.A2(n_895),
.B1(n_901),
.B2(n_894),
.Y(n_1521)
);

OAI221xp5_ASAP7_75t_L g1522 ( 
.A1(n_1239),
.A2(n_901),
.B1(n_924),
.B2(n_895),
.C(n_894),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_1348),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1189),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1180),
.B(n_35),
.Y(n_1525)
);

AO22x2_ASAP7_75t_L g1526 ( 
.A1(n_1363),
.A2(n_40),
.B1(n_36),
.B2(n_39),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1184),
.B(n_39),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1313),
.Y(n_1528)
);

OAI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1184),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_1529)
);

AOI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1268),
.A2(n_895),
.B1(n_901),
.B2(n_894),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1240),
.B(n_42),
.Y(n_1531)
);

OAI221xp5_ASAP7_75t_L g1532 ( 
.A1(n_1217),
.A2(n_924),
.B1(n_931),
.B2(n_901),
.C(n_895),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1266),
.Y(n_1533)
);

INVx4_ASAP7_75t_SL g1534 ( 
.A(n_1281),
.Y(n_1534)
);

AND2x4_ASAP7_75t_L g1535 ( 
.A(n_1357),
.B(n_43),
.Y(n_1535)
);

NAND2xp33_ASAP7_75t_L g1536 ( 
.A(n_1293),
.B(n_924),
.Y(n_1536)
);

INVxp67_ASAP7_75t_L g1537 ( 
.A(n_1201),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1177),
.B(n_43),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1266),
.Y(n_1539)
);

AO22x2_ASAP7_75t_L g1540 ( 
.A1(n_1370),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1304),
.Y(n_1541)
);

AO22x2_ASAP7_75t_L g1542 ( 
.A1(n_1372),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1304),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1289),
.Y(n_1544)
);

BUFx6f_ASAP7_75t_L g1545 ( 
.A(n_1293),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1291),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1321),
.B(n_47),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1300),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1329),
.B(n_47),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1351),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1337),
.B(n_48),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_SL g1552 ( 
.A(n_1293),
.B(n_924),
.Y(n_1552)
);

NAND2x1p5_ASAP7_75t_L g1553 ( 
.A(n_1297),
.B(n_1307),
.Y(n_1553)
);

AO22x2_ASAP7_75t_L g1554 ( 
.A1(n_1364),
.A2(n_1196),
.B1(n_1178),
.B2(n_1352),
.Y(n_1554)
);

NOR2x1_ASAP7_75t_L g1555 ( 
.A(n_1249),
.B(n_924),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1306),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1306),
.Y(n_1557)
);

BUFx2_ASAP7_75t_L g1558 ( 
.A(n_1297),
.Y(n_1558)
);

AO22x2_ASAP7_75t_L g1559 ( 
.A1(n_1301),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1341),
.Y(n_1560)
);

AO22x2_ASAP7_75t_L g1561 ( 
.A1(n_1308),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1341),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1319),
.Y(n_1563)
);

AO22x2_ASAP7_75t_L g1564 ( 
.A1(n_1271),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1325),
.Y(n_1565)
);

AO22x2_ASAP7_75t_L g1566 ( 
.A1(n_1358),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_1566)
);

INVxp67_ASAP7_75t_L g1567 ( 
.A(n_1317),
.Y(n_1567)
);

AOI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1328),
.A2(n_931),
.B1(n_58),
.B2(n_55),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1326),
.B(n_57),
.Y(n_1569)
);

NAND2x1p5_ASAP7_75t_L g1570 ( 
.A(n_1297),
.B(n_931),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1331),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1255),
.B(n_58),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_SL g1573 ( 
.A(n_1284),
.B(n_931),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1343),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1347),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1349),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1307),
.Y(n_1577)
);

INVxp67_ASAP7_75t_L g1578 ( 
.A(n_1335),
.Y(n_1578)
);

OAI221xp5_ASAP7_75t_L g1579 ( 
.A1(n_1316),
.A2(n_931),
.B1(n_61),
.B2(n_59),
.C(n_60),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1298),
.B(n_59),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1365),
.Y(n_1581)
);

INVx4_ASAP7_75t_L g1582 ( 
.A(n_1391),
.Y(n_1582)
);

O2A1O1Ixp33_ASAP7_75t_L g1583 ( 
.A1(n_1506),
.A2(n_1261),
.B(n_1336),
.C(n_1327),
.Y(n_1583)
);

AOI21xp5_ASAP7_75t_L g1584 ( 
.A1(n_1469),
.A2(n_1360),
.B(n_1368),
.Y(n_1584)
);

O2A1O1Ixp33_ASAP7_75t_L g1585 ( 
.A1(n_1425),
.A2(n_1374),
.B(n_1344),
.C(n_1338),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1383),
.B(n_1299),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1463),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1392),
.B(n_1385),
.Y(n_1588)
);

BUFx4f_ASAP7_75t_L g1589 ( 
.A(n_1485),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1435),
.B(n_1312),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1518),
.B(n_1314),
.Y(n_1591)
);

AOI21xp5_ASAP7_75t_L g1592 ( 
.A1(n_1476),
.A2(n_1368),
.B(n_1365),
.Y(n_1592)
);

AOI21x1_ASAP7_75t_L g1593 ( 
.A1(n_1492),
.A2(n_1330),
.B(n_1273),
.Y(n_1593)
);

NOR3xp33_ASAP7_75t_L g1594 ( 
.A(n_1477),
.B(n_1346),
.C(n_60),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1519),
.B(n_1307),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1520),
.B(n_1238),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1439),
.B(n_1406),
.Y(n_1597)
);

BUFx3_ASAP7_75t_L g1598 ( 
.A(n_1493),
.Y(n_1598)
);

AOI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1483),
.A2(n_1238),
.B(n_347),
.Y(n_1599)
);

A2O1A1Ixp33_ASAP7_75t_L g1600 ( 
.A1(n_1480),
.A2(n_1238),
.B(n_64),
.C(n_62),
.Y(n_1600)
);

AOI21xp5_ASAP7_75t_L g1601 ( 
.A1(n_1491),
.A2(n_1238),
.B(n_348),
.Y(n_1601)
);

INVx2_ASAP7_75t_SL g1602 ( 
.A(n_1402),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1524),
.B(n_1238),
.Y(n_1603)
);

OAI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1427),
.A2(n_62),
.B(n_63),
.Y(n_1604)
);

OAI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1481),
.A2(n_1497),
.B1(n_1500),
.B2(n_1494),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_SL g1606 ( 
.A(n_1462),
.B(n_63),
.Y(n_1606)
);

AOI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1505),
.A2(n_349),
.B(n_346),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1437),
.B(n_64),
.Y(n_1608)
);

AOI21xp5_ASAP7_75t_L g1609 ( 
.A1(n_1508),
.A2(n_353),
.B(n_351),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1537),
.B(n_65),
.Y(n_1610)
);

BUFx3_ASAP7_75t_L g1611 ( 
.A(n_1465),
.Y(n_1611)
);

A2O1A1Ixp33_ASAP7_75t_L g1612 ( 
.A1(n_1547),
.A2(n_1549),
.B(n_1471),
.C(n_1556),
.Y(n_1612)
);

AOI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1512),
.A2(n_357),
.B(n_355),
.Y(n_1613)
);

BUFx6f_ASAP7_75t_L g1614 ( 
.A(n_1456),
.Y(n_1614)
);

OAI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1513),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_1615)
);

BUFx6f_ASAP7_75t_L g1616 ( 
.A(n_1456),
.Y(n_1616)
);

AOI21x1_ASAP7_75t_L g1617 ( 
.A1(n_1492),
.A2(n_359),
.B(n_358),
.Y(n_1617)
);

AOI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1516),
.A2(n_363),
.B(n_360),
.Y(n_1618)
);

NOR2xp67_ASAP7_75t_L g1619 ( 
.A(n_1376),
.B(n_364),
.Y(n_1619)
);

BUFx6f_ASAP7_75t_L g1620 ( 
.A(n_1545),
.Y(n_1620)
);

OAI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1453),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_1621)
);

INVxp67_ASAP7_75t_L g1622 ( 
.A(n_1447),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1533),
.B(n_69),
.Y(n_1623)
);

AOI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1387),
.A2(n_372),
.B(n_367),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1404),
.B(n_69),
.Y(n_1625)
);

A2O1A1Ixp33_ASAP7_75t_L g1626 ( 
.A1(n_1557),
.A2(n_72),
.B(n_70),
.C(n_71),
.Y(n_1626)
);

NOR2xp33_ASAP7_75t_L g1627 ( 
.A(n_1389),
.B(n_70),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1539),
.B(n_71),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1394),
.Y(n_1629)
);

AOI21xp5_ASAP7_75t_L g1630 ( 
.A1(n_1511),
.A2(n_374),
.B(n_373),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1525),
.A2(n_379),
.B(n_376),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1378),
.Y(n_1632)
);

AOI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1496),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_SL g1634 ( 
.A(n_1457),
.B(n_380),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1390),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1541),
.B(n_75),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1395),
.Y(n_1637)
);

AOI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1527),
.A2(n_382),
.B(n_381),
.Y(n_1638)
);

OAI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1503),
.A2(n_76),
.B(n_77),
.Y(n_1639)
);

OAI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1551),
.A2(n_77),
.B(n_78),
.Y(n_1640)
);

AOI21xp5_ASAP7_75t_L g1641 ( 
.A1(n_1560),
.A2(n_388),
.B(n_386),
.Y(n_1641)
);

AOI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1562),
.A2(n_392),
.B(n_389),
.Y(n_1642)
);

AOI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1507),
.A2(n_394),
.B(n_393),
.Y(n_1643)
);

INVx3_ASAP7_75t_L g1644 ( 
.A(n_1545),
.Y(n_1644)
);

AOI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1536),
.A2(n_1543),
.B(n_1452),
.Y(n_1645)
);

AND2x6_ASAP7_75t_L g1646 ( 
.A(n_1443),
.B(n_396),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_SL g1647 ( 
.A(n_1535),
.B(n_78),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1461),
.B(n_79),
.Y(n_1648)
);

AO21x1_ASAP7_75t_L g1649 ( 
.A1(n_1384),
.A2(n_1490),
.B(n_1397),
.Y(n_1649)
);

BUFx6f_ASAP7_75t_L g1650 ( 
.A(n_1558),
.Y(n_1650)
);

AOI21x1_ASAP7_75t_L g1651 ( 
.A1(n_1554),
.A2(n_399),
.B(n_398),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1485),
.B(n_80),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1390),
.A2(n_1401),
.B1(n_1414),
.B2(n_1467),
.Y(n_1653)
);

OAI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1495),
.A2(n_83),
.B1(n_80),
.B2(n_81),
.Y(n_1654)
);

AOI21x1_ASAP7_75t_L g1655 ( 
.A1(n_1554),
.A2(n_403),
.B(n_402),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1464),
.B(n_81),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_SL g1657 ( 
.A(n_1509),
.B(n_84),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1401),
.B(n_84),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_SL g1659 ( 
.A(n_1514),
.B(n_1501),
.Y(n_1659)
);

AOI21xp5_ASAP7_75t_L g1660 ( 
.A1(n_1573),
.A2(n_408),
.B(n_404),
.Y(n_1660)
);

AOI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1552),
.A2(n_1421),
.B(n_1580),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1405),
.Y(n_1662)
);

BUFx4f_ASAP7_75t_L g1663 ( 
.A(n_1379),
.Y(n_1663)
);

OAI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1460),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.Y(n_1664)
);

AOI21x1_ASAP7_75t_L g1665 ( 
.A1(n_1424),
.A2(n_411),
.B(n_410),
.Y(n_1665)
);

AOI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1555),
.A2(n_413),
.B(n_412),
.Y(n_1666)
);

NAND2x1p5_ASAP7_75t_L g1667 ( 
.A(n_1451),
.B(n_414),
.Y(n_1667)
);

AOI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1412),
.A2(n_416),
.B(n_415),
.Y(n_1668)
);

BUFx6f_ASAP7_75t_L g1669 ( 
.A(n_1558),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1454),
.B(n_85),
.Y(n_1670)
);

OAI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1489),
.A2(n_86),
.B(n_87),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1522),
.A2(n_421),
.B(n_420),
.Y(n_1672)
);

OAI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1488),
.A2(n_88),
.B(n_89),
.Y(n_1673)
);

AOI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1532),
.A2(n_424),
.B(n_423),
.Y(n_1674)
);

AOI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1441),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1581),
.B(n_90),
.Y(n_1676)
);

AOI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1424),
.A2(n_430),
.B(n_428),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1434),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1407),
.B(n_91),
.Y(n_1679)
);

AOI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1521),
.A2(n_432),
.B(n_431),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1455),
.B(n_93),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1408),
.Y(n_1682)
);

INVx4_ASAP7_75t_L g1683 ( 
.A(n_1534),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1409),
.B(n_93),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1410),
.B(n_94),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1396),
.Y(n_1686)
);

INVx3_ASAP7_75t_L g1687 ( 
.A(n_1553),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1413),
.B(n_94),
.Y(n_1688)
);

OAI21xp5_ASAP7_75t_L g1689 ( 
.A1(n_1430),
.A2(n_95),
.B(n_96),
.Y(n_1689)
);

A2O1A1Ixp33_ASAP7_75t_L g1690 ( 
.A1(n_1442),
.A2(n_97),
.B(n_95),
.C(n_96),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1419),
.B(n_97),
.Y(n_1691)
);

NOR2xp33_ASAP7_75t_L g1692 ( 
.A(n_1567),
.B(n_98),
.Y(n_1692)
);

AOI21xp5_ASAP7_75t_L g1693 ( 
.A1(n_1411),
.A2(n_437),
.B(n_434),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1578),
.B(n_99),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1420),
.Y(n_1695)
);

OA22x2_ASAP7_75t_L g1696 ( 
.A1(n_1459),
.A2(n_103),
.B1(n_101),
.B2(n_102),
.Y(n_1696)
);

AOI21xp5_ASAP7_75t_L g1697 ( 
.A1(n_1569),
.A2(n_1444),
.B(n_1530),
.Y(n_1697)
);

INVx3_ASAP7_75t_L g1698 ( 
.A(n_1380),
.Y(n_1698)
);

AOI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1445),
.A2(n_440),
.B(n_438),
.Y(n_1699)
);

O2A1O1Ixp33_ASAP7_75t_SL g1700 ( 
.A1(n_1529),
.A2(n_103),
.B(n_101),
.C(n_102),
.Y(n_1700)
);

OAI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1498),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.Y(n_1701)
);

AOI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1570),
.A2(n_442),
.B(n_441),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1398),
.B(n_105),
.Y(n_1703)
);

AOI21xp5_ASAP7_75t_L g1704 ( 
.A1(n_1504),
.A2(n_444),
.B(n_443),
.Y(n_1704)
);

AOI21xp5_ASAP7_75t_L g1705 ( 
.A1(n_1478),
.A2(n_449),
.B(n_447),
.Y(n_1705)
);

A2O1A1Ixp33_ASAP7_75t_L g1706 ( 
.A1(n_1568),
.A2(n_108),
.B(n_106),
.C(n_107),
.Y(n_1706)
);

OAI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1450),
.A2(n_1517),
.B(n_1479),
.Y(n_1707)
);

O2A1O1Ixp5_ASAP7_75t_L g1708 ( 
.A1(n_1449),
.A2(n_109),
.B(n_107),
.C(n_108),
.Y(n_1708)
);

O2A1O1Ixp5_ASAP7_75t_L g1709 ( 
.A1(n_1458),
.A2(n_111),
.B(n_109),
.C(n_110),
.Y(n_1709)
);

OAI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1579),
.A2(n_110),
.B(n_111),
.Y(n_1710)
);

AOI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1478),
.A2(n_451),
.B(n_450),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1398),
.B(n_112),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1382),
.B(n_112),
.Y(n_1713)
);

BUFx2_ASAP7_75t_L g1714 ( 
.A(n_1502),
.Y(n_1714)
);

AOI33xp33_ASAP7_75t_L g1715 ( 
.A1(n_1538),
.A2(n_113),
.A3(n_114),
.B1(n_115),
.B2(n_116),
.B3(n_117),
.Y(n_1715)
);

AO22x1_ASAP7_75t_L g1716 ( 
.A1(n_1523),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.Y(n_1716)
);

INVx3_ASAP7_75t_L g1717 ( 
.A(n_1577),
.Y(n_1717)
);

OAI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1475),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_1718)
);

AOI21xp5_ASAP7_75t_L g1719 ( 
.A1(n_1422),
.A2(n_455),
.B(n_453),
.Y(n_1719)
);

A2O1A1Ixp33_ASAP7_75t_L g1720 ( 
.A1(n_1572),
.A2(n_121),
.B(n_118),
.C(n_120),
.Y(n_1720)
);

OAI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1475),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1467),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.Y(n_1722)
);

O2A1O1Ixp33_ASAP7_75t_L g1723 ( 
.A1(n_1400),
.A2(n_126),
.B(n_123),
.C(n_125),
.Y(n_1723)
);

AOI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1531),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_1724)
);

NOR2x1_ASAP7_75t_R g1725 ( 
.A(n_1377),
.B(n_128),
.Y(n_1725)
);

BUFx4f_ASAP7_75t_L g1726 ( 
.A(n_1482),
.Y(n_1726)
);

OAI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1448),
.A2(n_132),
.B1(n_130),
.B2(n_131),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1426),
.Y(n_1728)
);

AOI21xp5_ASAP7_75t_L g1729 ( 
.A1(n_1428),
.A2(n_457),
.B(n_456),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1399),
.Y(n_1730)
);

AOI22xp5_ASAP7_75t_L g1731 ( 
.A1(n_1388),
.A2(n_134),
.B1(n_130),
.B2(n_133),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1382),
.B(n_133),
.Y(n_1732)
);

INVxp67_ASAP7_75t_SL g1733 ( 
.A(n_1574),
.Y(n_1733)
);

AOI21xp5_ASAP7_75t_L g1734 ( 
.A1(n_1431),
.A2(n_460),
.B(n_458),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1403),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1381),
.B(n_134),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1433),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1550),
.B(n_135),
.Y(n_1738)
);

HB1xp67_ASAP7_75t_L g1739 ( 
.A(n_1534),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_SL g1740 ( 
.A(n_1486),
.B(n_135),
.Y(n_1740)
);

AOI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1414),
.A2(n_1561),
.B1(n_1564),
.B2(n_1559),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1386),
.A2(n_138),
.B1(n_136),
.B2(n_137),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1528),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1386),
.B(n_136),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1544),
.B(n_137),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1418),
.Y(n_1746)
);

INVx5_ASAP7_75t_L g1747 ( 
.A(n_1440),
.Y(n_1747)
);

OAI321xp33_ASAP7_75t_L g1748 ( 
.A1(n_1448),
.A2(n_138),
.A3(n_139),
.B1(n_140),
.B2(n_141),
.C(n_142),
.Y(n_1748)
);

AOI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1515),
.A2(n_463),
.B(n_461),
.Y(n_1749)
);

AOI21xp5_ASAP7_75t_L g1750 ( 
.A1(n_1515),
.A2(n_466),
.B(n_464),
.Y(n_1750)
);

AOI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1559),
.A2(n_141),
.B1(n_139),
.B2(n_140),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1546),
.B(n_143),
.Y(n_1752)
);

AOI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1526),
.A2(n_1542),
.B(n_1540),
.Y(n_1753)
);

NOR2xp33_ASAP7_75t_L g1754 ( 
.A(n_1563),
.B(n_144),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1548),
.B(n_144),
.Y(n_1755)
);

AOI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1526),
.A2(n_469),
.B(n_467),
.Y(n_1756)
);

NOR2xp33_ASAP7_75t_L g1757 ( 
.A(n_1565),
.B(n_145),
.Y(n_1757)
);

A2O1A1Ixp33_ASAP7_75t_L g1758 ( 
.A1(n_1571),
.A2(n_147),
.B(n_145),
.C(n_146),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1575),
.Y(n_1759)
);

BUFx6f_ASAP7_75t_L g1760 ( 
.A(n_1415),
.Y(n_1760)
);

AOI22xp33_ASAP7_75t_L g1761 ( 
.A1(n_1561),
.A2(n_149),
.B1(n_147),
.B2(n_148),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1576),
.Y(n_1762)
);

AOI21x1_ASAP7_75t_L g1763 ( 
.A1(n_1393),
.A2(n_473),
.B(n_470),
.Y(n_1763)
);

O2A1O1Ixp33_ASAP7_75t_L g1764 ( 
.A1(n_1564),
.A2(n_151),
.B(n_149),
.C(n_150),
.Y(n_1764)
);

HB1xp67_ASAP7_75t_L g1765 ( 
.A(n_1466),
.Y(n_1765)
);

AOI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1540),
.A2(n_475),
.B(n_474),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1393),
.B(n_151),
.Y(n_1767)
);

BUFx3_ASAP7_75t_L g1768 ( 
.A(n_1436),
.Y(n_1768)
);

INVx3_ASAP7_75t_L g1769 ( 
.A(n_1470),
.Y(n_1769)
);

AOI21x1_ASAP7_75t_L g1770 ( 
.A1(n_1416),
.A2(n_477),
.B(n_476),
.Y(n_1770)
);

NOR2xp33_ASAP7_75t_L g1771 ( 
.A(n_1446),
.B(n_152),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1468),
.B(n_1484),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1681),
.B(n_1472),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1632),
.Y(n_1774)
);

AOI21xp5_ASAP7_75t_L g1775 ( 
.A1(n_1599),
.A2(n_1542),
.B(n_1423),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_SL g1776 ( 
.A(n_1597),
.B(n_1487),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_R g1777 ( 
.A(n_1598),
.B(n_1440),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1714),
.B(n_152),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1662),
.Y(n_1779)
);

AOI21xp5_ASAP7_75t_L g1780 ( 
.A1(n_1601),
.A2(n_1423),
.B(n_1417),
.Y(n_1780)
);

BUFx6f_ASAP7_75t_L g1781 ( 
.A(n_1683),
.Y(n_1781)
);

O2A1O1Ixp33_ASAP7_75t_L g1782 ( 
.A1(n_1689),
.A2(n_1438),
.B(n_1473),
.C(n_1566),
.Y(n_1782)
);

O2A1O1Ixp33_ASAP7_75t_L g1783 ( 
.A1(n_1671),
.A2(n_1438),
.B(n_1473),
.C(n_1566),
.Y(n_1783)
);

AOI21x1_ASAP7_75t_L g1784 ( 
.A1(n_1593),
.A2(n_1416),
.B(n_1474),
.Y(n_1784)
);

INVx2_ASAP7_75t_SL g1785 ( 
.A(n_1663),
.Y(n_1785)
);

AOI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1605),
.A2(n_1697),
.B(n_1603),
.Y(n_1786)
);

A2O1A1Ixp33_ASAP7_75t_L g1787 ( 
.A1(n_1639),
.A2(n_1474),
.B(n_1472),
.C(n_1429),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_L g1788 ( 
.A(n_1725),
.B(n_153),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1587),
.B(n_153),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1682),
.Y(n_1790)
);

AOI21xp5_ASAP7_75t_L g1791 ( 
.A1(n_1596),
.A2(n_1429),
.B(n_1417),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1633),
.A2(n_1432),
.B1(n_1510),
.B2(n_1499),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_SL g1793 ( 
.A(n_1588),
.B(n_1432),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1695),
.B(n_154),
.Y(n_1794)
);

CKINVDCx14_ASAP7_75t_R g1795 ( 
.A(n_1663),
.Y(n_1795)
);

INVx4_ASAP7_75t_L g1796 ( 
.A(n_1683),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1728),
.Y(n_1797)
);

AOI21xp5_ASAP7_75t_L g1798 ( 
.A1(n_1645),
.A2(n_1440),
.B(n_155),
.Y(n_1798)
);

NOR2xp33_ASAP7_75t_L g1799 ( 
.A(n_1670),
.B(n_155),
.Y(n_1799)
);

BUFx6f_ASAP7_75t_L g1800 ( 
.A(n_1589),
.Y(n_1800)
);

OAI22xp5_ASAP7_75t_L g1801 ( 
.A1(n_1741),
.A2(n_158),
.B1(n_156),
.B2(n_157),
.Y(n_1801)
);

NOR2xp33_ASAP7_75t_SL g1802 ( 
.A(n_1747),
.B(n_157),
.Y(n_1802)
);

BUFx3_ASAP7_75t_L g1803 ( 
.A(n_1611),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_SL g1804 ( 
.A(n_1707),
.B(n_158),
.Y(n_1804)
);

AOI21xp5_ASAP7_75t_L g1805 ( 
.A1(n_1584),
.A2(n_159),
.B(n_160),
.Y(n_1805)
);

AOI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1661),
.A2(n_160),
.B(n_161),
.Y(n_1806)
);

O2A1O1Ixp33_ASAP7_75t_L g1807 ( 
.A1(n_1720),
.A2(n_163),
.B(n_161),
.C(n_162),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_SL g1808 ( 
.A(n_1589),
.B(n_163),
.Y(n_1808)
);

AOI21xp5_ASAP7_75t_L g1809 ( 
.A1(n_1612),
.A2(n_164),
.B(n_165),
.Y(n_1809)
);

AOI22xp5_ASAP7_75t_L g1810 ( 
.A1(n_1647),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.Y(n_1810)
);

BUFx2_ASAP7_75t_L g1811 ( 
.A(n_1614),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1737),
.Y(n_1812)
);

BUFx3_ASAP7_75t_L g1813 ( 
.A(n_1602),
.Y(n_1813)
);

AOI21xp5_ASAP7_75t_L g1814 ( 
.A1(n_1592),
.A2(n_166),
.B(n_167),
.Y(n_1814)
);

BUFx2_ASAP7_75t_L g1815 ( 
.A(n_1614),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1629),
.Y(n_1816)
);

BUFx12f_ASAP7_75t_L g1817 ( 
.A(n_1582),
.Y(n_1817)
);

AOI22xp5_ASAP7_75t_L g1818 ( 
.A1(n_1736),
.A2(n_169),
.B1(n_167),
.B2(n_168),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_L g1819 ( 
.A(n_1582),
.B(n_168),
.Y(n_1819)
);

BUFx12f_ASAP7_75t_L g1820 ( 
.A(n_1614),
.Y(n_1820)
);

NOR3xp33_ASAP7_75t_SL g1821 ( 
.A(n_1627),
.B(n_169),
.C(n_170),
.Y(n_1821)
);

O2A1O1Ixp33_ASAP7_75t_L g1822 ( 
.A1(n_1723),
.A2(n_173),
.B(n_171),
.C(n_172),
.Y(n_1822)
);

OAI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1675),
.A2(n_177),
.B1(n_174),
.B2(n_176),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1678),
.B(n_176),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1743),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1759),
.Y(n_1826)
);

BUFx2_ASAP7_75t_L g1827 ( 
.A(n_1616),
.Y(n_1827)
);

AOI21xp5_ASAP7_75t_L g1828 ( 
.A1(n_1680),
.A2(n_177),
.B(n_178),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1762),
.Y(n_1829)
);

NOR2xp33_ASAP7_75t_L g1830 ( 
.A(n_1657),
.B(n_178),
.Y(n_1830)
);

AOI21xp5_ASAP7_75t_L g1831 ( 
.A1(n_1672),
.A2(n_1674),
.B(n_1591),
.Y(n_1831)
);

INVx3_ASAP7_75t_L g1832 ( 
.A(n_1620),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_SL g1833 ( 
.A(n_1650),
.B(n_179),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1608),
.B(n_179),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1765),
.Y(n_1835)
);

NOR2xp67_ASAP7_75t_L g1836 ( 
.A(n_1739),
.B(n_478),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1590),
.B(n_180),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1637),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_SL g1839 ( 
.A(n_1650),
.B(n_180),
.Y(n_1839)
);

O2A1O1Ixp33_ASAP7_75t_SL g1840 ( 
.A1(n_1600),
.A2(n_183),
.B(n_181),
.C(n_182),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1686),
.Y(n_1841)
);

AOI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1694),
.A2(n_184),
.B1(n_181),
.B2(n_183),
.Y(n_1842)
);

OR2x2_ASAP7_75t_L g1843 ( 
.A(n_1622),
.B(n_184),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1653),
.B(n_185),
.Y(n_1844)
);

INVx5_ASAP7_75t_L g1845 ( 
.A(n_1646),
.Y(n_1845)
);

A2O1A1Ixp33_ASAP7_75t_L g1846 ( 
.A1(n_1583),
.A2(n_187),
.B(n_185),
.C(n_186),
.Y(n_1846)
);

A2O1A1Ixp33_ASAP7_75t_L g1847 ( 
.A1(n_1710),
.A2(n_188),
.B(n_186),
.C(n_187),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1730),
.Y(n_1848)
);

NAND3xp33_ASAP7_75t_L g1849 ( 
.A(n_1673),
.B(n_188),
.C(n_189),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1648),
.B(n_189),
.Y(n_1850)
);

A2O1A1Ixp33_ASAP7_75t_L g1851 ( 
.A1(n_1753),
.A2(n_192),
.B(n_190),
.C(n_191),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_SL g1852 ( 
.A(n_1650),
.B(n_190),
.Y(n_1852)
);

NOR2xp33_ASAP7_75t_L g1853 ( 
.A(n_1625),
.B(n_192),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1656),
.B(n_193),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1735),
.Y(n_1855)
);

AOI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1643),
.A2(n_194),
.B(n_195),
.Y(n_1856)
);

AOI21xp5_ASAP7_75t_L g1857 ( 
.A1(n_1586),
.A2(n_195),
.B(n_196),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_SL g1858 ( 
.A(n_1669),
.B(n_198),
.Y(n_1858)
);

AOI21xp5_ASAP7_75t_L g1859 ( 
.A1(n_1699),
.A2(n_198),
.B(n_199),
.Y(n_1859)
);

NOR2xp33_ASAP7_75t_L g1860 ( 
.A(n_1740),
.B(n_199),
.Y(n_1860)
);

HB1xp67_ASAP7_75t_L g1861 ( 
.A(n_1669),
.Y(n_1861)
);

NOR3xp33_ASAP7_75t_SL g1862 ( 
.A(n_1654),
.B(n_200),
.C(n_201),
.Y(n_1862)
);

OAI22xp5_ASAP7_75t_L g1863 ( 
.A1(n_1724),
.A2(n_203),
.B1(n_200),
.B2(n_201),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1715),
.B(n_203),
.Y(n_1864)
);

AOI21xp5_ASAP7_75t_L g1865 ( 
.A1(n_1630),
.A2(n_204),
.B(n_205),
.Y(n_1865)
);

AOI21xp5_ASAP7_75t_L g1866 ( 
.A1(n_1631),
.A2(n_1638),
.B(n_1649),
.Y(n_1866)
);

BUFx6f_ASAP7_75t_L g1867 ( 
.A(n_1669),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1746),
.Y(n_1868)
);

AOI21xp5_ASAP7_75t_L g1869 ( 
.A1(n_1607),
.A2(n_206),
.B(n_207),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1717),
.Y(n_1870)
);

NOR2xp33_ASAP7_75t_L g1871 ( 
.A(n_1644),
.B(n_208),
.Y(n_1871)
);

CKINVDCx5p33_ASAP7_75t_R g1872 ( 
.A(n_1616),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1772),
.Y(n_1873)
);

INVxp67_ASAP7_75t_L g1874 ( 
.A(n_1659),
.Y(n_1874)
);

BUFx2_ASAP7_75t_L g1875 ( 
.A(n_1616),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1733),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1717),
.Y(n_1877)
);

OAI22xp33_ASAP7_75t_L g1878 ( 
.A1(n_1696),
.A2(n_210),
.B1(n_208),
.B2(n_209),
.Y(n_1878)
);

AOI22xp33_ASAP7_75t_L g1879 ( 
.A1(n_1718),
.A2(n_212),
.B1(n_209),
.B2(n_211),
.Y(n_1879)
);

O2A1O1Ixp33_ASAP7_75t_L g1880 ( 
.A1(n_1722),
.A2(n_215),
.B(n_212),
.C(n_214),
.Y(n_1880)
);

AOI21xp5_ASAP7_75t_L g1881 ( 
.A1(n_1609),
.A2(n_215),
.B(n_216),
.Y(n_1881)
);

AOI21xp5_ASAP7_75t_L g1882 ( 
.A1(n_1613),
.A2(n_216),
.B(n_217),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1623),
.B(n_217),
.Y(n_1883)
);

NOR2xp33_ASAP7_75t_SL g1884 ( 
.A(n_1747),
.B(n_218),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1628),
.B(n_218),
.Y(n_1885)
);

NOR2xp33_ASAP7_75t_L g1886 ( 
.A(n_1644),
.B(n_219),
.Y(n_1886)
);

OAI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1751),
.A2(n_219),
.B1(n_220),
.B2(n_222),
.Y(n_1887)
);

O2A1O1Ixp33_ASAP7_75t_L g1888 ( 
.A1(n_1721),
.A2(n_223),
.B(n_224),
.C(n_225),
.Y(n_1888)
);

OA22x2_ASAP7_75t_L g1889 ( 
.A1(n_1731),
.A2(n_223),
.B1(n_224),
.B2(n_226),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1745),
.Y(n_1890)
);

INVxp67_ASAP7_75t_L g1891 ( 
.A(n_1692),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1752),
.Y(n_1892)
);

AOI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1618),
.A2(n_227),
.B(n_228),
.Y(n_1893)
);

AOI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1624),
.A2(n_227),
.B(n_228),
.Y(n_1894)
);

AOI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1641),
.A2(n_229),
.B(n_230),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1755),
.Y(n_1896)
);

BUFx2_ASAP7_75t_L g1897 ( 
.A(n_1620),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_SL g1898 ( 
.A(n_1747),
.B(n_230),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1713),
.Y(n_1899)
);

OR2x6_ASAP7_75t_L g1900 ( 
.A(n_1749),
.B(n_479),
.Y(n_1900)
);

OAI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1761),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_1901)
);

BUFx3_ASAP7_75t_L g1902 ( 
.A(n_1620),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1636),
.B(n_232),
.Y(n_1903)
);

AND2x4_ASAP7_75t_L g1904 ( 
.A(n_1768),
.B(n_234),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_SL g1905 ( 
.A(n_1760),
.B(n_1698),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1676),
.B(n_234),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1754),
.B(n_1757),
.Y(n_1907)
);

INVx1_ASAP7_75t_SL g1908 ( 
.A(n_1595),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1687),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1658),
.B(n_235),
.Y(n_1910)
);

AOI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1642),
.A2(n_236),
.B(n_237),
.Y(n_1911)
);

AOI22xp5_ASAP7_75t_L g1912 ( 
.A1(n_1652),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_1912)
);

NOR3xp33_ASAP7_75t_SL g1913 ( 
.A(n_1727),
.B(n_239),
.C(n_240),
.Y(n_1913)
);

BUFx6f_ASAP7_75t_SL g1914 ( 
.A(n_1646),
.Y(n_1914)
);

OAI22xp5_ASAP7_75t_L g1915 ( 
.A1(n_1635),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1738),
.B(n_242),
.Y(n_1916)
);

AOI21xp5_ASAP7_75t_L g1917 ( 
.A1(n_1585),
.A2(n_243),
.B(n_244),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1679),
.B(n_244),
.Y(n_1918)
);

AOI21xp5_ASAP7_75t_L g1919 ( 
.A1(n_1666),
.A2(n_245),
.B(n_246),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_SL g1920 ( 
.A(n_1760),
.B(n_245),
.Y(n_1920)
);

AOI21xp5_ASAP7_75t_L g1921 ( 
.A1(n_1719),
.A2(n_1734),
.B(n_1729),
.Y(n_1921)
);

AOI21xp5_ASAP7_75t_L g1922 ( 
.A1(n_1693),
.A2(n_247),
.B(n_248),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_R g1923 ( 
.A(n_1726),
.B(n_569),
.Y(n_1923)
);

INVxp67_ASAP7_75t_L g1924 ( 
.A(n_1610),
.Y(n_1924)
);

AOI21xp5_ASAP7_75t_L g1925 ( 
.A1(n_1640),
.A2(n_249),
.B(n_250),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1716),
.B(n_249),
.Y(n_1926)
);

OAI22xp5_ASAP7_75t_L g1927 ( 
.A1(n_1604),
.A2(n_250),
.B1(n_251),
.B2(n_252),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1684),
.B(n_251),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1732),
.B(n_252),
.Y(n_1929)
);

HB1xp67_ASAP7_75t_L g1930 ( 
.A(n_1744),
.Y(n_1930)
);

NOR2x1_ASAP7_75t_L g1931 ( 
.A(n_1703),
.B(n_253),
.Y(n_1931)
);

HB1xp67_ASAP7_75t_L g1932 ( 
.A(n_1712),
.Y(n_1932)
);

HB1xp67_ASAP7_75t_L g1933 ( 
.A(n_1767),
.Y(n_1933)
);

OAI22xp33_ASAP7_75t_L g1934 ( 
.A1(n_1748),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_1934)
);

INVx3_ASAP7_75t_L g1935 ( 
.A(n_1687),
.Y(n_1935)
);

AOI21xp5_ASAP7_75t_L g1936 ( 
.A1(n_1677),
.A2(n_254),
.B(n_255),
.Y(n_1936)
);

BUFx2_ASAP7_75t_L g1937 ( 
.A(n_1698),
.Y(n_1937)
);

AOI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1705),
.A2(n_1711),
.B(n_1660),
.Y(n_1938)
);

OAI21xp5_ASAP7_75t_L g1939 ( 
.A1(n_1849),
.A2(n_1756),
.B(n_1750),
.Y(n_1939)
);

CKINVDCx5p33_ASAP7_75t_R g1940 ( 
.A(n_1803),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1774),
.Y(n_1941)
);

CKINVDCx20_ASAP7_75t_R g1942 ( 
.A(n_1795),
.Y(n_1942)
);

A2O1A1Ixp33_ASAP7_75t_L g1943 ( 
.A1(n_1782),
.A2(n_1764),
.B(n_1766),
.C(n_1706),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1779),
.Y(n_1944)
);

AOI21xp5_ASAP7_75t_L g1945 ( 
.A1(n_1921),
.A2(n_1594),
.B(n_1700),
.Y(n_1945)
);

BUFx10_ASAP7_75t_L g1946 ( 
.A(n_1819),
.Y(n_1946)
);

AOI21xp5_ASAP7_75t_L g1947 ( 
.A1(n_1786),
.A2(n_1866),
.B(n_1831),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_SL g1948 ( 
.A(n_1845),
.B(n_1634),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1790),
.Y(n_1949)
);

OAI21x1_ASAP7_75t_L g1950 ( 
.A1(n_1938),
.A2(n_1665),
.B(n_1617),
.Y(n_1950)
);

AOI221x1_ASAP7_75t_L g1951 ( 
.A1(n_1801),
.A2(n_1887),
.B1(n_1787),
.B2(n_1925),
.C(n_1927),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1899),
.B(n_1685),
.Y(n_1952)
);

OAI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1891),
.A2(n_1742),
.B1(n_1690),
.B2(n_1626),
.Y(n_1953)
);

AOI21xp5_ASAP7_75t_L g1954 ( 
.A1(n_1780),
.A2(n_1668),
.B(n_1704),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1797),
.Y(n_1955)
);

AOI21xp5_ASAP7_75t_L g1956 ( 
.A1(n_1775),
.A2(n_1702),
.B(n_1701),
.Y(n_1956)
);

OR2x6_ASAP7_75t_L g1957 ( 
.A(n_1800),
.B(n_1667),
.Y(n_1957)
);

INVxp67_ASAP7_75t_L g1958 ( 
.A(n_1835),
.Y(n_1958)
);

BUFx3_ASAP7_75t_L g1959 ( 
.A(n_1813),
.Y(n_1959)
);

AOI21xp33_ASAP7_75t_L g1960 ( 
.A1(n_1783),
.A2(n_1621),
.B(n_1664),
.Y(n_1960)
);

INVx1_ASAP7_75t_SL g1961 ( 
.A(n_1872),
.Y(n_1961)
);

OAI21x1_ASAP7_75t_L g1962 ( 
.A1(n_1798),
.A2(n_1655),
.B(n_1651),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1773),
.B(n_1771),
.Y(n_1963)
);

AOI22xp5_ASAP7_75t_L g1964 ( 
.A1(n_1907),
.A2(n_1606),
.B1(n_1646),
.B2(n_1615),
.Y(n_1964)
);

AO21x1_ASAP7_75t_L g1965 ( 
.A1(n_1801),
.A2(n_1770),
.B(n_1691),
.Y(n_1965)
);

CKINVDCx11_ASAP7_75t_R g1966 ( 
.A(n_1817),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1930),
.B(n_1688),
.Y(n_1967)
);

HB1xp67_ASAP7_75t_L g1968 ( 
.A(n_1932),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1812),
.Y(n_1969)
);

AND2x4_ASAP7_75t_L g1970 ( 
.A(n_1867),
.B(n_1760),
.Y(n_1970)
);

OA21x2_ASAP7_75t_L g1971 ( 
.A1(n_1791),
.A2(n_1763),
.B(n_1709),
.Y(n_1971)
);

OAI21x1_ASAP7_75t_L g1972 ( 
.A1(n_1805),
.A2(n_1708),
.B(n_1769),
.Y(n_1972)
);

BUFx6f_ASAP7_75t_L g1973 ( 
.A(n_1800),
.Y(n_1973)
);

NOR2xp33_ASAP7_75t_SL g1974 ( 
.A(n_1800),
.B(n_1726),
.Y(n_1974)
);

AOI21xp5_ASAP7_75t_L g1975 ( 
.A1(n_1845),
.A2(n_1900),
.B(n_1849),
.Y(n_1975)
);

AOI21xp5_ASAP7_75t_L g1976 ( 
.A1(n_1845),
.A2(n_1900),
.B(n_1828),
.Y(n_1976)
);

AOI21xp5_ASAP7_75t_L g1977 ( 
.A1(n_1900),
.A2(n_1758),
.B(n_1646),
.Y(n_1977)
);

NOR2xp33_ASAP7_75t_L g1978 ( 
.A(n_1799),
.B(n_256),
.Y(n_1978)
);

AO31x2_ASAP7_75t_L g1979 ( 
.A1(n_1792),
.A2(n_1619),
.A3(n_568),
.B(n_567),
.Y(n_1979)
);

AOI21xp5_ASAP7_75t_L g1980 ( 
.A1(n_1856),
.A2(n_257),
.B(n_258),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1825),
.Y(n_1981)
);

BUFx3_ASAP7_75t_L g1982 ( 
.A(n_1820),
.Y(n_1982)
);

INVx2_ASAP7_75t_SL g1983 ( 
.A(n_1902),
.Y(n_1983)
);

AOI21xp5_ASAP7_75t_L g1984 ( 
.A1(n_1804),
.A2(n_258),
.B(n_259),
.Y(n_1984)
);

CKINVDCx20_ASAP7_75t_R g1985 ( 
.A(n_1861),
.Y(n_1985)
);

AO32x2_ASAP7_75t_L g1986 ( 
.A1(n_1887),
.A2(n_259),
.A3(n_260),
.B1(n_261),
.B2(n_262),
.Y(n_1986)
);

OAI21xp5_ASAP7_75t_L g1987 ( 
.A1(n_1847),
.A2(n_263),
.B(n_264),
.Y(n_1987)
);

NAND2x1p5_ASAP7_75t_L g1988 ( 
.A(n_1796),
.B(n_481),
.Y(n_1988)
);

BUFx2_ASAP7_75t_L g1989 ( 
.A(n_1867),
.Y(n_1989)
);

AO32x2_ASAP7_75t_L g1990 ( 
.A1(n_1823),
.A2(n_263),
.A3(n_264),
.B1(n_265),
.B2(n_266),
.Y(n_1990)
);

AOI21x1_ASAP7_75t_SL g1991 ( 
.A1(n_1864),
.A2(n_265),
.B(n_266),
.Y(n_1991)
);

NOR2xp67_ASAP7_75t_L g1992 ( 
.A(n_1796),
.B(n_1933),
.Y(n_1992)
);

AO22x2_ASAP7_75t_L g1993 ( 
.A1(n_1793),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_1993)
);

BUFx6f_ASAP7_75t_L g1994 ( 
.A(n_1781),
.Y(n_1994)
);

OAI21xp5_ASAP7_75t_L g1995 ( 
.A1(n_1846),
.A2(n_268),
.B(n_270),
.Y(n_1995)
);

OAI21x1_ASAP7_75t_L g1996 ( 
.A1(n_1936),
.A2(n_483),
.B(n_482),
.Y(n_1996)
);

AOI21x1_ASAP7_75t_L g1997 ( 
.A1(n_1784),
.A2(n_1917),
.B(n_1806),
.Y(n_1997)
);

OAI22xp5_ASAP7_75t_L g1998 ( 
.A1(n_1842),
.A2(n_271),
.B1(n_272),
.B2(n_273),
.Y(n_1998)
);

AOI221x1_ASAP7_75t_L g1999 ( 
.A1(n_1809),
.A2(n_273),
.B1(n_274),
.B2(n_275),
.C(n_276),
.Y(n_1999)
);

A2O1A1Ixp33_ASAP7_75t_L g2000 ( 
.A1(n_1822),
.A2(n_274),
.B(n_275),
.C(n_277),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1873),
.B(n_277),
.Y(n_2001)
);

NAND3xp33_ASAP7_75t_SL g2002 ( 
.A(n_1818),
.B(n_278),
.C(n_279),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1890),
.B(n_278),
.Y(n_2003)
);

O2A1O1Ixp5_ASAP7_75t_SL g2004 ( 
.A1(n_1892),
.A2(n_279),
.B(n_280),
.C(n_281),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_SL g2005 ( 
.A(n_1802),
.B(n_484),
.Y(n_2005)
);

AO32x2_ASAP7_75t_L g2006 ( 
.A1(n_1901),
.A2(n_1863),
.A3(n_1915),
.B1(n_1908),
.B2(n_1785),
.Y(n_2006)
);

OAI21x1_ASAP7_75t_L g2007 ( 
.A1(n_1859),
.A2(n_487),
.B(n_565),
.Y(n_2007)
);

AND2x4_ASAP7_75t_L g2008 ( 
.A(n_1908),
.B(n_488),
.Y(n_2008)
);

INVx1_ASAP7_75t_SL g2009 ( 
.A(n_1811),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_SL g2010 ( 
.A(n_1802),
.B(n_489),
.Y(n_2010)
);

AOI21x1_ASAP7_75t_L g2011 ( 
.A1(n_1814),
.A2(n_1896),
.B(n_1910),
.Y(n_2011)
);

O2A1O1Ixp5_ASAP7_75t_L g2012 ( 
.A1(n_1934),
.A2(n_280),
.B(n_282),
.C(n_283),
.Y(n_2012)
);

OAI21xp5_ASAP7_75t_L g2013 ( 
.A1(n_1869),
.A2(n_282),
.B(n_284),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1826),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1829),
.B(n_284),
.Y(n_2015)
);

AOI21xp5_ASAP7_75t_L g2016 ( 
.A1(n_1881),
.A2(n_285),
.B(n_286),
.Y(n_2016)
);

CKINVDCx5p33_ASAP7_75t_R g2017 ( 
.A(n_1815),
.Y(n_2017)
);

OAI21x1_ASAP7_75t_L g2018 ( 
.A1(n_1919),
.A2(n_492),
.B(n_563),
.Y(n_2018)
);

OAI21x1_ASAP7_75t_L g2019 ( 
.A1(n_1894),
.A2(n_491),
.B(n_562),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1924),
.B(n_287),
.Y(n_2020)
);

AOI21xp5_ASAP7_75t_L g2021 ( 
.A1(n_1882),
.A2(n_287),
.B(n_288),
.Y(n_2021)
);

AOI211x1_ASAP7_75t_L g2022 ( 
.A1(n_1878),
.A2(n_289),
.B(n_290),
.C(n_291),
.Y(n_2022)
);

OAI21x1_ASAP7_75t_SL g2023 ( 
.A1(n_1807),
.A2(n_289),
.B(n_290),
.Y(n_2023)
);

OAI21xp5_ASAP7_75t_L g2024 ( 
.A1(n_1893),
.A2(n_291),
.B(n_292),
.Y(n_2024)
);

AOI21xp33_ASAP7_75t_L g2025 ( 
.A1(n_1888),
.A2(n_293),
.B(n_294),
.Y(n_2025)
);

CKINVDCx8_ASAP7_75t_R g2026 ( 
.A(n_1781),
.Y(n_2026)
);

AOI21xp5_ASAP7_75t_L g2027 ( 
.A1(n_1895),
.A2(n_293),
.B(n_294),
.Y(n_2027)
);

OAI22x1_ASAP7_75t_L g2028 ( 
.A1(n_1926),
.A2(n_295),
.B1(n_296),
.B2(n_297),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1929),
.B(n_296),
.Y(n_2029)
);

HB1xp67_ASAP7_75t_L g2030 ( 
.A(n_1937),
.Y(n_2030)
);

AND2x4_ASAP7_75t_L g2031 ( 
.A(n_1827),
.B(n_493),
.Y(n_2031)
);

AND2x4_ASAP7_75t_L g2032 ( 
.A(n_1875),
.B(n_494),
.Y(n_2032)
);

OAI22xp5_ASAP7_75t_L g2033 ( 
.A1(n_1912),
.A2(n_297),
.B1(n_300),
.B2(n_301),
.Y(n_2033)
);

AOI221x1_ASAP7_75t_L g2034 ( 
.A1(n_1851),
.A2(n_1857),
.B1(n_1844),
.B2(n_1865),
.C(n_1911),
.Y(n_2034)
);

BUFx4f_ASAP7_75t_L g2035 ( 
.A(n_1781),
.Y(n_2035)
);

NOR2xp33_ASAP7_75t_L g2036 ( 
.A(n_1874),
.B(n_1853),
.Y(n_2036)
);

BUFx3_ASAP7_75t_L g2037 ( 
.A(n_1897),
.Y(n_2037)
);

INVx1_ASAP7_75t_SL g2038 ( 
.A(n_1923),
.Y(n_2038)
);

A2O1A1Ixp33_ASAP7_75t_L g2039 ( 
.A1(n_1880),
.A2(n_1860),
.B(n_1862),
.C(n_1830),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1941),
.Y(n_2040)
);

BUFx10_ASAP7_75t_L g2041 ( 
.A(n_1994),
.Y(n_2041)
);

INVx1_ASAP7_75t_SL g2042 ( 
.A(n_1959),
.Y(n_2042)
);

OAI21x1_ASAP7_75t_L g2043 ( 
.A1(n_1950),
.A2(n_1922),
.B(n_1877),
.Y(n_2043)
);

AOI22xp33_ASAP7_75t_L g2044 ( 
.A1(n_1993),
.A2(n_1889),
.B1(n_1914),
.B2(n_1931),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1968),
.B(n_1789),
.Y(n_2045)
);

OAI22xp33_ASAP7_75t_L g2046 ( 
.A1(n_1951),
.A2(n_1884),
.B1(n_1810),
.B2(n_1794),
.Y(n_2046)
);

OAI21x1_ASAP7_75t_L g2047 ( 
.A1(n_1947),
.A2(n_1962),
.B(n_1976),
.Y(n_2047)
);

OAI222xp33_ASAP7_75t_L g2048 ( 
.A1(n_1964),
.A2(n_1855),
.B1(n_1841),
.B2(n_1848),
.C1(n_1876),
.C2(n_1879),
.Y(n_2048)
);

OAI21x1_ASAP7_75t_SL g2049 ( 
.A1(n_1975),
.A2(n_1854),
.B(n_1850),
.Y(n_2049)
);

BUFx2_ASAP7_75t_L g2050 ( 
.A(n_2030),
.Y(n_2050)
);

OAI22xp33_ASAP7_75t_L g2051 ( 
.A1(n_1987),
.A2(n_1884),
.B1(n_1885),
.B2(n_1906),
.Y(n_2051)
);

BUFx10_ASAP7_75t_L g2052 ( 
.A(n_1994),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1944),
.Y(n_2053)
);

INVx3_ASAP7_75t_L g2054 ( 
.A(n_1971),
.Y(n_2054)
);

OA21x2_ASAP7_75t_L g2055 ( 
.A1(n_1939),
.A2(n_1870),
.B(n_1913),
.Y(n_2055)
);

AOI22xp33_ASAP7_75t_L g2056 ( 
.A1(n_1993),
.A2(n_1914),
.B1(n_1788),
.B2(n_1776),
.Y(n_2056)
);

AOI21xp5_ASAP7_75t_SL g2057 ( 
.A1(n_1977),
.A2(n_1948),
.B(n_1943),
.Y(n_2057)
);

OAI21x1_ASAP7_75t_L g2058 ( 
.A1(n_1954),
.A2(n_1898),
.B(n_1935),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1949),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1955),
.Y(n_2060)
);

OAI21x1_ASAP7_75t_L g2061 ( 
.A1(n_1945),
.A2(n_1935),
.B(n_1832),
.Y(n_2061)
);

OR2x2_ASAP7_75t_L g2062 ( 
.A(n_1958),
.B(n_1824),
.Y(n_2062)
);

OAI21x1_ASAP7_75t_L g2063 ( 
.A1(n_1997),
.A2(n_1832),
.B(n_1905),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1969),
.Y(n_2064)
);

OAI21x1_ASAP7_75t_L g2065 ( 
.A1(n_1956),
.A2(n_1839),
.B(n_1852),
.Y(n_2065)
);

AO21x2_ASAP7_75t_L g2066 ( 
.A1(n_1965),
.A2(n_1840),
.B(n_1837),
.Y(n_2066)
);

OAI21x1_ASAP7_75t_L g2067 ( 
.A1(n_2011),
.A2(n_1858),
.B(n_1833),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_1981),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2014),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1967),
.Y(n_2070)
);

INVx4_ASAP7_75t_L g2071 ( 
.A(n_1994),
.Y(n_2071)
);

AOI22xp33_ASAP7_75t_L g2072 ( 
.A1(n_1995),
.A2(n_1868),
.B1(n_1816),
.B2(n_1838),
.Y(n_2072)
);

OAI21xp5_ASAP7_75t_L g2073 ( 
.A1(n_2039),
.A2(n_1821),
.B(n_1883),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1952),
.Y(n_2074)
);

OAI21x1_ASAP7_75t_L g2075 ( 
.A1(n_1971),
.A2(n_1909),
.B(n_1903),
.Y(n_2075)
);

OAI21x1_ASAP7_75t_L g2076 ( 
.A1(n_1972),
.A2(n_1928),
.B(n_1918),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2015),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_1979),
.Y(n_2078)
);

AOI22xp33_ASAP7_75t_L g2079 ( 
.A1(n_1978),
.A2(n_1960),
.B1(n_2002),
.B2(n_1953),
.Y(n_2079)
);

OAI21x1_ASAP7_75t_L g2080 ( 
.A1(n_1991),
.A2(n_1836),
.B(n_1920),
.Y(n_2080)
);

OAI21x1_ASAP7_75t_L g2081 ( 
.A1(n_1996),
.A2(n_1916),
.B(n_1808),
.Y(n_2081)
);

OAI21x1_ASAP7_75t_L g2082 ( 
.A1(n_2007),
.A2(n_1843),
.B(n_1886),
.Y(n_2082)
);

OAI21x1_ASAP7_75t_L g2083 ( 
.A1(n_2018),
.A2(n_1871),
.B(n_1834),
.Y(n_2083)
);

AOI21xp5_ASAP7_75t_L g2084 ( 
.A1(n_2005),
.A2(n_1904),
.B(n_1778),
.Y(n_2084)
);

OR2x2_ASAP7_75t_L g2085 ( 
.A(n_1963),
.B(n_1904),
.Y(n_2085)
);

BUFx6f_ASAP7_75t_L g2086 ( 
.A(n_1973),
.Y(n_2086)
);

HB1xp67_ASAP7_75t_L g2087 ( 
.A(n_1992),
.Y(n_2087)
);

AOI221xp5_ASAP7_75t_L g2088 ( 
.A1(n_2028),
.A2(n_1777),
.B1(n_302),
.B2(n_303),
.C(n_304),
.Y(n_2088)
);

AND2x4_ASAP7_75t_L g2089 ( 
.A(n_1989),
.B(n_301),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2009),
.Y(n_2090)
);

BUFx6f_ASAP7_75t_L g2091 ( 
.A(n_2026),
.Y(n_2091)
);

OAI21x1_ASAP7_75t_L g2092 ( 
.A1(n_2019),
.A2(n_502),
.B(n_560),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2037),
.Y(n_2093)
);

OAI21xp5_ASAP7_75t_L g2094 ( 
.A1(n_2012),
.A2(n_2000),
.B(n_2016),
.Y(n_2094)
);

OA21x2_ASAP7_75t_L g2095 ( 
.A1(n_2034),
.A2(n_302),
.B(n_303),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2003),
.Y(n_2096)
);

NOR2xp33_ASAP7_75t_L g2097 ( 
.A(n_1961),
.B(n_304),
.Y(n_2097)
);

OAI21xp33_ASAP7_75t_L g2098 ( 
.A1(n_2079),
.A2(n_2024),
.B(n_2013),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_2054),
.Y(n_2099)
);

OA21x2_ASAP7_75t_L g2100 ( 
.A1(n_2047),
.A2(n_1999),
.B(n_2008),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_2054),
.Y(n_2101)
);

INVx8_ASAP7_75t_L g2102 ( 
.A(n_2091),
.Y(n_2102)
);

AND2x2_ASAP7_75t_L g2103 ( 
.A(n_2054),
.B(n_1986),
.Y(n_2103)
);

CKINVDCx5p33_ASAP7_75t_R g2104 ( 
.A(n_2042),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_2078),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2068),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2068),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_2050),
.B(n_1986),
.Y(n_2108)
);

INVx3_ASAP7_75t_L g2109 ( 
.A(n_2047),
.Y(n_2109)
);

BUFx3_ASAP7_75t_L g2110 ( 
.A(n_2049),
.Y(n_2110)
);

BUFx2_ASAP7_75t_L g2111 ( 
.A(n_2087),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_SL g2112 ( 
.A(n_2049),
.B(n_1946),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_2075),
.Y(n_2113)
);

AOI22xp33_ASAP7_75t_SL g2114 ( 
.A1(n_2066),
.A2(n_1946),
.B1(n_2036),
.B2(n_2008),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_2050),
.B(n_1986),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_2075),
.Y(n_2116)
);

AOI22xp33_ASAP7_75t_L g2117 ( 
.A1(n_2051),
.A2(n_1998),
.B1(n_2033),
.B2(n_2025),
.Y(n_2117)
);

INVx2_ASAP7_75t_SL g2118 ( 
.A(n_2040),
.Y(n_2118)
);

BUFx3_ASAP7_75t_L g2119 ( 
.A(n_2091),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_2043),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2053),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_2043),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_2059),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2060),
.Y(n_2124)
);

INVx1_ASAP7_75t_SL g2125 ( 
.A(n_2062),
.Y(n_2125)
);

BUFx2_ASAP7_75t_R g2126 ( 
.A(n_2085),
.Y(n_2126)
);

INVx6_ASAP7_75t_L g2127 ( 
.A(n_2041),
.Y(n_2127)
);

AOI22xp33_ASAP7_75t_L g2128 ( 
.A1(n_2046),
.A2(n_2023),
.B1(n_2029),
.B2(n_1984),
.Y(n_2128)
);

INVx3_ASAP7_75t_L g2129 ( 
.A(n_2061),
.Y(n_2129)
);

AOI22xp33_ASAP7_75t_SL g2130 ( 
.A1(n_2066),
.A2(n_2006),
.B1(n_1990),
.B2(n_2038),
.Y(n_2130)
);

AOI22xp33_ASAP7_75t_SL g2131 ( 
.A1(n_2108),
.A2(n_2066),
.B1(n_2095),
.B2(n_2055),
.Y(n_2131)
);

OAI22xp5_ASAP7_75t_L g2132 ( 
.A1(n_2098),
.A2(n_2057),
.B1(n_2044),
.B2(n_2084),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_2105),
.Y(n_2133)
);

OAI21xp33_ASAP7_75t_L g2134 ( 
.A1(n_2098),
.A2(n_2073),
.B(n_2094),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2123),
.Y(n_2135)
);

AOI22xp33_ASAP7_75t_L g2136 ( 
.A1(n_2130),
.A2(n_2095),
.B1(n_2088),
.B2(n_2072),
.Y(n_2136)
);

AOI22xp33_ASAP7_75t_L g2137 ( 
.A1(n_2130),
.A2(n_2095),
.B1(n_2056),
.B2(n_2055),
.Y(n_2137)
);

CKINVDCx5p33_ASAP7_75t_R g2138 ( 
.A(n_2104),
.Y(n_2138)
);

INVx3_ASAP7_75t_L g2139 ( 
.A(n_2110),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2123),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2123),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_2105),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_2108),
.B(n_2077),
.Y(n_2143)
);

AOI22xp33_ASAP7_75t_L g2144 ( 
.A1(n_2114),
.A2(n_2055),
.B1(n_2096),
.B2(n_1980),
.Y(n_2144)
);

AOI22xp33_ASAP7_75t_L g2145 ( 
.A1(n_2114),
.A2(n_2027),
.B1(n_2021),
.B2(n_2070),
.Y(n_2145)
);

OAI21xp5_ASAP7_75t_SL g2146 ( 
.A1(n_2117),
.A2(n_2097),
.B(n_2089),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_2111),
.B(n_2090),
.Y(n_2147)
);

OAI22xp5_ASAP7_75t_L g2148 ( 
.A1(n_2117),
.A2(n_2057),
.B1(n_2089),
.B2(n_2045),
.Y(n_2148)
);

AOI22xp33_ASAP7_75t_SL g2149 ( 
.A1(n_2108),
.A2(n_2083),
.B1(n_2089),
.B2(n_2082),
.Y(n_2149)
);

BUFx3_ASAP7_75t_R g2150 ( 
.A(n_2111),
.Y(n_2150)
);

AOI22xp33_ASAP7_75t_L g2151 ( 
.A1(n_2115),
.A2(n_2083),
.B1(n_2076),
.B2(n_2010),
.Y(n_2151)
);

AOI22xp33_ASAP7_75t_L g2152 ( 
.A1(n_2115),
.A2(n_2076),
.B1(n_2074),
.B2(n_2082),
.Y(n_2152)
);

NAND2xp33_ASAP7_75t_R g2153 ( 
.A(n_2138),
.B(n_2111),
.Y(n_2153)
);

AND2x4_ASAP7_75t_L g2154 ( 
.A(n_2139),
.B(n_2110),
.Y(n_2154)
);

AND2x4_ASAP7_75t_L g2155 ( 
.A(n_2139),
.B(n_2110),
.Y(n_2155)
);

NAND2xp33_ASAP7_75t_R g2156 ( 
.A(n_2138),
.B(n_2115),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_2134),
.B(n_2125),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_2134),
.B(n_2125),
.Y(n_2158)
);

AND2x4_ASAP7_75t_L g2159 ( 
.A(n_2139),
.B(n_2110),
.Y(n_2159)
);

NAND2x1p5_ASAP7_75t_L g2160 ( 
.A(n_2147),
.B(n_2091),
.Y(n_2160)
);

BUFx10_ASAP7_75t_L g2161 ( 
.A(n_2150),
.Y(n_2161)
);

CKINVDCx5p33_ASAP7_75t_R g2162 ( 
.A(n_2132),
.Y(n_2162)
);

AND2x2_ASAP7_75t_L g2163 ( 
.A(n_2161),
.B(n_2147),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_2157),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2158),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_2162),
.B(n_2143),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_2160),
.Y(n_2167)
);

AND2x2_ASAP7_75t_L g2168 ( 
.A(n_2159),
.B(n_2149),
.Y(n_2168)
);

INVxp67_ASAP7_75t_SL g2169 ( 
.A(n_2166),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2164),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_2163),
.B(n_2154),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_2164),
.Y(n_2172)
);

INVx1_ASAP7_75t_SL g2173 ( 
.A(n_2166),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2165),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_2168),
.B(n_2154),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_2167),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2164),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_2163),
.B(n_2155),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_SL g2179 ( 
.A(n_2173),
.B(n_2155),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_SL g2180 ( 
.A(n_2169),
.B(n_2159),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2174),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_2174),
.B(n_2146),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_2175),
.B(n_2118),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_2175),
.B(n_2118),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_2176),
.B(n_2152),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_2171),
.B(n_2118),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2171),
.B(n_2178),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2170),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2170),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2181),
.Y(n_2190)
);

AND2x4_ASAP7_75t_L g2191 ( 
.A(n_2187),
.B(n_2178),
.Y(n_2191)
);

OR2x2_ASAP7_75t_L g2192 ( 
.A(n_2182),
.B(n_2176),
.Y(n_2192)
);

AND2x2_ASAP7_75t_L g2193 ( 
.A(n_2184),
.B(n_1966),
.Y(n_2193)
);

OR2x2_ASAP7_75t_L g2194 ( 
.A(n_2180),
.B(n_2177),
.Y(n_2194)
);

HB1xp67_ASAP7_75t_L g2195 ( 
.A(n_2180),
.Y(n_2195)
);

OR2x2_ASAP7_75t_L g2196 ( 
.A(n_2179),
.B(n_2177),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2188),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2195),
.Y(n_2198)
);

INVxp67_ASAP7_75t_SL g2199 ( 
.A(n_2192),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2190),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_2191),
.B(n_2184),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_2201),
.B(n_2191),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_2199),
.B(n_2194),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2198),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_2201),
.B(n_2196),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2203),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2202),
.B(n_2198),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_2205),
.Y(n_2208)
);

AOI21xp5_ASAP7_75t_L g2209 ( 
.A1(n_2204),
.A2(n_2179),
.B(n_2193),
.Y(n_2209)
);

AOI22xp5_ASAP7_75t_L g2210 ( 
.A1(n_2203),
.A2(n_2185),
.B1(n_2189),
.B2(n_2156),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2207),
.Y(n_2211)
);

AOI21xp5_ASAP7_75t_L g2212 ( 
.A1(n_2209),
.A2(n_2200),
.B(n_2197),
.Y(n_2212)
);

AOI21xp5_ASAP7_75t_L g2213 ( 
.A1(n_2208),
.A2(n_2183),
.B(n_2186),
.Y(n_2213)
);

INVx1_ASAP7_75t_SL g2214 ( 
.A(n_2206),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_2210),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_2208),
.B(n_2186),
.Y(n_2216)
);

OAI22xp33_ASAP7_75t_L g2217 ( 
.A1(n_2210),
.A2(n_2172),
.B1(n_2153),
.B2(n_2148),
.Y(n_2217)
);

OAI221xp5_ASAP7_75t_L g2218 ( 
.A1(n_2210),
.A2(n_2172),
.B1(n_2131),
.B2(n_2137),
.C(n_2136),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_2208),
.B(n_2062),
.Y(n_2219)
);

AOI22xp5_ASAP7_75t_L g2220 ( 
.A1(n_2210),
.A2(n_1942),
.B1(n_2112),
.B2(n_2128),
.Y(n_2220)
);

OAI22xp5_ASAP7_75t_L g2221 ( 
.A1(n_2212),
.A2(n_1940),
.B1(n_2128),
.B2(n_2144),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2216),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2211),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2219),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2214),
.Y(n_2225)
);

NOR2xp33_ASAP7_75t_L g2226 ( 
.A(n_2213),
.B(n_1982),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_2215),
.Y(n_2227)
);

OR2x2_ASAP7_75t_L g2228 ( 
.A(n_2220),
.B(n_2020),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2218),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_2217),
.B(n_2112),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2216),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2214),
.B(n_2001),
.Y(n_2232)
);

INVxp67_ASAP7_75t_L g2233 ( 
.A(n_2211),
.Y(n_2233)
);

NOR2xp33_ASAP7_75t_L g2234 ( 
.A(n_2225),
.B(n_2126),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2232),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2223),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_2233),
.B(n_2151),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2227),
.Y(n_2238)
);

NAND3x1_ASAP7_75t_L g2239 ( 
.A(n_2222),
.B(n_2150),
.C(n_2093),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2231),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_SL g2241 ( 
.A(n_2226),
.B(n_2035),
.Y(n_2241)
);

AOI221xp5_ASAP7_75t_L g2242 ( 
.A1(n_2221),
.A2(n_2022),
.B1(n_2103),
.B2(n_2145),
.C(n_2113),
.Y(n_2242)
);

AOI211xp5_ASAP7_75t_L g2243 ( 
.A1(n_2221),
.A2(n_1974),
.B(n_2103),
.C(n_2080),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_2224),
.B(n_2085),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_2229),
.B(n_2135),
.Y(n_2245)
);

NAND3xp33_ASAP7_75t_SL g2246 ( 
.A(n_2230),
.B(n_1988),
.C(n_1985),
.Y(n_2246)
);

AOI21xp5_ASAP7_75t_L g2247 ( 
.A1(n_2234),
.A2(n_2228),
.B(n_2109),
.Y(n_2247)
);

AOI21xp5_ASAP7_75t_L g2248 ( 
.A1(n_2236),
.A2(n_2109),
.B(n_2103),
.Y(n_2248)
);

NAND3xp33_ASAP7_75t_L g2249 ( 
.A(n_2238),
.B(n_2004),
.C(n_2031),
.Y(n_2249)
);

A2O1A1Ixp33_ASAP7_75t_L g2250 ( 
.A1(n_2237),
.A2(n_2080),
.B(n_2081),
.C(n_2067),
.Y(n_2250)
);

AOI31xp33_ASAP7_75t_L g2251 ( 
.A1(n_2240),
.A2(n_2235),
.A3(n_2241),
.B(n_2243),
.Y(n_2251)
);

NAND3xp33_ASAP7_75t_L g2252 ( 
.A(n_2245),
.B(n_2032),
.C(n_2031),
.Y(n_2252)
);

OAI21xp5_ASAP7_75t_SL g2253 ( 
.A1(n_2246),
.A2(n_2091),
.B(n_2032),
.Y(n_2253)
);

AOI221xp5_ASAP7_75t_L g2254 ( 
.A1(n_2242),
.A2(n_2113),
.B1(n_2116),
.B2(n_2140),
.C(n_2135),
.Y(n_2254)
);

O2A1O1Ixp33_ASAP7_75t_L g2255 ( 
.A1(n_2244),
.A2(n_1957),
.B(n_1990),
.C(n_2100),
.Y(n_2255)
);

NOR2x1_ASAP7_75t_L g2256 ( 
.A(n_2239),
.B(n_305),
.Y(n_2256)
);

NOR4xp25_ASAP7_75t_L g2257 ( 
.A(n_2238),
.B(n_2140),
.C(n_2141),
.D(n_2116),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_2238),
.B(n_2141),
.Y(n_2258)
);

AND2x2_ASAP7_75t_L g2259 ( 
.A(n_2256),
.B(n_2126),
.Y(n_2259)
);

AOI21xp5_ASAP7_75t_L g2260 ( 
.A1(n_2251),
.A2(n_305),
.B(n_307),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_2252),
.B(n_1983),
.Y(n_2261)
);

AND2x2_ASAP7_75t_L g2262 ( 
.A(n_2247),
.B(n_2119),
.Y(n_2262)
);

AOI21xp5_ASAP7_75t_L g2263 ( 
.A1(n_2258),
.A2(n_307),
.B(n_308),
.Y(n_2263)
);

NOR2xp33_ASAP7_75t_L g2264 ( 
.A(n_2253),
.B(n_1957),
.Y(n_2264)
);

AOI221xp5_ASAP7_75t_SL g2265 ( 
.A1(n_2248),
.A2(n_2099),
.B1(n_2101),
.B2(n_2109),
.C(n_2121),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_2257),
.B(n_2119),
.Y(n_2266)
);

OAI21xp33_ASAP7_75t_L g2267 ( 
.A1(n_2249),
.A2(n_2017),
.B(n_2119),
.Y(n_2267)
);

AOI21xp33_ASAP7_75t_L g2268 ( 
.A1(n_2255),
.A2(n_308),
.B(n_309),
.Y(n_2268)
);

AND4x1_ASAP7_75t_L g2269 ( 
.A(n_2254),
.B(n_309),
.C(n_310),
.D(n_311),
.Y(n_2269)
);

O2A1O1Ixp5_ASAP7_75t_L g2270 ( 
.A1(n_2250),
.A2(n_2109),
.B(n_2129),
.C(n_2101),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2256),
.Y(n_2271)
);

AOI211xp5_ASAP7_75t_L g2272 ( 
.A1(n_2247),
.A2(n_2081),
.B(n_2092),
.C(n_1973),
.Y(n_2272)
);

OAI211xp5_ASAP7_75t_L g2273 ( 
.A1(n_2256),
.A2(n_310),
.B(n_311),
.C(n_312),
.Y(n_2273)
);

AOI21xp33_ASAP7_75t_SL g2274 ( 
.A1(n_2271),
.A2(n_312),
.B(n_313),
.Y(n_2274)
);

AOI21xp33_ASAP7_75t_L g2275 ( 
.A1(n_2273),
.A2(n_313),
.B(n_314),
.Y(n_2275)
);

AOI222xp33_ASAP7_75t_L g2276 ( 
.A1(n_2259),
.A2(n_1990),
.B1(n_2048),
.B2(n_2116),
.C1(n_2113),
.C2(n_2092),
.Y(n_2276)
);

NAND4xp25_ASAP7_75t_L g2277 ( 
.A(n_2260),
.B(n_2119),
.C(n_315),
.D(n_316),
.Y(n_2277)
);

NAND3xp33_ASAP7_75t_L g2278 ( 
.A(n_2263),
.B(n_1973),
.C(n_2113),
.Y(n_2278)
);

AOI211xp5_ASAP7_75t_L g2279 ( 
.A1(n_2267),
.A2(n_314),
.B(n_316),
.C(n_317),
.Y(n_2279)
);

AOI21xp33_ASAP7_75t_SL g2280 ( 
.A1(n_2268),
.A2(n_317),
.B(n_318),
.Y(n_2280)
);

AOI321xp33_ASAP7_75t_L g2281 ( 
.A1(n_2262),
.A2(n_2116),
.A3(n_2099),
.B1(n_2101),
.B2(n_2109),
.C(n_2122),
.Y(n_2281)
);

AOI221xp5_ASAP7_75t_L g2282 ( 
.A1(n_2266),
.A2(n_2270),
.B1(n_2264),
.B2(n_2261),
.C(n_2272),
.Y(n_2282)
);

AOI222xp33_ASAP7_75t_L g2283 ( 
.A1(n_2269),
.A2(n_2142),
.B1(n_2133),
.B2(n_2067),
.C1(n_2121),
.C2(n_2124),
.Y(n_2283)
);

NOR2x1_ASAP7_75t_L g2284 ( 
.A(n_2265),
.B(n_319),
.Y(n_2284)
);

AOI31xp33_ASAP7_75t_L g2285 ( 
.A1(n_2260),
.A2(n_319),
.A3(n_320),
.B(n_321),
.Y(n_2285)
);

AOI221xp5_ASAP7_75t_L g2286 ( 
.A1(n_2267),
.A2(n_2124),
.B1(n_2064),
.B2(n_2069),
.C(n_2120),
.Y(n_2286)
);

OAI211xp5_ASAP7_75t_L g2287 ( 
.A1(n_2260),
.A2(n_320),
.B(n_321),
.C(n_322),
.Y(n_2287)
);

OAI221xp5_ASAP7_75t_L g2288 ( 
.A1(n_2267),
.A2(n_2100),
.B1(n_2129),
.B2(n_2099),
.C(n_2101),
.Y(n_2288)
);

OAI21xp33_ASAP7_75t_L g2289 ( 
.A1(n_2259),
.A2(n_2099),
.B(n_2129),
.Y(n_2289)
);

AND2x2_ASAP7_75t_SL g2290 ( 
.A(n_2271),
.B(n_2071),
.Y(n_2290)
);

OAI211xp5_ASAP7_75t_SL g2291 ( 
.A1(n_2271),
.A2(n_322),
.B(n_323),
.C(n_324),
.Y(n_2291)
);

AOI21xp33_ASAP7_75t_L g2292 ( 
.A1(n_2271),
.A2(n_323),
.B(n_324),
.Y(n_2292)
);

NOR2xp33_ASAP7_75t_R g2293 ( 
.A(n_2271),
.B(n_325),
.Y(n_2293)
);

NAND3xp33_ASAP7_75t_SL g2294 ( 
.A(n_2271),
.B(n_325),
.C(n_326),
.Y(n_2294)
);

O2A1O1Ixp33_ASAP7_75t_L g2295 ( 
.A1(n_2271),
.A2(n_326),
.B(n_328),
.C(n_329),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2274),
.B(n_328),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_2285),
.B(n_329),
.Y(n_2297)
);

OAI21xp33_ASAP7_75t_L g2298 ( 
.A1(n_2277),
.A2(n_2129),
.B(n_2123),
.Y(n_2298)
);

NOR3xp33_ASAP7_75t_L g2299 ( 
.A(n_2294),
.B(n_330),
.C(n_331),
.Y(n_2299)
);

NOR2xp33_ASAP7_75t_L g2300 ( 
.A(n_2291),
.B(n_330),
.Y(n_2300)
);

NOR3xp33_ASAP7_75t_L g2301 ( 
.A(n_2292),
.B(n_331),
.C(n_332),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2284),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_2293),
.B(n_332),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_2280),
.B(n_333),
.Y(n_2304)
);

AND2x2_ASAP7_75t_L g2305 ( 
.A(n_2290),
.B(n_2279),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2295),
.Y(n_2306)
);

NAND4xp75_ASAP7_75t_L g2307 ( 
.A(n_2275),
.B(n_334),
.C(n_335),
.D(n_336),
.Y(n_2307)
);

HB1xp67_ASAP7_75t_L g2308 ( 
.A(n_2287),
.Y(n_2308)
);

NOR2x1_ASAP7_75t_L g2309 ( 
.A(n_2278),
.B(n_335),
.Y(n_2309)
);

AOI22xp33_ASAP7_75t_L g2310 ( 
.A1(n_2282),
.A2(n_2100),
.B1(n_2142),
.B2(n_2133),
.Y(n_2310)
);

AOI21xp5_ASAP7_75t_L g2311 ( 
.A1(n_2289),
.A2(n_336),
.B(n_337),
.Y(n_2311)
);

AND2x2_ASAP7_75t_L g2312 ( 
.A(n_2283),
.B(n_2129),
.Y(n_2312)
);

OA21x2_ASAP7_75t_L g2313 ( 
.A1(n_2303),
.A2(n_2286),
.B(n_2288),
.Y(n_2313)
);

NAND3xp33_ASAP7_75t_L g2314 ( 
.A(n_2302),
.B(n_2281),
.C(n_2276),
.Y(n_2314)
);

AOI21xp5_ASAP7_75t_L g2315 ( 
.A1(n_2296),
.A2(n_2297),
.B(n_2305),
.Y(n_2315)
);

NOR2xp33_ASAP7_75t_L g2316 ( 
.A(n_2308),
.B(n_337),
.Y(n_2316)
);

NOR3xp33_ASAP7_75t_SL g2317 ( 
.A(n_2306),
.B(n_338),
.C(n_339),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2300),
.B(n_338),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2304),
.Y(n_2319)
);

NOR3xp33_ASAP7_75t_L g2320 ( 
.A(n_2301),
.B(n_339),
.C(n_340),
.Y(n_2320)
);

AND3x4_ASAP7_75t_L g2321 ( 
.A(n_2299),
.B(n_341),
.C(n_342),
.Y(n_2321)
);

NOR2x1_ASAP7_75t_L g2322 ( 
.A(n_2307),
.B(n_341),
.Y(n_2322)
);

NOR2x1_ASAP7_75t_L g2323 ( 
.A(n_2309),
.B(n_343),
.Y(n_2323)
);

NOR3xp33_ASAP7_75t_L g2324 ( 
.A(n_2311),
.B(n_343),
.C(n_344),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_2298),
.B(n_2100),
.Y(n_2325)
);

NOR2xp33_ASAP7_75t_L g2326 ( 
.A(n_2312),
.B(n_344),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2310),
.Y(n_2327)
);

NOR2xp33_ASAP7_75t_L g2328 ( 
.A(n_2302),
.B(n_345),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2302),
.Y(n_2329)
);

NOR3xp33_ASAP7_75t_L g2330 ( 
.A(n_2303),
.B(n_345),
.C(n_495),
.Y(n_2330)
);

NAND4xp75_ASAP7_75t_L g2331 ( 
.A(n_2329),
.B(n_2100),
.C(n_498),
.D(n_500),
.Y(n_2331)
);

OAI322xp33_ASAP7_75t_L g2332 ( 
.A1(n_2326),
.A2(n_2122),
.A3(n_2120),
.B1(n_2086),
.B2(n_2071),
.C1(n_2106),
.C2(n_2107),
.Y(n_2332)
);

AND2x4_ASAP7_75t_L g2333 ( 
.A(n_2315),
.B(n_2071),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2323),
.B(n_1979),
.Y(n_2334)
);

INVx2_ASAP7_75t_SL g2335 ( 
.A(n_2322),
.Y(n_2335)
);

AOI221xp5_ASAP7_75t_L g2336 ( 
.A1(n_2314),
.A2(n_2122),
.B1(n_2120),
.B2(n_2086),
.C(n_2102),
.Y(n_2336)
);

BUFx3_ASAP7_75t_L g2337 ( 
.A(n_2328),
.Y(n_2337)
);

NOR4xp25_ASAP7_75t_L g2338 ( 
.A(n_2319),
.B(n_2122),
.C(n_2120),
.D(n_504),
.Y(n_2338)
);

OAI22xp5_ASAP7_75t_L g2339 ( 
.A1(n_2316),
.A2(n_2127),
.B1(n_2100),
.B2(n_2102),
.Y(n_2339)
);

NAND3xp33_ASAP7_75t_L g2340 ( 
.A(n_2317),
.B(n_2086),
.C(n_501),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2321),
.Y(n_2341)
);

NOR3xp33_ASAP7_75t_L g2342 ( 
.A(n_2318),
.B(n_496),
.C(n_505),
.Y(n_2342)
);

AND2x2_ASAP7_75t_L g2343 ( 
.A(n_2320),
.B(n_2127),
.Y(n_2343)
);

AOI211xp5_ASAP7_75t_L g2344 ( 
.A1(n_2327),
.A2(n_2086),
.B(n_2065),
.C(n_2063),
.Y(n_2344)
);

NOR2xp33_ASAP7_75t_R g2345 ( 
.A(n_2335),
.B(n_2324),
.Y(n_2345)
);

XNOR2xp5_ASAP7_75t_L g2346 ( 
.A(n_2341),
.B(n_2330),
.Y(n_2346)
);

NAND2xp33_ASAP7_75t_SL g2347 ( 
.A(n_2333),
.B(n_2325),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_SL g2348 ( 
.A(n_2340),
.B(n_2313),
.Y(n_2348)
);

NOR2xp33_ASAP7_75t_R g2349 ( 
.A(n_2337),
.B(n_2313),
.Y(n_2349)
);

NOR2xp33_ASAP7_75t_R g2350 ( 
.A(n_2343),
.B(n_506),
.Y(n_2350)
);

AND4x1_ASAP7_75t_L g2351 ( 
.A(n_2342),
.B(n_507),
.C(n_509),
.D(n_511),
.Y(n_2351)
);

NAND2xp33_ASAP7_75t_SL g2352 ( 
.A(n_2334),
.B(n_2086),
.Y(n_2352)
);

NAND3xp33_ASAP7_75t_L g2353 ( 
.A(n_2338),
.B(n_516),
.C(n_517),
.Y(n_2353)
);

NOR2xp33_ASAP7_75t_R g2354 ( 
.A(n_2331),
.B(n_518),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_2336),
.B(n_1979),
.Y(n_2355)
);

NOR3xp33_ASAP7_75t_SL g2356 ( 
.A(n_2332),
.B(n_2339),
.C(n_2344),
.Y(n_2356)
);

NOR2xp33_ASAP7_75t_R g2357 ( 
.A(n_2335),
.B(n_520),
.Y(n_2357)
);

XNOR2xp5_ASAP7_75t_L g2358 ( 
.A(n_2341),
.B(n_522),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2349),
.Y(n_2359)
);

INVx3_ASAP7_75t_L g2360 ( 
.A(n_2351),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2353),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2348),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2358),
.Y(n_2363)
);

AOI22xp5_ASAP7_75t_L g2364 ( 
.A1(n_2347),
.A2(n_2065),
.B1(n_2102),
.B2(n_2127),
.Y(n_2364)
);

INVxp67_ASAP7_75t_SL g2365 ( 
.A(n_2346),
.Y(n_2365)
);

AND2x2_ASAP7_75t_L g2366 ( 
.A(n_2354),
.B(n_2127),
.Y(n_2366)
);

INVx3_ASAP7_75t_L g2367 ( 
.A(n_2357),
.Y(n_2367)
);

BUFx2_ASAP7_75t_L g2368 ( 
.A(n_2359),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2362),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2367),
.Y(n_2370)
);

XNOR2xp5_ASAP7_75t_L g2371 ( 
.A(n_2365),
.B(n_2356),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2367),
.Y(n_2372)
);

OAI22xp5_ASAP7_75t_L g2373 ( 
.A1(n_2366),
.A2(n_2355),
.B1(n_2345),
.B2(n_2352),
.Y(n_2373)
);

XOR2xp5_ASAP7_75t_L g2374 ( 
.A(n_2363),
.B(n_2350),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2360),
.Y(n_2375)
);

OAI22xp5_ASAP7_75t_L g2376 ( 
.A1(n_2369),
.A2(n_2361),
.B1(n_2364),
.B2(n_2127),
.Y(n_2376)
);

CKINVDCx20_ASAP7_75t_R g2377 ( 
.A(n_2371),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_SL g2378 ( 
.A(n_2368),
.B(n_1970),
.Y(n_2378)
);

OAI21xp5_ASAP7_75t_L g2379 ( 
.A1(n_2375),
.A2(n_2063),
.B(n_2058),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2374),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_2377),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_2380),
.Y(n_2382)
);

OAI22xp5_ASAP7_75t_SL g2383 ( 
.A1(n_2376),
.A2(n_2372),
.B1(n_2370),
.B2(n_2373),
.Y(n_2383)
);

OAI22xp5_ASAP7_75t_SL g2384 ( 
.A1(n_2381),
.A2(n_2378),
.B1(n_2379),
.B2(n_2127),
.Y(n_2384)
);

AO21x2_ASAP7_75t_L g2385 ( 
.A1(n_2384),
.A2(n_2382),
.B(n_2383),
.Y(n_2385)
);

XNOR2xp5_ASAP7_75t_L g2386 ( 
.A(n_2385),
.B(n_523),
.Y(n_2386)
);

AOI22xp5_ASAP7_75t_L g2387 ( 
.A1(n_2385),
.A2(n_2102),
.B1(n_2052),
.B2(n_2041),
.Y(n_2387)
);

NAND3xp33_ASAP7_75t_L g2388 ( 
.A(n_2386),
.B(n_524),
.C(n_525),
.Y(n_2388)
);

OAI21xp5_ASAP7_75t_L g2389 ( 
.A1(n_2387),
.A2(n_527),
.B(n_528),
.Y(n_2389)
);

AOI21xp5_ASAP7_75t_L g2390 ( 
.A1(n_2388),
.A2(n_530),
.B(n_534),
.Y(n_2390)
);

AOI22x1_ASAP7_75t_L g2391 ( 
.A1(n_2390),
.A2(n_2389),
.B1(n_537),
.B2(n_538),
.Y(n_2391)
);

AOI221xp5_ASAP7_75t_L g2392 ( 
.A1(n_2391),
.A2(n_535),
.B1(n_544),
.B2(n_546),
.C(n_548),
.Y(n_2392)
);

AOI21xp5_ASAP7_75t_L g2393 ( 
.A1(n_2392),
.A2(n_549),
.B(n_551),
.Y(n_2393)
);

AOI22xp33_ASAP7_75t_SL g2394 ( 
.A1(n_2393),
.A2(n_2102),
.B1(n_553),
.B2(n_554),
.Y(n_2394)
);


endmodule