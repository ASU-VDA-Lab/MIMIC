module fake_netlist_6_270_n_852 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_852);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_852;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_222;
wire n_300;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_272;
wire n_526;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_722;
wire n_688;
wire n_351;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_817;
wire n_701;
wire n_629;
wire n_388;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_508;
wire n_361;
wire n_663;
wire n_379;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_664;
wire n_678;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g200 ( 
.A(n_51),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_89),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_195),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_110),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g204 ( 
.A(n_29),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_176),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_46),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_77),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_100),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_141),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_101),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_0),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_153),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_166),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_93),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_136),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_105),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_146),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_54),
.Y(n_218)
);

NOR2xp67_ASAP7_75t_L g219 ( 
.A(n_115),
.B(n_130),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_124),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_120),
.Y(n_221)
);

BUFx5_ASAP7_75t_L g222 ( 
.A(n_111),
.Y(n_222)
);

NOR2xp67_ASAP7_75t_L g223 ( 
.A(n_64),
.B(n_155),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_104),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_38),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_139),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_70),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_13),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_126),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_161),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_42),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_88),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_87),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_169),
.Y(n_234)
);

NOR2xp67_ASAP7_75t_L g235 ( 
.A(n_148),
.B(n_66),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_31),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_196),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_83),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_106),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_2),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_18),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_52),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_67),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_192),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_154),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_114),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_49),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_84),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_150),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_44),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_159),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_99),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_48),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_103),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_164),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_73),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_185),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_171),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_98),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_183),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_47),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_129),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_79),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_39),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_119),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_157),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_61),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_102),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_68),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_187),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_144),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_190),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_147),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_15),
.B(n_82),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_156),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_199),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_74),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_28),
.Y(n_278)
);

BUFx12f_ASAP7_75t_L g279 ( 
.A(n_270),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_236),
.B(n_0),
.Y(n_280)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_273),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_273),
.Y(n_282)
);

BUFx12f_ASAP7_75t_L g283 ( 
.A(n_228),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_240),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_216),
.Y(n_285)
);

BUFx8_ASAP7_75t_L g286 ( 
.A(n_274),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_241),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_211),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_204),
.Y(n_289)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_273),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_204),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_200),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_204),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_249),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_201),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_204),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_215),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_204),
.Y(n_298)
);

OAI22x1_ASAP7_75t_R g299 ( 
.A1(n_211),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_273),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g301 ( 
.A(n_278),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_202),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_207),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_203),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_229),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_231),
.B(n_272),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_215),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_230),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_204),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_222),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_222),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_210),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_243),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_212),
.Y(n_314)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_205),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_213),
.Y(n_316)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_206),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_224),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_260),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_238),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_266),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_222),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_242),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_237),
.B(n_4),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_246),
.Y(n_325)
);

AND2x4_ASAP7_75t_L g326 ( 
.A(n_251),
.B(n_23),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_222),
.B(n_5),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_255),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_257),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_222),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_304),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_315),
.B(n_317),
.Y(n_332)
);

AOI21x1_ASAP7_75t_L g333 ( 
.A1(n_327),
.A2(n_261),
.B(n_259),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_301),
.B(n_208),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_285),
.B(n_209),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_282),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_282),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_282),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_282),
.Y(n_339)
);

BUFx6f_ASAP7_75t_SL g340 ( 
.A(n_326),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_300),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_300),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_300),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_300),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_304),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_315),
.B(n_263),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_306),
.B(n_214),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_304),
.Y(n_348)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_304),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_308),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_285),
.B(n_277),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_324),
.A2(n_225),
.B1(n_239),
.B2(n_252),
.Y(n_352)
);

AOI21x1_ASAP7_75t_L g353 ( 
.A1(n_289),
.A2(n_271),
.B(n_264),
.Y(n_353)
);

AOI21x1_ASAP7_75t_L g354 ( 
.A1(n_289),
.A2(n_293),
.B(n_291),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_301),
.B(n_217),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_306),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_285),
.B(n_218),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_308),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_315),
.B(n_275),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_308),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_308),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_313),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_313),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_313),
.Y(n_364)
);

INVx2_ASAP7_75t_SL g365 ( 
.A(n_294),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_286),
.B(n_220),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_313),
.Y(n_367)
);

INVx8_ASAP7_75t_L g368 ( 
.A(n_281),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_294),
.B(n_295),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_319),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_319),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_319),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_319),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_321),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_321),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_321),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_317),
.B(n_276),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_321),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_326),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_323),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_284),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_326),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_379),
.B(n_330),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_360),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_379),
.B(n_330),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_349),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_349),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_379),
.B(n_291),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_382),
.B(n_293),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_360),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_382),
.B(n_296),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_382),
.B(n_296),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_365),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_356),
.B(n_317),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_331),
.Y(n_395)
);

AO221x1_ASAP7_75t_L g396 ( 
.A1(n_349),
.A2(n_329),
.B1(n_294),
.B2(n_325),
.C(n_323),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_331),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_357),
.B(n_281),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_357),
.B(n_281),
.Y(n_399)
);

OAI221xp5_ASAP7_75t_L g400 ( 
.A1(n_381),
.A2(n_305),
.B1(n_280),
.B2(n_292),
.C(n_302),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_371),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_356),
.B(n_286),
.Y(n_402)
);

O2A1O1Ixp33_ASAP7_75t_L g403 ( 
.A1(n_381),
.A2(n_316),
.B(n_312),
.C(n_314),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_369),
.B(n_334),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_371),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_331),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_371),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_352),
.B(n_286),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_345),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_R g410 ( 
.A(n_333),
.B(n_297),
.Y(n_410)
);

NAND2xp33_ASAP7_75t_SL g411 ( 
.A(n_340),
.B(n_297),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_370),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_345),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_370),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_334),
.B(n_279),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_355),
.B(n_279),
.Y(n_416)
);

NAND2xp33_ASAP7_75t_L g417 ( 
.A(n_355),
.B(n_222),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_335),
.B(n_290),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_348),
.Y(n_419)
);

INVxp33_ASAP7_75t_L g420 ( 
.A(n_369),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_332),
.B(n_280),
.Y(n_421)
);

OR2x2_ASAP7_75t_L g422 ( 
.A(n_335),
.B(n_288),
.Y(n_422)
);

NOR3xp33_ASAP7_75t_L g423 ( 
.A(n_347),
.B(n_307),
.C(n_303),
.Y(n_423)
);

OR2x2_ASAP7_75t_L g424 ( 
.A(n_351),
.B(n_307),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_359),
.B(n_283),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_366),
.A2(n_283),
.B1(n_221),
.B2(n_226),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_351),
.B(n_290),
.Y(n_427)
);

NOR2x1p5_ASAP7_75t_L g428 ( 
.A(n_346),
.B(n_287),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_377),
.B(n_227),
.Y(n_429)
);

BUFx5_ASAP7_75t_L g430 ( 
.A(n_338),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_348),
.B(n_318),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_372),
.B(n_290),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_333),
.B(n_232),
.Y(n_433)
);

NAND3xp33_ASAP7_75t_L g434 ( 
.A(n_373),
.B(n_320),
.C(n_323),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_380),
.B(n_233),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_380),
.B(n_234),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_340),
.A2(n_262),
.B1(n_244),
.B2(n_245),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_374),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_350),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_350),
.B(n_247),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_358),
.B(n_248),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_374),
.B(n_298),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_358),
.B(n_329),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_375),
.B(n_298),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_375),
.B(n_378),
.Y(n_445)
);

A2O1A1Ixp33_ASAP7_75t_L g446 ( 
.A1(n_404),
.A2(n_219),
.B(n_223),
.C(n_235),
.Y(n_446)
);

AOI33xp33_ASAP7_75t_L g447 ( 
.A1(n_394),
.A2(n_299),
.A3(n_309),
.B1(n_310),
.B2(n_311),
.B3(n_322),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_422),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_421),
.B(n_378),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_420),
.B(n_250),
.Y(n_450)
);

OAI21xp33_ASAP7_75t_L g451 ( 
.A1(n_400),
.A2(n_254),
.B(n_253),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_424),
.B(n_256),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_383),
.A2(n_354),
.B(n_353),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_393),
.B(n_340),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_383),
.B(n_361),
.Y(n_455)
);

OAI321xp33_ASAP7_75t_L g456 ( 
.A1(n_426),
.A2(n_353),
.A3(n_354),
.B1(n_328),
.B2(n_323),
.C(n_325),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_385),
.B(n_362),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_385),
.A2(n_368),
.B(n_363),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_388),
.B(n_362),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_428),
.A2(n_258),
.B1(n_265),
.B2(n_267),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_415),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_388),
.B(n_363),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_389),
.A2(n_368),
.B(n_376),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_389),
.B(n_364),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_395),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_443),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_391),
.A2(n_368),
.B(n_376),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_425),
.B(n_437),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_391),
.A2(n_367),
.B(n_364),
.Y(n_469)
);

AOI21x1_ASAP7_75t_L g470 ( 
.A1(n_433),
.A2(n_339),
.B(n_338),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_445),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_392),
.B(n_367),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_392),
.B(n_336),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_398),
.A2(n_368),
.B(n_337),
.Y(n_474)
);

AOI22xp33_ASAP7_75t_L g475 ( 
.A1(n_417),
.A2(n_328),
.B1(n_325),
.B2(n_310),
.Y(n_475)
);

OAI21xp33_ASAP7_75t_L g476 ( 
.A1(n_408),
.A2(n_269),
.B(n_268),
.Y(n_476)
);

INVx5_ASAP7_75t_L g477 ( 
.A(n_395),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_410),
.B(n_325),
.Y(n_478)
);

AND2x2_ASAP7_75t_SL g479 ( 
.A(n_423),
.B(n_431),
.Y(n_479)
);

O2A1O1Ixp33_ASAP7_75t_SL g480 ( 
.A1(n_399),
.A2(n_309),
.B(n_311),
.C(n_322),
.Y(n_480)
);

OAI21xp33_ASAP7_75t_L g481 ( 
.A1(n_416),
.A2(n_328),
.B(n_339),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_418),
.A2(n_368),
.B(n_337),
.Y(n_482)
);

OAI321xp33_ASAP7_75t_L g483 ( 
.A1(n_437),
.A2(n_328),
.A3(n_342),
.B1(n_341),
.B2(n_336),
.C(n_344),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_427),
.A2(n_342),
.B(n_341),
.Y(n_484)
);

CKINVDCx6p67_ASAP7_75t_R g485 ( 
.A(n_402),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_445),
.A2(n_444),
.B(n_442),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_384),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_442),
.A2(n_344),
.B(n_343),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_390),
.B(n_343),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_412),
.B(n_343),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_411),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_409),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_444),
.Y(n_493)
);

INVx2_ASAP7_75t_SL g494 ( 
.A(n_440),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_441),
.A2(n_344),
.B(n_107),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_414),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_429),
.B(n_395),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_438),
.B(n_24),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_397),
.B(n_5),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_397),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_L g501 ( 
.A1(n_396),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_413),
.A2(n_108),
.B(n_197),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_435),
.B(n_6),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_436),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_419),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_397),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_439),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_406),
.Y(n_508)
);

AO21x1_ASAP7_75t_L g509 ( 
.A1(n_386),
.A2(n_387),
.B(n_401),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_406),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_486),
.A2(n_432),
.B(n_406),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_453),
.A2(n_407),
.B(n_405),
.Y(n_512)
);

O2A1O1Ixp5_ASAP7_75t_L g513 ( 
.A1(n_509),
.A2(n_468),
.B(n_449),
.C(n_478),
.Y(n_513)
);

OA22x2_ASAP7_75t_L g514 ( 
.A1(n_448),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_514)
);

OAI21x1_ASAP7_75t_L g515 ( 
.A1(n_470),
.A2(n_434),
.B(n_403),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_487),
.B(n_25),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_455),
.A2(n_430),
.B(n_112),
.Y(n_517)
);

OAI21x1_ASAP7_75t_L g518 ( 
.A1(n_469),
.A2(n_463),
.B(n_458),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_479),
.B(n_430),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_SL g520 ( 
.A1(n_502),
.A2(n_430),
.B(n_113),
.Y(n_520)
);

A2O1A1Ixp33_ASAP7_75t_L g521 ( 
.A1(n_471),
.A2(n_430),
.B(n_10),
.C(n_11),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_496),
.Y(n_522)
);

OAI21x1_ASAP7_75t_L g523 ( 
.A1(n_467),
.A2(n_430),
.B(n_109),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_493),
.B(n_9),
.Y(n_524)
);

O2A1O1Ixp5_ASAP7_75t_L g525 ( 
.A1(n_497),
.A2(n_116),
.B(n_194),
.C(n_193),
.Y(n_525)
);

AO21x1_ASAP7_75t_L g526 ( 
.A1(n_503),
.A2(n_498),
.B(n_459),
.Y(n_526)
);

OAI21x1_ASAP7_75t_L g527 ( 
.A1(n_484),
.A2(n_198),
.B(n_96),
.Y(n_527)
);

AND2x6_ASAP7_75t_L g528 ( 
.A(n_454),
.B(n_26),
.Y(n_528)
);

AOI221x1_ASAP7_75t_L g529 ( 
.A1(n_446),
.A2(n_97),
.B1(n_189),
.B2(n_188),
.C(n_186),
.Y(n_529)
);

OAI21x1_ASAP7_75t_L g530 ( 
.A1(n_474),
.A2(n_94),
.B(n_184),
.Y(n_530)
);

OAI21x1_ASAP7_75t_L g531 ( 
.A1(n_473),
.A2(n_462),
.B(n_457),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_466),
.B(n_10),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g533 ( 
.A1(n_464),
.A2(n_191),
.B(n_92),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_472),
.A2(n_91),
.B(n_181),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_461),
.B(n_27),
.Y(n_535)
);

AOI21xp33_ASAP7_75t_L g536 ( 
.A1(n_451),
.A2(n_11),
.B(n_12),
.Y(n_536)
);

OAI21x1_ASAP7_75t_L g537 ( 
.A1(n_482),
.A2(n_182),
.B(n_95),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_485),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_494),
.B(n_30),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_500),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_505),
.Y(n_541)
);

OAI21x1_ASAP7_75t_L g542 ( 
.A1(n_488),
.A2(n_117),
.B(n_179),
.Y(n_542)
);

AO31x2_ASAP7_75t_L g543 ( 
.A1(n_495),
.A2(n_12),
.A3(n_13),
.B(n_14),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_507),
.B(n_14),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_492),
.Y(n_545)
);

AOI21x1_ASAP7_75t_L g546 ( 
.A1(n_489),
.A2(n_490),
.B(n_450),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_452),
.B(n_15),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_491),
.Y(n_548)
);

CKINVDCx8_ASAP7_75t_R g549 ( 
.A(n_500),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_465),
.B(n_16),
.Y(n_550)
);

OA21x2_ASAP7_75t_L g551 ( 
.A1(n_456),
.A2(n_121),
.B(n_178),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_465),
.B(n_16),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_504),
.B(n_17),
.Y(n_553)
);

INVxp67_ASAP7_75t_SL g554 ( 
.A(n_500),
.Y(n_554)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_477),
.A2(n_118),
.B(n_177),
.Y(n_555)
);

OAI21x1_ASAP7_75t_L g556 ( 
.A1(n_475),
.A2(n_180),
.B(n_90),
.Y(n_556)
);

OAI21x1_ASAP7_75t_SL g557 ( 
.A1(n_501),
.A2(n_86),
.B(n_175),
.Y(n_557)
);

OAI21x1_ASAP7_75t_SL g558 ( 
.A1(n_460),
.A2(n_85),
.B(n_174),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_506),
.B(n_17),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_510),
.B(n_32),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_506),
.Y(n_561)
);

AOI21x1_ASAP7_75t_SL g562 ( 
.A1(n_483),
.A2(n_18),
.B(n_19),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_460),
.B(n_33),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_L g564 ( 
.A1(n_476),
.A2(n_123),
.B(n_173),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_506),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_477),
.A2(n_122),
.B(n_172),
.Y(n_566)
);

OAI21x1_ASAP7_75t_L g567 ( 
.A1(n_523),
.A2(n_499),
.B(n_481),
.Y(n_567)
);

AO21x2_ASAP7_75t_L g568 ( 
.A1(n_526),
.A2(n_480),
.B(n_508),
.Y(n_568)
);

OA21x2_ASAP7_75t_L g569 ( 
.A1(n_518),
.A2(n_512),
.B(n_531),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_536),
.A2(n_508),
.B1(n_447),
.B2(n_477),
.Y(n_570)
);

INVx2_ASAP7_75t_SL g571 ( 
.A(n_541),
.Y(n_571)
);

NAND3xp33_ASAP7_75t_L g572 ( 
.A(n_547),
.B(n_508),
.C(n_20),
.Y(n_572)
);

OAI21x1_ASAP7_75t_L g573 ( 
.A1(n_511),
.A2(n_81),
.B(n_170),
.Y(n_573)
);

OAI21x1_ASAP7_75t_L g574 ( 
.A1(n_546),
.A2(n_80),
.B(n_168),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_538),
.Y(n_575)
);

AOI22x1_ASAP7_75t_L g576 ( 
.A1(n_517),
.A2(n_78),
.B1(n_167),
.B2(n_165),
.Y(n_576)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_548),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g578 ( 
.A(n_553),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_522),
.Y(n_579)
);

OAI21x1_ASAP7_75t_SL g580 ( 
.A1(n_557),
.A2(n_76),
.B(n_163),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_L g581 ( 
.A1(n_513),
.A2(n_75),
.B(n_162),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_545),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_545),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_R g584 ( 
.A(n_549),
.B(n_72),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g585 ( 
.A(n_540),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_520),
.A2(n_71),
.B(n_160),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_563),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_587)
);

OAI21x1_ASAP7_75t_L g588 ( 
.A1(n_515),
.A2(n_125),
.B(n_158),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_524),
.B(n_21),
.Y(n_589)
);

OAI21x1_ASAP7_75t_L g590 ( 
.A1(n_530),
.A2(n_127),
.B(n_34),
.Y(n_590)
);

OAI21x1_ASAP7_75t_L g591 ( 
.A1(n_542),
.A2(n_128),
.B(n_35),
.Y(n_591)
);

OA21x2_ASAP7_75t_L g592 ( 
.A1(n_527),
.A2(n_131),
.B(n_36),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_540),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_519),
.B(n_132),
.Y(n_594)
);

AOI21xp33_ASAP7_75t_L g595 ( 
.A1(n_532),
.A2(n_22),
.B(n_37),
.Y(n_595)
);

OAI21x1_ASAP7_75t_L g596 ( 
.A1(n_537),
.A2(n_133),
.B(n_40),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_561),
.Y(n_597)
);

AO21x2_ASAP7_75t_L g598 ( 
.A1(n_564),
.A2(n_134),
.B(n_41),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_565),
.Y(n_599)
);

OAI21x1_ASAP7_75t_L g600 ( 
.A1(n_562),
.A2(n_135),
.B(n_43),
.Y(n_600)
);

OAI21x1_ASAP7_75t_L g601 ( 
.A1(n_556),
.A2(n_533),
.B(n_525),
.Y(n_601)
);

OA21x2_ASAP7_75t_L g602 ( 
.A1(n_529),
.A2(n_137),
.B(n_45),
.Y(n_602)
);

OAI21x1_ASAP7_75t_L g603 ( 
.A1(n_550),
.A2(n_138),
.B(n_50),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_544),
.Y(n_604)
);

OAI21xp5_ASAP7_75t_L g605 ( 
.A1(n_552),
.A2(n_140),
.B(n_53),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_516),
.B(n_22),
.Y(n_606)
);

OAI21x1_ASAP7_75t_L g607 ( 
.A1(n_558),
.A2(n_55),
.B(n_56),
.Y(n_607)
);

BUFx8_ASAP7_75t_L g608 ( 
.A(n_528),
.Y(n_608)
);

OAI21x1_ASAP7_75t_L g609 ( 
.A1(n_551),
.A2(n_57),
.B(n_58),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_559),
.Y(n_610)
);

BUFx2_ASAP7_75t_SL g611 ( 
.A(n_516),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_593),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_579),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_583),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_583),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_582),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_597),
.Y(n_617)
);

OA21x2_ASAP7_75t_L g618 ( 
.A1(n_581),
.A2(n_521),
.B(n_534),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_573),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_597),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_577),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_599),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_600),
.Y(n_623)
);

AO21x1_ASAP7_75t_SL g624 ( 
.A1(n_605),
.A2(n_528),
.B(n_551),
.Y(n_624)
);

OAI21x1_ASAP7_75t_L g625 ( 
.A1(n_574),
.A2(n_566),
.B(n_555),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_571),
.Y(n_626)
);

BUFx2_ASAP7_75t_L g627 ( 
.A(n_593),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_600),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_568),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_568),
.Y(n_630)
);

BUFx2_ASAP7_75t_L g631 ( 
.A(n_585),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_610),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_606),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_604),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_611),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_570),
.B(n_589),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_609),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_589),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_572),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_570),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_609),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_594),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_594),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_578),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_573),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_587),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_567),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_587),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_567),
.Y(n_649)
);

NAND2x1p5_ASAP7_75t_L g650 ( 
.A(n_607),
.B(n_588),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_SL g651 ( 
.A1(n_608),
.A2(n_528),
.B1(n_514),
.B2(n_560),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_603),
.Y(n_652)
);

INVxp67_ASAP7_75t_SL g653 ( 
.A(n_644),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_615),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_631),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_636),
.B(n_543),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_615),
.B(n_607),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_638),
.B(n_560),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_636),
.B(n_543),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_612),
.Y(n_660)
);

HB1xp67_ASAP7_75t_L g661 ( 
.A(n_621),
.Y(n_661)
);

HB1xp67_ASAP7_75t_L g662 ( 
.A(n_626),
.Y(n_662)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_646),
.B(n_569),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_626),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_614),
.B(n_640),
.Y(n_665)
);

BUFx2_ASAP7_75t_L g666 ( 
.A(n_631),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_629),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_620),
.B(n_543),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_620),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_617),
.B(n_602),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_634),
.B(n_535),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_629),
.Y(n_672)
);

HB1xp67_ASAP7_75t_L g673 ( 
.A(n_627),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_616),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_613),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_630),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_642),
.B(n_591),
.Y(n_677)
);

OR2x2_ASAP7_75t_L g678 ( 
.A(n_648),
.B(n_569),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_632),
.B(n_528),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_639),
.B(n_602),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g681 ( 
.A(n_627),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_643),
.A2(n_595),
.B1(n_598),
.B2(n_539),
.Y(n_682)
);

INVx4_ASAP7_75t_L g683 ( 
.A(n_612),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_622),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_SL g685 ( 
.A1(n_618),
.A2(n_598),
.B(n_602),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_637),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_633),
.B(n_603),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_630),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_612),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_651),
.B(n_596),
.Y(n_690)
);

OR2x2_ASAP7_75t_L g691 ( 
.A(n_652),
.B(n_569),
.Y(n_691)
);

AND2x4_ASAP7_75t_L g692 ( 
.A(n_635),
.B(n_554),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_623),
.B(n_596),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_623),
.B(n_592),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_628),
.B(n_592),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_612),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_628),
.B(n_592),
.Y(n_697)
);

HB1xp67_ASAP7_75t_L g698 ( 
.A(n_612),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_689),
.B(n_641),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_673),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_689),
.B(n_641),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_660),
.Y(n_702)
);

OAI22xp5_ASAP7_75t_L g703 ( 
.A1(n_658),
.A2(n_575),
.B1(n_618),
.B2(n_586),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_656),
.B(n_649),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_653),
.B(n_575),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_671),
.B(n_608),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_686),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_656),
.B(n_649),
.Y(n_708)
);

NOR2xp67_ASAP7_75t_L g709 ( 
.A(n_661),
.B(n_619),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_660),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_662),
.B(n_608),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_667),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_667),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_672),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_682),
.A2(n_618),
.B1(n_624),
.B2(n_576),
.Y(n_715)
);

OR2x2_ASAP7_75t_L g716 ( 
.A(n_655),
.B(n_666),
.Y(n_716)
);

INVx2_ASAP7_75t_SL g717 ( 
.A(n_681),
.Y(n_717)
);

OR2x2_ASAP7_75t_L g718 ( 
.A(n_655),
.B(n_647),
.Y(n_718)
);

OR2x2_ASAP7_75t_L g719 ( 
.A(n_666),
.B(n_647),
.Y(n_719)
);

INVxp67_ASAP7_75t_SL g720 ( 
.A(n_664),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_686),
.Y(n_721)
);

INVxp67_ASAP7_75t_SL g722 ( 
.A(n_669),
.Y(n_722)
);

BUFx2_ASAP7_75t_L g723 ( 
.A(n_660),
.Y(n_723)
);

HB1xp67_ASAP7_75t_L g724 ( 
.A(n_698),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_659),
.B(n_645),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_675),
.B(n_584),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_672),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_675),
.B(n_584),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_659),
.B(n_645),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_674),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_660),
.Y(n_731)
);

INVx4_ASAP7_75t_L g732 ( 
.A(n_660),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_674),
.Y(n_733)
);

INVxp67_ASAP7_75t_SL g734 ( 
.A(n_669),
.Y(n_734)
);

INVxp67_ASAP7_75t_L g735 ( 
.A(n_684),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_668),
.B(n_687),
.Y(n_736)
);

OR2x6_ASAP7_75t_L g737 ( 
.A(n_703),
.B(n_685),
.Y(n_737)
);

HB1xp67_ASAP7_75t_L g738 ( 
.A(n_712),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_720),
.B(n_684),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_713),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_736),
.B(n_687),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_736),
.B(n_668),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_714),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_727),
.Y(n_744)
);

OR2x2_ASAP7_75t_L g745 ( 
.A(n_716),
.B(n_678),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_707),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_725),
.B(n_678),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_730),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_724),
.B(n_690),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_735),
.B(n_665),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_733),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_718),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_719),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_725),
.B(n_663),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_729),
.B(n_663),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_700),
.B(n_690),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_729),
.B(n_680),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_707),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_704),
.B(n_680),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_721),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_704),
.B(n_691),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_705),
.Y(n_762)
);

NAND2x1p5_ASAP7_75t_SL g763 ( 
.A(n_700),
.B(n_670),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_721),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_741),
.B(n_717),
.Y(n_765)
);

OR2x2_ASAP7_75t_L g766 ( 
.A(n_741),
.B(n_717),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_738),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_746),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_738),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_740),
.Y(n_770)
);

OR2x2_ASAP7_75t_L g771 ( 
.A(n_745),
.B(n_708),
.Y(n_771)
);

OR2x2_ASAP7_75t_L g772 ( 
.A(n_752),
.B(n_708),
.Y(n_772)
);

O2A1O1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_762),
.A2(n_726),
.B(n_728),
.C(n_706),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_753),
.B(n_734),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_743),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_742),
.B(n_731),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_737),
.A2(n_706),
.B1(n_715),
.B2(n_679),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_746),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_777),
.A2(n_737),
.B1(n_756),
.B2(n_749),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_770),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_775),
.Y(n_781)
);

AOI211x1_ASAP7_75t_L g782 ( 
.A1(n_774),
.A2(n_711),
.B(n_739),
.C(n_750),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_767),
.Y(n_783)
);

OAI22xp33_ASAP7_75t_SL g784 ( 
.A1(n_777),
.A2(n_737),
.B1(n_744),
.B2(n_748),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_769),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_768),
.Y(n_786)
);

AOI32xp33_ASAP7_75t_L g787 ( 
.A1(n_776),
.A2(n_742),
.A3(n_774),
.B1(n_759),
.B2(n_757),
.Y(n_787)
);

INVxp67_ASAP7_75t_L g788 ( 
.A(n_765),
.Y(n_788)
);

NOR2x1_ASAP7_75t_SL g789 ( 
.A(n_780),
.B(n_766),
.Y(n_789)
);

AOI221xp5_ASAP7_75t_L g790 ( 
.A1(n_782),
.A2(n_773),
.B1(n_763),
.B2(n_751),
.C(n_715),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_787),
.B(n_772),
.Y(n_791)
);

OAI22xp5_ASAP7_75t_L g792 ( 
.A1(n_779),
.A2(n_771),
.B1(n_709),
.B2(n_732),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_784),
.A2(n_755),
.B1(n_747),
.B2(n_754),
.Y(n_793)
);

NAND3xp33_ASAP7_75t_L g794 ( 
.A(n_790),
.B(n_785),
.C(n_783),
.Y(n_794)
);

OA21x2_ASAP7_75t_L g795 ( 
.A1(n_791),
.A2(n_781),
.B(n_786),
.Y(n_795)
);

OAI221xp5_ASAP7_75t_L g796 ( 
.A1(n_793),
.A2(n_784),
.B1(n_788),
.B2(n_778),
.C(n_764),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_789),
.Y(n_797)
);

AOI221xp5_ASAP7_75t_L g798 ( 
.A1(n_792),
.A2(n_763),
.B1(n_685),
.B2(n_692),
.C(n_758),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_790),
.A2(n_760),
.B(n_692),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_794),
.Y(n_800)
);

NOR2xp67_ASAP7_75t_L g801 ( 
.A(n_797),
.B(n_732),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_796),
.B(n_692),
.Y(n_802)
);

OAI21xp33_ASAP7_75t_L g803 ( 
.A1(n_798),
.A2(n_761),
.B(n_755),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_800),
.A2(n_795),
.B(n_799),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_802),
.Y(n_805)
);

OAI322xp33_ASAP7_75t_L g806 ( 
.A1(n_803),
.A2(n_759),
.A3(n_757),
.B1(n_761),
.B2(n_754),
.C1(n_747),
.C2(n_654),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_806),
.Y(n_807)
);

NAND3xp33_ASAP7_75t_L g808 ( 
.A(n_804),
.B(n_801),
.C(n_683),
.Y(n_808)
);

NAND4xp75_ASAP7_75t_L g809 ( 
.A(n_805),
.B(n_665),
.C(n_654),
.D(n_693),
.Y(n_809)
);

NAND4xp75_ASAP7_75t_L g810 ( 
.A(n_804),
.B(n_693),
.C(n_670),
.D(n_695),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_807),
.B(n_689),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_809),
.Y(n_812)
);

A2O1A1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_808),
.A2(n_710),
.B(n_696),
.C(n_590),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_810),
.B(n_723),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_808),
.B(n_696),
.Y(n_815)
);

AO22x2_ASAP7_75t_L g816 ( 
.A1(n_807),
.A2(n_683),
.B1(n_580),
.B2(n_732),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_807),
.B(n_710),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_811),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_817),
.A2(n_696),
.B1(n_683),
.B2(n_702),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_812),
.A2(n_702),
.B1(n_677),
.B2(n_701),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_816),
.B(n_702),
.Y(n_821)
);

NAND2xp33_ASAP7_75t_L g822 ( 
.A(n_814),
.B(n_702),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_SL g823 ( 
.A1(n_815),
.A2(n_650),
.B1(n_540),
.B2(n_722),
.Y(n_823)
);

NOR2x1_ASAP7_75t_L g824 ( 
.A(n_813),
.B(n_816),
.Y(n_824)
);

NAND4xp75_ASAP7_75t_L g825 ( 
.A(n_817),
.B(n_694),
.C(n_695),
.D(n_697),
.Y(n_825)
);

AO22x2_ASAP7_75t_L g826 ( 
.A1(n_818),
.A2(n_677),
.B1(n_699),
.B2(n_701),
.Y(n_826)
);

XNOR2xp5_ASAP7_75t_L g827 ( 
.A(n_819),
.B(n_59),
.Y(n_827)
);

OAI22xp5_ASAP7_75t_L g828 ( 
.A1(n_820),
.A2(n_701),
.B1(n_699),
.B2(n_677),
.Y(n_828)
);

OAI22x1_ASAP7_75t_SL g829 ( 
.A1(n_822),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_824),
.A2(n_677),
.B1(n_699),
.B2(n_657),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_821),
.Y(n_831)
);

NAND3xp33_ASAP7_75t_L g832 ( 
.A(n_823),
.B(n_657),
.C(n_619),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_825),
.Y(n_833)
);

AOI31xp33_ASAP7_75t_L g834 ( 
.A1(n_831),
.A2(n_650),
.A3(n_657),
.B(n_142),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_833),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_829),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_827),
.Y(n_837)
);

OR2x2_ASAP7_75t_L g838 ( 
.A(n_830),
.B(n_65),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_832),
.A2(n_657),
.B1(n_676),
.B2(n_688),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_836),
.B(n_826),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_835),
.A2(n_828),
.B1(n_624),
.B2(n_676),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_837),
.A2(n_838),
.B1(n_839),
.B2(n_834),
.Y(n_842)
);

OAI22xp5_ASAP7_75t_L g843 ( 
.A1(n_836),
.A2(n_688),
.B1(n_691),
.B2(n_650),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_836),
.A2(n_619),
.B1(n_694),
.B2(n_697),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_842),
.B(n_69),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_840),
.A2(n_625),
.B(n_601),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_843),
.A2(n_625),
.B(n_637),
.Y(n_847)
);

AOI22xp5_ASAP7_75t_L g848 ( 
.A1(n_845),
.A2(n_844),
.B1(n_841),
.B2(n_149),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_846),
.Y(n_849)
);

NAND2x1_ASAP7_75t_L g850 ( 
.A(n_848),
.B(n_847),
.Y(n_850)
);

AOI21x1_ASAP7_75t_L g851 ( 
.A1(n_850),
.A2(n_849),
.B(n_145),
.Y(n_851)
);

AOI31xp33_ASAP7_75t_L g852 ( 
.A1(n_851),
.A2(n_143),
.A3(n_151),
.B(n_152),
.Y(n_852)
);


endmodule