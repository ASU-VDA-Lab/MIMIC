module fake_jpeg_30936_n_470 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_470);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_470;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx2_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx6f_ASAP7_75t_SL g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_52),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_54),
.Y(n_120)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

AOI21xp33_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_15),
.B(n_2),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_58),
.B(n_86),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_59),
.Y(n_139)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_60),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_61),
.Y(n_150)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_63),
.Y(n_141)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_7),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_66),
.B(n_49),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_68),
.Y(n_135)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_69),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_71),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_74),
.Y(n_160)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_78),
.Y(n_140)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_16),
.Y(n_80)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_81),
.Y(n_162)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_82),
.Y(n_145)
);

BUFx10_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_83),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_84),
.Y(n_153)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_39),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_89),
.Y(n_159)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_19),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_90),
.Y(n_152)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_16),
.Y(n_91)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_93),
.Y(n_111)
);

BUFx12_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_23),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_17),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_95),
.Y(n_161)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_24),
.B(n_9),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_99),
.Y(n_125)
);

BUFx10_ASAP7_75t_L g98 ( 
.A(n_23),
.Y(n_98)
);

INVx6_ASAP7_75t_SL g113 ( 
.A(n_98),
.Y(n_113)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_27),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_24),
.B(n_9),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_100),
.B(n_37),
.Y(n_146)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_27),
.Y(n_101)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_27),
.Y(n_102)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_73),
.A2(n_29),
.B1(n_35),
.B2(n_31),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_107),
.A2(n_83),
.B1(n_0),
.B2(n_3),
.Y(n_204)
);

INVx6_ASAP7_75t_SL g122 ( 
.A(n_94),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_122),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_126),
.B(n_158),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_81),
.A2(n_34),
.B1(n_30),
.B2(n_41),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_133),
.A2(n_40),
.B1(n_30),
.B2(n_31),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_74),
.A2(n_29),
.B1(n_35),
.B2(n_49),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_134),
.A2(n_154),
.B1(n_113),
.B2(n_116),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_146),
.B(n_26),
.Y(n_171)
);

INVx6_ASAP7_75t_SL g151 ( 
.A(n_102),
.Y(n_151)
);

INVx13_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_84),
.A2(n_29),
.B1(n_35),
.B2(n_43),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_97),
.B(n_34),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_36),
.Y(n_173)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_100),
.Y(n_157)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_157),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_64),
.A2(n_41),
.B1(n_40),
.B2(n_37),
.Y(n_158)
);

A2O1A1Ixp33_ASAP7_75t_SL g233 ( 
.A1(n_163),
.A2(n_195),
.B(n_202),
.C(n_203),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_164),
.A2(n_189),
.B1(n_206),
.B2(n_107),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_165),
.Y(n_213)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_167),
.Y(n_225)
);

AOI32xp33_ASAP7_75t_L g168 ( 
.A1(n_105),
.A2(n_89),
.A3(n_88),
.B1(n_36),
.B2(n_43),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_168),
.B(n_183),
.Y(n_241)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_114),
.Y(n_169)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_169),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_109),
.Y(n_170)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_170),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_171),
.B(n_173),
.Y(n_227)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_124),
.Y(n_172)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_172),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_146),
.B(n_32),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_174),
.B(n_180),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_109),
.Y(n_176)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_176),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_126),
.B(n_26),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_185),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_117),
.Y(n_179)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_179),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_156),
.B(n_32),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_119),
.Y(n_182)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_182),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_105),
.B(n_17),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_129),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_184),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_125),
.B(n_54),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_130),
.Y(n_186)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_186),
.Y(n_236)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_142),
.Y(n_187)
);

INVx4_ASAP7_75t_SL g216 ( 
.A(n_187),
.Y(n_216)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_123),
.Y(n_188)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_188),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_144),
.A2(n_53),
.B1(n_51),
.B2(n_59),
.Y(n_189)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_141),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_190),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_118),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_191),
.Y(n_223)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_143),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_192),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_160),
.A2(n_85),
.B1(n_77),
.B2(n_29),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

INVx11_ASAP7_75t_L g194 ( 
.A(n_132),
.Y(n_194)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_194),
.Y(n_248)
);

OAI21xp33_ASAP7_75t_L g195 ( 
.A1(n_125),
.A2(n_92),
.B(n_35),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_160),
.A2(n_72),
.B1(n_67),
.B2(n_68),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_196),
.Y(n_232)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_121),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_197),
.Y(n_246)
);

FAx1_ASAP7_75t_SL g198 ( 
.A(n_131),
.B(n_98),
.CI(n_93),
.CON(n_198),
.SN(n_198)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_199),
.Y(n_229)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_149),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_140),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_208),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_L g201 ( 
.A1(n_162),
.A2(n_61),
.B1(n_103),
.B2(n_98),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_201),
.A2(n_204),
.B1(n_110),
.B2(n_137),
.Y(n_217)
);

AO22x1_ASAP7_75t_SL g202 ( 
.A1(n_145),
.A2(n_83),
.B1(n_0),
.B2(n_3),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_147),
.Y(n_203)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_123),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_205),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_112),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_206)
);

A2O1A1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_111),
.A2(n_2),
.B(n_5),
.C(n_10),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_207),
.A2(n_134),
.B(n_154),
.Y(n_230)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_152),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_161),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_111),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_104),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_215),
.A2(n_244),
.B1(n_201),
.B2(n_172),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_217),
.A2(n_206),
.B1(n_164),
.B2(n_177),
.Y(n_254)
);

AOI22x1_ASAP7_75t_L g218 ( 
.A1(n_195),
.A2(n_128),
.B1(n_148),
.B2(n_159),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_218),
.B(n_155),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_181),
.A2(n_136),
.B(n_152),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_220),
.A2(n_247),
.B(n_203),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_181),
.A2(n_135),
.B1(n_106),
.B2(n_137),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_224),
.A2(n_228),
.B1(n_243),
.B2(n_153),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_204),
.A2(n_135),
.B1(n_106),
.B2(n_139),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_230),
.B(n_202),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_181),
.A2(n_150),
.B1(n_139),
.B2(n_120),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_L g244 ( 
.A1(n_185),
.A2(n_150),
.B1(n_120),
.B2(n_115),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_173),
.B(n_115),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_202),
.Y(n_255)
);

NOR2xp67_ASAP7_75t_SL g247 ( 
.A(n_166),
.B(n_108),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_182),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_250),
.B(n_261),
.Y(n_304)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_212),
.Y(n_251)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_251),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_252),
.A2(n_268),
.B(n_233),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_214),
.B(n_178),
.C(n_198),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_253),
.B(n_218),
.C(n_233),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_254),
.A2(n_270),
.B1(n_274),
.B2(n_276),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_255),
.B(n_258),
.Y(n_288)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_222),
.Y(n_256)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_256),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_257),
.A2(n_273),
.B1(n_278),
.B2(n_219),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_184),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_214),
.B(n_207),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_259),
.B(n_263),
.Y(n_291)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_212),
.Y(n_260)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_260),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_227),
.B(n_177),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_226),
.Y(n_262)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_262),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_220),
.B(n_198),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_226),
.Y(n_264)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_264),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_229),
.B(n_169),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_265),
.B(n_266),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_229),
.B(n_200),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_267),
.Y(n_303)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_216),
.Y(n_269)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_269),
.Y(n_305)
);

OAI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_232),
.A2(n_205),
.B1(n_188),
.B2(n_197),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_216),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_271),
.B(n_275),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_229),
.B(n_175),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_272),
.B(n_280),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_215),
.A2(n_187),
.B1(n_192),
.B2(n_170),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_237),
.B(n_241),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_232),
.A2(n_190),
.B1(n_191),
.B2(n_199),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_277),
.A2(n_221),
.B1(n_223),
.B2(n_217),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_244),
.A2(n_176),
.B1(n_194),
.B2(n_175),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_225),
.B(n_224),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_219),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_237),
.B(n_2),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_268),
.A2(n_230),
.B(n_221),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_282),
.A2(n_293),
.B(n_306),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_256),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_284),
.B(n_271),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_243),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_285),
.B(n_292),
.C(n_296),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_236),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_295),
.A2(n_282),
.B(n_306),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_259),
.B(n_233),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_297),
.B(n_274),
.Y(n_312)
);

CKINVDCx14_ASAP7_75t_R g326 ( 
.A(n_299),
.Y(n_326)
);

OA21x2_ASAP7_75t_L g300 ( 
.A1(n_265),
.A2(n_233),
.B(n_218),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_274),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_302),
.A2(n_276),
.B1(n_279),
.B2(n_273),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_266),
.A2(n_233),
.B(n_246),
.Y(n_306)
);

AO21x2_ASAP7_75t_L g307 ( 
.A1(n_255),
.A2(n_231),
.B(n_246),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_307),
.A2(n_278),
.B1(n_257),
.B2(n_262),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_253),
.B(n_242),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_308),
.B(n_251),
.C(n_269),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_281),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_309),
.B(n_314),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_310),
.A2(n_318),
.B(n_319),
.Y(n_339)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_281),
.Y(n_311)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_311),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_312),
.B(n_301),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_291),
.B(n_264),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_313),
.B(n_327),
.C(n_291),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_286),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_304),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_315),
.Y(n_354)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_286),
.Y(n_316)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_316),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_295),
.A2(n_280),
.B(n_275),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_320),
.A2(n_334),
.B1(n_302),
.B2(n_293),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_288),
.B(n_258),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_321),
.B(n_322),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_297),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_323),
.A2(n_294),
.B1(n_290),
.B2(n_287),
.Y(n_347)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_305),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_324),
.B(n_325),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_288),
.B(n_260),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_328),
.B(n_330),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_294),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_329),
.Y(n_338)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_305),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_283),
.Y(n_331)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_331),
.Y(n_353)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_303),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_333),
.B(n_284),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_289),
.A2(n_231),
.B1(n_240),
.B2(n_238),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_287),
.B(n_213),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_335),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_317),
.B(n_296),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_336),
.B(n_340),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_326),
.A2(n_289),
.B1(n_298),
.B2(n_290),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_337),
.A2(n_351),
.B1(n_335),
.B2(n_311),
.Y(n_385)
);

XNOR2x1_ASAP7_75t_L g341 ( 
.A(n_317),
.B(n_285),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_341),
.B(n_348),
.Y(n_376)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_343),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_317),
.B(n_308),
.C(n_292),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_344),
.B(n_352),
.C(n_360),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_345),
.A2(n_355),
.B1(n_323),
.B2(n_329),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_347),
.A2(n_362),
.B1(n_330),
.B2(n_324),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_327),
.B(n_301),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_350),
.B(n_356),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_326),
.A2(n_298),
.B1(n_307),
.B2(n_300),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_327),
.B(n_303),
.C(n_307),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_320),
.A2(n_307),
.B1(n_300),
.B2(n_283),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_313),
.B(n_307),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_313),
.B(n_248),
.C(n_234),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_319),
.A2(n_238),
.B1(n_240),
.B2(n_249),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_363),
.A2(n_347),
.B1(n_338),
.B2(n_356),
.Y(n_390)
);

XOR2x2_ASAP7_75t_L g365 ( 
.A(n_336),
.B(n_339),
.Y(n_365)
);

XNOR2x1_ASAP7_75t_L g398 ( 
.A(n_365),
.B(n_358),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_354),
.B(n_315),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_367),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_341),
.B(n_312),
.C(n_318),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_368),
.B(n_371),
.C(n_372),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_354),
.A2(n_332),
.B1(n_334),
.B2(n_310),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_369),
.A2(n_381),
.B1(n_385),
.B2(n_355),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_359),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_370),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_340),
.B(n_348),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_344),
.B(n_312),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_346),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_374),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_346),
.Y(n_377)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_377),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_342),
.B(n_328),
.Y(n_378)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_378),
.Y(n_399)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_361),
.Y(n_379)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_379),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_360),
.B(n_332),
.C(n_325),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_380),
.B(n_382),
.C(n_345),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_352),
.B(n_321),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_359),
.Y(n_383)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_383),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_357),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_384),
.B(n_361),
.Y(n_403)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_357),
.Y(n_386)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_386),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_388),
.B(n_392),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_390),
.A2(n_368),
.B1(n_364),
.B2(n_331),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_372),
.B(n_350),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_369),
.A2(n_339),
.B(n_349),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_393),
.A2(n_380),
.B(n_381),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_373),
.B(n_349),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_397),
.B(n_398),
.C(n_405),
.Y(n_408)
);

BUFx24_ASAP7_75t_SL g401 ( 
.A(n_375),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_401),
.B(n_366),
.Y(n_410)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_403),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_404),
.B(n_382),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_366),
.B(n_353),
.C(n_333),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_406),
.B(n_410),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_407),
.A2(n_364),
.B(n_392),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_387),
.B(n_377),
.Y(n_409)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_409),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_405),
.B(n_404),
.C(n_397),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_411),
.B(n_414),
.C(n_417),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_395),
.A2(n_374),
.B1(n_309),
.B2(n_314),
.Y(n_412)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_412),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_394),
.B(n_373),
.C(n_371),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_391),
.B(n_362),
.Y(n_415)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_415),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_399),
.B(n_316),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_416),
.B(n_420),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_394),
.B(n_365),
.C(n_376),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_393),
.A2(n_390),
.B1(n_391),
.B2(n_396),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_419),
.B(n_388),
.Y(n_424)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_424),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_413),
.A2(n_403),
.B1(n_396),
.B2(n_389),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_425),
.A2(n_10),
.B1(n_11),
.B2(n_14),
.Y(n_446)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_415),
.Y(n_426)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_426),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_407),
.A2(n_389),
.B1(n_400),
.B2(n_402),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_429),
.B(n_433),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_L g430 ( 
.A1(n_420),
.A2(n_398),
.B1(n_213),
.B2(n_222),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_430),
.B(n_408),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_411),
.B(n_418),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_432),
.B(n_434),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_414),
.B(n_376),
.C(n_239),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_SL g436 ( 
.A(n_434),
.B(n_417),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_436),
.B(n_443),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_423),
.A2(n_418),
.B(n_408),
.Y(n_437)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_437),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_440),
.B(n_427),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_425),
.B(n_239),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_442),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_427),
.B(n_5),
.C(n_10),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_429),
.B(n_5),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_444),
.B(n_422),
.Y(n_451)
);

OAI21x1_ASAP7_75t_L g445 ( 
.A1(n_431),
.A2(n_5),
.B(n_10),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_445),
.B(n_446),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_449),
.B(n_451),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_438),
.B(n_424),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_452),
.B(n_454),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_435),
.B(n_428),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_441),
.B(n_421),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_455),
.A2(n_439),
.B(n_426),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_457),
.B(n_458),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_448),
.A2(n_439),
.B1(n_421),
.B2(n_444),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_450),
.A2(n_442),
.B(n_433),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_460),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_447),
.B(n_448),
.C(n_453),
.Y(n_461)
);

A2O1A1Ixp33_ASAP7_75t_SL g463 ( 
.A1(n_461),
.A2(n_453),
.B(n_14),
.C(n_15),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_463),
.B(n_459),
.C(n_456),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_465),
.A2(n_466),
.B(n_462),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_464),
.B(n_459),
.C(n_14),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_467),
.B(n_15),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_468),
.B(n_11),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_469),
.B(n_14),
.Y(n_470)
);


endmodule