module fake_jpeg_9162_n_104 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_104);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_104;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_25),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_20),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_31),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_39),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_15),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_49),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_60),
.Y(n_73)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_53),
.Y(n_64)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_66),
.A2(n_71),
.B1(n_61),
.B2(n_59),
.Y(n_75)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_68),
.Y(n_78)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_72),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_75),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_72),
.A2(n_55),
.B1(n_54),
.B2(n_47),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_76),
.A2(n_79),
.B1(n_83),
.B2(n_8),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_0),
.Y(n_77)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_77),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_72),
.A2(n_46),
.B1(n_42),
.B2(n_43),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_72),
.A2(n_48),
.B1(n_3),
.B2(n_5),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_80),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_88),
.B(n_89),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_90),
.B(n_85),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_92),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_93),
.A2(n_84),
.B(n_91),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_78),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_74),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_96),
.B(n_81),
.Y(n_97)
);

AOI21x1_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_16),
.B(n_17),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_98),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_27),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_100),
.B(n_29),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_33),
.C(n_34),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_35),
.C(n_36),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_38),
.Y(n_104)
);


endmodule