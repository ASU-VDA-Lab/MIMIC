module fake_aes_8347_n_748 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_748);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_748;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_622;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_695;
wire n_625;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g83 ( .A(n_8), .Y(n_83) );
NOR2xp67_ASAP7_75t_L g84 ( .A(n_79), .B(n_49), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_8), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_64), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_37), .Y(n_87) );
CKINVDCx20_ASAP7_75t_R g88 ( .A(n_5), .Y(n_88) );
INVxp67_ASAP7_75t_SL g89 ( .A(n_22), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_15), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_34), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_12), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_41), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_43), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_27), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_58), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_14), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_20), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_28), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_19), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_73), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_62), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_40), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_57), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g105 ( .A(n_55), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_4), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_48), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_13), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_32), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_5), .Y(n_110) );
INVxp33_ASAP7_75t_L g111 ( .A(n_52), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_9), .Y(n_112) );
INVx1_ASAP7_75t_SL g113 ( .A(n_76), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_11), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_59), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_6), .Y(n_116) );
CKINVDCx16_ASAP7_75t_R g117 ( .A(n_16), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_25), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_61), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_1), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_24), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_71), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_70), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_31), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_56), .Y(n_125) );
BUFx3_ASAP7_75t_L g126 ( .A(n_51), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_80), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_39), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_74), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_45), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_53), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_68), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_63), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_94), .Y(n_134) );
INVxp67_ASAP7_75t_L g135 ( .A(n_85), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_126), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_117), .B(n_0), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_83), .B(n_0), .Y(n_138) );
OA21x2_ASAP7_75t_L g139 ( .A1(n_91), .A2(n_33), .B(n_81), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_91), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_94), .B(n_1), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_126), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_111), .B(n_2), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_93), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_109), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_109), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_121), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_121), .Y(n_148) );
AND2x4_ASAP7_75t_L g149 ( .A(n_83), .B(n_2), .Y(n_149) );
BUFx8_ASAP7_75t_L g150 ( .A(n_130), .Y(n_150) );
OAI22xp5_ASAP7_75t_SL g151 ( .A1(n_88), .A2(n_3), .B1(n_4), .B2(n_6), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_130), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_93), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_96), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_96), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_99), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_99), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_100), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_90), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_90), .B(n_3), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_106), .B(n_7), .Y(n_161) );
OAI22xp5_ASAP7_75t_L g162 ( .A1(n_97), .A2(n_7), .B1(n_9), .B2(n_10), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_100), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_122), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_122), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_92), .Y(n_166) );
INVx3_ASAP7_75t_L g167 ( .A(n_92), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_112), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_112), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_86), .Y(n_170) );
AND2x2_ASAP7_75t_SL g171 ( .A(n_105), .B(n_82), .Y(n_171) );
OAI22xp5_ASAP7_75t_SL g172 ( .A1(n_106), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_87), .B(n_13), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_101), .Y(n_174) );
INVx3_ASAP7_75t_L g175 ( .A(n_97), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_102), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_104), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_107), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_110), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_179) );
OAI22xp33_ASAP7_75t_L g180 ( .A1(n_179), .A2(n_110), .B1(n_114), .B2(n_108), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_140), .B(n_119), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_136), .Y(n_182) );
AOI22xp33_ASAP7_75t_L g183 ( .A1(n_138), .A2(n_114), .B1(n_116), .B2(n_120), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_170), .B(n_133), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_170), .B(n_133), .Y(n_185) );
NAND2x1p5_ASAP7_75t_L g186 ( .A(n_143), .B(n_115), .Y(n_186) );
BUFx10_ASAP7_75t_L g187 ( .A(n_171), .Y(n_187) );
INVx2_ASAP7_75t_SL g188 ( .A(n_150), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_138), .Y(n_189) );
OAI22xp33_ASAP7_75t_L g190 ( .A1(n_179), .A2(n_129), .B1(n_95), .B2(n_132), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_136), .Y(n_191) );
NAND3xp33_ASAP7_75t_L g192 ( .A(n_143), .B(n_132), .C(n_95), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_135), .B(n_118), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_136), .Y(n_194) );
OR2x2_ASAP7_75t_L g195 ( .A(n_137), .B(n_118), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_176), .B(n_131), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g197 ( .A1(n_138), .A2(n_123), .B1(n_124), .B2(n_125), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_140), .B(n_128), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_176), .B(n_128), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_138), .Y(n_200) );
INVx4_ASAP7_75t_SL g201 ( .A(n_136), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_171), .Y(n_202) );
INVxp67_ASAP7_75t_L g203 ( .A(n_137), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_136), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_149), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_144), .B(n_103), .Y(n_206) );
BUFx3_ASAP7_75t_L g207 ( .A(n_142), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_144), .B(n_127), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_154), .B(n_103), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_154), .B(n_127), .Y(n_210) );
AOI22xp33_ASAP7_75t_L g211 ( .A1(n_149), .A2(n_98), .B1(n_89), .B2(n_113), .Y(n_211) );
INVx1_ASAP7_75t_SL g212 ( .A(n_161), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_155), .B(n_98), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_136), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_149), .B(n_84), .Y(n_215) );
AND3x2_ASAP7_75t_L g216 ( .A(n_149), .B(n_17), .C(n_18), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_160), .Y(n_217) );
AND2x6_ASAP7_75t_L g218 ( .A(n_160), .B(n_78), .Y(n_218) );
BUFx2_ASAP7_75t_L g219 ( .A(n_171), .Y(n_219) );
BUFx8_ASAP7_75t_SL g220 ( .A(n_160), .Y(n_220) );
BUFx4f_ASAP7_75t_L g221 ( .A(n_160), .Y(n_221) );
AND2x2_ASAP7_75t_L g222 ( .A(n_155), .B(n_21), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_175), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_163), .B(n_23), .Y(n_224) );
AOI22xp5_ASAP7_75t_SL g225 ( .A1(n_162), .A2(n_26), .B1(n_29), .B2(n_30), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_175), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_156), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_150), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_175), .Y(n_229) );
INVx4_ASAP7_75t_L g230 ( .A(n_175), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g231 ( .A1(n_163), .A2(n_35), .B1(n_36), .B2(n_38), .Y(n_231) );
CKINVDCx11_ASAP7_75t_R g232 ( .A(n_174), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_156), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_150), .B(n_42), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_153), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_153), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_156), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_158), .Y(n_238) );
BUFx3_ASAP7_75t_L g239 ( .A(n_142), .Y(n_239) );
INVx5_ASAP7_75t_L g240 ( .A(n_142), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_156), .Y(n_241) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_142), .Y(n_242) );
BUFx8_ASAP7_75t_SL g243 ( .A(n_174), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_156), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_177), .B(n_77), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_158), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_206), .B(n_150), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_209), .B(n_210), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_213), .B(n_178), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_230), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g251 ( .A1(n_202), .A2(n_172), .B1(n_178), .B2(n_177), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_230), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_193), .B(n_165), .Y(n_253) );
AOI221xp5_ASAP7_75t_SL g254 ( .A1(n_183), .A2(n_197), .B1(n_189), .B2(n_205), .C(n_200), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_192), .B(n_173), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_184), .B(n_164), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_188), .B(n_164), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_185), .B(n_165), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_199), .B(n_167), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_230), .B(n_167), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_217), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_212), .B(n_167), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_217), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_218), .A2(n_156), .B1(n_157), .B2(n_145), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_195), .B(n_141), .Y(n_265) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_188), .Y(n_266) );
BUFx6f_ASAP7_75t_L g267 ( .A(n_218), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_198), .B(n_169), .Y(n_268) );
AND2x4_ASAP7_75t_L g269 ( .A(n_215), .B(n_169), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_198), .B(n_168), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_208), .B(n_159), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_208), .B(n_159), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_215), .B(n_159), .Y(n_273) );
INVx4_ASAP7_75t_L g274 ( .A(n_228), .Y(n_274) );
BUFx6f_ASAP7_75t_L g275 ( .A(n_218), .Y(n_275) );
INVxp67_ASAP7_75t_L g276 ( .A(n_243), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_215), .B(n_159), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g278 ( .A1(n_218), .A2(n_157), .B1(n_134), .B2(n_145), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_218), .A2(n_157), .B1(n_152), .B2(n_134), .Y(n_279) );
BUFx2_ASAP7_75t_L g280 ( .A(n_243), .Y(n_280) );
AND2x2_ASAP7_75t_SL g281 ( .A(n_221), .B(n_139), .Y(n_281) );
INVx1_ASAP7_75t_SL g282 ( .A(n_232), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_228), .B(n_157), .Y(n_283) );
NOR2x2_ASAP7_75t_L g284 ( .A(n_232), .B(n_151), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_186), .B(n_167), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_217), .Y(n_286) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_220), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_186), .B(n_166), .Y(n_288) );
BUFx5_ASAP7_75t_L g289 ( .A(n_218), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_207), .Y(n_290) );
NAND2xp33_ASAP7_75t_L g291 ( .A(n_222), .B(n_157), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_203), .B(n_166), .Y(n_292) );
BUFx3_ASAP7_75t_L g293 ( .A(n_220), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_211), .B(n_168), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_221), .B(n_148), .Y(n_295) );
NOR2xp67_ASAP7_75t_L g296 ( .A(n_196), .B(n_152), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_207), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_221), .B(n_147), .Y(n_298) );
INVx3_ASAP7_75t_L g299 ( .A(n_235), .Y(n_299) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_187), .B(n_157), .Y(n_300) );
NAND2xp5_ASAP7_75t_SL g301 ( .A(n_187), .B(n_148), .Y(n_301) );
AND2x4_ASAP7_75t_L g302 ( .A(n_219), .B(n_147), .Y(n_302) );
OAI22xp5_ASAP7_75t_SL g303 ( .A1(n_202), .A2(n_151), .B1(n_172), .B2(n_139), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_239), .Y(n_304) );
INVx4_ASAP7_75t_L g305 ( .A(n_216), .Y(n_305) );
NOR3xp33_ASAP7_75t_L g306 ( .A(n_180), .B(n_146), .C(n_139), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_236), .B(n_146), .Y(n_307) );
AND2x6_ASAP7_75t_SL g308 ( .A(n_190), .B(n_139), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_238), .B(n_142), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_246), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_239), .Y(n_311) );
OAI22xp5_ASAP7_75t_L g312 ( .A1(n_223), .A2(n_44), .B1(n_46), .B2(n_47), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_226), .B(n_50), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g314 ( .A1(n_229), .A2(n_54), .B1(n_60), .B2(n_65), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_227), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_181), .B(n_66), .Y(n_316) );
INVx8_ASAP7_75t_L g317 ( .A(n_245), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_181), .B(n_67), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_187), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_299), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_248), .B(n_225), .Y(n_321) );
INVx3_ASAP7_75t_L g322 ( .A(n_299), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_280), .Y(n_323) );
NAND2xp5_ASAP7_75t_SL g324 ( .A(n_266), .B(n_274), .Y(n_324) );
AOI22xp33_ASAP7_75t_L g325 ( .A1(n_303), .A2(n_234), .B1(n_224), .B2(n_231), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_247), .A2(n_224), .B(n_241), .Y(n_326) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_257), .A2(n_244), .B(n_241), .Y(n_327) );
OAI22x1_ASAP7_75t_L g328 ( .A1(n_282), .A2(n_240), .B1(n_204), .B2(n_214), .Y(n_328) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_291), .A2(n_244), .B(n_237), .Y(n_329) );
AO22x1_ASAP7_75t_L g330 ( .A1(n_287), .A2(n_240), .B1(n_233), .B2(n_237), .Y(n_330) );
OAI21xp33_ASAP7_75t_SL g331 ( .A1(n_288), .A2(n_233), .B(n_227), .Y(n_331) );
BUFx2_ASAP7_75t_L g332 ( .A(n_276), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_285), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_278), .A2(n_240), .B1(n_194), .B2(n_214), .Y(n_334) );
NOR2xp33_ASAP7_75t_R g335 ( .A(n_293), .B(n_69), .Y(n_335) );
NAND2xp5_ASAP7_75t_SL g336 ( .A(n_266), .B(n_240), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_250), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_261), .Y(n_338) );
O2A1O1Ixp33_ASAP7_75t_L g339 ( .A1(n_251), .A2(n_194), .B(n_182), .C(n_204), .Y(n_339) );
BUFx12f_ASAP7_75t_L g340 ( .A(n_305), .Y(n_340) );
AOI21xp5_ASAP7_75t_L g341 ( .A1(n_256), .A2(n_182), .B(n_191), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_265), .B(n_319), .Y(n_342) );
AOI21xp5_ASAP7_75t_L g343 ( .A1(n_258), .A2(n_191), .B(n_242), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_252), .A2(n_191), .B(n_242), .Y(n_344) );
NAND2xp5_ASAP7_75t_SL g345 ( .A(n_266), .B(n_240), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_260), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_263), .Y(n_347) );
NAND2xp5_ASAP7_75t_SL g348 ( .A(n_266), .B(n_201), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_292), .B(n_201), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_273), .Y(n_350) );
O2A1O1Ixp33_ASAP7_75t_L g351 ( .A1(n_294), .A2(n_201), .B(n_242), .C(n_191), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_278), .A2(n_242), .B1(n_72), .B2(n_75), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_286), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_262), .Y(n_354) );
AOI21xp5_ASAP7_75t_L g355 ( .A1(n_281), .A2(n_300), .B(n_253), .Y(n_355) );
AOI21xp5_ASAP7_75t_L g356 ( .A1(n_281), .A2(n_249), .B(n_295), .Y(n_356) );
BUFx6f_ASAP7_75t_L g357 ( .A(n_267), .Y(n_357) );
OAI22xp5_ASAP7_75t_L g358 ( .A1(n_279), .A2(n_264), .B1(n_317), .B2(n_267), .Y(n_358) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_276), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_277), .Y(n_360) );
AND2x4_ASAP7_75t_L g361 ( .A(n_274), .B(n_269), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_269), .Y(n_362) );
INVx3_ASAP7_75t_L g363 ( .A(n_267), .Y(n_363) );
AOI22xp5_ASAP7_75t_L g364 ( .A1(n_255), .A2(n_317), .B1(n_302), .B2(n_254), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_310), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_317), .B(n_268), .Y(n_366) );
INVx4_ASAP7_75t_L g367 ( .A(n_267), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_279), .A2(n_264), .B1(n_275), .B2(n_259), .Y(n_368) );
INVx4_ASAP7_75t_L g369 ( .A(n_275), .Y(n_369) );
AOI22xp5_ASAP7_75t_L g370 ( .A1(n_255), .A2(n_302), .B1(n_305), .B2(n_268), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_287), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_308), .Y(n_372) );
O2A1O1Ixp33_ASAP7_75t_SL g373 ( .A1(n_316), .A2(n_318), .B(n_313), .C(n_283), .Y(n_373) );
AOI21xp5_ASAP7_75t_L g374 ( .A1(n_298), .A2(n_301), .B(n_271), .Y(n_374) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_272), .A2(n_270), .B(n_306), .Y(n_375) );
AO21x1_ASAP7_75t_L g376 ( .A1(n_306), .A2(n_312), .B(n_309), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_275), .A2(n_270), .B1(n_307), .B2(n_296), .Y(n_377) );
O2A1O1Ixp5_ASAP7_75t_L g378 ( .A1(n_376), .A2(n_297), .B(n_311), .C(n_304), .Y(n_378) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_354), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_365), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_321), .B(n_275), .Y(n_381) );
AOI22x1_ASAP7_75t_L g382 ( .A1(n_375), .A2(n_290), .B1(n_289), .B2(n_315), .Y(n_382) );
OAI21xp5_ASAP7_75t_L g383 ( .A1(n_356), .A2(n_314), .B(n_289), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_321), .A2(n_289), .B1(n_284), .B2(n_314), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_364), .A2(n_289), .B1(n_370), .B2(n_366), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_333), .A2(n_289), .B1(n_342), .B2(n_362), .Y(n_386) );
A2O1A1Ixp33_ASAP7_75t_L g387 ( .A1(n_339), .A2(n_289), .B(n_375), .C(n_355), .Y(n_387) );
NAND3xp33_ASAP7_75t_L g388 ( .A(n_325), .B(n_331), .C(n_372), .Y(n_388) );
BUFx3_ASAP7_75t_L g389 ( .A(n_340), .Y(n_389) );
NOR2xp67_ASAP7_75t_SL g390 ( .A(n_357), .B(n_369), .Y(n_390) );
AOI21xp5_ASAP7_75t_L g391 ( .A1(n_373), .A2(n_326), .B(n_343), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_350), .B(n_360), .Y(n_392) );
AOI22xp33_ASAP7_75t_SL g393 ( .A1(n_335), .A2(n_361), .B1(n_332), .B2(n_371), .Y(n_393) );
NOR3xp33_ASAP7_75t_SL g394 ( .A(n_323), .B(n_366), .C(n_324), .Y(n_394) );
OAI21x1_ASAP7_75t_L g395 ( .A1(n_351), .A2(n_344), .B(n_377), .Y(n_395) );
BUFx3_ASAP7_75t_L g396 ( .A(n_361), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_346), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_338), .Y(n_398) );
O2A1O1Ixp5_ASAP7_75t_L g399 ( .A1(n_330), .A2(n_377), .B(n_336), .C(n_345), .Y(n_399) );
BUFx3_ASAP7_75t_L g400 ( .A(n_357), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_357), .Y(n_401) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_359), .Y(n_402) );
A2O1A1Ixp33_ASAP7_75t_L g403 ( .A1(n_374), .A2(n_353), .B(n_347), .C(n_320), .Y(n_403) );
AOI21xp5_ASAP7_75t_L g404 ( .A1(n_341), .A2(n_368), .B(n_327), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_320), .B(n_322), .Y(n_405) );
AND2x4_ASAP7_75t_L g406 ( .A(n_322), .B(n_369), .Y(n_406) );
AND2x4_ASAP7_75t_L g407 ( .A(n_367), .B(n_349), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_337), .B(n_358), .Y(n_408) );
AOI21xp5_ASAP7_75t_L g409 ( .A1(n_368), .A2(n_329), .B(n_358), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_363), .Y(n_410) );
AOI221xp5_ASAP7_75t_SL g411 ( .A1(n_328), .A2(n_334), .B1(n_352), .B2(n_348), .C(n_363), .Y(n_411) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_367), .A2(n_202), .B1(n_232), .B2(n_321), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_352), .Y(n_413) );
NOR2xp67_ASAP7_75t_L g414 ( .A(n_379), .B(n_334), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_397), .B(n_392), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_402), .Y(n_416) );
AND2x4_ASAP7_75t_L g417 ( .A(n_397), .B(n_380), .Y(n_417) );
OAI21xp5_ASAP7_75t_L g418 ( .A1(n_387), .A2(n_378), .B(n_381), .Y(n_418) );
AOI21xp5_ASAP7_75t_L g419 ( .A1(n_391), .A2(n_404), .B(n_383), .Y(n_419) );
AOI21xp5_ASAP7_75t_L g420 ( .A1(n_409), .A2(n_413), .B(n_403), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_398), .B(n_380), .Y(n_421) );
OR2x6_ASAP7_75t_L g422 ( .A(n_396), .B(n_407), .Y(n_422) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_400), .Y(n_423) );
AOI21xp5_ASAP7_75t_L g424 ( .A1(n_413), .A2(n_382), .B(n_385), .Y(n_424) );
CKINVDCx11_ASAP7_75t_R g425 ( .A(n_389), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_398), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_384), .B(n_396), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_412), .B(n_393), .Y(n_428) );
XNOR2xp5_ASAP7_75t_L g429 ( .A(n_388), .B(n_394), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_401), .Y(n_430) );
OA21x2_ASAP7_75t_L g431 ( .A1(n_395), .A2(n_411), .B(n_382), .Y(n_431) );
AO21x2_ASAP7_75t_L g432 ( .A1(n_408), .A2(n_395), .B(n_410), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_405), .B(n_407), .Y(n_433) );
OA21x2_ASAP7_75t_L g434 ( .A1(n_399), .A2(n_410), .B(n_401), .Y(n_434) );
A2O1A1Ixp33_ASAP7_75t_L g435 ( .A1(n_386), .A2(n_405), .B(n_406), .C(n_407), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_406), .Y(n_436) );
O2A1O1Ixp5_ASAP7_75t_L g437 ( .A1(n_390), .A2(n_406), .B(n_400), .C(n_389), .Y(n_437) );
BUFx2_ASAP7_75t_L g438 ( .A(n_390), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_380), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_380), .Y(n_440) );
A2O1A1Ixp33_ASAP7_75t_L g441 ( .A1(n_381), .A2(n_375), .B(n_321), .C(n_409), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_384), .A2(n_232), .B1(n_303), .B2(n_220), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_384), .A2(n_232), .B1(n_282), .B2(n_202), .Y(n_443) );
OR2x6_ASAP7_75t_L g444 ( .A(n_435), .B(n_424), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_439), .Y(n_445) );
BUFx2_ASAP7_75t_L g446 ( .A(n_434), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_432), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_417), .B(n_421), .Y(n_448) );
INVx3_ASAP7_75t_L g449 ( .A(n_423), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_421), .B(n_415), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_442), .A2(n_427), .B1(n_428), .B2(n_417), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_425), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_417), .B(n_427), .Y(n_453) );
INVx3_ASAP7_75t_SL g454 ( .A(n_422), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_440), .B(n_441), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_419), .A2(n_420), .B(n_441), .Y(n_456) );
BUFx2_ASAP7_75t_L g457 ( .A(n_434), .Y(n_457) );
AO21x2_ASAP7_75t_L g458 ( .A1(n_418), .A2(n_435), .B(n_432), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_426), .B(n_430), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_432), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_430), .Y(n_461) );
AND2x4_ASAP7_75t_L g462 ( .A(n_423), .B(n_436), .Y(n_462) );
AND2x4_ASAP7_75t_L g463 ( .A(n_423), .B(n_422), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_433), .B(n_414), .Y(n_464) );
NAND4xp25_ASAP7_75t_SL g465 ( .A(n_443), .B(n_425), .C(n_429), .D(n_422), .Y(n_465) );
OA21x2_ASAP7_75t_L g466 ( .A1(n_437), .A2(n_431), .B(n_438), .Y(n_466) );
INVx2_ASAP7_75t_SL g467 ( .A(n_423), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_434), .B(n_422), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_431), .B(n_429), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_431), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_416), .B(n_417), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_421), .B(n_415), .Y(n_472) );
OA21x2_ASAP7_75t_L g473 ( .A1(n_419), .A2(n_424), .B(n_420), .Y(n_473) );
AO21x2_ASAP7_75t_L g474 ( .A1(n_424), .A2(n_419), .B(n_420), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_432), .Y(n_475) );
INVx2_ASAP7_75t_SL g476 ( .A(n_423), .Y(n_476) );
INVx3_ASAP7_75t_L g477 ( .A(n_423), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_417), .B(n_421), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_417), .B(n_421), .Y(n_479) );
OA21x2_ASAP7_75t_L g480 ( .A1(n_419), .A2(n_424), .B(n_420), .Y(n_480) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_461), .Y(n_481) );
INVx3_ASAP7_75t_L g482 ( .A(n_466), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_453), .B(n_469), .Y(n_483) );
BUFx2_ASAP7_75t_L g484 ( .A(n_468), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_453), .B(n_469), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_453), .B(n_469), .Y(n_486) );
INVx1_ASAP7_75t_SL g487 ( .A(n_471), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_455), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_447), .Y(n_489) );
BUFx2_ASAP7_75t_L g490 ( .A(n_468), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_444), .B(n_458), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_445), .B(n_472), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_455), .Y(n_493) );
INVx2_ASAP7_75t_SL g494 ( .A(n_463), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_448), .B(n_479), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_448), .B(n_479), .Y(n_496) );
AO21x2_ASAP7_75t_L g497 ( .A1(n_456), .A2(n_474), .B(n_460), .Y(n_497) );
NAND2x1_ASAP7_75t_L g498 ( .A(n_461), .B(n_468), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_450), .B(n_472), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_445), .Y(n_500) );
AND2x4_ASAP7_75t_L g501 ( .A(n_463), .B(n_444), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_459), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_444), .B(n_458), .Y(n_503) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_471), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_459), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_448), .B(n_479), .Y(n_506) );
INVx4_ASAP7_75t_L g507 ( .A(n_454), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_444), .B(n_458), .Y(n_508) );
INVx4_ASAP7_75t_L g509 ( .A(n_454), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_459), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_444), .B(n_458), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_444), .B(n_458), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_444), .B(n_478), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_478), .B(n_475), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_446), .Y(n_515) );
AO21x2_ASAP7_75t_L g516 ( .A1(n_456), .A2(n_474), .B(n_470), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_470), .Y(n_517) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_471), .Y(n_518) );
AND2x4_ASAP7_75t_L g519 ( .A(n_463), .B(n_449), .Y(n_519) );
NAND2x1_ASAP7_75t_L g520 ( .A(n_449), .B(n_477), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_446), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_450), .B(n_472), .Y(n_522) );
INVx5_ASAP7_75t_L g523 ( .A(n_449), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_470), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_446), .Y(n_525) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_474), .A2(n_464), .B(n_478), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_499), .B(n_450), .Y(n_527) );
INVx6_ASAP7_75t_L g528 ( .A(n_507), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_500), .Y(n_529) );
OR2x6_ASAP7_75t_L g530 ( .A(n_498), .B(n_457), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_483), .B(n_457), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_500), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_483), .B(n_457), .Y(n_533) );
INVxp67_ASAP7_75t_SL g534 ( .A(n_481), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_499), .Y(n_535) );
AOI21xp33_ASAP7_75t_L g536 ( .A1(n_526), .A2(n_451), .B(n_464), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_522), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_483), .B(n_474), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_522), .B(n_454), .Y(n_539) );
AND2x4_ASAP7_75t_SL g540 ( .A(n_507), .B(n_463), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_492), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_485), .B(n_474), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_492), .Y(n_543) );
OR2x2_ASAP7_75t_L g544 ( .A(n_504), .B(n_454), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_485), .B(n_480), .Y(n_545) );
NOR2x1_ASAP7_75t_L g546 ( .A(n_507), .B(n_452), .Y(n_546) );
NAND2x1p5_ASAP7_75t_L g547 ( .A(n_507), .B(n_463), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_481), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_509), .B(n_476), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_504), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_495), .B(n_451), .Y(n_551) );
INVxp67_ASAP7_75t_SL g552 ( .A(n_489), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_518), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_485), .B(n_480), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_486), .B(n_514), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_517), .Y(n_556) );
AOI31xp33_ASAP7_75t_L g557 ( .A1(n_518), .A2(n_452), .A3(n_465), .B(n_467), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_517), .Y(n_558) );
NAND2x1_ASAP7_75t_L g559 ( .A(n_509), .B(n_449), .Y(n_559) );
OAI21xp33_ASAP7_75t_SL g560 ( .A1(n_509), .A2(n_465), .B(n_467), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_526), .A2(n_462), .B1(n_473), .B2(n_480), .Y(n_561) );
NOR2x1_ASAP7_75t_L g562 ( .A(n_509), .B(n_449), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_486), .B(n_473), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_517), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_486), .B(n_473), .Y(n_565) );
NAND2x1p5_ASAP7_75t_L g566 ( .A(n_523), .B(n_477), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_495), .B(n_462), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_514), .B(n_473), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_487), .B(n_467), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_502), .Y(n_570) );
INVx2_ASAP7_75t_SL g571 ( .A(n_523), .Y(n_571) );
AND2x4_ASAP7_75t_L g572 ( .A(n_501), .B(n_477), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_502), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_524), .Y(n_574) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_487), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_496), .B(n_462), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_514), .B(n_473), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_496), .B(n_476), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_524), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_513), .B(n_473), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_513), .B(n_480), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_513), .B(n_480), .Y(n_582) );
NOR3xp33_ASAP7_75t_SL g583 ( .A(n_488), .B(n_462), .C(n_476), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_526), .B(n_480), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_526), .B(n_466), .Y(n_585) );
AND2x4_ASAP7_75t_L g586 ( .A(n_501), .B(n_477), .Y(n_586) );
OAI32xp33_ASAP7_75t_L g587 ( .A1(n_560), .A2(n_510), .A3(n_505), .B1(n_511), .B2(n_503), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_556), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_541), .B(n_506), .Y(n_589) );
NOR2x1_ASAP7_75t_L g590 ( .A(n_546), .B(n_498), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_529), .Y(n_591) );
NOR2xp33_ASAP7_75t_SL g592 ( .A(n_528), .B(n_523), .Y(n_592) );
INVx1_ASAP7_75t_SL g593 ( .A(n_578), .Y(n_593) );
INVx3_ASAP7_75t_SL g594 ( .A(n_528), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_555), .B(n_484), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_535), .B(n_537), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_556), .Y(n_597) );
NAND2x1p5_ASAP7_75t_L g598 ( .A(n_559), .B(n_523), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_538), .B(n_491), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_543), .B(n_506), .Y(n_600) );
INVxp67_ASAP7_75t_L g601 ( .A(n_575), .Y(n_601) );
INVx2_ASAP7_75t_SL g602 ( .A(n_528), .Y(n_602) );
INVx2_ASAP7_75t_L g603 ( .A(n_558), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_538), .B(n_491), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_550), .B(n_505), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_558), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_532), .Y(n_607) );
INVx1_ASAP7_75t_SL g608 ( .A(n_569), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_555), .B(n_542), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_564), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_542), .B(n_511), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_548), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_545), .B(n_511), .Y(n_613) );
INVx1_ASAP7_75t_SL g614 ( .A(n_540), .Y(n_614) );
NOR2xp67_ASAP7_75t_L g615 ( .A(n_571), .B(n_482), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_531), .B(n_484), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_564), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_574), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_553), .Y(n_619) );
AOI32xp33_ASAP7_75t_L g620 ( .A1(n_545), .A2(n_490), .A3(n_503), .B1(n_508), .B2(n_491), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_531), .B(n_490), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_570), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_573), .Y(n_623) );
OR2x2_ASAP7_75t_L g624 ( .A(n_533), .B(n_510), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_574), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_554), .B(n_512), .Y(n_626) );
INVx1_ASAP7_75t_SL g627 ( .A(n_540), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_534), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_554), .B(n_563), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_527), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_563), .B(n_512), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_567), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_533), .B(n_494), .Y(n_633) );
OR2x2_ASAP7_75t_L g634 ( .A(n_576), .B(n_494), .Y(n_634) );
OR2x2_ASAP7_75t_L g635 ( .A(n_565), .B(n_525), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_551), .B(n_493), .Y(n_636) );
AOI21xp33_ASAP7_75t_SL g637 ( .A1(n_557), .A2(n_494), .B(n_501), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_565), .B(n_512), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_580), .B(n_508), .Y(n_639) );
INVx1_ASAP7_75t_SL g640 ( .A(n_539), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_568), .B(n_488), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_580), .B(n_508), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_632), .B(n_568), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_612), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_622), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_630), .B(n_577), .Y(n_646) );
INVx2_ASAP7_75t_SL g647 ( .A(n_594), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_629), .B(n_582), .Y(n_648) );
INVx1_ASAP7_75t_SL g649 ( .A(n_594), .Y(n_649) );
NAND3xp33_ASAP7_75t_L g650 ( .A(n_620), .B(n_536), .C(n_561), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_623), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_596), .A2(n_501), .B1(n_581), .B2(n_582), .Y(n_652) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_637), .B(n_583), .Y(n_653) );
AOI21xp33_ASAP7_75t_SL g654 ( .A1(n_587), .A2(n_547), .B(n_549), .Y(n_654) );
OAI22xp33_ASAP7_75t_L g655 ( .A1(n_592), .A2(n_530), .B1(n_544), .B2(n_547), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_629), .B(n_581), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_591), .Y(n_657) );
NOR2xp33_ASAP7_75t_SL g658 ( .A(n_614), .B(n_571), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_613), .B(n_577), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_636), .B(n_493), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_588), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_607), .Y(n_662) );
OR2x2_ASAP7_75t_L g663 ( .A(n_609), .B(n_552), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_613), .B(n_503), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_609), .B(n_586), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_619), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_628), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_635), .Y(n_668) );
O2A1O1Ixp33_ASAP7_75t_SL g669 ( .A1(n_627), .A2(n_549), .B(n_520), .C(n_584), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_635), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_599), .B(n_525), .Y(n_671) );
OA21x2_ASAP7_75t_L g672 ( .A1(n_615), .A2(n_561), .B(n_585), .Y(n_672) );
OR2x2_ASAP7_75t_L g673 ( .A(n_595), .B(n_521), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_626), .B(n_585), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_624), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_599), .B(n_515), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_604), .B(n_515), .Y(n_677) );
OR2x2_ASAP7_75t_L g678 ( .A(n_621), .B(n_521), .Y(n_678) );
INVx1_ASAP7_75t_SL g679 ( .A(n_593), .Y(n_679) );
OR2x2_ASAP7_75t_L g680 ( .A(n_621), .B(n_579), .Y(n_680) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_601), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_626), .B(n_530), .Y(n_682) );
INVx1_ASAP7_75t_SL g683 ( .A(n_649), .Y(n_683) );
AOI211xp5_ASAP7_75t_L g684 ( .A1(n_653), .A2(n_602), .B(n_640), .C(n_596), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_668), .B(n_611), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_681), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_679), .B(n_608), .Y(n_687) );
INVxp67_ASAP7_75t_L g688 ( .A(n_681), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_670), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_645), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_674), .B(n_604), .Y(n_691) );
INVxp33_ASAP7_75t_L g692 ( .A(n_658), .Y(n_692) );
OAI211xp5_ASAP7_75t_L g693 ( .A1(n_653), .A2(n_590), .B(n_602), .C(n_641), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_651), .Y(n_694) );
AO22x2_ASAP7_75t_L g695 ( .A1(n_650), .A2(n_616), .B1(n_605), .B2(n_634), .Y(n_695) );
OAI222xp33_ASAP7_75t_L g696 ( .A1(n_647), .A2(n_530), .B1(n_611), .B2(n_639), .C1(n_642), .C2(n_638), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_657), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_674), .B(n_638), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_662), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_644), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_652), .A2(n_530), .B1(n_598), .B2(n_633), .Y(n_701) );
AND2x4_ASAP7_75t_L g702 ( .A(n_647), .B(n_631), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_666), .Y(n_703) );
INVx2_ASAP7_75t_L g704 ( .A(n_663), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_661), .Y(n_705) );
AOI22xp5_ASAP7_75t_SL g706 ( .A1(n_682), .A2(n_598), .B1(n_600), .B2(n_589), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_675), .B(n_631), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_683), .A2(n_682), .B1(n_655), .B2(n_672), .Y(n_708) );
AOI322xp5_ASAP7_75t_L g709 ( .A1(n_683), .A2(n_648), .A3(n_656), .B1(n_659), .B2(n_664), .C1(n_655), .C2(n_642), .Y(n_709) );
A2O1A1Ixp33_ASAP7_75t_L g710 ( .A1(n_684), .A2(n_654), .B(n_656), .C(n_648), .Y(n_710) );
AOI211x1_ASAP7_75t_L g711 ( .A1(n_696), .A2(n_659), .B(n_665), .C(n_664), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_686), .Y(n_712) );
OAI322xp33_ASAP7_75t_L g713 ( .A1(n_688), .A2(n_673), .A3(n_678), .B1(n_646), .B2(n_667), .C1(n_643), .C2(n_660), .Y(n_713) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_702), .Y(n_714) );
O2A1O1Ixp33_ASAP7_75t_L g715 ( .A1(n_693), .A2(n_669), .B(n_584), .C(n_672), .Y(n_715) );
AOI21xp33_ASAP7_75t_L g716 ( .A1(n_695), .A2(n_672), .B(n_497), .Y(n_716) );
AOI222xp33_ASAP7_75t_L g717 ( .A1(n_695), .A2(n_639), .B1(n_677), .B2(n_676), .C1(n_671), .C2(n_661), .Y(n_717) );
OAI22xp33_ASAP7_75t_L g718 ( .A1(n_692), .A2(n_680), .B1(n_669), .B2(n_562), .Y(n_718) );
NOR3xp33_ASAP7_75t_L g719 ( .A(n_701), .B(n_477), .C(n_482), .Y(n_719) );
OAI222xp33_ASAP7_75t_L g720 ( .A1(n_706), .A2(n_572), .B1(n_586), .B2(n_566), .C1(n_519), .C2(n_610), .Y(n_720) );
NOR2x1_ASAP7_75t_L g721 ( .A(n_701), .B(n_520), .Y(n_721) );
AOI221xp5_ASAP7_75t_L g722 ( .A1(n_689), .A2(n_707), .B1(n_694), .B2(n_690), .C(n_703), .Y(n_722) );
A2O1A1Ixp33_ASAP7_75t_L g723 ( .A1(n_710), .A2(n_687), .B(n_702), .C(n_685), .Y(n_723) );
NAND2xp5_ASAP7_75t_SL g724 ( .A(n_718), .B(n_704), .Y(n_724) );
AOI22xp5_ASAP7_75t_L g725 ( .A1(n_708), .A2(n_697), .B1(n_700), .B2(n_699), .Y(n_725) );
NAND3xp33_ASAP7_75t_SL g726 ( .A(n_715), .B(n_698), .C(n_691), .Y(n_726) );
OAI222xp33_ASAP7_75t_L g727 ( .A1(n_721), .A2(n_685), .B1(n_705), .B2(n_586), .C1(n_572), .C2(n_566), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_722), .B(n_625), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_717), .B(n_625), .Y(n_729) );
AOI321xp33_ASAP7_75t_L g730 ( .A1(n_719), .A2(n_572), .A3(n_519), .B1(n_618), .B2(n_597), .C(n_617), .Y(n_730) );
AOI211xp5_ASAP7_75t_L g731 ( .A1(n_720), .A2(n_519), .B(n_617), .C(n_610), .Y(n_731) );
AOI221xp5_ASAP7_75t_SL g732 ( .A1(n_723), .A2(n_713), .B1(n_716), .B2(n_711), .C(n_712), .Y(n_732) );
OAI211xp5_ASAP7_75t_SL g733 ( .A1(n_731), .A2(n_709), .B(n_714), .C(n_482), .Y(n_733) );
NAND3xp33_ASAP7_75t_SL g734 ( .A(n_725), .B(n_618), .C(n_606), .Y(n_734) );
NOR4xp25_ASAP7_75t_L g735 ( .A(n_726), .B(n_482), .C(n_603), .D(n_606), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_724), .A2(n_519), .B1(n_597), .B2(n_588), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_736), .Y(n_737) );
NOR2x1_ASAP7_75t_L g738 ( .A(n_734), .B(n_727), .Y(n_738) );
NOR2x1_ASAP7_75t_L g739 ( .A(n_733), .B(n_728), .Y(n_739) );
INVx2_ASAP7_75t_L g740 ( .A(n_737), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_738), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_740), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_740), .Y(n_743) );
BUFx4f_ASAP7_75t_SL g744 ( .A(n_742), .Y(n_744) );
OAI22x1_ASAP7_75t_SL g745 ( .A1(n_744), .A2(n_743), .B1(n_741), .B2(n_732), .Y(n_745) );
NAND3xp33_ASAP7_75t_L g746 ( .A(n_745), .B(n_739), .C(n_735), .Y(n_746) );
AO21x2_ASAP7_75t_L g747 ( .A1(n_746), .A2(n_729), .B(n_730), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_747), .A2(n_497), .B1(n_603), .B2(n_516), .Y(n_748) );
endmodule