module fake_ariane_542_n_760 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_760);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_760;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_679;
wire n_643;
wire n_226;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_151;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_733;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_455;
wire n_365;
wire n_429;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;
wire n_675;

INVx2_ASAP7_75t_SL g150 ( 
.A(n_20),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_31),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_70),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_86),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_26),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_145),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_63),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_6),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_51),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_47),
.B(n_54),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_88),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_44),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_106),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_123),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_75),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_33),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_11),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_108),
.Y(n_171)
);

INVxp67_ASAP7_75t_SL g172 ( 
.A(n_133),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_65),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_10),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_28),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_125),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_115),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_97),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_24),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_111),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_112),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_55),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_36),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_67),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_128),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_80),
.Y(n_189)
);

NOR2xp67_ASAP7_75t_L g190 ( 
.A(n_143),
.B(n_56),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_62),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_147),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_76),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_109),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_29),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_49),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_69),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_119),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_52),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_15),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_95),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_107),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_0),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_174),
.Y(n_205)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_196),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_199),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_199),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_153),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_161),
.Y(n_210)
);

BUFx12f_ASAP7_75t_L g211 ( 
.A(n_150),
.Y(n_211)
);

AND2x6_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_16),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_168),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_170),
.Y(n_214)
);

BUFx12f_ASAP7_75t_L g215 ( 
.A(n_152),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_151),
.Y(n_216)
);

AND2x4_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_1),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_154),
.Y(n_218)
);

NOR2x1_ASAP7_75t_L g219 ( 
.A(n_156),
.B(n_17),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_162),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_164),
.B(n_2),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_175),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_178),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_153),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_179),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_155),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_181),
.B(n_3),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_182),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_183),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_184),
.B(n_3),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_196),
.Y(n_231)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_196),
.Y(n_232)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_196),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_194),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_200),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_155),
.Y(n_236)
);

AND2x6_ASAP7_75t_L g237 ( 
.A(n_165),
.B(n_18),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_165),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_198),
.Y(n_239)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_157),
.Y(n_240)
);

BUFx12f_ASAP7_75t_L g241 ( 
.A(n_158),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_198),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_231),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_231),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_231),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_209),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_236),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_217),
.B(n_204),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_214),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_236),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_236),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_241),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_236),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_215),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_214),
.B(n_195),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_207),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_215),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_224),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_239),
.Y(n_259)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_207),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_R g261 ( 
.A(n_203),
.B(n_173),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_224),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_205),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_240),
.Y(n_264)
);

NOR2xp67_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_163),
.Y(n_265)
);

NOR2xp67_ASAP7_75t_L g266 ( 
.A(n_211),
.B(n_159),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_239),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_211),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_R g269 ( 
.A(n_203),
.B(n_166),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_205),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_216),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_216),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_223),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_223),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_234),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_234),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_208),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_231),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_210),
.B(n_186),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_208),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_239),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_220),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_226),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_R g284 ( 
.A(n_225),
.B(n_167),
.Y(n_284)
);

AND3x2_ASAP7_75t_L g285 ( 
.A(n_217),
.B(n_172),
.C(n_186),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_239),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_213),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_242),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_242),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_218),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_286),
.Y(n_291)
);

NAND2xp33_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_212),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_256),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_273),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_218),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_256),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_275),
.B(n_222),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_248),
.B(n_222),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_265),
.B(n_282),
.Y(n_299)
);

A2O1A1Ixp33_ASAP7_75t_L g300 ( 
.A1(n_248),
.A2(n_221),
.B(n_230),
.C(n_227),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_260),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_260),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_255),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_277),
.B(n_228),
.Y(n_304)
);

NAND3xp33_ASAP7_75t_L g305 ( 
.A(n_283),
.B(n_221),
.C(n_235),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_280),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_228),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_286),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_280),
.B(n_229),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_261),
.B(n_229),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_261),
.B(n_235),
.Y(n_311)
);

INVx2_ASAP7_75t_SL g312 ( 
.A(n_271),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_269),
.B(n_238),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_249),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_247),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_276),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_250),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_251),
.Y(n_318)
);

NAND3xp33_ASAP7_75t_L g319 ( 
.A(n_279),
.B(n_242),
.C(n_219),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_284),
.B(n_238),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_253),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_259),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_268),
.B(n_242),
.Y(n_323)
);

NOR3xp33_ASAP7_75t_L g324 ( 
.A(n_258),
.B(n_262),
.C(n_246),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_267),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_281),
.A2(n_212),
.B1(n_237),
.B2(n_197),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_289),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_243),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_252),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_284),
.B(n_212),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_243),
.Y(n_331)
);

OR2x6_ASAP7_75t_L g332 ( 
.A(n_266),
.B(n_190),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_244),
.B(n_212),
.Y(n_333)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_244),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_245),
.B(n_212),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_245),
.B(n_206),
.Y(n_336)
);

OR2x6_ASAP7_75t_L g337 ( 
.A(n_285),
.B(n_232),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_278),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_278),
.B(n_206),
.Y(n_339)
);

NAND2x1_ASAP7_75t_L g340 ( 
.A(n_254),
.B(n_237),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g341 ( 
.A(n_257),
.Y(n_341)
);

NOR2xp67_ASAP7_75t_L g342 ( 
.A(n_263),
.B(n_206),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_270),
.B(n_169),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_287),
.B(n_206),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_249),
.B(n_232),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_256),
.Y(n_346)
);

AND2x4_ASAP7_75t_L g347 ( 
.A(n_272),
.B(n_237),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_272),
.B(n_233),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_256),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_286),
.Y(n_350)
);

NOR2xp67_ASAP7_75t_L g351 ( 
.A(n_252),
.B(n_233),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_272),
.B(n_171),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_286),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_309),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_314),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_293),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_301),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_299),
.B(n_303),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_346),
.Y(n_359)
);

INVx5_ASAP7_75t_L g360 ( 
.A(n_347),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_349),
.Y(n_361)
);

NAND2xp33_ASAP7_75t_L g362 ( 
.A(n_330),
.B(n_237),
.Y(n_362)
);

NAND3xp33_ASAP7_75t_SL g363 ( 
.A(n_324),
.B(n_202),
.C(n_177),
.Y(n_363)
);

INVx4_ASAP7_75t_L g364 ( 
.A(n_347),
.Y(n_364)
);

AND2x4_ASAP7_75t_L g365 ( 
.A(n_342),
.B(n_237),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_298),
.B(n_176),
.Y(n_366)
);

INVx2_ASAP7_75t_SL g367 ( 
.A(n_345),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_300),
.B(n_180),
.Y(n_368)
);

NOR3xp33_ASAP7_75t_SL g369 ( 
.A(n_343),
.B(n_187),
.C(n_188),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_294),
.B(n_189),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_312),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_316),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_296),
.Y(n_373)
);

BUFx4f_ASAP7_75t_L g374 ( 
.A(n_341),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_302),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_290),
.B(n_191),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_329),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_310),
.B(n_311),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_306),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_313),
.B(n_192),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_318),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_337),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_304),
.B(n_193),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_R g384 ( 
.A(n_292),
.B(n_201),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_325),
.Y(n_385)
);

NOR3xp33_ASAP7_75t_SL g386 ( 
.A(n_305),
.B(n_4),
.C(n_5),
.Y(n_386)
);

AND2x6_ASAP7_75t_SL g387 ( 
.A(n_332),
.B(n_337),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_350),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_332),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_350),
.Y(n_390)
);

INVx5_ASAP7_75t_L g391 ( 
.A(n_291),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_353),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_L g393 ( 
.A1(n_319),
.A2(n_232),
.B1(n_233),
.B2(n_9),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_315),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_315),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_351),
.B(n_7),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_344),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_295),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_297),
.B(n_233),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_321),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_320),
.B(n_7),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_327),
.Y(n_402)
);

OR2x6_ASAP7_75t_L g403 ( 
.A(n_323),
.B(n_8),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_307),
.B(n_8),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_348),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_353),
.B(n_9),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_334),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_352),
.B(n_10),
.Y(n_408)
);

NAND2xp33_ASAP7_75t_L g409 ( 
.A(n_326),
.B(n_11),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_334),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_328),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_331),
.B(n_12),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_338),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_317),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_340),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_317),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_317),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_322),
.B(n_13),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_291),
.B(n_14),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_322),
.Y(n_420)
);

AOI21xp33_ASAP7_75t_L g421 ( 
.A1(n_409),
.A2(n_335),
.B(n_333),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_362),
.A2(n_339),
.B(n_336),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_398),
.B(n_322),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_397),
.B(n_291),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_355),
.B(n_308),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_388),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_358),
.B(n_308),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_390),
.Y(n_428)
);

O2A1O1Ixp33_ASAP7_75t_L g429 ( 
.A1(n_376),
.A2(n_308),
.B(n_21),
.C(n_22),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_354),
.B(n_19),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_394),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_377),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_399),
.A2(n_23),
.B(n_25),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_383),
.B(n_27),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_383),
.B(n_30),
.Y(n_435)
);

INVx4_ASAP7_75t_L g436 ( 
.A(n_360),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_360),
.B(n_32),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_372),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_395),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_400),
.Y(n_440)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_360),
.Y(n_441)
);

O2A1O1Ixp33_ASAP7_75t_L g442 ( 
.A1(n_368),
.A2(n_34),
.B(n_35),
.C(n_37),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_382),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_420),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_364),
.B(n_374),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_366),
.B(n_38),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_399),
.A2(n_39),
.B(n_40),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_367),
.B(n_41),
.Y(n_448)
);

A2O1A1Ixp33_ASAP7_75t_L g449 ( 
.A1(n_408),
.A2(n_42),
.B(n_43),
.C(n_45),
.Y(n_449)
);

A2O1A1Ixp33_ASAP7_75t_L g450 ( 
.A1(n_408),
.A2(n_46),
.B(n_48),
.C(n_50),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_366),
.B(n_53),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_371),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_404),
.B(n_57),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_402),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_380),
.B(n_58),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_391),
.Y(n_456)
);

A2O1A1Ixp33_ASAP7_75t_L g457 ( 
.A1(n_368),
.A2(n_59),
.B(n_60),
.C(n_61),
.Y(n_457)
);

NOR2x1_ASAP7_75t_L g458 ( 
.A(n_363),
.B(n_364),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_380),
.B(n_64),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_378),
.A2(n_66),
.B(n_68),
.Y(n_460)
);

A2O1A1Ixp33_ASAP7_75t_L g461 ( 
.A1(n_401),
.A2(n_71),
.B(n_72),
.C(n_73),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_374),
.B(n_74),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_403),
.B(n_386),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_405),
.B(n_77),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_370),
.B(n_149),
.Y(n_465)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_403),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_396),
.B(n_78),
.Y(n_467)
);

O2A1O1Ixp5_ASAP7_75t_L g468 ( 
.A1(n_406),
.A2(n_412),
.B(n_419),
.C(n_373),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_375),
.A2(n_79),
.B(n_81),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_392),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_379),
.B(n_82),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_L g472 ( 
.A1(n_411),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_R g473 ( 
.A(n_387),
.B(n_87),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_359),
.B(n_89),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_387),
.B(n_148),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_391),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_356),
.B(n_90),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_456),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_446),
.A2(n_412),
.B(n_419),
.Y(n_479)
);

BUFx2_ASAP7_75t_R g480 ( 
.A(n_432),
.Y(n_480)
);

INVx2_ASAP7_75t_SL g481 ( 
.A(n_438),
.Y(n_481)
);

OAI21x1_ASAP7_75t_L g482 ( 
.A1(n_422),
.A2(n_413),
.B(n_417),
.Y(n_482)
);

OAI21x1_ASAP7_75t_L g483 ( 
.A1(n_468),
.A2(n_474),
.B(n_477),
.Y(n_483)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_443),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_440),
.Y(n_485)
);

AOI22x1_ASAP7_75t_L g486 ( 
.A1(n_431),
.A2(n_407),
.B1(n_361),
.B2(n_357),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_473),
.Y(n_487)
);

OAI21x1_ASAP7_75t_L g488 ( 
.A1(n_471),
.A2(n_416),
.B(n_414),
.Y(n_488)
);

INVx5_ASAP7_75t_L g489 ( 
.A(n_456),
.Y(n_489)
);

BUFx4f_ASAP7_75t_SL g490 ( 
.A(n_452),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_425),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_436),
.Y(n_492)
);

BUFx12f_ASAP7_75t_L g493 ( 
.A(n_476),
.Y(n_493)
);

OA21x2_ASAP7_75t_L g494 ( 
.A1(n_451),
.A2(n_418),
.B(n_381),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_444),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_434),
.A2(n_415),
.B(n_369),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_439),
.B(n_385),
.Y(n_497)
);

OAI21x1_ASAP7_75t_L g498 ( 
.A1(n_455),
.A2(n_415),
.B(n_393),
.Y(n_498)
);

INVx8_ASAP7_75t_L g499 ( 
.A(n_456),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_454),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_436),
.Y(n_501)
);

NAND2x1p5_ASAP7_75t_L g502 ( 
.A(n_441),
.B(n_391),
.Y(n_502)
);

INVx5_ASAP7_75t_L g503 ( 
.A(n_476),
.Y(n_503)
);

BUFx12f_ASAP7_75t_L g504 ( 
.A(n_476),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_426),
.B(n_410),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_444),
.Y(n_506)
);

OAI21x1_ASAP7_75t_L g507 ( 
.A1(n_459),
.A2(n_430),
.B(n_447),
.Y(n_507)
);

AOI22x1_ASAP7_75t_L g508 ( 
.A1(n_433),
.A2(n_396),
.B1(n_365),
.B2(n_384),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_444),
.Y(n_509)
);

NAND2x1p5_ASAP7_75t_L g510 ( 
.A(n_441),
.B(n_365),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_428),
.Y(n_511)
);

OAI21x1_ASAP7_75t_L g512 ( 
.A1(n_435),
.A2(n_403),
.B(n_93),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_421),
.A2(n_389),
.B(n_94),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_424),
.Y(n_514)
);

NAND2x1p5_ASAP7_75t_L g515 ( 
.A(n_445),
.B(n_389),
.Y(n_515)
);

BUFx2_ASAP7_75t_SL g516 ( 
.A(n_462),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_470),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_423),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_466),
.Y(n_519)
);

CKINVDCx16_ASAP7_75t_R g520 ( 
.A(n_463),
.Y(n_520)
);

BUFx4f_ASAP7_75t_L g521 ( 
.A(n_458),
.Y(n_521)
);

INVx1_ASAP7_75t_SL g522 ( 
.A(n_427),
.Y(n_522)
);

INVx5_ASAP7_75t_L g523 ( 
.A(n_449),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_491),
.B(n_475),
.Y(n_524)
);

CKINVDCx6p67_ASAP7_75t_R g525 ( 
.A(n_493),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_490),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_SL g527 ( 
.A1(n_513),
.A2(n_464),
.B1(n_465),
.B2(n_453),
.Y(n_527)
);

NAND2x1p5_ASAP7_75t_L g528 ( 
.A(n_489),
.B(n_467),
.Y(n_528)
);

AO21x1_ASAP7_75t_L g529 ( 
.A1(n_513),
.A2(n_429),
.B(n_442),
.Y(n_529)
);

AO21x1_ASAP7_75t_SL g530 ( 
.A1(n_496),
.A2(n_472),
.B(n_421),
.Y(n_530)
);

BUFx2_ASAP7_75t_SL g531 ( 
.A(n_489),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_485),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_504),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_514),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_L g535 ( 
.A1(n_496),
.A2(n_448),
.B1(n_437),
.B2(n_469),
.Y(n_535)
);

NAND2x1_ASAP7_75t_L g536 ( 
.A(n_492),
.B(n_460),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_SL g537 ( 
.A1(n_515),
.A2(n_450),
.B1(n_457),
.B2(n_461),
.Y(n_537)
);

BUFx2_ASAP7_75t_R g538 ( 
.A(n_487),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_500),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_510),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_511),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_499),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_510),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_509),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_SL g545 ( 
.A1(n_515),
.A2(n_523),
.B1(n_522),
.B2(n_520),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_517),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_478),
.Y(n_547)
);

INVx6_ASAP7_75t_L g548 ( 
.A(n_489),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_499),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_SL g550 ( 
.A1(n_523),
.A2(n_91),
.B1(n_96),
.B2(n_98),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_497),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_482),
.Y(n_552)
);

CKINVDCx11_ASAP7_75t_R g553 ( 
.A(n_484),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_497),
.Y(n_554)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_479),
.A2(n_99),
.B(n_100),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_518),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_SL g557 ( 
.A1(n_523),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_557)
);

AOI21x1_ASAP7_75t_L g558 ( 
.A1(n_479),
.A2(n_104),
.B(n_105),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_505),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_505),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_486),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_495),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_481),
.Y(n_563)
);

BUFx2_ASAP7_75t_R g564 ( 
.A(n_516),
.Y(n_564)
);

NAND2x1p5_ASAP7_75t_L g565 ( 
.A(n_503),
.B(n_110),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_548),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_541),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_548),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_551),
.B(n_522),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_532),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_546),
.Y(n_571)
);

NAND2xp33_ASAP7_75t_R g572 ( 
.A(n_561),
.B(n_494),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_534),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_554),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_539),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_525),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_527),
.A2(n_521),
.B1(n_480),
.B2(n_508),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_524),
.B(n_519),
.Y(n_578)
);

O2A1O1Ixp33_ASAP7_75t_L g579 ( 
.A1(n_529),
.A2(n_492),
.B(n_501),
.C(n_506),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_563),
.B(n_519),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_526),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_563),
.B(n_503),
.Y(n_582)
);

NAND2xp33_ASAP7_75t_R g583 ( 
.A(n_527),
.B(n_494),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_562),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_544),
.B(n_480),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_556),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_544),
.B(n_503),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_552),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_559),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_560),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_545),
.A2(n_498),
.B1(n_521),
.B2(n_512),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_547),
.Y(n_592)
);

NOR2x1p5_ASAP7_75t_L g593 ( 
.A(n_533),
.B(n_478),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_553),
.B(n_545),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_547),
.B(n_478),
.Y(n_595)
);

INVxp67_ASAP7_75t_L g596 ( 
.A(n_531),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_548),
.Y(n_597)
);

NAND2xp33_ASAP7_75t_SL g598 ( 
.A(n_535),
.B(n_501),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_526),
.Y(n_599)
);

AND2x4_ASAP7_75t_L g600 ( 
.A(n_540),
.B(n_488),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_537),
.A2(n_499),
.B1(n_507),
.B2(n_502),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_R g602 ( 
.A(n_533),
.B(n_502),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_536),
.Y(n_603)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_540),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_553),
.B(n_483),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_565),
.Y(n_606)
);

OR2x6_ASAP7_75t_L g607 ( 
.A(n_528),
.B(n_565),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_542),
.B(n_113),
.Y(n_608)
);

OAI21x1_ASAP7_75t_SL g609 ( 
.A1(n_535),
.A2(n_114),
.B(n_116),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_558),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_543),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_543),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_570),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_577),
.A2(n_537),
.B1(n_530),
.B2(n_550),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_575),
.B(n_557),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_603),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_586),
.B(n_557),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_589),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_574),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_574),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_569),
.B(n_549),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_588),
.B(n_550),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_567),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_588),
.B(n_528),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_578),
.B(n_564),
.Y(n_625)
);

OR2x2_ASAP7_75t_L g626 ( 
.A(n_605),
.B(n_584),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_567),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_571),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_590),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_580),
.B(n_555),
.Y(n_630)
);

NOR2x1_ASAP7_75t_SL g631 ( 
.A(n_607),
.B(n_538),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_600),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_604),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_600),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_612),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_612),
.Y(n_636)
);

OR2x2_ASAP7_75t_L g637 ( 
.A(n_573),
.B(n_117),
.Y(n_637)
);

NOR2x1_ASAP7_75t_L g638 ( 
.A(n_582),
.B(n_118),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_610),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_610),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_594),
.A2(n_121),
.B1(n_122),
.B2(n_124),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_611),
.Y(n_642)
);

OAI21x1_ASAP7_75t_L g643 ( 
.A1(n_591),
.A2(n_126),
.B(n_129),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_603),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_604),
.B(n_130),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_601),
.A2(n_132),
.B1(n_134),
.B2(n_135),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_632),
.B(n_591),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_618),
.B(n_613),
.Y(n_648)
);

INVxp67_ASAP7_75t_SL g649 ( 
.A(n_633),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_632),
.B(n_607),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_619),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_620),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_635),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_628),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_629),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_634),
.B(n_624),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_634),
.B(n_626),
.Y(n_657)
);

OAI21xp5_ASAP7_75t_L g658 ( 
.A1(n_614),
.A2(n_598),
.B(n_579),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_626),
.B(n_592),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_644),
.Y(n_660)
);

NAND2x1p5_ASAP7_75t_L g661 ( 
.A(n_645),
.B(n_606),
.Y(n_661)
);

HB1xp67_ASAP7_75t_L g662 ( 
.A(n_636),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_615),
.B(n_617),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_615),
.B(n_596),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_622),
.B(n_601),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_622),
.B(n_585),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_644),
.B(n_581),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_616),
.B(n_581),
.Y(n_668)
);

HB1xp67_ASAP7_75t_L g669 ( 
.A(n_616),
.Y(n_669)
);

AND2x4_ASAP7_75t_SL g670 ( 
.A(n_624),
.B(n_607),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_617),
.B(n_587),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_660),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_667),
.B(n_639),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_653),
.Y(n_674)
);

HB1xp67_ASAP7_75t_L g675 ( 
.A(n_669),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_662),
.Y(n_676)
);

BUFx2_ASAP7_75t_L g677 ( 
.A(n_649),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_648),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_660),
.Y(n_679)
);

INVx2_ASAP7_75t_SL g680 ( 
.A(n_668),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_663),
.B(n_642),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_667),
.B(n_639),
.Y(n_682)
);

OR2x2_ASAP7_75t_L g683 ( 
.A(n_657),
.B(n_640),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_668),
.B(n_640),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_657),
.B(n_642),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_655),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_651),
.Y(n_687)
);

NOR3xp33_ASAP7_75t_L g688 ( 
.A(n_674),
.B(n_658),
.C(n_676),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_678),
.A2(n_665),
.B1(n_583),
.B2(n_666),
.Y(n_689)
);

AOI211xp5_ASAP7_75t_L g690 ( 
.A1(n_687),
.A2(n_665),
.B(n_664),
.C(n_666),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_686),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_675),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_677),
.Y(n_693)
);

NAND2x1p5_ASAP7_75t_L g694 ( 
.A(n_680),
.B(n_645),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_680),
.B(n_684),
.Y(n_695)
);

OR2x2_ASAP7_75t_L g696 ( 
.A(n_681),
.B(n_671),
.Y(n_696)
);

NAND5xp2_ASAP7_75t_L g697 ( 
.A(n_684),
.B(n_661),
.C(n_630),
.D(n_625),
.E(n_641),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_685),
.Y(n_698)
);

AOI21xp33_ASAP7_75t_L g699 ( 
.A1(n_689),
.A2(n_691),
.B(n_693),
.Y(n_699)
);

AOI21xp33_ASAP7_75t_SL g700 ( 
.A1(n_688),
.A2(n_599),
.B(n_661),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_692),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_698),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_689),
.A2(n_583),
.B1(n_647),
.B2(n_673),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_702),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_701),
.B(n_695),
.Y(n_705)
);

AND2x2_ASAP7_75t_SL g706 ( 
.A(n_703),
.B(n_625),
.Y(n_706)
);

AOI22xp5_ASAP7_75t_L g707 ( 
.A1(n_699),
.A2(n_690),
.B1(n_647),
.B2(n_659),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_700),
.Y(n_708)
);

INVx1_ASAP7_75t_SL g709 ( 
.A(n_708),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_705),
.B(n_576),
.Y(n_710)
);

NOR3x1_ASAP7_75t_L g711 ( 
.A(n_704),
.B(n_637),
.C(n_621),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_707),
.B(n_659),
.Y(n_712)
);

AOI211xp5_ASAP7_75t_L g713 ( 
.A1(n_709),
.A2(n_697),
.B(n_704),
.C(n_637),
.Y(n_713)
);

OAI21xp33_ASAP7_75t_L g714 ( 
.A1(n_712),
.A2(n_710),
.B(n_706),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_711),
.A2(n_631),
.B(n_576),
.Y(n_715)
);

O2A1O1Ixp33_ASAP7_75t_L g716 ( 
.A1(n_713),
.A2(n_646),
.B(n_609),
.C(n_661),
.Y(n_716)
);

NAND2xp33_ASAP7_75t_SL g717 ( 
.A(n_714),
.B(n_602),
.Y(n_717)
);

NAND4xp25_ASAP7_75t_L g718 ( 
.A(n_715),
.B(n_638),
.C(n_598),
.D(n_679),
.Y(n_718)
);

AOI322xp5_ASAP7_75t_L g719 ( 
.A1(n_714),
.A2(n_685),
.A3(n_682),
.B1(n_673),
.B2(n_631),
.C1(n_656),
.C2(n_651),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_719),
.Y(n_720)
);

OAI211xp5_ASAP7_75t_L g721 ( 
.A1(n_717),
.A2(n_602),
.B(n_679),
.C(n_672),
.Y(n_721)
);

NOR2x1_ASAP7_75t_L g722 ( 
.A(n_718),
.B(n_593),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_716),
.B(n_694),
.Y(n_723)
);

NOR2x1_ASAP7_75t_L g724 ( 
.A(n_718),
.B(n_672),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_717),
.Y(n_725)
);

NOR2x1_ASAP7_75t_L g726 ( 
.A(n_718),
.B(n_672),
.Y(n_726)
);

AOI22x1_ASAP7_75t_L g727 ( 
.A1(n_725),
.A2(n_679),
.B1(n_608),
.B2(n_597),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_720),
.Y(n_728)
);

AOI221xp5_ASAP7_75t_SL g729 ( 
.A1(n_723),
.A2(n_696),
.B1(n_652),
.B2(n_595),
.C(n_660),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_722),
.Y(n_730)
);

AND3x2_ASAP7_75t_L g731 ( 
.A(n_721),
.B(n_682),
.C(n_650),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_724),
.A2(n_572),
.B1(n_643),
.B2(n_652),
.Y(n_732)
);

NOR2x1_ASAP7_75t_L g733 ( 
.A(n_726),
.B(n_568),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_730),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_728),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_727),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_732),
.Y(n_737)
);

BUFx2_ASAP7_75t_L g738 ( 
.A(n_733),
.Y(n_738)
);

INVx1_ASAP7_75t_SL g739 ( 
.A(n_731),
.Y(n_739)
);

INVx1_ASAP7_75t_SL g740 ( 
.A(n_729),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_728),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_735),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_735),
.B(n_597),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_734),
.Y(n_744)
);

XOR2xp5_ASAP7_75t_L g745 ( 
.A(n_741),
.B(n_597),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_740),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_739),
.B(n_597),
.Y(n_747)
);

AOI22xp5_ASAP7_75t_L g748 ( 
.A1(n_746),
.A2(n_737),
.B1(n_736),
.B2(n_738),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_747),
.A2(n_629),
.B1(n_643),
.B2(n_566),
.Y(n_749)
);

INVx5_ASAP7_75t_L g750 ( 
.A(n_744),
.Y(n_750)
);

AO22x2_ASAP7_75t_L g751 ( 
.A1(n_742),
.A2(n_568),
.B1(n_683),
.B2(n_650),
.Y(n_751)
);

OAI22x1_ASAP7_75t_L g752 ( 
.A1(n_748),
.A2(n_745),
.B1(n_743),
.B2(n_650),
.Y(n_752)
);

OAI22x1_ASAP7_75t_SL g753 ( 
.A1(n_750),
.A2(n_566),
.B1(n_138),
.B2(n_139),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_751),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_SL g755 ( 
.A1(n_754),
.A2(n_749),
.B1(n_566),
.B2(n_670),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_752),
.A2(n_572),
.B1(n_566),
.B2(n_670),
.Y(n_756)
);

AOI21xp33_ASAP7_75t_SL g757 ( 
.A1(n_756),
.A2(n_753),
.B(n_140),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_757),
.A2(n_755),
.B1(n_656),
.B2(n_654),
.Y(n_758)
);

AOI221xp5_ASAP7_75t_L g759 ( 
.A1(n_758),
.A2(n_623),
.B1(n_627),
.B2(n_628),
.C(n_654),
.Y(n_759)
);

AOI211xp5_ASAP7_75t_L g760 ( 
.A1(n_759),
.A2(n_136),
.B(n_141),
.C(n_142),
.Y(n_760)
);


endmodule