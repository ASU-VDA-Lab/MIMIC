module fake_netlist_1_8056_n_37 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_37);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_37;
wire n_20;
wire n_36;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_30;
wire n_13;
wire n_26;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_3), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_2), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_10), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_4), .Y(n_14) );
INVx1_ASAP7_75t_SL g15 ( .A(n_10), .Y(n_15) );
NAND2xp5_ASAP7_75t_SL g16 ( .A(n_4), .B(n_9), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_8), .Y(n_17) );
AOI22xp5_ASAP7_75t_L g18 ( .A1(n_13), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_18) );
NOR2xp33_ASAP7_75t_L g19 ( .A(n_17), .B(n_0), .Y(n_19) );
AOI21x1_ASAP7_75t_L g20 ( .A1(n_13), .A2(n_1), .B(n_3), .Y(n_20) );
INVx4_ASAP7_75t_L g21 ( .A(n_13), .Y(n_21) );
AOI221xp5_ASAP7_75t_L g22 ( .A1(n_14), .A2(n_5), .B1(n_6), .B2(n_7), .C(n_8), .Y(n_22) );
AO31x2_ASAP7_75t_L g23 ( .A1(n_21), .A2(n_14), .A3(n_16), .B(n_15), .Y(n_23) );
CKINVDCx16_ASAP7_75t_R g24 ( .A(n_18), .Y(n_24) );
AO21x2_ASAP7_75t_L g25 ( .A1(n_20), .A2(n_16), .B(n_11), .Y(n_25) );
INVx2_ASAP7_75t_SL g26 ( .A(n_25), .Y(n_26) );
NAND2xp5_ASAP7_75t_L g27 ( .A(n_23), .B(n_21), .Y(n_27) );
NAND2xp5_ASAP7_75t_L g28 ( .A(n_23), .B(n_19), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_28), .B(n_23), .Y(n_29) );
AOI22xp33_ASAP7_75t_L g30 ( .A1(n_27), .A2(n_25), .B1(n_24), .B2(n_22), .Y(n_30) );
OAI211xp5_ASAP7_75t_SL g31 ( .A1(n_30), .A2(n_15), .B(n_26), .C(n_12), .Y(n_31) );
AOI221x1_ASAP7_75t_L g32 ( .A1(n_29), .A2(n_26), .B1(n_23), .B2(n_25), .C(n_9), .Y(n_32) );
INVx1_ASAP7_75t_SL g33 ( .A(n_31), .Y(n_33) );
INVx5_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
CKINVDCx5p33_ASAP7_75t_R g35 ( .A(n_31), .Y(n_35) );
OAI22xp5_ASAP7_75t_SL g36 ( .A1(n_35), .A2(n_23), .B1(n_6), .B2(n_7), .Y(n_36) );
AOI22xp5_ASAP7_75t_L g37 ( .A1(n_36), .A2(n_33), .B1(n_34), .B2(n_5), .Y(n_37) );
endmodule