module fake_jpeg_8819_n_46 (n_3, n_2, n_1, n_0, n_4, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

INVx6_ASAP7_75t_SL g8 ( 
.A(n_0),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx16f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_14),
.A2(n_7),
.B1(n_11),
.B2(n_8),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_9),
.B(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_17),
.A2(n_18),
.B1(n_11),
.B2(n_8),
.Y(n_22)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_3),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_SL g25 ( 
.A(n_19),
.B(n_20),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_7),
.B(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_14),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_27),
.A2(n_6),
.B(n_10),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_16),
.C(n_18),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_8),
.C(n_26),
.Y(n_33)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_30),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_20),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_31),
.A2(n_24),
.B1(n_25),
.B2(n_17),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_13),
.B1(n_6),
.B2(n_29),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_6),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_6),
.B(n_26),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_28),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_39),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_10),
.C(n_4),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_41),
.Y(n_44)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

AOI321xp33_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_4),
.A3(n_5),
.B1(n_10),
.B2(n_38),
.C(n_44),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_43),
.C(n_10),
.Y(n_46)
);


endmodule