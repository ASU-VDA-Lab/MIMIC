module fake_jpeg_9112_n_342 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_41),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_23),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_40),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_8),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_43),
.Y(n_53)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_49),
.Y(n_99)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_57),
.Y(n_75)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_46),
.B(n_19),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_58),
.B(n_56),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_63),
.Y(n_78)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_65),
.Y(n_81)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_39),
.A2(n_29),
.B1(n_20),
.B2(n_33),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_67),
.A2(n_39),
.B1(n_43),
.B2(n_34),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_73),
.B(n_94),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_61),
.B(n_48),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_74),
.B(n_79),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_50),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_84),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_22),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_52),
.A2(n_20),
.B1(n_29),
.B2(n_33),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_85),
.B1(n_90),
.B2(n_25),
.Y(n_101)
);

CKINVDCx12_ASAP7_75t_R g84 ( 
.A(n_49),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_71),
.A2(n_29),
.B1(n_20),
.B2(n_22),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_86),
.A2(n_91),
.B1(n_93),
.B2(n_95),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_59),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_92),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_55),
.B(n_32),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_98),
.B(n_17),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_71),
.A2(n_25),
.B1(n_32),
.B2(n_30),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_59),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_97),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_62),
.B(n_30),
.Y(n_98)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_100),
.B(n_104),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_101),
.Y(n_142)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

MAJx2_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_62),
.C(n_45),
.Y(n_106)
);

MAJx2_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_111),
.C(n_115),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_75),
.A2(n_70),
.B1(n_69),
.B2(n_51),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_107),
.A2(n_120),
.B1(n_121),
.B2(n_125),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_109),
.B(n_122),
.Y(n_136)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_110),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_26),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx4_ASAP7_75t_SL g145 ( 
.A(n_112),
.Y(n_145)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_113),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_87),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_114),
.B(n_118),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_26),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_87),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g120 ( 
.A1(n_86),
.A2(n_65),
.B1(n_69),
.B2(n_70),
.Y(n_120)
);

AO21x2_ASAP7_75t_L g121 ( 
.A1(n_76),
.A2(n_44),
.B(n_51),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_81),
.Y(n_122)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_124),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_75),
.A2(n_37),
.B1(n_26),
.B2(n_44),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_79),
.B(n_68),
.C(n_26),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_93),
.Y(n_140)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_129),
.Y(n_132)
);

NAND2x1_ASAP7_75t_SL g130 ( 
.A(n_121),
.B(n_18),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_130),
.A2(n_133),
.B(n_103),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_121),
.A2(n_94),
.B(n_80),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_140),
.B(n_152),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_115),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_156),
.Y(n_158)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_148),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_107),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_151),
.Y(n_183)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_125),
.A2(n_98),
.B(n_89),
.Y(n_152)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

AND2x6_ASAP7_75t_L g155 ( 
.A(n_106),
.B(n_7),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_155),
.Y(n_163)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_108),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_142),
.A2(n_120),
.B1(n_119),
.B2(n_126),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_157),
.Y(n_187)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_160),
.Y(n_189)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_149),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_132),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_164),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_128),
.Y(n_162)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_162),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_151),
.A2(n_142),
.B1(n_150),
.B2(n_140),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_165),
.A2(n_167),
.B1(n_168),
.B2(n_170),
.Y(n_202)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_166),
.B(n_173),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_146),
.A2(n_120),
.B1(n_116),
.B2(n_129),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_130),
.A2(n_76),
.B1(n_95),
.B2(n_80),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_130),
.A2(n_146),
.B1(n_155),
.B2(n_136),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_176),
.Y(n_191)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_134),
.Y(n_173)
);

AO21x2_ASAP7_75t_L g174 ( 
.A1(n_138),
.A2(n_123),
.B(n_110),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_174),
.A2(n_137),
.B1(n_134),
.B2(n_147),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_156),
.B(n_73),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_175),
.Y(n_188)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_135),
.A2(n_109),
.B(n_17),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_182),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_152),
.A2(n_91),
.B1(n_143),
.B2(n_138),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_179),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_135),
.A2(n_91),
.B1(n_102),
.B2(n_96),
.Y(n_181)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_181),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_84),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_144),
.A2(n_19),
.B(n_92),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_153),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_169),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_190),
.B(n_197),
.Y(n_233)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_195),
.Y(n_217)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_174),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_158),
.B(n_131),
.Y(n_198)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_198),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_158),
.B(n_131),
.Y(n_199)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_199),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_200),
.A2(n_201),
.B1(n_173),
.B2(n_171),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_163),
.A2(n_137),
.B1(n_154),
.B2(n_99),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_184),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_206),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_153),
.Y(n_205)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_205),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_165),
.Y(n_206)
);

INVx13_ASAP7_75t_L g208 ( 
.A(n_174),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_209),
.Y(n_223)
);

INVx13_ASAP7_75t_L g209 ( 
.A(n_174),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_167),
.B(n_0),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_211),
.Y(n_227)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_168),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_113),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_180),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_226),
.C(n_228),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_182),
.Y(n_214)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_193),
.B(n_180),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_216),
.B(n_221),
.Y(n_240)
);

AO21x2_ASAP7_75t_L g220 ( 
.A1(n_208),
.A2(n_176),
.B(n_170),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_220),
.A2(n_208),
.B1(n_209),
.B2(n_195),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_194),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_205),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_232),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_189),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_230),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_162),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_191),
.B(n_178),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_160),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_238),
.C(n_196),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_188),
.B(n_159),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_188),
.B(n_172),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_235),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_207),
.Y(n_232)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_196),
.Y(n_234)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_234),
.Y(n_242)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_189),
.Y(n_235)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_236),
.Y(n_245)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_198),
.Y(n_237)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_237),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_202),
.B(n_99),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_239),
.A2(n_233),
.B(n_232),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_243),
.A2(n_259),
.B1(n_214),
.B2(n_112),
.Y(n_278)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_244),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_220),
.A2(n_185),
.B1(n_212),
.B2(n_203),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_246),
.A2(n_251),
.B1(n_262),
.B2(n_24),
.Y(n_281)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_234),
.Y(n_247)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_220),
.A2(n_185),
.B1(n_192),
.B2(n_187),
.Y(n_248)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_248),
.Y(n_267)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_217),
.Y(n_249)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_249),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_220),
.A2(n_206),
.B1(n_211),
.B2(n_186),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_222),
.Y(n_254)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_254),
.Y(n_273)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_224),
.Y(n_256)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_256),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_227),
.A2(n_201),
.B1(n_200),
.B2(n_204),
.Y(n_257)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_257),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_223),
.A2(n_186),
.B1(n_199),
.B2(n_197),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_227),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_260),
.A2(n_145),
.B1(n_132),
.B2(n_24),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_216),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_215),
.A2(n_210),
.B1(n_190),
.B2(n_171),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_226),
.C(n_229),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_268),
.C(n_270),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_266),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_218),
.C(n_228),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_238),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_245),
.A2(n_210),
.B1(n_219),
.B2(n_214),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_271),
.A2(n_281),
.B1(n_249),
.B2(n_243),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_241),
.C(n_240),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_275),
.C(n_263),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_258),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_274),
.B(n_273),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_213),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_259),
.Y(n_282)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_278),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_255),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_282),
.B(n_297),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_269),
.A2(n_241),
.B(n_244),
.Y(n_283)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_283),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_276),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_285),
.B(n_287),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_286),
.A2(n_295),
.B1(n_285),
.B2(n_267),
.Y(n_299)
);

NAND3xp33_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_262),
.C(n_246),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_288),
.A2(n_291),
.B(n_294),
.Y(n_306)
);

AO22x1_ASAP7_75t_L g290 ( 
.A1(n_281),
.A2(n_252),
.B1(n_250),
.B2(n_242),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_290),
.A2(n_12),
.B(n_16),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_31),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_0),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_268),
.A2(n_11),
.B(n_16),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_279),
.A2(n_35),
.B1(n_28),
.B2(n_24),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_12),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_296),
.B(n_272),
.C(n_264),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_304),
.C(n_307),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_299),
.A2(n_301),
.B1(n_310),
.B2(n_302),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_297),
.A2(n_265),
.B(n_275),
.Y(n_300)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_300),
.Y(n_316)
);

AO21x1_ASAP7_75t_L g319 ( 
.A1(n_302),
.A2(n_9),
.B(n_2),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_293),
.A2(n_35),
.B1(n_28),
.B2(n_24),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_303),
.A2(n_35),
.B1(n_28),
.B2(n_31),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_31),
.C(n_18),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_288),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_10),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_290),
.A2(n_284),
.B1(n_282),
.B2(n_289),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_31),
.C(n_0),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_309),
.A2(n_1),
.B(n_31),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_311),
.B(n_0),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_312),
.A2(n_321),
.B(n_309),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_313),
.B(n_315),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_306),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_319),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_320),
.Y(n_329)
);

OAI21x1_ASAP7_75t_L g321 ( 
.A1(n_308),
.A2(n_31),
.B(n_2),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_308),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_323),
.B(n_12),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_298),
.C(n_304),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_324),
.A2(n_326),
.B(n_328),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_9),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_1),
.C(n_3),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_9),
.C(n_3),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_330),
.B(n_333),
.Y(n_336)
);

OAI21x1_ASAP7_75t_L g331 ( 
.A1(n_323),
.A2(n_6),
.B(n_3),
.Y(n_331)
);

OAI21x1_ASAP7_75t_SL g335 ( 
.A1(n_331),
.A2(n_334),
.B(n_326),
.Y(n_335)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_329),
.Y(n_333)
);

NOR3xp33_ASAP7_75t_L g337 ( 
.A(n_335),
.B(n_332),
.C(n_327),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_322),
.B(n_336),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_4),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_4),
.B(n_5),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_5),
.B1(n_6),
.B2(n_14),
.Y(n_341)
);

A2O1A1Ixp33_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_15),
.B(n_16),
.C(n_1),
.Y(n_342)
);


endmodule