module real_aes_4220_n_234 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_234);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_234;
wire n_480;
wire n_476;
wire n_758;
wire n_887;
wire n_436;
wire n_599;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_254;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_857;
wire n_461;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_884;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_763;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_892;
wire n_372;
wire n_528;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_875;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_898;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_598;
wire n_756;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_899;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_888;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_279;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_849;
wire n_554;
wire n_475;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
wire n_862;
HB1xp67_ASAP7_75t_L g245 ( .A(n_0), .Y(n_245) );
AND2x4_ASAP7_75t_L g668 ( .A(n_0), .B(n_224), .Y(n_668) );
AND2x4_ASAP7_75t_L g673 ( .A(n_0), .B(n_674), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_1), .A2(n_39), .B1(n_406), .B2(n_408), .Y(n_405) );
INVx1_ASAP7_75t_L g570 ( .A(n_2), .Y(n_570) );
AO22x1_ASAP7_75t_L g706 ( .A1(n_2), .A2(n_6), .B1(n_669), .B2(n_679), .Y(n_706) );
INVx1_ASAP7_75t_L g876 ( .A(n_3), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_4), .A2(n_65), .B1(n_308), .B2(n_312), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_5), .A2(n_164), .B1(n_672), .B2(n_675), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_7), .A2(n_15), .B1(n_606), .B2(n_607), .Y(n_605) );
XNOR2x2_ASAP7_75t_L g600 ( .A(n_8), .B(n_601), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_9), .A2(n_77), .B1(n_501), .B2(n_502), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_10), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_11), .A2(n_63), .B1(n_349), .B2(n_351), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g868 ( .A1(n_12), .A2(n_23), .B1(n_338), .B2(n_520), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_13), .A2(n_18), .B1(n_484), .B2(n_879), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_14), .A2(n_127), .B1(n_498), .B2(n_499), .Y(n_882) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_16), .A2(n_181), .B1(n_561), .B2(n_592), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_17), .A2(n_103), .B1(n_493), .B2(n_502), .Y(n_543) );
INVx1_ASAP7_75t_L g628 ( .A(n_19), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_20), .A2(n_167), .B1(n_561), .B2(n_636), .Y(n_635) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_21), .A2(n_97), .B1(n_696), .B2(n_704), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_22), .A2(n_182), .B1(n_419), .B2(n_422), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g564 ( .A1(n_24), .A2(n_29), .B1(n_382), .B2(n_565), .C(n_568), .Y(n_564) );
INVx1_ASAP7_75t_L g363 ( .A(n_25), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_26), .A2(n_67), .B1(n_411), .B2(n_412), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_27), .A2(n_173), .B1(n_338), .B2(n_578), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_28), .A2(n_141), .B1(n_498), .B2(n_499), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g583 ( .A1(n_30), .A2(n_481), .B(n_584), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_31), .A2(n_114), .B1(n_481), .B2(n_485), .Y(n_524) );
XNOR2x1_ASAP7_75t_L g355 ( .A(n_32), .B(n_356), .Y(n_355) );
AOI21xp5_ASAP7_75t_L g874 ( .A1(n_33), .A2(n_565), .B(n_875), .Y(n_874) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_34), .B(n_169), .Y(n_243) );
INVx1_ASAP7_75t_L g280 ( .A(n_34), .Y(n_280) );
INVxp67_ASAP7_75t_L g293 ( .A(n_34), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_35), .A2(n_101), .B1(n_481), .B2(n_495), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_36), .A2(n_130), .B1(n_333), .B2(n_554), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_37), .A2(n_69), .B1(n_362), .B2(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_38), .B(n_638), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_40), .A2(n_139), .B1(n_326), .B2(n_604), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_41), .A2(n_59), .B1(n_492), .B2(n_493), .Y(n_523) );
XNOR2x1_ASAP7_75t_L g573 ( .A(n_42), .B(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_43), .B(n_265), .Y(n_276) );
INVx1_ASAP7_75t_L g516 ( .A(n_44), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_45), .A2(n_210), .B1(n_610), .B2(n_611), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g414 ( .A1(n_46), .A2(n_113), .B1(n_415), .B2(n_416), .Y(n_414) );
CKINVDCx20_ASAP7_75t_R g427 ( .A(n_47), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_48), .A2(n_213), .B1(n_484), .B2(n_485), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_49), .A2(n_185), .B1(n_482), .B2(n_484), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_50), .A2(n_191), .B1(n_373), .B2(n_375), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_51), .A2(n_199), .B1(n_620), .B2(n_622), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_52), .A2(n_85), .B1(n_495), .B2(n_496), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_53), .A2(n_138), .B1(n_665), .B2(n_669), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_54), .A2(n_145), .B1(n_351), .B2(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g569 ( .A(n_55), .Y(n_569) );
INVx2_ASAP7_75t_L g240 ( .A(n_56), .Y(n_240) );
INVx1_ASAP7_75t_L g667 ( .A(n_57), .Y(n_667) );
AND2x4_ASAP7_75t_L g670 ( .A(n_57), .B(n_240), .Y(n_670) );
INVx1_ASAP7_75t_SL g702 ( .A(n_57), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_58), .A2(n_155), .B1(n_338), .B2(n_520), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_60), .A2(n_258), .B(n_283), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_61), .A2(n_151), .B1(n_679), .B2(n_686), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_62), .A2(n_195), .B1(n_482), .B2(n_485), .Y(n_880) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_64), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_66), .A2(n_211), .B1(n_443), .B2(n_444), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_68), .A2(n_171), .B1(n_498), .B2(n_499), .Y(n_497) );
INVx1_ASAP7_75t_L g385 ( .A(n_70), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_71), .A2(n_230), .B1(n_496), .B2(n_501), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g869 ( .A1(n_72), .A2(n_165), .B1(n_373), .B2(n_870), .Y(n_869) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_73), .A2(n_131), .B1(n_672), .B2(n_694), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_74), .A2(n_75), .B1(n_485), .B2(n_492), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_76), .A2(n_160), .B1(n_665), .B2(n_669), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_78), .A2(n_142), .B1(n_669), .B2(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g266 ( .A(n_79), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_79), .B(n_168), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_80), .A2(n_214), .B1(n_349), .B2(n_375), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_81), .A2(n_122), .B1(n_346), .B2(n_417), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g325 ( .A1(n_82), .A2(n_187), .B1(n_326), .B2(n_330), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_83), .A2(n_146), .B1(n_417), .B2(n_440), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_84), .A2(n_112), .B1(n_438), .B2(n_439), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_86), .A2(n_137), .B1(n_672), .B2(n_683), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_87), .A2(n_176), .B1(n_481), .B2(n_482), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_88), .A2(n_124), .B1(n_362), .B2(n_621), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_89), .A2(n_205), .B1(n_419), .B2(n_446), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_90), .A2(n_93), .B1(n_672), .B2(n_675), .Y(n_680) );
XNOR2x1_ASAP7_75t_L g530 ( .A(n_91), .B(n_531), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_92), .A2(n_194), .B1(n_438), .B2(n_614), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_94), .A2(n_170), .B1(n_683), .B2(n_761), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_95), .A2(n_116), .B1(n_333), .B2(n_338), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_96), .A2(n_178), .B1(n_367), .B2(n_398), .Y(n_397) );
XNOR2x1_ASAP7_75t_L g865 ( .A(n_97), .B(n_866), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_97), .A2(n_890), .B1(n_894), .B2(n_896), .Y(n_889) );
AOI22xp5_ASAP7_75t_L g690 ( .A1(n_98), .A2(n_212), .B1(n_672), .B2(n_675), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_99), .A2(n_133), .B1(n_349), .B2(n_351), .Y(n_348) );
INVx1_ASAP7_75t_L g872 ( .A(n_100), .Y(n_872) );
AOI21xp33_ASAP7_75t_L g536 ( .A1(n_102), .A2(n_487), .B(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g538 ( .A(n_104), .Y(n_538) );
INVx1_ASAP7_75t_L g365 ( .A(n_105), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_106), .A2(n_223), .B1(n_492), .B2(n_493), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_107), .A2(n_132), .B1(n_554), .B2(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_108), .B(n_402), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_109), .A2(n_140), .B1(n_343), .B2(n_346), .Y(n_342) );
XOR2x2_ASAP7_75t_L g510 ( .A(n_110), .B(n_511), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g640 ( .A1(n_111), .A2(n_367), .B(n_641), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_115), .A2(n_117), .B1(n_333), .B2(n_375), .Y(n_374) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_118), .A2(n_209), .B1(n_675), .B2(n_701), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_119), .A2(n_159), .B1(n_362), .B2(n_394), .Y(n_588) );
INVx1_ASAP7_75t_L g632 ( .A(n_120), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_121), .B(n_404), .Y(n_533) );
INVx1_ASAP7_75t_L g585 ( .A(n_123), .Y(n_585) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_125), .Y(n_458) );
AOI22xp33_ASAP7_75t_SL g317 ( .A1(n_126), .A2(n_190), .B1(n_318), .B2(n_322), .Y(n_317) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_128), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_129), .B(n_296), .Y(n_295) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_134), .A2(n_175), .B1(n_343), .B2(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g475 ( .A(n_135), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_135), .A2(n_177), .B1(n_665), .B2(n_696), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_136), .A2(n_208), .B1(n_326), .B2(n_581), .Y(n_580) );
XNOR2x2_ASAP7_75t_L g435 ( .A(n_138), .B(n_436), .Y(n_435) );
AO221x2_ASAP7_75t_L g705 ( .A1(n_143), .A2(n_192), .B1(n_672), .B2(n_694), .C(n_706), .Y(n_705) );
OA22x2_ASAP7_75t_L g270 ( .A1(n_144), .A2(n_169), .B1(n_265), .B2(n_269), .Y(n_270) );
INVx1_ASAP7_75t_L g306 ( .A(n_144), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_147), .A2(n_232), .B1(n_346), .B2(n_380), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_148), .A2(n_188), .B1(n_326), .B2(n_330), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_149), .A2(n_193), .B1(n_411), .B2(n_426), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_150), .A2(n_162), .B1(n_469), .B2(n_470), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_152), .A2(n_201), .B1(n_617), .B2(n_618), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_153), .A2(n_156), .B1(n_498), .B2(n_499), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_154), .A2(n_216), .B1(n_665), .B2(n_686), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_157), .A2(n_189), .B1(n_369), .B2(n_563), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_158), .A2(n_207), .B1(n_501), .B2(n_502), .Y(n_518) );
XNOR2x2_ASAP7_75t_L g254 ( .A(n_161), .B(n_255), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_163), .A2(n_184), .B1(n_482), .B2(n_484), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_166), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g282 ( .A(n_168), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_168), .B(n_303), .Y(n_302) );
OAI21xp33_ASAP7_75t_L g316 ( .A1(n_169), .A2(n_180), .B(n_294), .Y(n_316) );
INVx1_ASAP7_75t_L g360 ( .A(n_172), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_174), .A2(n_206), .B1(n_492), .B2(n_493), .Y(n_491) );
AOI221xp5_ASAP7_75t_L g512 ( .A1(n_179), .A2(n_229), .B1(n_513), .B2(n_514), .C(n_515), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_180), .B(n_215), .Y(n_244) );
INVx1_ASAP7_75t_L g268 ( .A(n_180), .Y(n_268) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_183), .Y(n_464) );
AOI221xp5_ASAP7_75t_L g381 ( .A1(n_186), .A2(n_219), .B1(n_382), .B2(n_383), .C(n_384), .Y(n_381) );
INVx1_ASAP7_75t_L g284 ( .A(n_196), .Y(n_284) );
INVx1_ASAP7_75t_L g642 ( .A(n_197), .Y(n_642) );
INVx1_ASAP7_75t_L g489 ( .A(n_198), .Y(n_489) );
AOI21xp33_ASAP7_75t_L g486 ( .A1(n_200), .A2(n_487), .B(n_488), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g645 ( .A1(n_202), .A2(n_226), .B1(n_646), .B2(n_647), .Y(n_645) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_203), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_204), .A2(n_217), .B1(n_393), .B2(n_395), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_215), .B(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_218), .B(n_590), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g890 ( .A1(n_220), .A2(n_891), .B1(n_892), .B2(n_893), .Y(n_890) );
CKINVDCx5p33_ASAP7_75t_R g892 ( .A(n_220), .Y(n_892) );
AOI221xp5_ASAP7_75t_L g623 ( .A1(n_221), .A2(n_225), .B1(n_406), .B2(n_624), .C(n_627), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_222), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g674 ( .A(n_224), .Y(n_674) );
HB1xp67_ASAP7_75t_L g899 ( .A(n_224), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_227), .A2(n_228), .B1(n_326), .B2(n_330), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_231), .A2(n_233), .B1(n_330), .B2(n_378), .Y(n_377) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_246), .B(n_653), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
BUFx4_ASAP7_75t_SL g236 ( .A(n_237), .Y(n_236) );
NAND3xp33_ASAP7_75t_L g237 ( .A(n_238), .B(n_241), .C(n_245), .Y(n_237) );
AND2x2_ASAP7_75t_L g886 ( .A(n_238), .B(n_887), .Y(n_886) );
AND2x2_ASAP7_75t_L g895 ( .A(n_238), .B(n_888), .Y(n_895) );
AOI21xp5_ASAP7_75t_L g900 ( .A1(n_238), .A2(n_245), .B(n_702), .Y(n_900) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AO21x1_ASAP7_75t_L g897 ( .A1(n_239), .A2(n_898), .B(n_900), .Y(n_897) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g666 ( .A(n_240), .B(n_667), .Y(n_666) );
AND3x4_ASAP7_75t_L g701 ( .A(n_240), .B(n_673), .C(n_702), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g887 ( .A(n_241), .B(n_888), .Y(n_887) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AO21x2_ASAP7_75t_L g299 ( .A1(n_242), .A2(n_300), .B(n_301), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
INVx1_ASAP7_75t_L g888 ( .A(n_245), .Y(n_888) );
OAI22xp5_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_248), .B1(n_430), .B2(n_652), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OAI22x1_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_388), .B1(n_428), .B2(n_429), .Y(n_251) );
INVx1_ASAP7_75t_L g428 ( .A(n_252), .Y(n_428) );
OA22x2_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_254), .B1(n_354), .B2(n_387), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_324), .Y(n_255) );
NAND3xp33_ASAP7_75t_L g256 ( .A(n_257), .B(n_307), .C(n_317), .Y(n_256) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g383 ( .A(n_259), .Y(n_383) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g479 ( .A(n_260), .Y(n_479) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
BUFx3_ASAP7_75t_L g404 ( .A(n_261), .Y(n_404) );
INVx3_ASAP7_75t_L g467 ( .A(n_261), .Y(n_467) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_271), .Y(n_261) );
AND2x2_ASAP7_75t_L g323 ( .A(n_262), .B(n_321), .Y(n_323) );
AND2x2_ASAP7_75t_L g334 ( .A(n_262), .B(n_335), .Y(n_334) );
AND2x4_ASAP7_75t_L g339 ( .A(n_262), .B(n_340), .Y(n_339) );
AND2x4_ASAP7_75t_L g482 ( .A(n_262), .B(n_321), .Y(n_482) );
AND2x4_ASAP7_75t_L g495 ( .A(n_262), .B(n_335), .Y(n_495) );
AND2x4_ASAP7_75t_L g496 ( .A(n_262), .B(n_345), .Y(n_496) );
AND2x2_ASAP7_75t_L g521 ( .A(n_262), .B(n_335), .Y(n_521) );
AND2x2_ASAP7_75t_L g567 ( .A(n_262), .B(n_271), .Y(n_567) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_270), .Y(n_262) );
INVx1_ASAP7_75t_L g311 ( .A(n_263), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_267), .Y(n_263) );
NAND2xp33_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g269 ( .A(n_265), .Y(n_269) );
INVx3_ASAP7_75t_L g275 ( .A(n_265), .Y(n_275) );
NAND2xp33_ASAP7_75t_L g281 ( .A(n_265), .B(n_282), .Y(n_281) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_265), .Y(n_289) );
INVx1_ASAP7_75t_L g294 ( .A(n_265), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_266), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
OAI21xp5_ASAP7_75t_L g292 ( .A1(n_268), .A2(n_293), .B(n_294), .Y(n_292) );
AND2x2_ASAP7_75t_L g291 ( .A(n_270), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g310 ( .A(n_270), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g329 ( .A(n_270), .Y(n_329) );
AND2x4_ASAP7_75t_L g309 ( .A(n_271), .B(n_310), .Y(n_309) );
AND2x4_ASAP7_75t_L g314 ( .A(n_271), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g331 ( .A(n_271), .B(n_328), .Y(n_331) );
AND2x4_ASAP7_75t_L g485 ( .A(n_271), .B(n_315), .Y(n_485) );
AND2x2_ASAP7_75t_L g487 ( .A(n_271), .B(n_310), .Y(n_487) );
AND2x4_ASAP7_75t_L g499 ( .A(n_271), .B(n_328), .Y(n_499) );
AND2x4_ASAP7_75t_L g271 ( .A(n_272), .B(n_277), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g287 ( .A(n_273), .B(n_288), .Y(n_287) );
AND2x4_ASAP7_75t_L g321 ( .A(n_273), .B(n_277), .Y(n_321) );
AND2x4_ASAP7_75t_L g335 ( .A(n_273), .B(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g341 ( .A(n_273), .B(n_337), .Y(n_341) );
AND2x4_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_275), .B(n_280), .Y(n_279) );
INVxp67_ASAP7_75t_L g303 ( .A(n_275), .Y(n_303) );
NAND3xp33_ASAP7_75t_L g301 ( .A(n_276), .B(n_302), .C(n_304), .Y(n_301) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g337 ( .A(n_278), .Y(n_337) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
OAI21xp33_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_285), .B(n_295), .Y(n_283) );
INVx4_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x4_ASAP7_75t_L g286 ( .A(n_287), .B(n_291), .Y(n_286) );
AND2x4_ASAP7_75t_L g370 ( .A(n_287), .B(n_291), .Y(n_370) );
AND2x2_ASAP7_75t_L g484 ( .A(n_287), .B(n_291), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
INVx1_ASAP7_75t_L g300 ( .A(n_289), .Y(n_300) );
INVx2_ASAP7_75t_L g386 ( .A(n_296), .Y(n_386) );
INVx4_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g408 ( .A(n_297), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_297), .B(n_489), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_297), .B(n_516), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_297), .B(n_538), .Y(n_537) );
INVx4_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx3_ASAP7_75t_L g471 ( .A(n_298), .Y(n_471) );
INVx3_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_299), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_303), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g315 ( .A(n_304), .B(n_316), .Y(n_315) );
BUFx8_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
BUFx3_ASAP7_75t_L g382 ( .A(n_309), .Y(n_382) );
BUFx6f_ASAP7_75t_L g394 ( .A(n_309), .Y(n_394) );
BUFx6f_ASAP7_75t_L g621 ( .A(n_309), .Y(n_621) );
AND2x4_ASAP7_75t_L g320 ( .A(n_310), .B(n_321), .Y(n_320) );
AND2x4_ASAP7_75t_L g481 ( .A(n_310), .B(n_321), .Y(n_481) );
AND2x4_ASAP7_75t_L g328 ( .A(n_311), .B(n_329), .Y(n_328) );
INVx3_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g622 ( .A(n_313), .Y(n_622) );
INVx3_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_314), .Y(n_362) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_314), .Y(n_396) );
AND2x4_ASAP7_75t_L g347 ( .A(n_315), .B(n_345), .Y(n_347) );
AND2x4_ASAP7_75t_L g353 ( .A(n_315), .B(n_335), .Y(n_353) );
AND2x4_ASAP7_75t_L g493 ( .A(n_315), .B(n_345), .Y(n_493) );
AND2x4_ASAP7_75t_L g502 ( .A(n_315), .B(n_335), .Y(n_502) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g452 ( .A(n_319), .Y(n_452) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_320), .Y(n_367) );
BUFx3_ASAP7_75t_L g563 ( .A(n_320), .Y(n_563) );
BUFx3_ASAP7_75t_L g879 ( .A(n_320), .Y(n_879) );
AND2x4_ASAP7_75t_L g327 ( .A(n_321), .B(n_328), .Y(n_327) );
AND2x4_ASAP7_75t_L g498 ( .A(n_321), .B(n_328), .Y(n_498) );
INVx3_ASAP7_75t_L g359 ( .A(n_322), .Y(n_359) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g400 ( .A(n_323), .Y(n_400) );
BUFx3_ASAP7_75t_L g561 ( .A(n_323), .Y(n_561) );
NAND4xp25_ASAP7_75t_L g324 ( .A(n_325), .B(n_332), .C(n_342), .D(n_348), .Y(n_324) );
BUFx12f_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_327), .Y(n_378) );
INVx3_ASAP7_75t_L g421 ( .A(n_327), .Y(n_421) );
AND2x4_ASAP7_75t_L g344 ( .A(n_328), .B(n_345), .Y(n_344) );
AND2x4_ASAP7_75t_L g350 ( .A(n_328), .B(n_335), .Y(n_350) );
AND2x4_ASAP7_75t_L g492 ( .A(n_328), .B(n_340), .Y(n_492) );
AND2x4_ASAP7_75t_L g501 ( .A(n_328), .B(n_335), .Y(n_501) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g424 ( .A(n_331), .Y(n_424) );
BUFx5_ASAP7_75t_L g446 ( .A(n_331), .Y(n_446) );
BUFx3_ASAP7_75t_L g581 ( .A(n_331), .Y(n_581) );
BUFx3_ASAP7_75t_L g610 ( .A(n_333), .Y(n_610) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx8_ASAP7_75t_L g426 ( .A(n_334), .Y(n_426) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
BUFx12f_ASAP7_75t_L g380 ( .A(n_339), .Y(n_380) );
BUFx3_ASAP7_75t_L g411 ( .A(n_339), .Y(n_411) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_339), .Y(n_554) );
BUFx6f_ASAP7_75t_L g612 ( .A(n_339), .Y(n_612) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g345 ( .A(n_341), .Y(n_345) );
BUFx3_ASAP7_75t_L g438 ( .A(n_343), .Y(n_438) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_344), .Y(n_417) );
BUFx6f_ASAP7_75t_L g646 ( .A(n_344), .Y(n_646) );
BUFx3_ASAP7_75t_L g614 ( .A(n_346), .Y(n_614) );
BUFx12f_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx6_ASAP7_75t_L g413 ( .A(n_347), .Y(n_413) );
BUFx2_ASAP7_75t_SL g606 ( .A(n_349), .Y(n_606) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx12f_ASAP7_75t_L g373 ( .A(n_350), .Y(n_373) );
INVx4_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g375 ( .A(n_352), .Y(n_375) );
INVx4_ASAP7_75t_L g444 ( .A(n_352), .Y(n_444) );
INVx1_ASAP7_75t_L g870 ( .A(n_352), .Y(n_870) );
INVx8_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g387 ( .A(n_354), .Y(n_387) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND4xp75_ASAP7_75t_L g356 ( .A(n_357), .B(n_371), .C(n_376), .D(n_381), .Y(n_356) );
NOR2xp67_ASAP7_75t_L g357 ( .A(n_358), .B(n_364), .Y(n_357) );
OAI22xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_360), .B1(n_361), .B2(n_363), .Y(n_358) );
INVx3_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx3_ASAP7_75t_L g462 ( .A(n_362), .Y(n_462) );
OAI21xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_366), .B(n_368), .Y(n_364) );
INVx4_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx4f_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx5_ASAP7_75t_L g407 ( .A(n_370), .Y(n_407) );
BUFx2_ASAP7_75t_L g592 ( .A(n_370), .Y(n_592) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_373), .Y(n_415) );
BUFx12f_ASAP7_75t_L g443 ( .A(n_373), .Y(n_443) );
BUFx2_ASAP7_75t_SL g607 ( .A(n_375), .Y(n_607) );
AND2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_379), .Y(n_376) );
INVx2_ASAP7_75t_L g459 ( .A(n_382), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
INVx1_ASAP7_75t_L g429 ( .A(n_388), .Y(n_429) );
BUFx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
XOR2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_427), .Y(n_389) );
NOR2x1_ASAP7_75t_L g390 ( .A(n_391), .B(n_409), .Y(n_390) );
NAND4xp25_ASAP7_75t_L g391 ( .A(n_392), .B(n_397), .C(n_401), .D(n_405), .Y(n_391) );
BUFx3_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g873 ( .A(n_394), .Y(n_873) );
BUFx3_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g456 ( .A(n_400), .Y(n_456) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx3_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g469 ( .A(n_407), .Y(n_469) );
INVx2_ASAP7_75t_L g636 ( .A(n_407), .Y(n_636) );
NAND4xp25_ASAP7_75t_L g409 ( .A(n_410), .B(n_414), .C(n_418), .D(n_425), .Y(n_409) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx5_ASAP7_75t_L g440 ( .A(n_413), .Y(n_440) );
INVx2_ASAP7_75t_L g647 ( .A(n_413), .Y(n_647) );
BUFx3_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx4f_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g652 ( .A(n_430), .Y(n_652) );
XNOR2xp5_ASAP7_75t_L g430 ( .A(n_431), .B(n_546), .Y(n_430) );
AOI22xp33_ASAP7_75t_SL g431 ( .A1(n_432), .A2(n_433), .B1(n_505), .B2(n_506), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_435), .B1(n_472), .B2(n_503), .Y(n_433) );
INVx3_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NAND3xp33_ASAP7_75t_SL g436 ( .A(n_437), .B(n_441), .C(n_448), .Y(n_436) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AND3x1_ASAP7_75t_L g441 ( .A(n_442), .B(n_445), .C(n_447), .Y(n_441) );
BUFx3_ASAP7_75t_L g604 ( .A(n_446), .Y(n_604) );
NOR3xp33_ASAP7_75t_L g448 ( .A(n_449), .B(n_457), .C(n_463), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_451), .B1(n_453), .B2(n_454), .Y(n_449) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVxp67_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_459), .B1(n_460), .B2(n_461), .Y(n_457) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
OAI21xp33_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B(n_468), .Y(n_463) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx3_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g513 ( .A(n_467), .Y(n_513) );
INVx2_ASAP7_75t_L g590 ( .A(n_467), .Y(n_590) );
INVx2_ASAP7_75t_L g626 ( .A(n_467), .Y(n_626) );
INVx2_ASAP7_75t_L g638 ( .A(n_467), .Y(n_638) );
INVx4_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_471), .B(n_569), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_471), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx3_ASAP7_75t_L g504 ( .A(n_474), .Y(n_504) );
XNOR2x1_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
OR2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_490), .Y(n_476) );
NAND4xp25_ASAP7_75t_L g477 ( .A(n_478), .B(n_480), .C(n_483), .D(n_486), .Y(n_477) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_487), .Y(n_514) );
NAND4xp25_ASAP7_75t_L g490 ( .A(n_491), .B(n_494), .C(n_497), .D(n_500), .Y(n_490) );
INVx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B1(n_527), .B2(n_544), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NAND3x1_ASAP7_75t_L g511 ( .A(n_512), .B(n_517), .C(n_522), .Y(n_511) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
BUFx4f_ASAP7_75t_L g578 ( .A(n_521), .Y(n_578) );
AND4x1_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .C(n_525), .D(n_526), .Y(n_522) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_529), .Y(n_545) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
OR2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_539), .Y(n_531) );
NAND4xp25_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .C(n_535), .D(n_536), .Y(n_532) );
NAND4xp25_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .C(n_542), .D(n_543), .Y(n_539) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
XOR2xp5_ASAP7_75t_SL g546 ( .A(n_547), .B(n_599), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_571), .B1(n_593), .B2(n_595), .Y(n_547) );
CKINVDCx5p33_ASAP7_75t_R g548 ( .A(n_549), .Y(n_548) );
BUFx3_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g594 ( .A(n_550), .Y(n_594) );
XNOR2x1_ASAP7_75t_L g550 ( .A(n_551), .B(n_570), .Y(n_550) );
NAND4xp75_ASAP7_75t_L g551 ( .A(n_552), .B(n_556), .C(n_559), .D(n_564), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_555), .Y(n_552) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_562), .Y(n_559) );
BUFx2_ASAP7_75t_L g618 ( .A(n_561), .Y(n_618) );
BUFx2_ASAP7_75t_L g617 ( .A(n_563), .Y(n_617) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
HB1xp67_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g598 ( .A(n_573), .Y(n_598) );
NOR2x1_ASAP7_75t_L g574 ( .A(n_575), .B(n_582), .Y(n_574) );
NAND4xp25_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .C(n_579), .D(n_580), .Y(n_575) );
NAND4xp25_ASAP7_75t_SL g582 ( .A(n_583), .B(n_588), .C(n_589), .D(n_591), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g875 ( .A(n_586), .B(n_876), .Y(n_875) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
BUFx6f_ASAP7_75t_L g643 ( .A(n_587), .Y(n_643) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVxp67_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_629), .B1(n_630), .B2(n_651), .Y(n_599) );
INVx2_ASAP7_75t_SL g651 ( .A(n_600), .Y(n_651) );
NAND4xp75_ASAP7_75t_L g601 ( .A(n_602), .B(n_608), .C(n_615), .D(n_623), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_605), .Y(n_602) );
AND2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_613), .Y(n_608) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_619), .Y(n_615) );
BUFx3_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
XNOR2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
NOR2xp67_ASAP7_75t_L g633 ( .A(n_634), .B(n_644), .Y(n_633) );
NAND4xp25_ASAP7_75t_L g634 ( .A(n_635), .B(n_637), .C(n_639), .D(n_640), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
NAND4xp25_ASAP7_75t_SL g644 ( .A(n_645), .B(n_648), .C(n_649), .D(n_650), .Y(n_644) );
OAI221xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_860), .B1(n_862), .B2(n_884), .C(n_889), .Y(n_653) );
AND5x1_ASAP7_75t_L g654 ( .A(n_655), .B(n_797), .C(n_848), .D(n_853), .E(n_858), .Y(n_654) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_758), .B(n_764), .Y(n_655) );
NAND3xp33_ASAP7_75t_SL g656 ( .A(n_657), .B(n_718), .C(n_729), .Y(n_656) );
O2A1O1Ixp33_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_687), .B(n_691), .C(n_707), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_676), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_659), .B(n_851), .Y(n_850) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g722 ( .A(n_660), .Y(n_722) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g778 ( .A(n_661), .Y(n_778) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
OR2x2_ASAP7_75t_L g742 ( .A(n_662), .B(n_743), .Y(n_742) );
INVx2_ASAP7_75t_L g826 ( .A(n_662), .Y(n_826) );
INVx4_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_663), .B(n_688), .Y(n_687) );
OR2x2_ASAP7_75t_L g744 ( .A(n_663), .B(n_677), .Y(n_744) );
AND2x2_ASAP7_75t_L g754 ( .A(n_663), .B(n_743), .Y(n_754) );
OR2x2_ASAP7_75t_L g788 ( .A(n_663), .B(n_743), .Y(n_788) );
NOR2xp33_ASAP7_75t_L g837 ( .A(n_663), .B(n_767), .Y(n_837) );
AND2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_671), .Y(n_663) );
AND2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_668), .Y(n_665) );
AND2x4_ASAP7_75t_L g672 ( .A(n_666), .B(n_673), .Y(n_672) );
AND2x4_ASAP7_75t_L g679 ( .A(n_666), .B(n_668), .Y(n_679) );
AND2x2_ASAP7_75t_L g704 ( .A(n_666), .B(n_668), .Y(n_704) );
AND2x2_ASAP7_75t_L g669 ( .A(n_668), .B(n_670), .Y(n_669) );
AND2x4_ASAP7_75t_L g686 ( .A(n_668), .B(n_670), .Y(n_686) );
AND2x2_ASAP7_75t_L g696 ( .A(n_668), .B(n_670), .Y(n_696) );
AND2x4_ASAP7_75t_L g675 ( .A(n_670), .B(n_673), .Y(n_675) );
AND2x4_ASAP7_75t_L g694 ( .A(n_670), .B(n_673), .Y(n_694) );
INVx3_ASAP7_75t_L g762 ( .A(n_672), .Y(n_762) );
INVx2_ASAP7_75t_SL g684 ( .A(n_675), .Y(n_684) );
INVx1_ASAP7_75t_L g717 ( .A(n_676), .Y(n_717) );
AND2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_681), .Y(n_676) );
INVx2_ASAP7_75t_L g743 ( .A(n_677), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_680), .Y(n_677) );
BUFx2_ASAP7_75t_L g861 ( .A(n_679), .Y(n_861) );
INVx4_ASAP7_75t_L g756 ( .A(n_681), .Y(n_756) );
AND2x2_ASAP7_75t_L g768 ( .A(n_681), .B(n_741), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_681), .B(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g800 ( .A(n_681), .Y(n_800) );
AND2x2_ASAP7_75t_L g825 ( .A(n_681), .B(n_826), .Y(n_825) );
AND2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_685), .Y(n_681) );
INVx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g817 ( .A(n_687), .Y(n_817) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_688), .B(n_710), .Y(n_709) );
INVx3_ASAP7_75t_L g727 ( .A(n_688), .Y(n_727) );
INVx2_ASAP7_75t_L g740 ( .A(n_688), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_688), .B(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g767 ( .A(n_688), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_688), .B(n_756), .Y(n_796) );
AND2x2_ASAP7_75t_L g810 ( .A(n_688), .B(n_714), .Y(n_810) );
AND2x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
AND2x2_ASAP7_75t_L g845 ( .A(n_691), .B(n_740), .Y(n_845) );
AND2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_697), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_692), .B(n_705), .Y(n_710) );
CKINVDCx6p67_ASAP7_75t_R g714 ( .A(n_692), .Y(n_714) );
AND2x2_ASAP7_75t_L g732 ( .A(n_692), .B(n_726), .Y(n_732) );
AND2x2_ASAP7_75t_L g735 ( .A(n_692), .B(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_L g783 ( .A(n_692), .B(n_715), .Y(n_783) );
AND2x2_ASAP7_75t_L g784 ( .A(n_692), .B(n_699), .Y(n_784) );
NOR2xp33_ASAP7_75t_L g815 ( .A(n_692), .B(n_698), .Y(n_815) );
AND2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_695), .Y(n_692) );
INVx1_ASAP7_75t_L g752 ( .A(n_697), .Y(n_752) );
AND2x2_ASAP7_75t_L g802 ( .A(n_697), .B(n_714), .Y(n_802) );
AND2x2_ASAP7_75t_L g809 ( .A(n_697), .B(n_810), .Y(n_809) );
AND2x2_ASAP7_75t_L g697 ( .A(n_698), .B(n_705), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_698), .B(n_714), .Y(n_795) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AND2x2_ASAP7_75t_L g715 ( .A(n_699), .B(n_716), .Y(n_715) );
OR2x2_ASAP7_75t_L g728 ( .A(n_699), .B(n_705), .Y(n_728) );
AND2x2_ASAP7_75t_L g733 ( .A(n_699), .B(n_705), .Y(n_733) );
OAI22xp33_ASAP7_75t_L g745 ( .A1(n_699), .A2(n_746), .B1(n_749), .B2(n_753), .Y(n_745) );
AND2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_703), .Y(n_699) );
INVx1_ASAP7_75t_L g716 ( .A(n_705), .Y(n_716) );
AND2x2_ASAP7_75t_L g771 ( .A(n_705), .B(n_714), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_705), .B(n_732), .Y(n_829) );
AOI21xp5_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_711), .B(n_717), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
O2A1O1Ixp33_ASAP7_75t_L g791 ( .A1(n_709), .A2(n_783), .B(n_787), .C(n_792), .Y(n_791) );
OAI322xp33_ASAP7_75t_L g798 ( .A1(n_711), .A2(n_714), .A3(n_741), .B1(n_742), .B2(n_786), .C1(n_799), .C2(n_801), .Y(n_798) );
INVx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g757 ( .A(n_713), .B(n_738), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_714), .B(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g822 ( .A(n_714), .B(n_733), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_714), .B(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g751 ( .A(n_715), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_715), .B(n_726), .Y(n_832) );
OAI211xp5_ASAP7_75t_SL g811 ( .A1(n_716), .A2(n_812), .B(n_814), .C(n_827), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_719), .B(n_723), .Y(n_718) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g818 ( .A(n_720), .B(n_819), .Y(n_818) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g808 ( .A(n_722), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_723), .B(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g823 ( .A(n_725), .Y(n_823) );
O2A1O1Ixp33_ASAP7_75t_L g853 ( .A1(n_725), .A2(n_768), .B(n_854), .C(n_856), .Y(n_853) );
NOR2x1_ASAP7_75t_L g725 ( .A(n_726), .B(n_728), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_726), .B(n_747), .Y(n_746) );
AOI22xp5_ASAP7_75t_L g812 ( .A1(n_726), .A2(n_741), .B1(n_755), .B2(n_813), .Y(n_812) );
INVx3_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g844 ( .A(n_727), .B(n_733), .Y(n_844) );
INVx1_ASAP7_75t_L g736 ( .A(n_728), .Y(n_736) );
AOI211xp5_ASAP7_75t_SL g792 ( .A1(n_728), .A2(n_742), .B(n_793), .C(n_796), .Y(n_792) );
AOI221xp5_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_737), .B1(n_745), .B2(n_755), .C(n_757), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_731), .B(n_734), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
AND2x2_ASAP7_75t_L g851 ( .A(n_732), .B(n_736), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_733), .B(n_810), .Y(n_819) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g766 ( .A(n_735), .B(n_767), .Y(n_766) );
NAND3xp33_ASAP7_75t_L g836 ( .A(n_736), .B(n_774), .C(n_837), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_744), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g769 ( .A(n_740), .B(n_770), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_740), .B(n_783), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_740), .B(n_784), .Y(n_806) );
NOR2xp33_ASAP7_75t_L g813 ( .A(n_740), .B(n_744), .Y(n_813) );
NOR2xp33_ASAP7_75t_L g846 ( .A(n_740), .B(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g748 ( .A(n_743), .Y(n_748) );
INVxp67_ASAP7_75t_L g774 ( .A(n_743), .Y(n_774) );
AND2x2_ASAP7_75t_L g840 ( .A(n_743), .B(n_756), .Y(n_840) );
INVx1_ASAP7_75t_L g790 ( .A(n_744), .Y(n_790) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_744), .B(n_756), .Y(n_805) );
OAI22xp33_ASAP7_75t_L g856 ( .A1(n_744), .A2(n_806), .B1(n_834), .B2(n_857), .Y(n_856) );
OAI221xp5_ASAP7_75t_L g803 ( .A1(n_747), .A2(n_770), .B1(n_804), .B2(n_806), .C(n_807), .Y(n_803) );
INVx3_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_748), .B(n_756), .Y(n_834) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_751), .B(n_752), .Y(n_750) );
INVx1_ASAP7_75t_L g779 ( .A(n_754), .Y(n_779) );
NOR2xp33_ASAP7_75t_L g816 ( .A(n_755), .B(n_817), .Y(n_816) );
OAI21xp33_ASAP7_75t_L g848 ( .A1(n_755), .A2(n_849), .B(n_852), .Y(n_848) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
OR2x2_ASAP7_75t_L g773 ( .A(n_756), .B(n_774), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_756), .B(n_787), .Y(n_786) );
AND2x2_ASAP7_75t_L g830 ( .A(n_756), .B(n_826), .Y(n_830) );
INVx2_ASAP7_75t_L g780 ( .A(n_758), .Y(n_780) );
OAI21xp5_ASAP7_75t_L g838 ( .A1(n_758), .A2(n_839), .B(n_841), .Y(n_838) );
CKINVDCx5p33_ASAP7_75t_R g758 ( .A(n_759), .Y(n_758) );
OAI211xp5_ASAP7_75t_L g833 ( .A1(n_759), .A2(n_834), .B(n_835), .C(n_836), .Y(n_833) );
AND2x2_ASAP7_75t_L g759 ( .A(n_760), .B(n_763), .Y(n_759) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
NAND4xp25_ASAP7_75t_SL g764 ( .A(n_765), .B(n_775), .C(n_789), .D(n_791), .Y(n_764) );
OAI31xp33_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_768), .A3(n_769), .B(n_772), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g854 ( .A(n_767), .B(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
AOI22xp5_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_781), .B1(n_784), .B2(n_785), .Y(n_775) );
AOI21xp33_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_779), .B(n_780), .Y(n_776) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g847 ( .A(n_783), .Y(n_847) );
INVx1_ASAP7_75t_L g835 ( .A(n_784), .Y(n_835) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
AOI221xp5_ASAP7_75t_L g827 ( .A1(n_790), .A2(n_828), .B1(n_830), .B2(n_831), .C(n_833), .Y(n_827) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
OAI31xp33_ASAP7_75t_SL g797 ( .A1(n_798), .A2(n_803), .A3(n_811), .B(n_838), .Y(n_797) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
NOR2xp33_ASAP7_75t_L g859 ( .A(n_804), .B(n_821), .Y(n_859) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_808), .B(n_809), .Y(n_807) );
AOI211xp5_ASAP7_75t_L g814 ( .A1(n_815), .A2(n_816), .B(n_818), .C(n_820), .Y(n_814) );
INVx1_ASAP7_75t_L g855 ( .A(n_815), .Y(n_855) );
INVx1_ASAP7_75t_L g852 ( .A(n_819), .Y(n_852) );
AOI21xp33_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_823), .B(n_824), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
AOI211xp5_ASAP7_75t_L g841 ( .A1(n_826), .A2(n_842), .B(n_845), .C(n_846), .Y(n_841) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVxp33_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g857 ( .A(n_851), .Y(n_857) );
INVxp67_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
CKINVDCx5p33_ASAP7_75t_R g860 ( .A(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
HB1xp67_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
HB1xp67_ASAP7_75t_L g891 ( .A(n_866), .Y(n_891) );
NAND4xp75_ASAP7_75t_L g866 ( .A(n_867), .B(n_871), .C(n_877), .D(n_881), .Y(n_866) );
AND2x2_ASAP7_75t_L g867 ( .A(n_868), .B(n_869), .Y(n_867) );
OA21x2_ASAP7_75t_L g871 ( .A1(n_872), .A2(n_873), .B(n_874), .Y(n_871) );
AND2x2_ASAP7_75t_L g877 ( .A(n_878), .B(n_880), .Y(n_877) );
AND2x2_ASAP7_75t_L g881 ( .A(n_882), .B(n_883), .Y(n_881) );
INVx1_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
HB1xp67_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx1_ASAP7_75t_L g893 ( .A(n_891), .Y(n_893) );
BUFx3_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
BUFx3_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
CKINVDCx5p33_ASAP7_75t_R g898 ( .A(n_899), .Y(n_898) );
endmodule