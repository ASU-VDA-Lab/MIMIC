module fake_jpeg_2642_n_126 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_126);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_126;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_26),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_32),
.C(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_47),
.Y(n_53)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_48),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_44),
.Y(n_49)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_34),
.A2(n_28),
.B1(n_24),
.B2(n_23),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_50),
.A2(n_39),
.B1(n_41),
.B2(n_36),
.Y(n_56)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_49),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_61),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_49),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_41),
.B1(n_39),
.B2(n_42),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_57),
.A2(n_40),
.B1(n_35),
.B2(n_44),
.Y(n_67)
);

NAND3xp33_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_43),
.C(n_35),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_37),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_63),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_37),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_64),
.A2(n_73),
.B1(n_70),
.B2(n_68),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_38),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_66),
.Y(n_84)
);

NOR2x1_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_58),
.A2(n_0),
.B(n_1),
.Y(n_69)
);

FAx1_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_1),
.CI(n_2),
.CON(n_79),
.SN(n_79)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

NOR2xp67_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_46),
.Y(n_72)
);

NOR2xp67_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_22),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_64),
.A2(n_52),
.B1(n_60),
.B2(n_3),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_75),
.A2(n_85),
.B1(n_4),
.B2(n_5),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_71),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_77),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_52),
.Y(n_78)
);

XNOR2x1_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_70),
.Y(n_92)
);

NOR3xp33_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_81),
.C(n_83),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_60),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_74),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_89),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

AND2x6_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_73),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_98),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_84),
.A2(n_66),
.B(n_69),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_91),
.A2(n_94),
.B(n_84),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_96),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_85),
.A2(n_21),
.B1(n_20),
.B2(n_19),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_SL g102 ( 
.A1(n_93),
.A2(n_75),
.B(n_79),
.C(n_80),
.Y(n_102)
);

OAI22x1_ASAP7_75t_L g94 ( 
.A1(n_78),
.A2(n_18),
.B1(n_17),
.B2(n_5),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_97),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_3),
.C(n_4),
.Y(n_96)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_102),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_86),
.A2(n_79),
.B(n_7),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_105),
.Y(n_112)
);

NOR4xp25_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_6),
.C(n_7),
.D(n_8),
.Y(n_104)
);

BUFx24_ASAP7_75t_SL g113 ( 
.A(n_104),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_93),
.B(n_6),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_9),
.B(n_10),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_106),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_15),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_88),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_114),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_109),
.B(n_87),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_108),
.B1(n_105),
.B2(n_101),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_116),
.A2(n_102),
.B(n_113),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_100),
.C(n_111),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_119),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_102),
.C(n_12),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_120),
.B(n_117),
.C(n_12),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_121),
.Y(n_123)
);

OAI321xp33_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_11),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.C(n_121),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_13),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_125),
.Y(n_126)
);


endmodule