module fake_jpeg_26871_n_227 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_227);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_3),
.B(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_2),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_43),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_23),
.B(n_2),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_23),
.B(n_3),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_26),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_27),
.B(n_33),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_26),
.C(n_17),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_38),
.B(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_54),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_32),
.B1(n_29),
.B2(n_22),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_52),
.A2(n_19),
.B1(n_24),
.B2(n_18),
.Y(n_68)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_45),
.B(n_33),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_55),
.B(n_61),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_40),
.A2(n_25),
.B1(n_30),
.B2(n_23),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_57),
.A2(n_62),
.B1(n_44),
.B2(n_29),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_63),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_35),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_39),
.B(n_32),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_37),
.A2(n_25),
.B1(n_30),
.B2(n_23),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_35),
.B(n_22),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_64),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_99)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_70),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_19),
.B1(n_24),
.B2(n_18),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_67),
.A2(n_73),
.B1(n_77),
.B2(n_78),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_68),
.B(n_72),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_60),
.A2(n_44),
.B1(n_26),
.B2(n_17),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_54),
.A2(n_17),
.B1(n_36),
.B2(n_41),
.Y(n_73)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_53),
.A2(n_55),
.B1(n_47),
.B2(n_46),
.Y(n_77)
);

O2A1O1Ixp33_ASAP7_75t_SL g78 ( 
.A1(n_47),
.A2(n_46),
.B(n_50),
.C(n_57),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_35),
.B(n_36),
.C(n_41),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_79),
.A2(n_80),
.B1(n_6),
.B2(n_7),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_51),
.A2(n_20),
.B1(n_34),
.B2(n_28),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_34),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_53),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_85),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_86),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_60),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_6),
.Y(n_112)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_16),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_71),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_34),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_95),
.Y(n_115)
);

NAND2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_28),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_94),
.A2(n_65),
.B(n_78),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_28),
.Y(n_95)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_98),
.B(n_107),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_99),
.A2(n_109),
.B1(n_9),
.B2(n_10),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_4),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_106),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_5),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_6),
.Y(n_107)
);

NAND3xp33_ASAP7_75t_L g108 ( 
.A(n_66),
.B(n_15),
.C(n_14),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_111),
.Y(n_116)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_113),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_66),
.B(n_7),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_8),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_128),
.Y(n_139)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_119),
.B(n_121),
.Y(n_159)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_94),
.A2(n_84),
.B(n_68),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_124),
.A2(n_127),
.B(n_131),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_111),
.A2(n_72),
.B1(n_64),
.B2(n_70),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_125),
.A2(n_103),
.B1(n_109),
.B2(n_91),
.Y(n_145)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_130),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_SL g127 ( 
.A1(n_93),
.A2(n_85),
.B(n_87),
.C(n_86),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_74),
.C(n_89),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_107),
.Y(n_153)
);

INVxp33_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_101),
.A2(n_83),
.B(n_9),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_133),
.Y(n_146)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_137),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_92),
.B(n_76),
.Y(n_135)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_135),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_92),
.B(n_8),
.Y(n_136)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_118),
.A2(n_98),
.B1(n_93),
.B2(n_103),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_141),
.A2(n_147),
.B1(n_152),
.B2(n_158),
.Y(n_173)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_150),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_149),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_125),
.A2(n_106),
.B1(n_95),
.B2(n_96),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_113),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_122),
.A2(n_96),
.B1(n_104),
.B2(n_114),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_157),
.Y(n_170)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_155),
.Y(n_172)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_117),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_156),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_97),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_122),
.A2(n_105),
.B1(n_97),
.B2(n_11),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_146),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_161),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_151),
.A2(n_131),
.B(n_115),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_162),
.A2(n_163),
.B(n_165),
.Y(n_188)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_159),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_151),
.A2(n_127),
.B(n_141),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_158),
.Y(n_166)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_166),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_115),
.C(n_128),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_174),
.C(n_177),
.Y(n_178)
);

AO21x1_ASAP7_75t_L g171 ( 
.A1(n_140),
.A2(n_116),
.B(n_121),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_175),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_127),
.C(n_120),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_145),
.A2(n_119),
.B(n_127),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_155),
.Y(n_176)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_127),
.C(n_120),
.Y(n_177)
);

BUFx24_ASAP7_75t_SL g179 ( 
.A(n_164),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_189),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_153),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_182),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_170),
.B(n_147),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_152),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_184),
.C(n_163),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_164),
.B(n_148),
.C(n_143),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_137),
.Y(n_189)
);

OAI21xp33_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_133),
.B(n_138),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_190),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_144),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_162),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_187),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_196),
.Y(n_202)
);

OA21x2_ASAP7_75t_L g195 ( 
.A1(n_190),
.A2(n_172),
.B(n_166),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_182),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_180),
.B(n_160),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_198),
.C(n_199),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_169),
.C(n_175),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_173),
.C(n_172),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_183),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_205),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_195),
.A2(n_188),
.B(n_186),
.Y(n_204)
);

NOR3xp33_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_207),
.C(n_208),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_200),
.A2(n_176),
.B(n_185),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_195),
.A2(n_171),
.B(n_167),
.Y(n_207)
);

NAND4xp25_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_173),
.C(n_161),
.D(n_167),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_197),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_199),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_211),
.Y(n_218)
);

INVx11_ASAP7_75t_L g211 ( 
.A(n_202),
.Y(n_211)
);

NOR2x1_ASAP7_75t_SL g212 ( 
.A(n_209),
.B(n_198),
.Y(n_212)
);

AOI21x1_ASAP7_75t_L g219 ( 
.A1(n_212),
.A2(n_9),
.B(n_10),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_213),
.A2(n_194),
.B(n_138),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_214),
.A2(n_194),
.B(n_181),
.Y(n_216)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_216),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_217),
.Y(n_221)
);

AOI21x1_ASAP7_75t_L g222 ( 
.A1(n_219),
.A2(n_214),
.B(n_11),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_11),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_224),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_218),
.C(n_215),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_221),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_211),
.Y(n_227)
);


endmodule