module real_jpeg_23510_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_213;
wire n_167;
wire n_179;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx1_ASAP7_75t_L g132 ( 
.A(n_0),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_2),
.B(n_28),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_2),
.B(n_48),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_2),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_3),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_3),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_3),
.B(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_3),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_3),
.B(n_28),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_3),
.B(n_48),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_3),
.B(n_168),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_4),
.B(n_26),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_4),
.B(n_31),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_4),
.B(n_65),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_4),
.B(n_73),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_4),
.B(n_48),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_4),
.B(n_44),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_4),
.B(n_28),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_4),
.B(n_94),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx8_ASAP7_75t_SL g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_8),
.B(n_31),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_8),
.B(n_26),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_8),
.B(n_65),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_8),
.B(n_44),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_8),
.B(n_28),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_9),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_9),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_9),
.B(n_48),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_9),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_10),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_10),
.B(n_26),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_10),
.B(n_44),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_10),
.B(n_28),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_10),
.B(n_65),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_10),
.B(n_168),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_11),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_11),
.B(n_28),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_13),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_14),
.B(n_83),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_14),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_14),
.B(n_48),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_16),
.B(n_65),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_16),
.B(n_73),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_16),
.B(n_44),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_16),
.B(n_26),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_16),
.B(n_48),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_16),
.B(n_28),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_16),
.B(n_206),
.Y(n_205)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_17),
.Y(n_84)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_17),
.Y(n_109)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_17),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_146),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_111),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_77),
.C(n_99),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_21),
.A2(n_22),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_50),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_23),
.B(n_51),
.C(n_60),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_34),
.C(n_42),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_24),
.B(n_231),
.Y(n_230)
);

BUFx24_ASAP7_75t_SL g242 ( 
.A(n_24),
.Y(n_242)
);

FAx1_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_27),
.CI(n_30),
.CON(n_24),
.SN(n_24)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_25),
.B(n_27),
.C(n_30),
.Y(n_101)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_26),
.Y(n_120)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_28),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_32),
.B(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_34),
.A2(n_35),
.B1(n_42),
.B2(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_36),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_40),
.Y(n_131)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_42),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.C(n_47),
.Y(n_42)
);

FAx1_ASAP7_75t_SL g218 ( 
.A(n_43),
.B(n_46),
.CI(n_47),
.CON(n_218),
.SN(n_218)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx13_ASAP7_75t_L g202 ( 
.A(n_48),
.Y(n_202)
);

BUFx24_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_60),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_52),
.B(n_56),
.C(n_59),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_53),
.B(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_54),
.B(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_58),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_69),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_64),
.B2(n_68),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_62),
.B(n_68),
.C(n_69),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_64),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_75),
.C(n_76),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_71),
.B(n_202),
.Y(n_201)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_76),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_77),
.B(n_99),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_80),
.C(n_87),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_78),
.A2(n_80),
.B1(n_81),
.B2(n_235),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_78),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_85),
.B(n_86),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_85),
.Y(n_86)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_84),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_101),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_86),
.B(n_101),
.C(n_102),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_87),
.B(n_234),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_95),
.C(n_97),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_88),
.A2(n_89),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_92),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_90),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_95),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_102),
.Y(n_99)
);

CKINVDCx5p33_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_141),
.Y(n_140)
);

FAx1_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_107),
.CI(n_110),
.CON(n_103),
.SN(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_144),
.B2(n_145),
.Y(n_111)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_136),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_123),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_118),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_121),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_128),
.B2(n_135),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_126),
.Y(n_135)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_133),
.B2(n_134),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_236),
.C(n_237),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_224),
.C(n_225),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_212),
.C(n_213),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_174),
.C(n_185),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_164),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_159),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_152),
.B(n_159),
.C(n_164),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.C(n_157),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_153),
.A2(n_154),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_160),
.B(n_162),
.C(n_163),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_171),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_165),
.B(n_172),
.C(n_173),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_166),
.A2(n_167),
.B1(n_169),
.B2(n_170),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.C(n_184),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_178),
.A2(n_179),
.B1(n_184),
.B2(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_180),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_208),
.C(n_209),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_194),
.C(n_199),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_192),
.C(n_193),
.Y(n_208)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_197),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_195),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.C(n_203),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_219),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_220),
.C(n_223),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_218),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_217),
.C(n_218),
.Y(n_228)
);

BUFx24_ASAP7_75t_SL g240 ( 
.A(n_218),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_223),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_233),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_229),
.C(n_233),
.Y(n_236)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_238),
.Y(n_239)
);


endmodule