module real_jpeg_2881_n_7 (n_5, n_4, n_0, n_1, n_2, n_6, n_3, n_7);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_3;

output n_7;

wire n_17;
wire n_8;
wire n_57;
wire n_43;
wire n_37;
wire n_21;
wire n_54;
wire n_65;
wire n_38;
wire n_33;
wire n_50;
wire n_35;
wire n_29;
wire n_55;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_52;
wire n_58;
wire n_63;
wire n_12;
wire n_24;
wire n_66;
wire n_34;
wire n_28;
wire n_44;
wire n_60;
wire n_46;
wire n_62;
wire n_59;
wire n_64;
wire n_23;
wire n_11;
wire n_14;
wire n_47;
wire n_51;
wire n_45;
wire n_25;
wire n_61;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_39;
wire n_36;
wire n_40;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_56;
wire n_30;
wire n_48;
wire n_16;
wire n_15;
wire n_13;

INVx2_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_2),
.B(n_16),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_2),
.A2(n_12),
.B1(n_13),
.B2(n_25),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_2),
.B(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_2),
.A2(n_25),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_2),
.B(n_12),
.C(n_30),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_2),
.B(n_59),
.Y(n_58)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_4),
.A2(n_12),
.B1(n_13),
.B2(n_21),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_4),
.A2(n_21),
.B1(n_38),
.B2(n_39),
.Y(n_44)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_50),
.Y(n_7)
);

OAI21xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_33),
.B(n_49),
.Y(n_8)
);

AOI21xp5_ASAP7_75t_L g9 ( 
.A1(n_10),
.A2(n_26),
.B(n_32),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_17),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_15),
.Y(n_11)
);

AO22x1_ASAP7_75t_SL g29 ( 
.A1(n_12),
.A2(n_13),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_16),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_16),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_27)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

OA21x2_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B(n_22),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_24),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_28),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_27),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_30),
.A2(n_31),
.B1(n_38),
.B2(n_39),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_48),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_48),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_36),
.B1(n_45),
.B2(n_47),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_47),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_37),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_64)
);

AOI22x1_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_39),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_46),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_45),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_66),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_53),
.B(n_54),
.Y(n_66)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_57)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);


endmodule