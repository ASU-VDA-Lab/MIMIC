module fake_jpeg_25094_n_9 (n_3, n_2, n_1, n_0, n_4, n_9);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_9;

wire n_8;
wire n_6;
wire n_5;
wire n_7;

OAI22xp5_ASAP7_75t_L g5 ( 
.A1(n_3),
.A2(n_4),
.B1(n_2),
.B2(n_1),
.Y(n_5)
);

OAI32xp33_ASAP7_75t_L g6 ( 
.A1(n_2),
.A2(n_0),
.A3(n_1),
.B1(n_4),
.B2(n_3),
.Y(n_6)
);

NAND2xp5_ASAP7_75t_L g7 ( 
.A(n_0),
.B(n_1),
.Y(n_7)
);

AOI321xp33_ASAP7_75t_L g8 ( 
.A1(n_6),
.A2(n_0),
.A3(n_2),
.B1(n_5),
.B2(n_7),
.C(n_4),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_8),
.B(n_6),
.Y(n_9)
);


endmodule