module fake_ariane_2731_n_1995 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1995);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1995;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_727;
wire n_590;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_928;
wire n_253;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1904;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_784;
wire n_648;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_33),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_99),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_135),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_38),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_171),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_26),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_169),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_33),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_86),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_35),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_162),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_39),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_80),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_77),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_72),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_54),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_150),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_128),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_113),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_114),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_74),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_6),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_75),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_10),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_19),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_190),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_67),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_70),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_43),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_173),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_51),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_22),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_64),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_76),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_28),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_194),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_172),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_54),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_161),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_131),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_23),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_94),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_0),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_3),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_43),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_107),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_23),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_180),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_164),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_101),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_83),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_37),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_111),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_183),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_28),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_155),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_67),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_87),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_35),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_1),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_174),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_89),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_30),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_182),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_178),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_167),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_157),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_12),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_118),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_140),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_134),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_1),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_39),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_191),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_129),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_56),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_175),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_123),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_13),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_188),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_60),
.Y(n_276)
);

BUFx10_ASAP7_75t_L g277 ( 
.A(n_69),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_63),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_98),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_69),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_59),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_170),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_112),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_17),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_93),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_64),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_52),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_78),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_36),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_40),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_47),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_146),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_137),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_26),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_5),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_41),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_158),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_3),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_34),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_88),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_125),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_36),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_51),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_136),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_145),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_40),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_141),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_166),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_15),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_149),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_71),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_165),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_106),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_153),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_184),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_60),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_66),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_16),
.Y(n_318)
);

BUFx10_ASAP7_75t_L g319 ( 
.A(n_120),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_9),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_10),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_84),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_179),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_176),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_73),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_4),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_9),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_22),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_187),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_30),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_85),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_96),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_104),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_45),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_49),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_79),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_138),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_193),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_92),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_47),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_31),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_102),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_32),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_37),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_19),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_56),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_15),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_116),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_52),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_48),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_11),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_38),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_163),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_11),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_44),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_45),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_159),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_109),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_115),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_24),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_4),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_117),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_133),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_81),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_186),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_100),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_12),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_6),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_91),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_17),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_152),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_126),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_192),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_68),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_63),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_156),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_103),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_130),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_82),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_58),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_31),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_50),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_0),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_57),
.Y(n_384)
);

INVx2_ASAP7_75t_SL g385 ( 
.A(n_142),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_46),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_5),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_29),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_119),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_198),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_388),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_296),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_296),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_237),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_296),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_241),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_197),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_257),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_197),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_198),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_269),
.Y(n_401)
);

OR2x2_ASAP7_75t_L g402 ( 
.A(n_368),
.B(n_2),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_279),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_288),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_203),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_333),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_203),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_205),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_232),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_339),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_365),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_195),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_200),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_368),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_202),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_280),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_335),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_207),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_211),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_229),
.B(n_2),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_217),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_205),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_220),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_224),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_227),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_206),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_206),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_319),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_319),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_208),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_319),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_208),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_262),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_228),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_233),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_212),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_330),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_239),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_262),
.Y(n_439)
);

INVxp67_ASAP7_75t_SL g440 ( 
.A(n_302),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_240),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_272),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_242),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_212),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_214),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_250),
.Y(n_446)
);

BUFx2_ASAP7_75t_SL g447 ( 
.A(n_246),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_214),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_272),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_221),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_219),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_254),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_221),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_330),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_302),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_367),
.Y(n_456)
);

INVxp67_ASAP7_75t_SL g457 ( 
.A(n_367),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_310),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_219),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_225),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_225),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_255),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_267),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_268),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_271),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_231),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_231),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_235),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_277),
.B(n_7),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_310),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_235),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_312),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_312),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_243),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_277),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_274),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_277),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_243),
.Y(n_478)
);

INVxp33_ASAP7_75t_SL g479 ( 
.A(n_276),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_248),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_277),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_222),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g483 ( 
.A(n_330),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_248),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g485 ( 
.A(n_330),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_278),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_204),
.B(n_7),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_260),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_286),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_290),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_294),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_299),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_437),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_488),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_488),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_488),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_488),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_488),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_397),
.B(n_204),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_397),
.B(n_330),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_399),
.B(n_256),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_488),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_486),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_437),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_454),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_454),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_483),
.B(n_311),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_472),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_420),
.B(n_381),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_399),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_392),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_405),
.B(n_381),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_400),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_405),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_447),
.B(n_315),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_392),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_393),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_407),
.B(n_347),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_393),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_407),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_408),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_408),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_422),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_395),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_422),
.B(n_426),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_426),
.Y(n_526)
);

NAND2xp33_ASAP7_75t_L g527 ( 
.A(n_469),
.B(n_381),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_395),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_427),
.Y(n_529)
);

AND2x2_ASAP7_75t_SL g530 ( 
.A(n_487),
.B(n_218),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_427),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_430),
.B(n_432),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_430),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_472),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_432),
.B(n_347),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_436),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_436),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_444),
.Y(n_538)
);

AND2x6_ASAP7_75t_L g539 ( 
.A(n_487),
.B(n_210),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_444),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_445),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_445),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_448),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_448),
.B(n_450),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_450),
.Y(n_545)
);

INVxp67_ASAP7_75t_L g546 ( 
.A(n_489),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_453),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_453),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_460),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_394),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_460),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_461),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_461),
.B(n_256),
.Y(n_553)
);

AND2x2_ASAP7_75t_SL g554 ( 
.A(n_469),
.B(n_218),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_466),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_466),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_467),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_409),
.B(n_412),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_467),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_468),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_468),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_471),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_471),
.Y(n_563)
);

OA21x2_ASAP7_75t_L g564 ( 
.A1(n_474),
.A2(n_261),
.B(n_259),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_474),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_478),
.Y(n_566)
);

AND2x6_ASAP7_75t_L g567 ( 
.A(n_478),
.B(n_210),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_472),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_396),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_480),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_480),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_484),
.Y(n_572)
);

INVx1_ASAP7_75t_SL g573 ( 
.A(n_503),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_510),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_503),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_510),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_515),
.B(n_409),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_510),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_510),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_515),
.B(n_413),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_508),
.B(n_479),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_510),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_510),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_554),
.B(n_415),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_510),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_525),
.B(n_544),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_508),
.Y(n_587)
);

BUFx10_ASAP7_75t_L g588 ( 
.A(n_550),
.Y(n_588)
);

INVx1_ASAP7_75t_SL g589 ( 
.A(n_503),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_510),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_510),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_508),
.B(n_418),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_510),
.Y(n_593)
);

OAI21xp33_ASAP7_75t_SL g594 ( 
.A1(n_530),
.A2(n_402),
.B(n_484),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_531),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_531),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_554),
.B(n_421),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_550),
.Y(n_598)
);

AND2x6_ASAP7_75t_L g599 ( 
.A(n_525),
.B(n_259),
.Y(n_599)
);

INVx5_ASAP7_75t_L g600 ( 
.A(n_539),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_525),
.B(n_440),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_531),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_531),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_554),
.B(n_530),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_546),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_531),
.Y(n_606)
);

BUFx10_ASAP7_75t_L g607 ( 
.A(n_569),
.Y(n_607)
);

AND2x6_ASAP7_75t_L g608 ( 
.A(n_525),
.B(n_261),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_513),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_554),
.B(n_447),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_508),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_534),
.B(n_423),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_531),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_531),
.Y(n_614)
);

NAND2xp33_ASAP7_75t_L g615 ( 
.A(n_539),
.B(n_402),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_534),
.B(n_424),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_531),
.Y(n_617)
);

INVx4_ASAP7_75t_L g618 ( 
.A(n_539),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_544),
.B(n_457),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_531),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_531),
.Y(n_621)
);

AND2x4_ASAP7_75t_L g622 ( 
.A(n_544),
.B(n_451),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_554),
.B(n_485),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_543),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_544),
.B(n_455),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_530),
.A2(n_419),
.B1(n_390),
.B2(n_414),
.Y(n_626)
);

INVx4_ASAP7_75t_L g627 ( 
.A(n_539),
.Y(n_627)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_539),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_530),
.A2(n_419),
.B1(n_439),
.B2(n_433),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_543),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_530),
.B(n_425),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_543),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_543),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_543),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_513),
.B(n_398),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_534),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_543),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_543),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_543),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_499),
.B(n_456),
.Y(n_640)
);

BUFx10_ASAP7_75t_L g641 ( 
.A(n_569),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_543),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_543),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_563),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_563),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_499),
.B(n_459),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_563),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_563),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_539),
.A2(n_449),
.B1(n_458),
.B2(n_442),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_563),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_563),
.Y(n_651)
);

BUFx10_ASAP7_75t_L g652 ( 
.A(n_539),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_534),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_568),
.Y(n_654)
);

OAI22xp33_ASAP7_75t_SL g655 ( 
.A1(n_507),
.A2(n_482),
.B1(n_401),
.B2(n_404),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_568),
.B(n_434),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_563),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_499),
.B(n_435),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_546),
.B(n_438),
.Y(n_659)
);

INVxp33_ASAP7_75t_L g660 ( 
.A(n_558),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_563),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_539),
.A2(n_441),
.B1(n_446),
.B2(n_443),
.Y(n_662)
);

OAI22xp5_ASAP7_75t_L g663 ( 
.A1(n_558),
.A2(n_236),
.B1(n_309),
.B2(n_306),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_563),
.Y(n_664)
);

BUFx10_ASAP7_75t_L g665 ( 
.A(n_539),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_563),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_568),
.B(n_452),
.Y(n_667)
);

INVxp67_ASAP7_75t_L g668 ( 
.A(n_507),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_568),
.B(n_462),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_499),
.B(n_463),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_514),
.B(n_464),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_511),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_511),
.Y(n_673)
);

AND3x2_ASAP7_75t_L g674 ( 
.A(n_518),
.B(n_226),
.C(n_222),
.Y(n_674)
);

BUFx2_ASAP7_75t_L g675 ( 
.A(n_539),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_514),
.B(n_465),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_559),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_559),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_559),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_518),
.B(n_470),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_559),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_559),
.B(n_539),
.Y(n_682)
);

NOR2x1p5_ASAP7_75t_L g683 ( 
.A(n_532),
.B(n_391),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_532),
.B(n_476),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_532),
.B(n_491),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_559),
.B(n_473),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_514),
.B(n_428),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_520),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_520),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_520),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_528),
.Y(n_691)
);

AND2x6_ASAP7_75t_L g692 ( 
.A(n_500),
.B(n_266),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_521),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_528),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_521),
.B(n_490),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_521),
.B(n_522),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_511),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_539),
.A2(n_492),
.B1(n_230),
.B2(n_298),
.Y(n_698)
);

NAND3xp33_ASAP7_75t_SL g699 ( 
.A(n_501),
.B(n_406),
.C(n_403),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_516),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_522),
.Y(n_701)
);

INVx5_ASAP7_75t_L g702 ( 
.A(n_539),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_522),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_504),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_523),
.B(n_429),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_516),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_523),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_523),
.B(n_431),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_518),
.B(n_535),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_526),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_526),
.B(n_196),
.Y(n_711)
);

INVx5_ASAP7_75t_L g712 ( 
.A(n_567),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_526),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_529),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_518),
.B(n_226),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_529),
.B(n_313),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_527),
.A2(n_349),
.B1(n_317),
.B2(n_320),
.Y(n_717)
);

INVx5_ASAP7_75t_L g718 ( 
.A(n_567),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_529),
.B(n_321),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_533),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_533),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_528),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_533),
.Y(n_723)
);

OAI22xp5_ASAP7_75t_L g724 ( 
.A1(n_501),
.A2(n_345),
.B1(n_326),
.B2(n_327),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_693),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_672),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_587),
.Y(n_727)
);

NAND2xp33_ASAP7_75t_L g728 ( 
.A(n_599),
.B(n_567),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_693),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_672),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_575),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_618),
.B(n_538),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_668),
.B(n_538),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_673),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_671),
.B(n_538),
.Y(n_735)
);

INVxp67_ASAP7_75t_SL g736 ( 
.A(n_615),
.Y(n_736)
);

INVx8_ASAP7_75t_L g737 ( 
.A(n_599),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_L g738 ( 
.A1(n_604),
.A2(n_564),
.B1(n_567),
.B2(n_527),
.Y(n_738)
);

OAI22xp33_ASAP7_75t_L g739 ( 
.A1(n_698),
.A2(n_553),
.B1(n_501),
.B2(n_541),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_605),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_676),
.B(n_540),
.Y(n_741)
);

NAND2xp33_ASAP7_75t_L g742 ( 
.A(n_599),
.B(n_567),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_592),
.B(n_540),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_707),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_707),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_673),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_612),
.B(n_540),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_605),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_618),
.B(n_627),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_631),
.B(n_509),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_688),
.Y(n_751)
);

NOR3xp33_ASAP7_75t_L g752 ( 
.A(n_659),
.B(n_247),
.C(n_238),
.Y(n_752)
);

NAND2xp33_ASAP7_75t_L g753 ( 
.A(n_599),
.B(n_567),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_584),
.B(n_509),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_616),
.B(n_541),
.Y(n_755)
);

AND2x4_ASAP7_75t_L g756 ( 
.A(n_586),
.B(n_535),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_581),
.B(n_541),
.Y(n_757)
);

NOR2xp67_ASAP7_75t_L g758 ( 
.A(n_598),
.B(n_553),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_618),
.B(n_627),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_610),
.B(n_545),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_697),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_688),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_627),
.B(n_545),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_577),
.B(n_545),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_586),
.B(n_547),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_689),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_697),
.Y(n_767)
);

INVx2_ASAP7_75t_SL g768 ( 
.A(n_635),
.Y(n_768)
);

INVx4_ASAP7_75t_L g769 ( 
.A(n_600),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_597),
.B(n_547),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_586),
.B(n_547),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_689),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_628),
.B(n_549),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_690),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_700),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_711),
.B(n_549),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_652),
.Y(n_777)
);

OAI221xp5_ASAP7_75t_L g778 ( 
.A1(n_594),
.A2(n_284),
.B1(n_281),
.B2(n_287),
.C(n_289),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_700),
.Y(n_779)
);

NOR2x1p5_ASAP7_75t_L g780 ( 
.A(n_598),
.B(n_553),
.Y(n_780)
);

NAND2xp33_ASAP7_75t_L g781 ( 
.A(n_599),
.B(n_567),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_716),
.B(n_549),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_690),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_601),
.B(n_551),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_601),
.B(n_551),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_619),
.B(n_551),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_701),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_615),
.A2(n_556),
.B1(n_561),
.B2(n_552),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_686),
.B(n_552),
.Y(n_789)
);

NOR3xp33_ASAP7_75t_L g790 ( 
.A(n_687),
.B(n_247),
.C(n_238),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_619),
.B(n_552),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_599),
.A2(n_561),
.B1(n_562),
.B2(n_556),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_608),
.B(n_556),
.Y(n_793)
);

NOR2x1p5_ASAP7_75t_L g794 ( 
.A(n_635),
.B(n_528),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_608),
.B(n_561),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_706),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_580),
.B(n_562),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_588),
.Y(n_798)
);

NAND2xp33_ASAP7_75t_L g799 ( 
.A(n_608),
.B(n_567),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_608),
.A2(n_565),
.B1(n_566),
.B2(n_562),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_684),
.B(n_565),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_628),
.B(n_565),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_656),
.A2(n_669),
.B(n_667),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_703),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_703),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_710),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_628),
.B(n_566),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_608),
.B(n_566),
.Y(n_808)
);

INVx4_ASAP7_75t_L g809 ( 
.A(n_600),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_710),
.Y(n_810)
);

NAND2xp33_ASAP7_75t_L g811 ( 
.A(n_608),
.B(n_567),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_675),
.B(n_571),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_629),
.B(n_658),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_706),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_713),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_713),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_714),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_714),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_720),
.Y(n_819)
);

O2A1O1Ixp5_ASAP7_75t_L g820 ( 
.A1(n_719),
.A2(n_571),
.B(n_528),
.C(n_537),
.Y(n_820)
);

INVxp67_ASAP7_75t_L g821 ( 
.A(n_705),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_675),
.A2(n_564),
.B1(n_567),
.B2(n_537),
.Y(n_822)
);

AND2x4_ASAP7_75t_L g823 ( 
.A(n_709),
.B(n_535),
.Y(n_823)
);

INVxp33_ASAP7_75t_L g824 ( 
.A(n_708),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_721),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_658),
.B(n_571),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_670),
.A2(n_567),
.B1(n_535),
.B2(n_537),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_680),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_723),
.Y(n_829)
);

OR2x2_ASAP7_75t_L g830 ( 
.A(n_573),
.B(n_410),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_600),
.B(n_528),
.Y(n_831)
);

O2A1O1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_685),
.A2(n_537),
.B(n_542),
.C(n_536),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_678),
.Y(n_833)
);

INVxp67_ASAP7_75t_L g834 ( 
.A(n_589),
.Y(n_834)
);

AND2x4_ASAP7_75t_L g835 ( 
.A(n_709),
.B(n_500),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_600),
.B(n_536),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_670),
.B(n_536),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_622),
.B(n_542),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_622),
.B(n_542),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_678),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_660),
.B(n_662),
.Y(n_841)
);

AO22x2_ASAP7_75t_L g842 ( 
.A1(n_680),
.A2(n_316),
.B1(n_352),
.B2(n_252),
.Y(n_842)
);

AOI22xp5_ASAP7_75t_L g843 ( 
.A1(n_623),
.A2(n_567),
.B1(n_570),
.B2(n_572),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_679),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_679),
.Y(n_845)
);

NAND2xp33_ASAP7_75t_L g846 ( 
.A(n_682),
.B(n_638),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_600),
.B(n_542),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_702),
.B(n_548),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_622),
.B(n_548),
.Y(n_849)
);

INVx4_ASAP7_75t_L g850 ( 
.A(n_702),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_681),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_681),
.Y(n_852)
);

OR2x2_ASAP7_75t_L g853 ( 
.A(n_609),
.B(n_411),
.Y(n_853)
);

NAND3xp33_ASAP7_75t_L g854 ( 
.A(n_626),
.B(n_555),
.C(n_548),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_677),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_677),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_702),
.B(n_555),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_680),
.Y(n_858)
);

AND2x4_ASAP7_75t_SL g859 ( 
.A(n_588),
.B(n_475),
.Y(n_859)
);

BUFx4_ASAP7_75t_L g860 ( 
.A(n_575),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_691),
.Y(n_861)
);

BUFx3_ASAP7_75t_L g862 ( 
.A(n_587),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_691),
.B(n_555),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_691),
.B(n_694),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_694),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_640),
.B(n_416),
.Y(n_866)
);

HB1xp67_ASAP7_75t_L g867 ( 
.A(n_625),
.Y(n_867)
);

BUFx3_ASAP7_75t_L g868 ( 
.A(n_611),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_694),
.B(n_555),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_722),
.B(n_557),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_722),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_696),
.A2(n_722),
.B1(n_646),
.B2(n_649),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_695),
.B(n_557),
.Y(n_873)
);

NAND3xp33_ASAP7_75t_L g874 ( 
.A(n_663),
.B(n_560),
.C(n_557),
.Y(n_874)
);

INVxp67_ASAP7_75t_L g875 ( 
.A(n_646),
.Y(n_875)
);

NOR2xp67_ASAP7_75t_L g876 ( 
.A(n_699),
.B(n_557),
.Y(n_876)
);

NOR2xp67_ASAP7_75t_L g877 ( 
.A(n_717),
.B(n_560),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_574),
.Y(n_878)
);

O2A1O1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_724),
.A2(n_570),
.B(n_560),
.C(n_572),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_702),
.B(n_560),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_625),
.B(n_570),
.Y(n_881)
);

AOI221xp5_ASAP7_75t_L g882 ( 
.A1(n_640),
.A2(n_352),
.B1(n_252),
.B2(n_258),
.C(n_263),
.Y(n_882)
);

AND2x4_ASAP7_75t_L g883 ( 
.A(n_715),
.B(n_500),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_702),
.B(n_570),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_715),
.B(n_417),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_683),
.A2(n_572),
.B1(n_328),
.B2(n_334),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_611),
.B(n_572),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_636),
.B(n_516),
.Y(n_888)
);

BUFx3_ASAP7_75t_L g889 ( 
.A(n_636),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_692),
.B(n_653),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_653),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_SL g892 ( 
.A(n_834),
.B(n_588),
.Y(n_892)
);

INVx4_ASAP7_75t_L g893 ( 
.A(n_737),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_830),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_803),
.A2(n_582),
.B(n_579),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_764),
.B(n_692),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_821),
.B(n_607),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_881),
.B(n_692),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_881),
.B(n_692),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_758),
.B(n_607),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_735),
.B(n_692),
.Y(n_901)
);

BUFx8_ASAP7_75t_L g902 ( 
.A(n_731),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_727),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_727),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_740),
.B(n_607),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_SL g906 ( 
.A(n_859),
.B(n_641),
.Y(n_906)
);

INVx3_ASAP7_75t_L g907 ( 
.A(n_862),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_824),
.B(n_641),
.Y(n_908)
);

O2A1O1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_872),
.A2(n_519),
.B(n_524),
.C(n_517),
.Y(n_909)
);

O2A1O1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_875),
.A2(n_741),
.B(n_757),
.C(n_826),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_736),
.B(n_652),
.Y(n_911)
);

AOI22xp5_ASAP7_75t_L g912 ( 
.A1(n_841),
.A2(n_692),
.B1(n_641),
.B2(n_665),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_737),
.B(n_815),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_733),
.B(n_654),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_837),
.B(n_654),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_748),
.B(n_477),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_784),
.B(n_785),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_823),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_743),
.A2(n_755),
.B(n_747),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_846),
.A2(n_582),
.B(n_579),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_862),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_786),
.B(n_481),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_864),
.A2(n_595),
.B(n_593),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_841),
.B(n_652),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_751),
.Y(n_925)
);

INVx1_ASAP7_75t_SL g926 ( 
.A(n_860),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_732),
.A2(n_595),
.B(n_593),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_791),
.B(n_674),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_789),
.B(n_517),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_789),
.B(n_517),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_762),
.Y(n_931)
);

OAI21xp5_ASAP7_75t_L g932 ( 
.A1(n_770),
.A2(n_602),
.B(n_596),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_732),
.A2(n_602),
.B(n_596),
.Y(n_933)
);

NAND2xp33_ASAP7_75t_L g934 ( 
.A(n_737),
.B(n_638),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_828),
.B(n_655),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_763),
.A2(n_606),
.B(n_603),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_858),
.B(n_665),
.Y(n_937)
);

HB1xp67_ASAP7_75t_L g938 ( 
.A(n_823),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_SL g939 ( 
.A(n_859),
.B(n_665),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_756),
.B(n_517),
.Y(n_940)
);

INVxp67_ASAP7_75t_SL g941 ( 
.A(n_822),
.Y(n_941)
);

A2O1A1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_797),
.A2(n_576),
.B(n_578),
.C(n_574),
.Y(n_942)
);

INVx4_ASAP7_75t_L g943 ( 
.A(n_835),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_763),
.A2(n_606),
.B(n_603),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_773),
.A2(n_620),
.B(n_614),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_773),
.A2(n_620),
.B(n_614),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_802),
.A2(n_632),
.B(n_630),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_813),
.B(n_630),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_756),
.B(n_519),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_L g950 ( 
.A1(n_792),
.A2(n_800),
.B1(n_766),
.B2(n_774),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_802),
.A2(n_633),
.B(n_632),
.Y(n_951)
);

OAI21xp5_ASAP7_75t_L g952 ( 
.A1(n_770),
.A2(n_634),
.B(n_633),
.Y(n_952)
);

O2A1O1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_790),
.A2(n_524),
.B(n_519),
.C(n_263),
.Y(n_953)
);

AOI21xp33_ASAP7_75t_L g954 ( 
.A1(n_739),
.A2(n_754),
.B(n_750),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_883),
.B(n_519),
.Y(n_955)
);

OAI21xp33_ASAP7_75t_L g956 ( 
.A1(n_801),
.A2(n_341),
.B(n_340),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_807),
.A2(n_642),
.B(n_634),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_807),
.A2(n_644),
.B(n_642),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_868),
.Y(n_959)
);

BUFx4f_ASAP7_75t_L g960 ( 
.A(n_768),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_797),
.A2(n_576),
.B(n_583),
.C(n_578),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_883),
.B(n_524),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_867),
.B(n_650),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_L g964 ( 
.A1(n_794),
.A2(n_567),
.B1(n_664),
.B2(n_661),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_838),
.B(n_524),
.Y(n_965)
);

NOR2xp67_ASAP7_75t_L g966 ( 
.A(n_798),
.B(n_500),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_863),
.A2(n_664),
.B(n_661),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_839),
.B(n_500),
.Y(n_968)
);

OAI21xp5_ASAP7_75t_L g969 ( 
.A1(n_760),
.A2(n_585),
.B(n_583),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_772),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_849),
.B(n_500),
.Y(n_971)
);

INVx1_ASAP7_75t_SL g972 ( 
.A(n_853),
.Y(n_972)
);

NAND2x1p5_ASAP7_75t_L g973 ( 
.A(n_868),
.B(n_712),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_801),
.B(n_500),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_815),
.B(n_638),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_889),
.B(n_712),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_889),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_783),
.A2(n_617),
.B1(n_591),
.B2(n_585),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_869),
.A2(n_591),
.B(n_590),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_765),
.B(n_712),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_870),
.A2(n_613),
.B(n_590),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_873),
.B(n_512),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_771),
.B(n_712),
.Y(n_983)
);

INVx4_ASAP7_75t_L g984 ( 
.A(n_835),
.Y(n_984)
);

NOR3xp33_ASAP7_75t_L g985 ( 
.A(n_778),
.B(n_281),
.C(n_258),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_835),
.B(n_718),
.Y(n_986)
);

OR2x2_ASAP7_75t_L g987 ( 
.A(n_866),
.B(n_885),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_776),
.B(n_512),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_782),
.B(n_512),
.Y(n_989)
);

O2A1O1Ixp5_ASAP7_75t_L g990 ( 
.A1(n_820),
.A2(n_647),
.B(n_613),
.C(n_617),
.Y(n_990)
);

OR2x2_ASAP7_75t_L g991 ( 
.A(n_780),
.B(n_512),
.Y(n_991)
);

OAI21xp5_ASAP7_75t_L g992 ( 
.A1(n_843),
.A2(n_624),
.B(n_621),
.Y(n_992)
);

A2O1A1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_750),
.A2(n_637),
.B(n_621),
.C(n_624),
.Y(n_993)
);

AO21x1_ASAP7_75t_L g994 ( 
.A1(n_754),
.A2(n_292),
.B(n_266),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_819),
.B(n_512),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_793),
.Y(n_996)
);

O2A1O1Ixp33_ASAP7_75t_SL g997 ( 
.A1(n_795),
.A2(n_637),
.B(n_651),
.C(n_648),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_812),
.B(n_639),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_842),
.B(n_564),
.Y(n_999)
);

INVx4_ASAP7_75t_L g1000 ( 
.A(n_769),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_749),
.A2(n_643),
.B(n_639),
.Y(n_1001)
);

AO21x2_ASAP7_75t_L g1002 ( 
.A1(n_808),
.A2(n_647),
.B(n_643),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_725),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_812),
.Y(n_1004)
);

O2A1O1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_787),
.A2(n_805),
.B(n_806),
.C(n_804),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_840),
.A2(n_651),
.B(n_648),
.Y(n_1006)
);

INVx2_ASAP7_75t_SL g1007 ( 
.A(n_842),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_769),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_825),
.B(n_564),
.Y(n_1009)
);

O2A1O1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_810),
.A2(n_289),
.B(n_355),
.C(n_351),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_840),
.B(n_638),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_844),
.B(n_638),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_729),
.B(n_657),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_829),
.B(n_564),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_749),
.A2(n_657),
.B(n_645),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_759),
.A2(n_666),
.B(n_645),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_816),
.B(n_564),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_817),
.B(n_564),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_759),
.A2(n_666),
.B(n_645),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_878),
.A2(n_666),
.B(n_645),
.Y(n_1020)
);

OAI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_827),
.A2(n_316),
.B1(n_343),
.B2(n_344),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_818),
.B(n_645),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_744),
.B(n_666),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_878),
.A2(n_666),
.B(n_704),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_745),
.B(n_704),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_844),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_833),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_855),
.B(n_704),
.Y(n_1028)
);

OR2x6_ASAP7_75t_L g1029 ( 
.A(n_842),
.B(n_284),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_788),
.B(n_704),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_876),
.B(n_718),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_877),
.A2(n_359),
.B(n_357),
.C(n_362),
.Y(n_1032)
);

INVx1_ASAP7_75t_SL g1033 ( 
.A(n_886),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_890),
.B(n_718),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_856),
.B(n_704),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_845),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_851),
.A2(n_287),
.B(n_291),
.C(n_384),
.Y(n_1037)
);

AND2x4_ASAP7_75t_SL g1038 ( 
.A(n_752),
.B(n_291),
.Y(n_1038)
);

A2O1A1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_832),
.A2(n_852),
.B(n_861),
.C(n_856),
.Y(n_1039)
);

AOI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_728),
.A2(n_348),
.B1(n_246),
.B2(n_385),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_861),
.B(n_718),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_871),
.B(n_295),
.Y(n_1042)
);

AOI22xp33_ASAP7_75t_SL g1043 ( 
.A1(n_854),
.A2(n_343),
.B1(n_303),
.B2(n_355),
.Y(n_1043)
);

A2O1A1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_871),
.A2(n_362),
.B(n_292),
.C(n_376),
.Y(n_1044)
);

NAND3xp33_ASAP7_75t_L g1045 ( 
.A(n_882),
.B(n_350),
.C(n_346),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_887),
.B(n_865),
.Y(n_1046)
);

NOR2xp67_ASAP7_75t_L g1047 ( 
.A(n_874),
.B(n_505),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_887),
.B(n_295),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_726),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_726),
.B(n_303),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_809),
.B(n_718),
.Y(n_1051)
);

NOR3xp33_ASAP7_75t_L g1052 ( 
.A(n_879),
.B(n_344),
.C(n_318),
.Y(n_1052)
);

INVxp67_ASAP7_75t_SL g1053 ( 
.A(n_822),
.Y(n_1053)
);

BUFx8_ASAP7_75t_L g1054 ( 
.A(n_891),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_888),
.B(n_318),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_831),
.A2(n_888),
.B(n_753),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_742),
.A2(n_351),
.B(n_384),
.C(n_364),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_831),
.A2(n_496),
.B(n_495),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_730),
.B(n_734),
.Y(n_1059)
);

A2O1A1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_781),
.A2(n_338),
.B(n_364),
.C(n_304),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_730),
.B(n_354),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_734),
.B(n_356),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_746),
.B(n_360),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_746),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_761),
.B(n_361),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_799),
.A2(n_496),
.B(n_495),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_761),
.Y(n_1067)
);

BUFx3_ASAP7_75t_L g1068 ( 
.A(n_767),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_767),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_775),
.B(n_370),
.Y(n_1070)
);

INVxp67_ASAP7_75t_L g1071 ( 
.A(n_836),
.Y(n_1071)
);

AOI211xp5_ASAP7_75t_L g1072 ( 
.A1(n_811),
.A2(n_374),
.B(n_375),
.C(n_380),
.Y(n_1072)
);

NOR3xp33_ASAP7_75t_L g1073 ( 
.A(n_836),
.B(n_383),
.C(n_382),
.Y(n_1073)
);

NOR2x1_ASAP7_75t_L g1074 ( 
.A(n_847),
.B(n_304),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_775),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_779),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_779),
.Y(n_1077)
);

OR2x2_ASAP7_75t_L g1078 ( 
.A(n_987),
.B(n_796),
.Y(n_1078)
);

OAI22x1_ASAP7_75t_L g1079 ( 
.A1(n_1007),
.A2(n_386),
.B1(n_796),
.B2(n_814),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_960),
.B(n_777),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_904),
.Y(n_1081)
);

A2O1A1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_954),
.A2(n_738),
.B(n_777),
.C(n_814),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_917),
.B(n_738),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_919),
.B(n_809),
.Y(n_1084)
);

O2A1O1Ixp5_ASAP7_75t_L g1085 ( 
.A1(n_994),
.A2(n_880),
.B(n_857),
.C(n_847),
.Y(n_1085)
);

AND2x2_ASAP7_75t_SL g1086 ( 
.A(n_906),
.B(n_939),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_925),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_892),
.B(n_850),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_904),
.Y(n_1089)
);

OAI21xp33_ASAP7_75t_L g1090 ( 
.A1(n_956),
.A2(n_387),
.B(n_381),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_929),
.A2(n_930),
.B(n_901),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_R g1092 ( 
.A(n_902),
.B(n_850),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_910),
.A2(n_884),
.B(n_880),
.C(n_857),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_904),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_931),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_985),
.A2(n_884),
.B(n_848),
.C(n_308),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_970),
.Y(n_1097)
);

NAND2x1p5_ASAP7_75t_L g1098 ( 
.A(n_893),
.B(n_848),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_902),
.Y(n_1099)
);

NOR2xp67_ASAP7_75t_L g1100 ( 
.A(n_908),
.B(n_505),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_896),
.A2(n_952),
.B(n_932),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_897),
.B(n_493),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_926),
.Y(n_1103)
);

BUFx8_ASAP7_75t_L g1104 ( 
.A(n_916),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_895),
.A2(n_496),
.B(n_495),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1024),
.A2(n_385),
.B(n_502),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_897),
.B(n_922),
.Y(n_1107)
);

INVx2_ASAP7_75t_SL g1108 ( 
.A(n_1054),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_948),
.B(n_308),
.Y(n_1109)
);

INVx6_ASAP7_75t_L g1110 ( 
.A(n_1054),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_918),
.B(n_493),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_972),
.A2(n_336),
.B1(n_337),
.B2(n_338),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_943),
.B(n_199),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_918),
.B(n_493),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_938),
.B(n_506),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_985),
.A2(n_337),
.B(n_359),
.C(n_357),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_938),
.B(n_506),
.Y(n_1117)
);

OR2x6_ASAP7_75t_L g1118 ( 
.A(n_1029),
.B(n_336),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_SL g1119 ( 
.A1(n_908),
.A2(n_498),
.B(n_497),
.C(n_505),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1033),
.B(n_506),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_894),
.B(n_505),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_905),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_963),
.B(n_505),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_915),
.A2(n_496),
.B(n_502),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_904),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_984),
.B(n_201),
.Y(n_1126)
);

AND2x4_ASAP7_75t_L g1127 ( 
.A(n_984),
.B(n_505),
.Y(n_1127)
);

O2A1O1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_1010),
.A2(n_376),
.B(n_210),
.C(n_358),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_1029),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1027),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1036),
.Y(n_1131)
);

BUFx8_ASAP7_75t_L g1132 ( 
.A(n_999),
.Y(n_1132)
);

O2A1O1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_900),
.A2(n_1037),
.B(n_953),
.C(n_1021),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_959),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1026),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_893),
.B(n_504),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_928),
.B(n_209),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_SL g1138 ( 
.A1(n_1029),
.A2(n_381),
.B1(n_387),
.B2(n_389),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1056),
.A2(n_502),
.B(n_495),
.Y(n_1139)
);

O2A1O1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_1021),
.A2(n_297),
.B(n_358),
.C(n_497),
.Y(n_1140)
);

NOR3xp33_ASAP7_75t_L g1141 ( 
.A(n_1045),
.B(n_297),
.C(n_497),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_963),
.B(n_387),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_935),
.B(n_213),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_935),
.B(n_215),
.Y(n_1144)
);

OAI21xp33_ASAP7_75t_SL g1145 ( 
.A1(n_941),
.A2(n_8),
.B(n_13),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1020),
.A2(n_502),
.B(n_497),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_1003),
.Y(n_1147)
);

XOR2xp5_ASAP7_75t_L g1148 ( 
.A(n_912),
.B(n_216),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1050),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1042),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1057),
.A2(n_1005),
.B(n_948),
.C(n_1032),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_991),
.B(n_223),
.Y(n_1152)
);

OAI21xp33_ASAP7_75t_L g1153 ( 
.A1(n_1052),
.A2(n_949),
.B(n_940),
.Y(n_1153)
);

AOI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1004),
.A2(n_322),
.B1(n_234),
.B2(n_244),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1015),
.A2(n_497),
.B(n_498),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1004),
.B(n_387),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_959),
.B(n_245),
.Y(n_1157)
);

A2O1A1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_898),
.A2(n_498),
.B(n_497),
.C(n_387),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_903),
.B(n_249),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1046),
.A2(n_498),
.B(n_324),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_941),
.B(n_498),
.Y(n_1161)
);

AOI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_966),
.A2(n_323),
.B1(n_253),
.B2(n_264),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1070),
.B(n_8),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_974),
.B(n_14),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_1038),
.B(n_1071),
.Y(n_1165)
);

INVx3_ASAP7_75t_L g1166 ( 
.A(n_1000),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1017),
.A2(n_498),
.B(n_329),
.Y(n_1167)
);

O2A1O1Ixp5_ASAP7_75t_L g1168 ( 
.A1(n_975),
.A2(n_14),
.B(n_16),
.C(n_18),
.Y(n_1168)
);

INVxp67_ASAP7_75t_L g1169 ( 
.A(n_1061),
.Y(n_1169)
);

INVxp67_ASAP7_75t_L g1170 ( 
.A(n_1062),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1018),
.A2(n_325),
.B(n_265),
.Y(n_1171)
);

AND2x4_ASAP7_75t_L g1172 ( 
.A(n_903),
.B(n_504),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_955),
.B(n_18),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1001),
.A2(n_331),
.B(n_270),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_907),
.B(n_921),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_996),
.B(n_20),
.Y(n_1176)
);

O2A1O1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_950),
.A2(n_20),
.B(n_21),
.C(n_24),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_907),
.B(n_504),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1053),
.B(n_504),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1035),
.A2(n_332),
.B(n_273),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1069),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_914),
.A2(n_342),
.B(n_275),
.Y(n_1182)
);

AOI221xp5_ASAP7_75t_L g1183 ( 
.A1(n_1043),
.A2(n_314),
.B1(n_379),
.B2(n_282),
.C(n_377),
.Y(n_1183)
);

AOI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1073),
.A2(n_353),
.B1(n_283),
.B2(n_293),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_962),
.B(n_21),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_979),
.A2(n_363),
.B(n_300),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_981),
.A2(n_251),
.B(n_307),
.Y(n_1187)
);

OR2x2_ASAP7_75t_L g1188 ( 
.A(n_1063),
.B(n_504),
.Y(n_1188)
);

AOI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1073),
.A2(n_937),
.B1(n_899),
.B2(n_924),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1053),
.B(n_504),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_988),
.A2(n_369),
.B1(n_301),
.B2(n_373),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_989),
.A2(n_305),
.B1(n_371),
.B2(n_372),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_921),
.B(n_504),
.Y(n_1193)
);

INVx4_ASAP7_75t_L g1194 ( 
.A(n_977),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_998),
.A2(n_504),
.B(n_378),
.C(n_366),
.Y(n_1195)
);

AOI221xp5_ASAP7_75t_L g1196 ( 
.A1(n_1043),
.A2(n_504),
.B1(n_378),
.B2(n_366),
.C(n_285),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_996),
.B(n_25),
.Y(n_1197)
);

O2A1O1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1052),
.A2(n_25),
.B(n_27),
.C(n_29),
.Y(n_1198)
);

BUFx2_ASAP7_75t_L g1199 ( 
.A(n_977),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1048),
.B(n_1055),
.Y(n_1200)
);

NOR2x1_ASAP7_75t_L g1201 ( 
.A(n_1000),
.B(n_378),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1016),
.A2(n_494),
.B(n_378),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1019),
.A2(n_494),
.B(n_378),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_1068),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_920),
.A2(n_494),
.B(n_366),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1077),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_965),
.B(n_27),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_1008),
.Y(n_1208)
);

OR2x2_ASAP7_75t_L g1209 ( 
.A(n_1065),
.B(n_32),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1049),
.Y(n_1210)
);

OAI21xp33_ASAP7_75t_L g1211 ( 
.A1(n_995),
.A2(n_260),
.B(n_285),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_982),
.B(n_34),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1071),
.B(n_41),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_923),
.A2(n_494),
.B(n_366),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1030),
.A2(n_494),
.B(n_366),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_1074),
.Y(n_1216)
);

INVx1_ASAP7_75t_SL g1217 ( 
.A(n_1023),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1064),
.Y(n_1218)
);

INVx4_ASAP7_75t_L g1219 ( 
.A(n_1008),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_SL g1220 ( 
.A1(n_1028),
.A2(n_42),
.B(n_44),
.C(n_46),
.Y(n_1220)
);

BUFx2_ASAP7_75t_SL g1221 ( 
.A(n_1051),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_968),
.B(n_42),
.Y(n_1222)
);

O2A1O1Ixp5_ASAP7_75t_L g1223 ( 
.A1(n_975),
.A2(n_48),
.B(n_49),
.C(n_50),
.Y(n_1223)
);

O2A1O1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1039),
.A2(n_1044),
.B(n_942),
.C(n_961),
.Y(n_1224)
);

INVx4_ASAP7_75t_L g1225 ( 
.A(n_1008),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_967),
.A2(n_494),
.B(n_285),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_971),
.B(n_53),
.Y(n_1227)
);

BUFx4f_ASAP7_75t_L g1228 ( 
.A(n_1008),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1067),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1075),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_998),
.B(n_53),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1076),
.B(n_55),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_969),
.A2(n_494),
.B(n_285),
.Y(n_1233)
);

OAI22x1_ASAP7_75t_L g1234 ( 
.A1(n_1143),
.A2(n_1040),
.B1(n_913),
.B2(n_964),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1105),
.A2(n_990),
.B(n_909),
.Y(n_1235)
);

INVxp67_ASAP7_75t_L g1236 ( 
.A(n_1147),
.Y(n_1236)
);

AOI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1144),
.A2(n_937),
.B1(n_1072),
.B2(n_1013),
.Y(n_1237)
);

AO21x2_ASAP7_75t_L g1238 ( 
.A1(n_1233),
.A2(n_1002),
.B(n_1047),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1118),
.A2(n_1009),
.B1(n_1014),
.B2(n_1022),
.Y(n_1239)
);

OAI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1101),
.A2(n_993),
.B(n_990),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1202),
.A2(n_1006),
.B(n_992),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1129),
.B(n_55),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1118),
.A2(n_1060),
.B1(n_978),
.B2(n_1013),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1087),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1091),
.A2(n_934),
.B(n_997),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1203),
.A2(n_1066),
.B(n_951),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1084),
.A2(n_1011),
.B(n_1012),
.Y(n_1247)
);

INVx4_ASAP7_75t_L g1248 ( 
.A(n_1228),
.Y(n_1248)
);

AOI221x1_ASAP7_75t_L g1249 ( 
.A1(n_1090),
.A2(n_1028),
.B1(n_1025),
.B2(n_1058),
.C(n_927),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1104),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1095),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1084),
.A2(n_1012),
.B(n_1011),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1200),
.A2(n_958),
.B(n_957),
.Y(n_1253)
);

AO32x2_ASAP7_75t_L g1254 ( 
.A1(n_1138),
.A2(n_1002),
.A3(n_1059),
.B1(n_946),
.B2(n_947),
.Y(n_1254)
);

OR2x2_ASAP7_75t_L g1255 ( 
.A(n_1078),
.B(n_986),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1215),
.A2(n_933),
.B(n_945),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1083),
.A2(n_1109),
.B(n_1151),
.Y(n_1257)
);

NAND3xp33_ASAP7_75t_L g1258 ( 
.A(n_1177),
.B(n_983),
.C(n_980),
.Y(n_1258)
);

BUFx3_ASAP7_75t_L g1259 ( 
.A(n_1099),
.Y(n_1259)
);

AO31x2_ASAP7_75t_L g1260 ( 
.A1(n_1195),
.A2(n_936),
.A3(n_944),
.B(n_911),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1139),
.A2(n_1034),
.B(n_1031),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1107),
.B(n_1051),
.Y(n_1262)
);

AOI221x1_ASAP7_75t_L g1263 ( 
.A1(n_1079),
.A2(n_1231),
.B1(n_1109),
.B2(n_1116),
.C(n_1153),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1149),
.B(n_973),
.Y(n_1264)
);

BUFx2_ASAP7_75t_L g1265 ( 
.A(n_1104),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1165),
.B(n_973),
.Y(n_1266)
);

A2O1A1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1133),
.A2(n_976),
.B(n_1041),
.C(n_260),
.Y(n_1267)
);

O2A1O1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1198),
.A2(n_57),
.B(n_58),
.C(n_59),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1083),
.A2(n_260),
.B(n_494),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1097),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_SL g1271 ( 
.A(n_1228),
.B(n_260),
.Y(n_1271)
);

INVx4_ASAP7_75t_L g1272 ( 
.A(n_1110),
.Y(n_1272)
);

A2O1A1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1163),
.A2(n_61),
.B(n_62),
.C(n_65),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1224),
.A2(n_1226),
.B(n_1214),
.Y(n_1274)
);

AND2x4_ASAP7_75t_L g1275 ( 
.A(n_1118),
.B(n_127),
.Y(n_1275)
);

INVx1_ASAP7_75t_SL g1276 ( 
.A(n_1122),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1130),
.Y(n_1277)
);

INVxp67_ASAP7_75t_L g1278 ( 
.A(n_1121),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1110),
.Y(n_1279)
);

AO31x2_ASAP7_75t_L g1280 ( 
.A1(n_1082),
.A2(n_124),
.A3(n_181),
.B(n_177),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1131),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1205),
.A2(n_122),
.B(n_168),
.Y(n_1282)
);

AO31x2_ASAP7_75t_L g1283 ( 
.A1(n_1167),
.A2(n_121),
.A3(n_160),
.B(n_154),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1169),
.B(n_61),
.Y(n_1284)
);

O2A1O1Ixp33_ASAP7_75t_SL g1285 ( 
.A1(n_1164),
.A2(n_62),
.B(n_65),
.C(n_66),
.Y(n_1285)
);

O2A1O1Ixp33_ASAP7_75t_SL g1286 ( 
.A1(n_1212),
.A2(n_68),
.B(n_90),
.C(n_95),
.Y(n_1286)
);

INVx3_ASAP7_75t_SL g1287 ( 
.A(n_1103),
.Y(n_1287)
);

AO31x2_ASAP7_75t_L g1288 ( 
.A1(n_1179),
.A2(n_97),
.A3(n_105),
.B(n_108),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1135),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1158),
.A2(n_110),
.B(n_132),
.Y(n_1290)
);

CKINVDCx20_ASAP7_75t_R g1291 ( 
.A(n_1092),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1209),
.A2(n_139),
.B1(n_143),
.B2(n_144),
.Y(n_1292)
);

NAND2xp33_ASAP7_75t_L g1293 ( 
.A(n_1166),
.B(n_147),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1181),
.Y(n_1294)
);

A2O1A1Ixp33_ASAP7_75t_L g1295 ( 
.A1(n_1170),
.A2(n_1128),
.B(n_1189),
.C(n_1150),
.Y(n_1295)
);

NOR2xp67_ASAP7_75t_L g1296 ( 
.A(n_1204),
.B(n_148),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_SL g1297 ( 
.A1(n_1176),
.A2(n_151),
.B(n_185),
.Y(n_1297)
);

INVxp67_ASAP7_75t_L g1298 ( 
.A(n_1199),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_SL g1299 ( 
.A1(n_1093),
.A2(n_1190),
.B(n_1179),
.Y(n_1299)
);

NOR2x1_ASAP7_75t_SL g1300 ( 
.A(n_1221),
.B(n_1081),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_1108),
.Y(n_1301)
);

AOI221x1_ASAP7_75t_L g1302 ( 
.A1(n_1211),
.A2(n_1106),
.B1(n_1141),
.B2(n_1207),
.C(n_1197),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1206),
.Y(n_1303)
);

NOR2xp67_ASAP7_75t_L g1304 ( 
.A(n_1219),
.B(n_1225),
.Y(n_1304)
);

AO31x2_ASAP7_75t_L g1305 ( 
.A1(n_1190),
.A2(n_1161),
.A3(n_1160),
.B(n_1142),
.Y(n_1305)
);

AO31x2_ASAP7_75t_L g1306 ( 
.A1(n_1161),
.A2(n_1124),
.A3(n_1232),
.B(n_1229),
.Y(n_1306)
);

OR2x2_ASAP7_75t_L g1307 ( 
.A(n_1213),
.B(n_1112),
.Y(n_1307)
);

O2A1O1Ixp33_ASAP7_75t_SL g1308 ( 
.A1(n_1222),
.A2(n_1227),
.B(n_1207),
.C(n_1119),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1081),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1152),
.B(n_1086),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1123),
.A2(n_1102),
.B(n_1155),
.Y(n_1311)
);

AOI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1148),
.A2(n_1185),
.B1(n_1173),
.B2(n_1145),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1146),
.A2(n_1193),
.B(n_1171),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1210),
.Y(n_1314)
);

AND2x2_ASAP7_75t_SL g1315 ( 
.A(n_1081),
.B(n_1125),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1218),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1175),
.A2(n_1100),
.B(n_1217),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1137),
.B(n_1217),
.Y(n_1318)
);

AO31x2_ASAP7_75t_L g1319 ( 
.A1(n_1232),
.A2(n_1230),
.A3(n_1156),
.B(n_1096),
.Y(n_1319)
);

O2A1O1Ixp33_ASAP7_75t_SL g1320 ( 
.A1(n_1080),
.A2(n_1220),
.B(n_1126),
.C(n_1113),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1172),
.A2(n_1178),
.B(n_1180),
.Y(n_1321)
);

AO21x1_ASAP7_75t_L g1322 ( 
.A1(n_1191),
.A2(n_1192),
.B(n_1120),
.Y(n_1322)
);

AND2x4_ASAP7_75t_L g1323 ( 
.A(n_1127),
.B(n_1166),
.Y(n_1323)
);

OAI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1085),
.A2(n_1188),
.B(n_1168),
.Y(n_1324)
);

NOR2xp67_ASAP7_75t_SL g1325 ( 
.A(n_1208),
.B(n_1194),
.Y(n_1325)
);

CKINVDCx20_ASAP7_75t_R g1326 ( 
.A(n_1132),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1172),
.A2(n_1178),
.B(n_1194),
.Y(n_1327)
);

AND2x4_ASAP7_75t_L g1328 ( 
.A(n_1127),
.B(n_1225),
.Y(n_1328)
);

AOI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1191),
.A2(n_1192),
.B1(n_1184),
.B2(n_1183),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1159),
.A2(n_1182),
.B(n_1088),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1111),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_1089),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1114),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1115),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_SL g1335 ( 
.A(n_1132),
.B(n_1219),
.Y(n_1335)
);

AOI221xp5_ASAP7_75t_SL g1336 ( 
.A1(n_1140),
.A2(n_1186),
.B1(n_1187),
.B2(n_1196),
.C(n_1174),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1136),
.A2(n_1157),
.B(n_1201),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1216),
.A2(n_1154),
.B1(n_1117),
.B2(n_1162),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1136),
.A2(n_1098),
.B(n_1208),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1098),
.A2(n_1208),
.B(n_1223),
.Y(n_1340)
);

NAND3xp33_ASAP7_75t_L g1341 ( 
.A(n_1089),
.B(n_1094),
.C(n_1125),
.Y(n_1341)
);

AO31x2_ASAP7_75t_L g1342 ( 
.A1(n_1089),
.A2(n_1094),
.A3(n_1125),
.B(n_1134),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_1094),
.Y(n_1343)
);

OAI22x1_ASAP7_75t_L g1344 ( 
.A1(n_1134),
.A2(n_1143),
.B1(n_1144),
.B2(n_1129),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1134),
.A2(n_919),
.B(n_1091),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1105),
.A2(n_1203),
.B(n_1202),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1107),
.B(n_821),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1105),
.A2(n_1203),
.B(n_1202),
.Y(n_1348)
);

AOI221xp5_ASAP7_75t_SL g1349 ( 
.A1(n_1177),
.A2(n_1198),
.B1(n_778),
.B2(n_910),
.C(n_1145),
.Y(n_1349)
);

AO21x1_ASAP7_75t_L g1350 ( 
.A1(n_1109),
.A2(n_954),
.B(n_1231),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1091),
.A2(n_919),
.B(n_1084),
.Y(n_1351)
);

OAI22x1_ASAP7_75t_L g1352 ( 
.A1(n_1143),
.A2(n_1144),
.B1(n_1129),
.B2(n_598),
.Y(n_1352)
);

O2A1O1Ixp5_ASAP7_75t_L g1353 ( 
.A1(n_1231),
.A2(n_954),
.B(n_824),
.C(n_1143),
.Y(n_1353)
);

A2O1A1Ixp33_ASAP7_75t_L g1354 ( 
.A1(n_1143),
.A2(n_954),
.B(n_841),
.C(n_577),
.Y(n_1354)
);

BUFx3_ASAP7_75t_L g1355 ( 
.A(n_1099),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1105),
.A2(n_1203),
.B(n_1202),
.Y(n_1356)
);

AOI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1143),
.A2(n_985),
.B1(n_821),
.B2(n_790),
.Y(n_1357)
);

NOR2xp67_ASAP7_75t_L g1358 ( 
.A(n_1169),
.B(n_834),
.Y(n_1358)
);

A2O1A1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1143),
.A2(n_954),
.B(n_841),
.C(n_577),
.Y(n_1359)
);

AOI31xp67_ASAP7_75t_L g1360 ( 
.A1(n_1084),
.A2(n_1189),
.A3(n_1142),
.B(n_975),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_SL g1361 ( 
.A(n_1107),
.B(n_960),
.Y(n_1361)
);

AOI31xp67_ASAP7_75t_L g1362 ( 
.A1(n_1084),
.A2(n_1189),
.A3(n_1142),
.B(n_975),
.Y(n_1362)
);

AO21x1_ASAP7_75t_L g1363 ( 
.A1(n_1109),
.A2(n_954),
.B(n_1231),
.Y(n_1363)
);

CKINVDCx20_ASAP7_75t_R g1364 ( 
.A(n_1103),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1107),
.B(n_821),
.Y(n_1365)
);

A2O1A1Ixp33_ASAP7_75t_L g1366 ( 
.A1(n_1143),
.A2(n_954),
.B(n_841),
.C(n_577),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1091),
.A2(n_919),
.B(n_1084),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1105),
.A2(n_1203),
.B(n_1202),
.Y(n_1368)
);

AO31x2_ASAP7_75t_L g1369 ( 
.A1(n_1233),
.A2(n_994),
.A3(n_1215),
.B(n_1101),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_SL g1370 ( 
.A(n_1107),
.B(n_960),
.Y(n_1370)
);

AOI221xp5_ASAP7_75t_SL g1371 ( 
.A1(n_1177),
.A2(n_1198),
.B1(n_778),
.B2(n_910),
.C(n_1145),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_1107),
.B(n_824),
.Y(n_1372)
);

INVx3_ASAP7_75t_L g1373 ( 
.A(n_1228),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1087),
.Y(n_1374)
);

BUFx6f_ASAP7_75t_L g1375 ( 
.A(n_1228),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1107),
.B(n_821),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1087),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1087),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1105),
.A2(n_1203),
.B(n_1202),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1107),
.B(n_821),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1118),
.A2(n_1109),
.B1(n_917),
.B2(n_1029),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1107),
.B(n_821),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1107),
.B(n_821),
.Y(n_1383)
);

OA21x2_ASAP7_75t_L g1384 ( 
.A1(n_1233),
.A2(n_1215),
.B(n_1101),
.Y(n_1384)
);

BUFx10_ASAP7_75t_L g1385 ( 
.A(n_1110),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1107),
.B(n_824),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1087),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1105),
.A2(n_1203),
.B(n_1202),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1087),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1105),
.A2(n_1203),
.B(n_1202),
.Y(n_1390)
);

AOI31xp67_ASAP7_75t_L g1391 ( 
.A1(n_1084),
.A2(n_1189),
.A3(n_1142),
.B(n_975),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1105),
.A2(n_1203),
.B(n_1202),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_1107),
.B(n_824),
.Y(n_1393)
);

AOI221x1_ASAP7_75t_L g1394 ( 
.A1(n_1090),
.A2(n_954),
.B1(n_1079),
.B2(n_790),
.C(n_1231),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1091),
.A2(n_919),
.B(n_1084),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_SL g1396 ( 
.A1(n_1381),
.A2(n_1307),
.B1(n_1275),
.B2(n_1310),
.Y(n_1396)
);

OAI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1357),
.A2(n_1329),
.B1(n_1312),
.B2(n_1381),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1357),
.A2(n_1366),
.B1(n_1359),
.B2(n_1354),
.Y(n_1398)
);

CKINVDCx11_ASAP7_75t_R g1399 ( 
.A(n_1364),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1244),
.Y(n_1400)
);

INVx6_ASAP7_75t_L g1401 ( 
.A(n_1385),
.Y(n_1401)
);

CKINVDCx11_ASAP7_75t_R g1402 ( 
.A(n_1287),
.Y(n_1402)
);

OAI21xp33_ASAP7_75t_L g1403 ( 
.A1(n_1347),
.A2(n_1376),
.B(n_1365),
.Y(n_1403)
);

INVxp67_ASAP7_75t_SL g1404 ( 
.A(n_1351),
.Y(n_1404)
);

BUFx12f_ASAP7_75t_L g1405 ( 
.A(n_1385),
.Y(n_1405)
);

AOI22x1_ASAP7_75t_SL g1406 ( 
.A1(n_1326),
.A2(n_1301),
.B1(n_1291),
.B2(n_1272),
.Y(n_1406)
);

BUFx10_ASAP7_75t_L g1407 ( 
.A(n_1372),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1329),
.A2(n_1382),
.B1(n_1380),
.B2(n_1383),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1251),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1312),
.A2(n_1363),
.B1(n_1350),
.B2(n_1322),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1270),
.Y(n_1411)
);

INVx6_ASAP7_75t_L g1412 ( 
.A(n_1375),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1386),
.A2(n_1393),
.B1(n_1237),
.B2(n_1262),
.Y(n_1413)
);

BUFx12f_ASAP7_75t_L g1414 ( 
.A(n_1250),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1275),
.A2(n_1352),
.B1(n_1344),
.B2(n_1257),
.Y(n_1415)
);

INVx5_ASAP7_75t_L g1416 ( 
.A(n_1248),
.Y(n_1416)
);

NAND2x1p5_ASAP7_75t_L g1417 ( 
.A(n_1315),
.B(n_1248),
.Y(n_1417)
);

CKINVDCx11_ASAP7_75t_R g1418 ( 
.A(n_1265),
.Y(n_1418)
);

BUFx3_ASAP7_75t_L g1419 ( 
.A(n_1279),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1242),
.B(n_1278),
.Y(n_1420)
);

BUFx2_ASAP7_75t_L g1421 ( 
.A(n_1343),
.Y(n_1421)
);

CKINVDCx11_ASAP7_75t_R g1422 ( 
.A(n_1259),
.Y(n_1422)
);

INVx1_ASAP7_75t_SL g1423 ( 
.A(n_1276),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1277),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1318),
.B(n_1333),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_SL g1426 ( 
.A1(n_1243),
.A2(n_1292),
.B1(n_1239),
.B2(n_1293),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_SL g1427 ( 
.A1(n_1284),
.A2(n_1272),
.B1(n_1355),
.B2(n_1292),
.Y(n_1427)
);

BUFx8_ASAP7_75t_L g1428 ( 
.A(n_1281),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1237),
.A2(n_1316),
.B1(n_1314),
.B2(n_1234),
.Y(n_1429)
);

OAI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1243),
.A2(n_1331),
.B1(n_1334),
.B2(n_1263),
.Y(n_1430)
);

INVx3_ASAP7_75t_L g1431 ( 
.A(n_1373),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_SL g1432 ( 
.A1(n_1239),
.A2(n_1290),
.B1(n_1377),
.B2(n_1374),
.Y(n_1432)
);

INVx3_ASAP7_75t_L g1433 ( 
.A(n_1373),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1338),
.A2(n_1255),
.B1(n_1389),
.B2(n_1387),
.Y(n_1434)
);

BUFx12f_ASAP7_75t_L g1435 ( 
.A(n_1328),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1361),
.A2(n_1370),
.B1(n_1295),
.B2(n_1236),
.Y(n_1436)
);

AOI21xp5_ASAP7_75t_SL g1437 ( 
.A1(n_1267),
.A2(n_1300),
.B(n_1268),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1378),
.A2(n_1303),
.B1(n_1289),
.B2(n_1294),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1264),
.A2(n_1258),
.B1(n_1358),
.B2(n_1290),
.Y(n_1439)
);

INVx1_ASAP7_75t_SL g1440 ( 
.A(n_1332),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1258),
.A2(n_1266),
.B1(n_1296),
.B2(n_1317),
.Y(n_1441)
);

AOI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1349),
.A2(n_1371),
.B1(n_1335),
.B2(n_1323),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1309),
.Y(n_1443)
);

OAI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1335),
.A2(n_1394),
.B1(n_1298),
.B2(n_1302),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_SL g1445 ( 
.A1(n_1353),
.A2(n_1371),
.B1(n_1349),
.B2(n_1324),
.Y(n_1445)
);

BUFx4_ASAP7_75t_R g1446 ( 
.A(n_1325),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1324),
.A2(n_1297),
.B1(n_1238),
.B2(n_1321),
.Y(n_1447)
);

OAI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1327),
.A2(n_1339),
.B1(n_1274),
.B2(n_1311),
.Y(n_1448)
);

OAI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1367),
.A2(n_1395),
.B1(n_1285),
.B2(n_1340),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1342),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1341),
.Y(n_1451)
);

INVx2_ASAP7_75t_SL g1452 ( 
.A(n_1341),
.Y(n_1452)
);

BUFx2_ASAP7_75t_L g1453 ( 
.A(n_1319),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_SL g1454 ( 
.A1(n_1240),
.A2(n_1273),
.B1(n_1238),
.B2(n_1299),
.Y(n_1454)
);

BUFx6f_ASAP7_75t_L g1455 ( 
.A(n_1271),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1330),
.A2(n_1337),
.B1(n_1252),
.B2(n_1247),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_SL g1457 ( 
.A1(n_1240),
.A2(n_1241),
.B1(n_1245),
.B2(n_1282),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1253),
.A2(n_1269),
.B1(n_1345),
.B2(n_1384),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1384),
.A2(n_1313),
.B1(n_1304),
.B2(n_1261),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1288),
.B(n_1254),
.Y(n_1460)
);

INVx6_ASAP7_75t_L g1461 ( 
.A(n_1320),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1288),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1308),
.B(n_1288),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1336),
.A2(n_1286),
.B1(n_1256),
.B2(n_1235),
.Y(n_1464)
);

CKINVDCx20_ASAP7_75t_R g1465 ( 
.A(n_1360),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1362),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1391),
.Y(n_1467)
);

BUFx12f_ASAP7_75t_L g1468 ( 
.A(n_1280),
.Y(n_1468)
);

BUFx2_ASAP7_75t_L g1469 ( 
.A(n_1254),
.Y(n_1469)
);

OAI21xp5_ASAP7_75t_SL g1470 ( 
.A1(n_1249),
.A2(n_1280),
.B(n_1336),
.Y(n_1470)
);

BUFx12f_ASAP7_75t_L g1471 ( 
.A(n_1280),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1246),
.A2(n_1368),
.B1(n_1390),
.B2(n_1388),
.Y(n_1472)
);

INVx6_ASAP7_75t_L g1473 ( 
.A(n_1283),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1346),
.A2(n_1356),
.B1(n_1379),
.B2(n_1392),
.Y(n_1474)
);

CKINVDCx11_ASAP7_75t_R g1475 ( 
.A(n_1283),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1305),
.Y(n_1476)
);

NAND2x1p5_ASAP7_75t_L g1477 ( 
.A(n_1348),
.B(n_1260),
.Y(n_1477)
);

OAI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1305),
.A2(n_1357),
.B1(n_1029),
.B2(n_1118),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1260),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1369),
.Y(n_1480)
);

OAI21xp5_ASAP7_75t_SL g1481 ( 
.A1(n_1369),
.A2(n_1357),
.B(n_1329),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1244),
.Y(n_1482)
);

BUFx8_ASAP7_75t_L g1483 ( 
.A(n_1250),
.Y(n_1483)
);

AOI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1357),
.A2(n_1359),
.B1(n_1366),
.B2(n_1354),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_SL g1485 ( 
.A1(n_1381),
.A2(n_1029),
.B1(n_842),
.B2(n_813),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1244),
.Y(n_1486)
);

INVx1_ASAP7_75t_SL g1487 ( 
.A(n_1287),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1357),
.A2(n_1359),
.B1(n_1366),
.B2(n_1354),
.Y(n_1488)
);

INVxp67_ASAP7_75t_SL g1489 ( 
.A(n_1351),
.Y(n_1489)
);

BUFx2_ASAP7_75t_SL g1490 ( 
.A(n_1291),
.Y(n_1490)
);

BUFx3_ASAP7_75t_L g1491 ( 
.A(n_1385),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1381),
.A2(n_1029),
.B1(n_813),
.B2(n_842),
.Y(n_1492)
);

BUFx3_ASAP7_75t_L g1493 ( 
.A(n_1385),
.Y(n_1493)
);

BUFx8_ASAP7_75t_SL g1494 ( 
.A(n_1364),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1244),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1381),
.A2(n_1029),
.B1(n_813),
.B2(n_842),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1244),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1372),
.B(n_1386),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_SL g1499 ( 
.A1(n_1381),
.A2(n_1029),
.B1(n_842),
.B2(n_813),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1381),
.A2(n_1029),
.B1(n_813),
.B2(n_842),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_1364),
.Y(n_1501)
);

INVx6_ASAP7_75t_L g1502 ( 
.A(n_1385),
.Y(n_1502)
);

BUFx8_ASAP7_75t_L g1503 ( 
.A(n_1250),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1381),
.A2(n_1029),
.B1(n_813),
.B2(n_842),
.Y(n_1504)
);

OAI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1357),
.A2(n_1029),
.B1(n_1118),
.B2(n_1329),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1244),
.Y(n_1506)
);

INVx1_ASAP7_75t_SL g1507 ( 
.A(n_1287),
.Y(n_1507)
);

BUFx3_ASAP7_75t_L g1508 ( 
.A(n_1385),
.Y(n_1508)
);

AO22x1_ASAP7_75t_L g1509 ( 
.A1(n_1275),
.A2(n_598),
.B1(n_1144),
.B2(n_1143),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1381),
.A2(n_1029),
.B1(n_813),
.B2(n_842),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1244),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1248),
.Y(n_1512)
);

BUFx2_ASAP7_75t_L g1513 ( 
.A(n_1343),
.Y(n_1513)
);

BUFx6f_ASAP7_75t_SL g1514 ( 
.A(n_1385),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1372),
.B(n_1386),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1381),
.A2(n_1029),
.B1(n_813),
.B2(n_842),
.Y(n_1516)
);

OAI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1357),
.A2(n_1029),
.B1(n_1118),
.B2(n_1329),
.Y(n_1517)
);

INVx6_ASAP7_75t_L g1518 ( 
.A(n_1385),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_1364),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1244),
.Y(n_1520)
);

BUFx8_ASAP7_75t_L g1521 ( 
.A(n_1250),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1381),
.A2(n_1029),
.B1(n_813),
.B2(n_842),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1306),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1244),
.Y(n_1524)
);

BUFx2_ASAP7_75t_SL g1525 ( 
.A(n_1291),
.Y(n_1525)
);

AOI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1351),
.A2(n_1395),
.B(n_1367),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1244),
.Y(n_1527)
);

OAI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1357),
.A2(n_1029),
.B1(n_1118),
.B2(n_1329),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1244),
.Y(n_1529)
);

AOI21x1_ASAP7_75t_L g1530 ( 
.A1(n_1463),
.A2(n_1467),
.B(n_1466),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1400),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1443),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1485),
.A2(n_1499),
.B1(n_1505),
.B2(n_1517),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1409),
.Y(n_1534)
);

NAND2x1p5_ASAP7_75t_L g1535 ( 
.A(n_1451),
.B(n_1452),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1411),
.Y(n_1536)
);

AO21x1_ASAP7_75t_SL g1537 ( 
.A1(n_1484),
.A2(n_1410),
.B(n_1447),
.Y(n_1537)
);

INVx2_ASAP7_75t_SL g1538 ( 
.A(n_1424),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1482),
.Y(n_1539)
);

INVx3_ASAP7_75t_L g1540 ( 
.A(n_1477),
.Y(n_1540)
);

CKINVDCx11_ASAP7_75t_R g1541 ( 
.A(n_1399),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1469),
.B(n_1481),
.Y(n_1542)
);

INVx2_ASAP7_75t_SL g1543 ( 
.A(n_1486),
.Y(n_1543)
);

OR2x6_ASAP7_75t_L g1544 ( 
.A(n_1468),
.B(n_1471),
.Y(n_1544)
);

AO21x2_ASAP7_75t_L g1545 ( 
.A1(n_1470),
.A2(n_1462),
.B(n_1430),
.Y(n_1545)
);

AOI21x1_ASAP7_75t_L g1546 ( 
.A1(n_1526),
.A2(n_1509),
.B(n_1480),
.Y(n_1546)
);

OR2x6_ASAP7_75t_L g1547 ( 
.A(n_1453),
.B(n_1437),
.Y(n_1547)
);

OR2x6_ASAP7_75t_L g1548 ( 
.A(n_1450),
.B(n_1473),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1523),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1523),
.Y(n_1550)
);

INVx6_ASAP7_75t_L g1551 ( 
.A(n_1435),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1476),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1476),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1529),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1495),
.Y(n_1555)
);

OA21x2_ASAP7_75t_L g1556 ( 
.A1(n_1458),
.A2(n_1472),
.B(n_1474),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1497),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1506),
.Y(n_1558)
);

OAI21x1_ASAP7_75t_L g1559 ( 
.A1(n_1477),
.A2(n_1472),
.B(n_1458),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1408),
.B(n_1403),
.Y(n_1560)
);

INVx2_ASAP7_75t_SL g1561 ( 
.A(n_1511),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1520),
.Y(n_1562)
);

INVx1_ASAP7_75t_SL g1563 ( 
.A(n_1421),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1485),
.A2(n_1499),
.B1(n_1528),
.B2(n_1505),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1524),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1527),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1479),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1460),
.B(n_1438),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1404),
.Y(n_1569)
);

OAI21xp5_ASAP7_75t_L g1570 ( 
.A1(n_1398),
.A2(n_1488),
.B(n_1426),
.Y(n_1570)
);

INVxp67_ASAP7_75t_L g1571 ( 
.A(n_1498),
.Y(n_1571)
);

BUFx3_ASAP7_75t_L g1572 ( 
.A(n_1401),
.Y(n_1572)
);

INVx3_ASAP7_75t_L g1573 ( 
.A(n_1461),
.Y(n_1573)
);

AOI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1517),
.A2(n_1528),
.B1(n_1397),
.B2(n_1426),
.Y(n_1574)
);

BUFx3_ASAP7_75t_L g1575 ( 
.A(n_1401),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1438),
.Y(n_1576)
);

HB1xp67_ASAP7_75t_L g1577 ( 
.A(n_1423),
.Y(n_1577)
);

OAI21x1_ASAP7_75t_L g1578 ( 
.A1(n_1459),
.A2(n_1464),
.B(n_1456),
.Y(n_1578)
);

OA21x2_ASAP7_75t_L g1579 ( 
.A1(n_1464),
.A2(n_1404),
.B(n_1489),
.Y(n_1579)
);

BUFx8_ASAP7_75t_SL g1580 ( 
.A(n_1494),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1425),
.Y(n_1581)
);

AO21x1_ASAP7_75t_L g1582 ( 
.A1(n_1397),
.A2(n_1478),
.B(n_1430),
.Y(n_1582)
);

OAI21x1_ASAP7_75t_L g1583 ( 
.A1(n_1459),
.A2(n_1447),
.B(n_1489),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1478),
.Y(n_1584)
);

BUFx2_ASAP7_75t_L g1585 ( 
.A(n_1465),
.Y(n_1585)
);

BUFx12f_ASAP7_75t_L g1586 ( 
.A(n_1422),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1432),
.B(n_1410),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1434),
.Y(n_1588)
);

CKINVDCx6p67_ASAP7_75t_R g1589 ( 
.A(n_1514),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1434),
.Y(n_1590)
);

OAI21x1_ASAP7_75t_L g1591 ( 
.A1(n_1441),
.A2(n_1429),
.B(n_1439),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1420),
.Y(n_1592)
);

INVxp67_ASAP7_75t_R g1593 ( 
.A(n_1427),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1442),
.Y(n_1594)
);

BUFx3_ASAP7_75t_L g1595 ( 
.A(n_1502),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1448),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1448),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1449),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1449),
.Y(n_1599)
);

OAI21x1_ASAP7_75t_L g1600 ( 
.A1(n_1439),
.A2(n_1415),
.B(n_1436),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1454),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1454),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1445),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1413),
.B(n_1515),
.Y(n_1604)
);

AO31x2_ASAP7_75t_L g1605 ( 
.A1(n_1432),
.A2(n_1475),
.A3(n_1457),
.B(n_1445),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1444),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1396),
.B(n_1407),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1396),
.B(n_1415),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1444),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1431),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1433),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1455),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1440),
.Y(n_1613)
);

BUFx3_ASAP7_75t_L g1614 ( 
.A(n_1502),
.Y(n_1614)
);

BUFx3_ASAP7_75t_L g1615 ( 
.A(n_1518),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1407),
.B(n_1492),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1428),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1492),
.B(n_1504),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1455),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1428),
.Y(n_1620)
);

OAI21x1_ASAP7_75t_L g1621 ( 
.A1(n_1512),
.A2(n_1417),
.B(n_1510),
.Y(n_1621)
);

CKINVDCx14_ASAP7_75t_R g1622 ( 
.A(n_1418),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1496),
.B(n_1500),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1416),
.B(n_1513),
.Y(n_1624)
);

A2O1A1Ixp33_ASAP7_75t_SL g1625 ( 
.A1(n_1446),
.A2(n_1496),
.B(n_1522),
.C(n_1504),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1500),
.B(n_1510),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1516),
.Y(n_1627)
);

BUFx8_ASAP7_75t_L g1628 ( 
.A(n_1514),
.Y(n_1628)
);

INVx4_ASAP7_75t_L g1629 ( 
.A(n_1518),
.Y(n_1629)
);

BUFx3_ASAP7_75t_L g1630 ( 
.A(n_1491),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1516),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1522),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1487),
.B(n_1507),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1585),
.B(n_1592),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1570),
.B(n_1406),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1585),
.B(n_1490),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1557),
.B(n_1525),
.Y(n_1637)
);

AO32x2_ASAP7_75t_L g1638 ( 
.A1(n_1538),
.A2(n_1483),
.A3(n_1503),
.B1(n_1521),
.B2(n_1414),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1538),
.B(n_1419),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1543),
.B(n_1493),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1569),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1543),
.B(n_1508),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1532),
.B(n_1402),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1571),
.B(n_1519),
.Y(n_1644)
);

OAI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1560),
.A2(n_1600),
.B(n_1574),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1604),
.B(n_1483),
.Y(n_1646)
);

AOI221xp5_ASAP7_75t_L g1647 ( 
.A1(n_1606),
.A2(n_1501),
.B1(n_1503),
.B2(n_1521),
.C(n_1412),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1563),
.B(n_1405),
.Y(n_1648)
);

NOR2xp33_ASAP7_75t_L g1649 ( 
.A(n_1603),
.B(n_1573),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1561),
.B(n_1547),
.Y(n_1650)
);

O2A1O1Ixp33_ASAP7_75t_SL g1651 ( 
.A1(n_1593),
.A2(n_1625),
.B(n_1617),
.C(n_1620),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1577),
.B(n_1587),
.Y(n_1652)
);

AND2x2_ASAP7_75t_SL g1653 ( 
.A(n_1608),
.B(n_1542),
.Y(n_1653)
);

OAI21xp5_ASAP7_75t_L g1654 ( 
.A1(n_1591),
.A2(n_1602),
.B(n_1601),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_1580),
.Y(n_1655)
);

A2O1A1Ixp33_ASAP7_75t_L g1656 ( 
.A1(n_1533),
.A2(n_1564),
.B(n_1608),
.C(n_1591),
.Y(n_1656)
);

OAI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1601),
.A2(n_1602),
.B(n_1609),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1554),
.Y(n_1658)
);

A2O1A1Ixp33_ASAP7_75t_L g1659 ( 
.A1(n_1606),
.A2(n_1609),
.B(n_1542),
.C(n_1607),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1568),
.B(n_1535),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1573),
.B(n_1629),
.Y(n_1661)
);

AND2x4_ASAP7_75t_L g1662 ( 
.A(n_1547),
.B(n_1544),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1554),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1555),
.Y(n_1664)
);

INVx3_ASAP7_75t_L g1665 ( 
.A(n_1624),
.Y(n_1665)
);

AOI221xp5_ASAP7_75t_L g1666 ( 
.A1(n_1582),
.A2(n_1594),
.B1(n_1576),
.B2(n_1616),
.C(n_1590),
.Y(n_1666)
);

NAND4xp25_ASAP7_75t_L g1667 ( 
.A(n_1633),
.B(n_1610),
.C(n_1611),
.D(n_1569),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1566),
.B(n_1555),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1535),
.B(n_1613),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_1580),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1558),
.B(n_1562),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1558),
.B(n_1562),
.Y(n_1672)
);

OA21x2_ASAP7_75t_L g1673 ( 
.A1(n_1583),
.A2(n_1578),
.B(n_1559),
.Y(n_1673)
);

OAI211xp5_ASAP7_75t_L g1674 ( 
.A1(n_1596),
.A2(n_1597),
.B(n_1599),
.C(n_1598),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1535),
.B(n_1531),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_SL g1676 ( 
.A1(n_1626),
.A2(n_1618),
.B1(n_1623),
.B2(n_1616),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1534),
.B(n_1536),
.Y(n_1677)
);

OA21x2_ASAP7_75t_L g1678 ( 
.A1(n_1578),
.A2(n_1559),
.B(n_1596),
.Y(n_1678)
);

INVxp67_ASAP7_75t_L g1679 ( 
.A(n_1619),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1549),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1539),
.B(n_1630),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1565),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1565),
.B(n_1581),
.Y(n_1683)
);

A2O1A1Ixp33_ASAP7_75t_L g1684 ( 
.A1(n_1623),
.A2(n_1626),
.B(n_1584),
.C(n_1582),
.Y(n_1684)
);

INVx1_ASAP7_75t_SL g1685 ( 
.A(n_1541),
.Y(n_1685)
);

OR2x6_ASAP7_75t_L g1686 ( 
.A(n_1621),
.B(n_1548),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_1541),
.Y(n_1687)
);

AO21x2_ASAP7_75t_L g1688 ( 
.A1(n_1530),
.A2(n_1545),
.B(n_1546),
.Y(n_1688)
);

A2O1A1Ixp33_ASAP7_75t_L g1689 ( 
.A1(n_1605),
.A2(n_1597),
.B(n_1537),
.C(n_1588),
.Y(n_1689)
);

OA21x2_ASAP7_75t_L g1690 ( 
.A1(n_1598),
.A2(n_1599),
.B(n_1553),
.Y(n_1690)
);

AND2x4_ASAP7_75t_L g1691 ( 
.A(n_1624),
.B(n_1612),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1572),
.B(n_1575),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1572),
.B(n_1575),
.Y(n_1693)
);

A2O1A1Ixp33_ASAP7_75t_L g1694 ( 
.A1(n_1605),
.A2(n_1627),
.B(n_1631),
.C(n_1632),
.Y(n_1694)
);

AND2x4_ASAP7_75t_L g1695 ( 
.A(n_1612),
.B(n_1540),
.Y(n_1695)
);

OA21x2_ASAP7_75t_L g1696 ( 
.A1(n_1552),
.A2(n_1553),
.B(n_1549),
.Y(n_1696)
);

INVx3_ASAP7_75t_L g1697 ( 
.A(n_1665),
.Y(n_1697)
);

BUFx3_ASAP7_75t_L g1698 ( 
.A(n_1691),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1680),
.Y(n_1699)
);

AOI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1666),
.A2(n_1545),
.B1(n_1551),
.B2(n_1621),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1641),
.B(n_1550),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1650),
.B(n_1605),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1652),
.B(n_1550),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1641),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1658),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1650),
.B(n_1605),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1696),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1660),
.B(n_1683),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1663),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1664),
.Y(n_1710)
);

NOR2x1p5_ASAP7_75t_L g1711 ( 
.A(n_1667),
.B(n_1586),
.Y(n_1711)
);

INVx2_ASAP7_75t_SL g1712 ( 
.A(n_1691),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1668),
.B(n_1552),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1682),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1677),
.B(n_1545),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1671),
.Y(n_1716)
);

INVxp67_ASAP7_75t_SL g1717 ( 
.A(n_1690),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1672),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1634),
.B(n_1579),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1678),
.B(n_1556),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1679),
.Y(n_1721)
);

HB1xp67_ASAP7_75t_L g1722 ( 
.A(n_1678),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1678),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1675),
.B(n_1556),
.Y(n_1724)
);

INVx2_ASAP7_75t_SL g1725 ( 
.A(n_1691),
.Y(n_1725)
);

INVxp67_ASAP7_75t_L g1726 ( 
.A(n_1669),
.Y(n_1726)
);

HB1xp67_ASAP7_75t_L g1727 ( 
.A(n_1688),
.Y(n_1727)
);

BUFx2_ASAP7_75t_L g1728 ( 
.A(n_1695),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1673),
.B(n_1556),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1659),
.B(n_1567),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1673),
.B(n_1540),
.Y(n_1731)
);

BUFx2_ASAP7_75t_L g1732 ( 
.A(n_1695),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1689),
.B(n_1653),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1688),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1704),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1704),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1719),
.B(n_1673),
.Y(n_1737)
);

HB1xp67_ASAP7_75t_L g1738 ( 
.A(n_1721),
.Y(n_1738)
);

INVxp67_ASAP7_75t_SL g1739 ( 
.A(n_1707),
.Y(n_1739)
);

OAI221xp5_ASAP7_75t_L g1740 ( 
.A1(n_1700),
.A2(n_1684),
.B1(n_1645),
.B2(n_1656),
.C(n_1635),
.Y(n_1740)
);

OAI21xp5_ASAP7_75t_SL g1741 ( 
.A1(n_1700),
.A2(n_1635),
.B(n_1684),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1707),
.Y(n_1742)
);

OAI31xp33_ASAP7_75t_L g1743 ( 
.A1(n_1733),
.A2(n_1656),
.A3(n_1689),
.B(n_1694),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1699),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1719),
.B(n_1681),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_SL g1746 ( 
.A(n_1715),
.B(n_1687),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1701),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1701),
.Y(n_1748)
);

INVxp67_ASAP7_75t_L g1749 ( 
.A(n_1721),
.Y(n_1749)
);

INVx4_ASAP7_75t_L g1750 ( 
.A(n_1697),
.Y(n_1750)
);

INVx5_ASAP7_75t_L g1751 ( 
.A(n_1729),
.Y(n_1751)
);

NOR3xp33_ASAP7_75t_L g1752 ( 
.A(n_1733),
.B(n_1651),
.C(n_1674),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1703),
.B(n_1637),
.Y(n_1753)
);

BUFx2_ASAP7_75t_L g1754 ( 
.A(n_1698),
.Y(n_1754)
);

OAI33xp33_ASAP7_75t_L g1755 ( 
.A1(n_1730),
.A2(n_1639),
.A3(n_1642),
.B1(n_1640),
.B2(n_1646),
.B3(n_1692),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1716),
.B(n_1694),
.Y(n_1756)
);

BUFx2_ASAP7_75t_L g1757 ( 
.A(n_1698),
.Y(n_1757)
);

AOI33xp33_ASAP7_75t_L g1758 ( 
.A1(n_1716),
.A2(n_1676),
.A3(n_1651),
.B1(n_1685),
.B2(n_1636),
.B3(n_1643),
.Y(n_1758)
);

A2O1A1Ixp33_ASAP7_75t_SL g1759 ( 
.A1(n_1697),
.A2(n_1622),
.B(n_1661),
.C(n_1693),
.Y(n_1759)
);

NAND2xp33_ASAP7_75t_SL g1760 ( 
.A(n_1711),
.B(n_1655),
.Y(n_1760)
);

AO21x2_ASAP7_75t_L g1761 ( 
.A1(n_1717),
.A2(n_1734),
.B(n_1727),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1718),
.B(n_1649),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1718),
.B(n_1715),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1705),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1705),
.Y(n_1765)
);

AND2x4_ASAP7_75t_L g1766 ( 
.A(n_1731),
.B(n_1686),
.Y(n_1766)
);

NOR3xp33_ASAP7_75t_L g1767 ( 
.A(n_1717),
.B(n_1647),
.C(n_1654),
.Y(n_1767)
);

BUFx2_ASAP7_75t_L g1768 ( 
.A(n_1728),
.Y(n_1768)
);

HB1xp67_ASAP7_75t_L g1769 ( 
.A(n_1722),
.Y(n_1769)
);

NOR2xp33_ASAP7_75t_L g1770 ( 
.A(n_1708),
.B(n_1586),
.Y(n_1770)
);

INVx2_ASAP7_75t_SL g1771 ( 
.A(n_1751),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1761),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1751),
.B(n_1732),
.Y(n_1773)
);

BUFx3_ASAP7_75t_L g1774 ( 
.A(n_1770),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1747),
.B(n_1709),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1747),
.B(n_1709),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1748),
.B(n_1710),
.Y(n_1777)
);

NAND2x1p5_ASAP7_75t_L g1778 ( 
.A(n_1751),
.B(n_1662),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1764),
.Y(n_1779)
);

NAND2x1_ASAP7_75t_L g1780 ( 
.A(n_1768),
.B(n_1732),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1748),
.B(n_1710),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1764),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1751),
.B(n_1712),
.Y(n_1783)
);

AND2x4_ASAP7_75t_L g1784 ( 
.A(n_1751),
.B(n_1750),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1768),
.B(n_1725),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1749),
.B(n_1714),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1765),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1749),
.B(n_1714),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1745),
.B(n_1725),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_SL g1790 ( 
.A(n_1752),
.B(n_1724),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1761),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1735),
.B(n_1713),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1745),
.B(n_1726),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1745),
.B(n_1726),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1763),
.B(n_1713),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1735),
.B(n_1722),
.Y(n_1796)
);

HB1xp67_ASAP7_75t_L g1797 ( 
.A(n_1761),
.Y(n_1797)
);

AND2x4_ASAP7_75t_L g1798 ( 
.A(n_1750),
.B(n_1702),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1765),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1736),
.B(n_1723),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1761),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1736),
.Y(n_1802)
);

INVxp67_ASAP7_75t_L g1803 ( 
.A(n_1738),
.Y(n_1803)
);

HB1xp67_ASAP7_75t_L g1804 ( 
.A(n_1744),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1762),
.B(n_1703),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1772),
.Y(n_1806)
);

OAI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1790),
.A2(n_1741),
.B(n_1752),
.Y(n_1807)
);

AOI21xp33_ASAP7_75t_SL g1808 ( 
.A1(n_1778),
.A2(n_1670),
.B(n_1655),
.Y(n_1808)
);

AOI32xp33_ASAP7_75t_L g1809 ( 
.A1(n_1774),
.A2(n_1740),
.A3(n_1767),
.B1(n_1741),
.B2(n_1737),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1772),
.Y(n_1810)
);

OAI22xp33_ASAP7_75t_L g1811 ( 
.A1(n_1805),
.A2(n_1740),
.B1(n_1756),
.B2(n_1730),
.Y(n_1811)
);

INVxp67_ASAP7_75t_L g1812 ( 
.A(n_1774),
.Y(n_1812)
);

INVxp33_ASAP7_75t_L g1813 ( 
.A(n_1774),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1805),
.B(n_1767),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1779),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1793),
.B(n_1754),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1793),
.B(n_1794),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1779),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1795),
.B(n_1762),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1803),
.B(n_1758),
.Y(n_1820)
);

NOR2x1_ASAP7_75t_L g1821 ( 
.A(n_1780),
.B(n_1784),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1772),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1803),
.B(n_1756),
.Y(n_1823)
);

BUFx3_ASAP7_75t_L g1824 ( 
.A(n_1780),
.Y(n_1824)
);

HB1xp67_ASAP7_75t_L g1825 ( 
.A(n_1786),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1782),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1793),
.B(n_1794),
.Y(n_1827)
);

BUFx6f_ASAP7_75t_L g1828 ( 
.A(n_1801),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1782),
.Y(n_1829)
);

AND2x4_ASAP7_75t_SL g1830 ( 
.A(n_1798),
.B(n_1784),
.Y(n_1830)
);

INVxp67_ASAP7_75t_SL g1831 ( 
.A(n_1804),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1787),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1795),
.B(n_1737),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1795),
.B(n_1737),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1794),
.B(n_1754),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1789),
.B(n_1757),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1787),
.Y(n_1837)
);

NOR2x1p5_ASAP7_75t_L g1838 ( 
.A(n_1784),
.B(n_1589),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1792),
.B(n_1753),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1801),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1789),
.B(n_1757),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1799),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1799),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1801),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1792),
.B(n_1753),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1791),
.Y(n_1846)
);

AOI22xp5_ASAP7_75t_L g1847 ( 
.A1(n_1791),
.A2(n_1755),
.B1(n_1711),
.B2(n_1657),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1786),
.B(n_1788),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1802),
.Y(n_1849)
);

AND2x4_ASAP7_75t_L g1850 ( 
.A(n_1798),
.B(n_1766),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1828),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1815),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_SL g1853 ( 
.A(n_1809),
.B(n_1784),
.Y(n_1853)
);

INVx2_ASAP7_75t_SL g1854 ( 
.A(n_1830),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1817),
.B(n_1798),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1809),
.B(n_1814),
.Y(n_1856)
);

NOR2xp33_ASAP7_75t_L g1857 ( 
.A(n_1813),
.B(n_1670),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1817),
.B(n_1798),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1811),
.B(n_1804),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1827),
.B(n_1798),
.Y(n_1860)
);

INVxp67_ASAP7_75t_L g1861 ( 
.A(n_1820),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1819),
.B(n_1788),
.Y(n_1862)
);

OR2x2_ASAP7_75t_L g1863 ( 
.A(n_1819),
.B(n_1775),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1815),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1827),
.B(n_1773),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1812),
.B(n_1755),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1816),
.B(n_1773),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1807),
.B(n_1775),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1818),
.Y(n_1869)
);

OR2x2_ASAP7_75t_L g1870 ( 
.A(n_1839),
.B(n_1776),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1845),
.B(n_1776),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1823),
.B(n_1777),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1825),
.B(n_1777),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1816),
.B(n_1773),
.Y(n_1874)
);

NAND2xp33_ASAP7_75t_SL g1875 ( 
.A(n_1838),
.B(n_1771),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1818),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1826),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1847),
.B(n_1781),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1828),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1826),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1829),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1848),
.B(n_1781),
.Y(n_1882)
);

OR2x2_ASAP7_75t_L g1883 ( 
.A(n_1833),
.B(n_1796),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1829),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1835),
.B(n_1783),
.Y(n_1885)
);

NOR2xp33_ASAP7_75t_L g1886 ( 
.A(n_1808),
.B(n_1589),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1847),
.B(n_1785),
.Y(n_1887)
);

NAND4xp25_ASAP7_75t_L g1888 ( 
.A(n_1824),
.B(n_1759),
.C(n_1760),
.D(n_1785),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1854),
.B(n_1835),
.Y(n_1889)
);

AOI22xp5_ASAP7_75t_L g1890 ( 
.A1(n_1866),
.A2(n_1729),
.B1(n_1720),
.B2(n_1706),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1856),
.B(n_1831),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1880),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1868),
.B(n_1836),
.Y(n_1893)
);

AOI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1853),
.A2(n_1821),
.B(n_1824),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1880),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1861),
.B(n_1836),
.Y(n_1896)
);

OAI22xp33_ASAP7_75t_L g1897 ( 
.A1(n_1887),
.A2(n_1797),
.B1(n_1824),
.B2(n_1834),
.Y(n_1897)
);

OAI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1859),
.A2(n_1778),
.B1(n_1821),
.B2(n_1830),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1852),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1872),
.B(n_1841),
.Y(n_1900)
);

NAND2x1p5_ASAP7_75t_L g1901 ( 
.A(n_1854),
.B(n_1838),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1855),
.B(n_1830),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1865),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1863),
.B(n_1841),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1864),
.Y(n_1905)
);

AOI22xp5_ASAP7_75t_L g1906 ( 
.A1(n_1878),
.A2(n_1729),
.B1(n_1720),
.B2(n_1706),
.Y(n_1906)
);

HB1xp67_ASAP7_75t_L g1907 ( 
.A(n_1869),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1865),
.Y(n_1908)
);

A2O1A1Ixp33_ASAP7_75t_L g1909 ( 
.A1(n_1888),
.A2(n_1743),
.B(n_1797),
.C(n_1808),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1863),
.B(n_1832),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1867),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1862),
.B(n_1832),
.Y(n_1912)
);

INVx2_ASAP7_75t_SL g1913 ( 
.A(n_1855),
.Y(n_1913)
);

INVxp67_ASAP7_75t_L g1914 ( 
.A(n_1857),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1862),
.B(n_1837),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1907),
.Y(n_1916)
);

INVxp67_ASAP7_75t_L g1917 ( 
.A(n_1891),
.Y(n_1917)
);

NAND4xp25_ASAP7_75t_L g1918 ( 
.A(n_1909),
.B(n_1875),
.C(n_1886),
.D(n_1874),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1907),
.Y(n_1919)
);

NAND3xp33_ASAP7_75t_L g1920 ( 
.A(n_1909),
.B(n_1879),
.C(n_1851),
.Y(n_1920)
);

OR2x2_ASAP7_75t_L g1921 ( 
.A(n_1911),
.B(n_1870),
.Y(n_1921)
);

INVx1_ASAP7_75t_SL g1922 ( 
.A(n_1889),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1892),
.Y(n_1923)
);

AOI22xp33_ASAP7_75t_L g1924 ( 
.A1(n_1890),
.A2(n_1743),
.B1(n_1906),
.B2(n_1897),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1895),
.Y(n_1925)
);

HB1xp67_ASAP7_75t_L g1926 ( 
.A(n_1911),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_SL g1927 ( 
.A(n_1897),
.B(n_1875),
.Y(n_1927)
);

AOI211xp5_ASAP7_75t_SL g1928 ( 
.A1(n_1894),
.A2(n_1858),
.B(n_1860),
.C(n_1851),
.Y(n_1928)
);

AO22x1_ASAP7_75t_L g1929 ( 
.A1(n_1896),
.A2(n_1628),
.B1(n_1879),
.B2(n_1881),
.Y(n_1929)
);

OAI222xp33_ASAP7_75t_L g1930 ( 
.A1(n_1893),
.A2(n_1883),
.B1(n_1882),
.B2(n_1870),
.C1(n_1871),
.C2(n_1873),
.Y(n_1930)
);

INVx3_ASAP7_75t_L g1931 ( 
.A(n_1903),
.Y(n_1931)
);

OAI332xp33_ASAP7_75t_L g1932 ( 
.A1(n_1898),
.A2(n_1846),
.A3(n_1883),
.B1(n_1876),
.B2(n_1884),
.B3(n_1877),
.C1(n_1882),
.C2(n_1871),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1899),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1903),
.B(n_1908),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1905),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1910),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1902),
.B(n_1908),
.Y(n_1937)
);

A2O1A1Ixp33_ASAP7_75t_L g1938 ( 
.A1(n_1928),
.A2(n_1915),
.B(n_1912),
.C(n_1900),
.Y(n_1938)
);

OR2x2_ASAP7_75t_L g1939 ( 
.A(n_1921),
.B(n_1904),
.Y(n_1939)
);

INVx1_ASAP7_75t_SL g1940 ( 
.A(n_1922),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1931),
.Y(n_1941)
);

OAI222xp33_ASAP7_75t_L g1942 ( 
.A1(n_1924),
.A2(n_1913),
.B1(n_1901),
.B2(n_1914),
.C1(n_1846),
.C2(n_1806),
.Y(n_1942)
);

NOR2xp33_ASAP7_75t_L g1943 ( 
.A(n_1932),
.B(n_1930),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1937),
.B(n_1913),
.Y(n_1944)
);

OR2x2_ASAP7_75t_L g1945 ( 
.A(n_1921),
.B(n_1867),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1926),
.Y(n_1946)
);

OR2x2_ASAP7_75t_L g1947 ( 
.A(n_1934),
.B(n_1874),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1931),
.B(n_1858),
.Y(n_1948)
);

NOR2x1_ASAP7_75t_L g1949 ( 
.A(n_1927),
.B(n_1860),
.Y(n_1949)
);

O2A1O1Ixp33_ASAP7_75t_L g1950 ( 
.A1(n_1942),
.A2(n_1927),
.B(n_1917),
.C(n_1916),
.Y(n_1950)
);

AOI21xp5_ASAP7_75t_L g1951 ( 
.A1(n_1949),
.A2(n_1916),
.B(n_1919),
.Y(n_1951)
);

AOI21xp5_ASAP7_75t_L g1952 ( 
.A1(n_1943),
.A2(n_1920),
.B(n_1918),
.Y(n_1952)
);

OAI21xp5_ASAP7_75t_SL g1953 ( 
.A1(n_1940),
.A2(n_1901),
.B(n_1937),
.Y(n_1953)
);

OAI21xp33_ASAP7_75t_L g1954 ( 
.A1(n_1944),
.A2(n_1940),
.B(n_1948),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1945),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1941),
.Y(n_1956)
);

INVx1_ASAP7_75t_SL g1957 ( 
.A(n_1939),
.Y(n_1957)
);

INVxp67_ASAP7_75t_SL g1958 ( 
.A(n_1946),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1947),
.Y(n_1959)
);

NAND4xp25_ASAP7_75t_L g1960 ( 
.A(n_1952),
.B(n_1938),
.C(n_1931),
.D(n_1936),
.Y(n_1960)
);

AOI211xp5_ASAP7_75t_L g1961 ( 
.A1(n_1950),
.A2(n_1929),
.B(n_1933),
.C(n_1935),
.Y(n_1961)
);

OAI222xp33_ASAP7_75t_L g1962 ( 
.A1(n_1951),
.A2(n_1925),
.B1(n_1923),
.B2(n_1846),
.C1(n_1929),
.C2(n_1822),
.Y(n_1962)
);

NOR2xp33_ASAP7_75t_R g1963 ( 
.A(n_1957),
.B(n_1959),
.Y(n_1963)
);

AOI222xp33_ASAP7_75t_L g1964 ( 
.A1(n_1958),
.A2(n_1828),
.B1(n_1822),
.B2(n_1844),
.C1(n_1810),
.C2(n_1840),
.Y(n_1964)
);

OAI211xp5_ASAP7_75t_L g1965 ( 
.A1(n_1951),
.A2(n_1885),
.B(n_1771),
.C(n_1739),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1961),
.B(n_1954),
.Y(n_1966)
);

INVx1_ASAP7_75t_SL g1967 ( 
.A(n_1963),
.Y(n_1967)
);

OAI21xp33_ASAP7_75t_SL g1968 ( 
.A1(n_1960),
.A2(n_1956),
.B(n_1955),
.Y(n_1968)
);

AND3x2_ASAP7_75t_L g1969 ( 
.A(n_1962),
.B(n_1953),
.C(n_1628),
.Y(n_1969)
);

AOI21xp5_ASAP7_75t_SL g1970 ( 
.A1(n_1965),
.A2(n_1771),
.B(n_1628),
.Y(n_1970)
);

AOI211xp5_ASAP7_75t_L g1971 ( 
.A1(n_1964),
.A2(n_1885),
.B(n_1850),
.C(n_1828),
.Y(n_1971)
);

AOI22xp33_ASAP7_75t_L g1972 ( 
.A1(n_1960),
.A2(n_1828),
.B1(n_1844),
.B2(n_1810),
.Y(n_1972)
);

CKINVDCx5p33_ASAP7_75t_R g1973 ( 
.A(n_1967),
.Y(n_1973)
);

CKINVDCx20_ASAP7_75t_R g1974 ( 
.A(n_1966),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1969),
.B(n_1837),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_L g1976 ( 
.A(n_1968),
.B(n_1648),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1970),
.Y(n_1977)
);

NOR2xp33_ASAP7_75t_L g1978 ( 
.A(n_1972),
.B(n_1842),
.Y(n_1978)
);

AOI322xp5_ASAP7_75t_L g1979 ( 
.A1(n_1974),
.A2(n_1810),
.A3(n_1822),
.B1(n_1844),
.B2(n_1806),
.C1(n_1840),
.C2(n_1828),
.Y(n_1979)
);

NOR4xp75_ASAP7_75t_L g1980 ( 
.A(n_1975),
.B(n_1971),
.C(n_1746),
.D(n_1800),
.Y(n_1980)
);

OR2x2_ASAP7_75t_L g1981 ( 
.A(n_1973),
.B(n_1842),
.Y(n_1981)
);

OAI21xp5_ASAP7_75t_L g1982 ( 
.A1(n_1976),
.A2(n_1977),
.B(n_1978),
.Y(n_1982)
);

OR2x2_ASAP7_75t_L g1983 ( 
.A(n_1981),
.B(n_1982),
.Y(n_1983)
);

AOI22xp5_ASAP7_75t_L g1984 ( 
.A1(n_1983),
.A2(n_1980),
.B1(n_1979),
.B2(n_1850),
.Y(n_1984)
);

HB1xp67_ASAP7_75t_L g1985 ( 
.A(n_1984),
.Y(n_1985)
);

OAI22xp5_ASAP7_75t_L g1986 ( 
.A1(n_1984),
.A2(n_1849),
.B1(n_1843),
.B2(n_1850),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1985),
.Y(n_1987)
);

OAI21xp5_ASAP7_75t_L g1988 ( 
.A1(n_1986),
.A2(n_1849),
.B(n_1843),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1987),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_SL g1990 ( 
.A(n_1988),
.B(n_1850),
.Y(n_1990)
);

AOI21xp5_ASAP7_75t_L g1991 ( 
.A1(n_1989),
.A2(n_1739),
.B(n_1796),
.Y(n_1991)
);

OR2x2_ASAP7_75t_L g1992 ( 
.A(n_1991),
.B(n_1990),
.Y(n_1992)
);

AOI21xp5_ASAP7_75t_L g1993 ( 
.A1(n_1992),
.A2(n_1644),
.B(n_1800),
.Y(n_1993)
);

OAI221xp5_ASAP7_75t_R g1994 ( 
.A1(n_1993),
.A2(n_1638),
.B1(n_1742),
.B2(n_1769),
.C(n_1784),
.Y(n_1994)
);

AOI211xp5_ASAP7_75t_L g1995 ( 
.A1(n_1994),
.A2(n_1615),
.B(n_1614),
.C(n_1595),
.Y(n_1995)
);


endmodule