module fake_jpeg_1022_n_491 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_491);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_491;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_17),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_5),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_5),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_56),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_57),
.Y(n_130)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_58),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_23),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_59),
.B(n_74),
.Y(n_169)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_62),
.Y(n_125)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_36),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_64),
.B(n_66),
.Y(n_148)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_65),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_32),
.B(n_10),
.Y(n_66)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_67),
.Y(n_194)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx3_ASAP7_75t_SL g127 ( 
.A(n_68),
.Y(n_127)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_69),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_40),
.Y(n_71)
);

NAND2xp33_ASAP7_75t_SL g199 ( 
.A(n_71),
.B(n_117),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_21),
.B(n_10),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_72),
.B(n_88),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_73),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_47),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_75),
.Y(n_140)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_76),
.Y(n_152)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_77),
.Y(n_165)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_78),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_79),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_80),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_47),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_81),
.B(n_91),
.Y(n_172)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_52),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_83),
.Y(n_196)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_84),
.Y(n_174)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_18),
.Y(n_85)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_85),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_86),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_87),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_24),
.B(n_11),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_24),
.B(n_17),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_89),
.B(n_93),
.Y(n_175)
);

BUFx12_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_30),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_31),
.B(n_36),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_95),
.Y(n_171)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_96),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_31),
.B(n_16),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_99),
.B(n_106),
.Y(n_191)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_35),
.Y(n_100)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_102),
.Y(n_151)
);

CKINVDCx12_ASAP7_75t_R g103 ( 
.A(n_25),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_103),
.B(n_111),
.Y(n_180)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_37),
.Y(n_105)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_105),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_28),
.B(n_14),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_25),
.Y(n_107)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_107),
.Y(n_155)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_28),
.Y(n_108)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_108),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_33),
.Y(n_109)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_109),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_26),
.Y(n_110)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_110),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_20),
.B(n_15),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_33),
.Y(n_112)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_112),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_19),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_113),
.B(n_115),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_34),
.Y(n_114)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_114),
.Y(n_164)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_37),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_34),
.Y(n_116)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_116),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_25),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_41),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_119),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_26),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_51),
.C(n_50),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_120),
.B(n_176),
.C(n_140),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_118),
.B(n_19),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_123),
.B(n_156),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_100),
.A2(n_22),
.B1(n_53),
.B2(n_49),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_173),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_83),
.A2(n_51),
.B1(n_50),
.B2(n_41),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_80),
.A2(n_55),
.B1(n_53),
.B2(n_49),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_86),
.A2(n_94),
.B1(n_95),
.B2(n_97),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_147),
.A2(n_158),
.B1(n_159),
.B2(n_167),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_60),
.A2(n_44),
.B(n_48),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_154),
.A2(n_179),
.B(n_167),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_63),
.B(n_55),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_102),
.A2(n_48),
.B1(n_46),
.B2(n_42),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_101),
.A2(n_46),
.B1(n_42),
.B2(n_22),
.Y(n_159)
);

NAND2x1_ASAP7_75t_L g161 ( 
.A(n_61),
.B(n_44),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_161),
.B(n_190),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_76),
.A2(n_20),
.B1(n_1),
.B2(n_2),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_163),
.A2(n_183),
.B1(n_194),
.B2(n_196),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_73),
.B(n_15),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_166),
.B(n_182),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_104),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_77),
.A2(n_12),
.B1(n_13),
.B2(n_4),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_70),
.B(n_12),
.C(n_3),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_98),
.A2(n_0),
.B1(n_4),
.B2(n_7),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_178),
.A2(n_197),
.B1(n_195),
.B2(n_155),
.Y(n_253)
);

OAI21xp33_ASAP7_75t_L g179 ( 
.A1(n_109),
.A2(n_0),
.B(n_4),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_57),
.B(n_7),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_96),
.A2(n_8),
.B1(n_56),
.B2(n_69),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_112),
.B(n_8),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_184),
.B(n_185),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_117),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_57),
.B(n_107),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_188),
.B(n_198),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_114),
.A2(n_116),
.B1(n_67),
.B2(n_68),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_107),
.A2(n_79),
.B1(n_58),
.B2(n_90),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_68),
.B(n_58),
.Y(n_198)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_186),
.Y(n_200)
);

INVxp67_ASAP7_75t_SL g309 ( 
.A(n_200),
.Y(n_309)
);

NAND3xp33_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_90),
.C(n_87),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_201),
.B(n_237),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_121),
.B(n_110),
.Y(n_202)
);

AO22x1_ASAP7_75t_L g270 ( 
.A1(n_202),
.A2(n_226),
.B1(n_227),
.B2(n_237),
.Y(n_270)
);

OA22x2_ASAP7_75t_L g281 ( 
.A1(n_203),
.A2(n_253),
.B1(n_200),
.B2(n_226),
.Y(n_281)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_138),
.Y(n_204)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_204),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_131),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_205),
.Y(n_304)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_142),
.Y(n_207)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_207),
.Y(n_274)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_177),
.Y(n_208)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_208),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_121),
.A2(n_119),
.B(n_159),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_209),
.A2(n_226),
.B(n_202),
.Y(n_279)
);

AND2x2_ASAP7_75t_SL g210 ( 
.A(n_125),
.B(n_137),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_210),
.B(n_232),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_124),
.A2(n_160),
.B1(n_126),
.B2(n_172),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_212),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_127),
.Y(n_214)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_214),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_148),
.B(n_180),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_215),
.B(n_220),
.Y(n_268)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_138),
.Y(n_216)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_216),
.Y(n_285)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_189),
.Y(n_217)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_217),
.Y(n_275)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_165),
.Y(n_218)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_218),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_131),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_219),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_162),
.B(n_175),
.Y(n_220)
);

BUFx12f_ASAP7_75t_L g221 ( 
.A(n_155),
.Y(n_221)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_221),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_181),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_222),
.B(n_229),
.Y(n_276)
);

AO22x1_ASAP7_75t_SL g223 ( 
.A1(n_178),
.A2(n_145),
.B1(n_143),
.B2(n_165),
.Y(n_223)
);

AO22x1_ASAP7_75t_SL g295 ( 
.A1(n_223),
.A2(n_227),
.B1(n_218),
.B2(n_210),
.Y(n_295)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_157),
.Y(n_225)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_225),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_161),
.B(n_199),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_128),
.Y(n_227)
);

INVx13_ASAP7_75t_L g228 ( 
.A(n_135),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_228),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_169),
.B(n_164),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_158),
.B(n_179),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_230),
.B(n_243),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_144),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_231),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_187),
.B(n_192),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_234),
.B(n_239),
.Y(n_271)
);

INVx8_ASAP7_75t_L g235 ( 
.A(n_168),
.Y(n_235)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_235),
.Y(n_284)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_152),
.Y(n_236)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_236),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_127),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_128),
.Y(n_238)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_238),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_129),
.B(n_151),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_135),
.B(n_141),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_240),
.B(n_244),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_149),
.B(n_151),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_241),
.B(n_262),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_141),
.Y(n_242)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_242),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_136),
.B(n_135),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_146),
.B(n_136),
.Y(n_244)
);

OAI211xp5_ASAP7_75t_L g287 ( 
.A1(n_245),
.A2(n_246),
.B(n_247),
.C(n_252),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_144),
.B(n_153),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_146),
.B(n_122),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_153),
.Y(n_248)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_248),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_140),
.Y(n_250)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_250),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_122),
.B(n_130),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_139),
.Y(n_254)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_254),
.Y(n_307)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_149),
.Y(n_255)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_255),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_152),
.Y(n_256)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_256),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_150),
.B(n_195),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_257),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_174),
.B(n_170),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_258),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_174),
.A2(n_170),
.B1(n_122),
.B2(n_183),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_259),
.A2(n_260),
.B1(n_263),
.B2(n_264),
.Y(n_300)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_171),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_163),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_261),
.A2(n_265),
.B1(n_214),
.B2(n_204),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_168),
.B(n_139),
.Y(n_262)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_171),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_147),
.Y(n_264)
);

NOR3xp33_ASAP7_75t_L g265 ( 
.A(n_191),
.B(n_162),
.C(n_175),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_213),
.A2(n_232),
.B1(n_261),
.B2(n_253),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_266),
.A2(n_294),
.B1(n_267),
.B2(n_284),
.Y(n_347)
);

AO22x2_ASAP7_75t_L g267 ( 
.A1(n_223),
.A2(n_209),
.B1(n_233),
.B2(n_224),
.Y(n_267)
);

A2O1A1Ixp33_ASAP7_75t_SL g315 ( 
.A1(n_267),
.A2(n_235),
.B(n_216),
.C(n_236),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_270),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_223),
.A2(n_213),
.B1(n_224),
.B2(n_239),
.Y(n_278)
);

INVxp33_ASAP7_75t_L g350 ( 
.A(n_278),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_279),
.A2(n_283),
.B(n_272),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_281),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_245),
.B(n_251),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_282),
.B(n_287),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_202),
.A2(n_234),
.B(n_227),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_249),
.A2(n_206),
.B1(n_211),
.B2(n_241),
.Y(n_294)
);

OA21x2_ASAP7_75t_L g334 ( 
.A1(n_295),
.A2(n_301),
.B(n_281),
.Y(n_334)
);

O2A1O1Ixp33_ASAP7_75t_L g297 ( 
.A1(n_250),
.A2(n_210),
.B(n_238),
.C(n_225),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_297),
.A2(n_302),
.B(n_283),
.Y(n_328)
);

OA22x2_ASAP7_75t_L g301 ( 
.A1(n_207),
.A2(n_255),
.B1(n_263),
.B2(n_260),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_310),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_315),
.B(n_316),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_271),
.B(n_205),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_271),
.B(n_219),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_317),
.B(n_319),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_298),
.B(n_231),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_297),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_320),
.B(n_321),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_248),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_311),
.Y(n_322)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_322),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_276),
.B(n_221),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_323),
.Y(n_379)
);

XNOR2x2_ASAP7_75t_L g324 ( 
.A(n_282),
.B(n_228),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_324),
.A2(n_328),
.B(n_336),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_273),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_325),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_268),
.B(n_221),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_326),
.B(n_327),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_308),
.B(n_305),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_289),
.B(n_288),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_329),
.B(n_332),
.Y(n_367)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_274),
.Y(n_330)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_330),
.Y(n_371)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_274),
.Y(n_331)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_331),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_306),
.B(n_269),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_306),
.B(n_302),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_333),
.B(n_335),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_334),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_302),
.B(n_266),
.Y(n_335)
);

AOI22x1_ASAP7_75t_SL g336 ( 
.A1(n_267),
.A2(n_279),
.B1(n_281),
.B2(n_270),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_273),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_338),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_339),
.B(n_292),
.C(n_314),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_301),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_341),
.A2(n_343),
.B1(n_349),
.B2(n_351),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_295),
.B(n_267),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_342),
.A2(n_347),
.B1(n_291),
.B2(n_285),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_301),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_281),
.B(n_275),
.Y(n_344)
);

BUFx24_ASAP7_75t_SL g373 ( 
.A(n_344),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_272),
.A2(n_300),
.B(n_295),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_345),
.A2(n_346),
.B(n_309),
.Y(n_355)
);

AO21x2_ASAP7_75t_L g348 ( 
.A1(n_301),
.A2(n_296),
.B(n_280),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_348),
.A2(n_307),
.B1(n_290),
.B2(n_291),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_293),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_293),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_353),
.B(n_319),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_355),
.A2(n_359),
.B(n_340),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_358),
.A2(n_361),
.B1(n_365),
.B2(n_375),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_328),
.A2(n_346),
.B(n_344),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_339),
.B(n_286),
.C(n_285),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_360),
.B(n_378),
.C(n_380),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_347),
.A2(n_318),
.B1(n_342),
.B2(n_350),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_363),
.B(n_376),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_318),
.A2(n_304),
.B1(n_312),
.B2(n_299),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_334),
.A2(n_304),
.B1(n_312),
.B2(n_299),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_366),
.A2(n_348),
.B1(n_334),
.B2(n_357),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_334),
.A2(n_277),
.B1(n_303),
.B2(n_341),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_372),
.A2(n_348),
.B1(n_315),
.B2(n_317),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_335),
.A2(n_277),
.B1(n_303),
.B2(n_343),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_337),
.A2(n_320),
.B1(n_345),
.B2(n_333),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_324),
.B(n_332),
.C(n_327),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_324),
.B(n_336),
.C(n_316),
.Y(n_380)
);

INVx4_ASAP7_75t_SL g382 ( 
.A(n_357),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_382),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_379),
.B(n_326),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_383),
.B(n_384),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_367),
.B(n_323),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_367),
.B(n_329),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_385),
.B(n_387),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_386),
.B(n_360),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_362),
.B(n_321),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_388),
.A2(n_391),
.B1(n_356),
.B2(n_364),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_389),
.Y(n_416)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_352),
.Y(n_390)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_390),
.Y(n_417)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_352),
.Y(n_392)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_392),
.Y(n_423)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_371),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_393),
.B(n_398),
.Y(n_409)
);

CKINVDCx14_ASAP7_75t_R g396 ( 
.A(n_362),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_396),
.B(n_404),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_381),
.B(n_322),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_397),
.B(n_381),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_369),
.B(n_315),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_371),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_399),
.B(n_400),
.Y(n_425)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_377),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_369),
.B(n_338),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_401),
.B(n_403),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_370),
.B(n_315),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_377),
.Y(n_404)
);

AO32x1_ASAP7_75t_L g405 ( 
.A1(n_373),
.A2(n_315),
.A3(n_348),
.B1(n_325),
.B2(n_349),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_405),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_370),
.B(n_351),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_406),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_408),
.B(n_418),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_395),
.B(n_378),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_410),
.B(n_413),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_SL g418 ( 
.A(n_397),
.B(n_381),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_395),
.B(n_353),
.C(n_354),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_419),
.B(n_422),
.C(n_406),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_421),
.A2(n_363),
.B1(n_411),
.B2(n_409),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_386),
.B(n_354),
.C(n_380),
.Y(n_422)
);

XNOR2x1_ASAP7_75t_L g424 ( 
.A(n_389),
.B(n_359),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_424),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_394),
.A2(n_356),
.B1(n_372),
.B2(n_364),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_427),
.A2(n_375),
.B1(n_391),
.B2(n_402),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_427),
.A2(n_388),
.B1(n_382),
.B2(n_361),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_428),
.A2(n_434),
.B1(n_436),
.B2(n_421),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_420),
.B(n_401),
.Y(n_429)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_429),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_416),
.A2(n_382),
.B1(n_376),
.B2(n_394),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_430),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_431),
.B(n_443),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_432),
.B(n_433),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_426),
.A2(n_398),
.B(n_403),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_414),
.A2(n_366),
.B1(n_365),
.B2(n_402),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_410),
.B(n_355),
.C(n_368),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_437),
.B(n_440),
.C(n_424),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_415),
.B(n_368),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_438),
.B(n_442),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_419),
.B(n_413),
.C(n_422),
.Y(n_440)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_425),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_408),
.B(n_374),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_443),
.B(n_418),
.Y(n_446)
);

MAJx2_ASAP7_75t_L g464 ( 
.A(n_446),
.B(n_452),
.C(n_439),
.Y(n_464)
);

OAI21xp33_ASAP7_75t_L g447 ( 
.A1(n_441),
.A2(n_416),
.B(n_426),
.Y(n_447)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_447),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_449),
.A2(n_374),
.B1(n_405),
.B2(n_423),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_441),
.A2(n_407),
.B(n_409),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_451),
.B(n_455),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_435),
.B(n_407),
.C(n_425),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_454),
.B(n_431),
.C(n_435),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_433),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_444),
.A2(n_428),
.B1(n_437),
.B2(n_405),
.Y(n_457)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_457),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_453),
.B(n_412),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_458),
.B(n_459),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_SL g460 ( 
.A(n_446),
.B(n_439),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_460),
.B(n_463),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_450),
.B(n_440),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_461),
.B(n_465),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_464),
.B(n_452),
.Y(n_468)
);

OAI221xp5_ASAP7_75t_L g465 ( 
.A1(n_448),
.A2(n_423),
.B1(n_417),
.B2(n_430),
.C(n_392),
.Y(n_465)
);

OR2x2_ASAP7_75t_L g478 ( 
.A(n_468),
.B(n_473),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_456),
.A2(n_445),
.B(n_447),
.Y(n_470)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_470),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_462),
.A2(n_449),
.B(n_450),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_472),
.B(n_460),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_459),
.B(n_454),
.C(n_404),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_471),
.B(n_457),
.C(n_464),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_474),
.B(n_476),
.Y(n_480)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_475),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_467),
.B(n_417),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_473),
.B(n_390),
.Y(n_479)
);

INVxp33_ASAP7_75t_L g481 ( 
.A(n_479),
.Y(n_481)
);

A2O1A1Ixp33_ASAP7_75t_L g482 ( 
.A1(n_477),
.A2(n_470),
.B(n_466),
.C(n_469),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_482),
.A2(n_475),
.B(n_469),
.Y(n_484)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_484),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_480),
.Y(n_485)
);

A2O1A1O1Ixp25_ASAP7_75t_L g486 ( 
.A1(n_485),
.A2(n_481),
.B(n_483),
.C(n_478),
.D(n_399),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_486),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_488),
.A2(n_487),
.B(n_393),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_489),
.A2(n_400),
.B(n_358),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_490),
.B(n_348),
.Y(n_491)
);


endmodule