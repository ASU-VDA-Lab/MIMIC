module real_jpeg_32624_n_9 (n_79, n_5, n_4, n_8, n_0, n_81, n_84, n_85, n_1, n_80, n_78, n_2, n_82, n_83, n_6, n_7, n_3, n_9);

input n_79;
input n_5;
input n_4;
input n_8;
input n_0;
input n_81;
input n_84;
input n_85;
input n_1;
input n_80;
input n_78;
input n_2;
input n_82;
input n_83;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_49;
wire n_10;
wire n_68;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_65;
wire n_33;
wire n_67;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_39;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_61;
wire n_70;
wire n_41;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_57;
wire n_43;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_16;

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_0),
.B(n_36),
.Y(n_35)
);

AOI221xp5_ASAP7_75t_L g33 ( 
.A1(n_1),
.A2(n_3),
.B1(n_34),
.B2(n_40),
.C(n_42),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_1),
.B(n_34),
.C(n_40),
.Y(n_45)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g10 ( 
.A1(n_4),
.A2(n_11),
.B1(n_12),
.B2(n_18),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_6),
.B(n_72),
.Y(n_71)
);

HAxp5_ASAP7_75t_SL g74 ( 
.A(n_6),
.B(n_75),
.CON(n_74),
.SN(n_74)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_7),
.B(n_64),
.Y(n_70)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_19),
.Y(n_9)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_14),
.Y(n_12)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_71),
.B(n_74),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_62),
.B(n_69),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_56),
.C(n_57),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_46),
.B(n_55),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_33),
.B1(n_44),
.B2(n_45),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_35),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_81),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_54),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_54),
.Y(n_55)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_68),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

BUFx24_ASAP7_75t_SL g77 ( 
.A(n_74),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_78),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_79),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_80),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_82),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_83),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_84),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_85),
.Y(n_73)
);


endmodule