module fake_jpeg_11829_n_28 (n_3, n_2, n_1, n_0, n_4, n_5, n_28);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_28;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

AOI22xp33_ASAP7_75t_SL g6 ( 
.A1(n_5),
.A2(n_1),
.B1(n_4),
.B2(n_3),
.Y(n_6)
);

OAI22xp33_ASAP7_75t_L g7 ( 
.A1(n_3),
.A2(n_5),
.B1(n_4),
.B2(n_2),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_0),
.B(n_3),
.Y(n_8)
);

INVx6_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

OAI22xp5_ASAP7_75t_SL g12 ( 
.A1(n_6),
.A2(n_0),
.B1(n_1),
.B2(n_9),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_12),
.A2(n_15),
.B1(n_17),
.B2(n_11),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_8),
.B(n_1),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g15 ( 
.A1(n_6),
.A2(n_8),
.B(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_16),
.A2(n_9),
.B1(n_11),
.B2(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_18),
.A2(n_20),
.B(n_17),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_15),
.A2(n_9),
.B1(n_7),
.B2(n_11),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_22),
.B(n_9),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_24),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_12),
.C(n_19),
.Y(n_25)
);

NOR2xp67_ASAP7_75t_SL g26 ( 
.A(n_25),
.B(n_19),
.Y(n_26)
);

OAI21x1_ASAP7_75t_L g28 ( 
.A1(n_26),
.A2(n_21),
.B(n_27),
.Y(n_28)
);


endmodule