module fake_jpeg_296_n_125 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_125);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_9),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_6),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_6),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_7),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_41),
.Y(n_52)
);

HAxp5_ASAP7_75t_SL g41 ( 
.A(n_21),
.B(n_0),
.CON(n_41),
.SN(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_44),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_15),
.B1(n_19),
.B2(n_27),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_47),
.A2(n_57),
.B1(n_61),
.B2(n_39),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_34),
.A2(n_37),
.B1(n_42),
.B2(n_36),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_58),
.A2(n_60),
.B1(n_55),
.B2(n_31),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_30),
.A2(n_27),
.B1(n_24),
.B2(n_22),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_44),
.A2(n_24),
.B1(n_16),
.B2(n_1),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_50),
.A2(n_35),
.B1(n_41),
.B2(n_39),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_53),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_16),
.C(n_32),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_67),
.C(n_74),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_68),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_51),
.B(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_69),
.Y(n_78)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_31),
.C(n_23),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_70),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_72),
.Y(n_81)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

NOR3xp33_ASAP7_75t_SL g88 ( 
.A(n_73),
.B(n_75),
.C(n_2),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_57),
.A2(n_54),
.B(n_61),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_53),
.A2(n_23),
.B1(n_4),
.B2(n_5),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_59),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_77),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_54),
.B(n_2),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_64),
.A2(n_59),
.B1(n_45),
.B2(n_7),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_80),
.A2(n_66),
.B1(n_70),
.B2(n_68),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_45),
.C(n_4),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_62),
.C(n_11),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_11),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_85),
.A2(n_76),
.B(n_74),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_89),
.A2(n_87),
.B(n_79),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_75),
.B1(n_63),
.B2(n_62),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_93),
.B1(n_80),
.B2(n_84),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_78),
.B(n_9),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_96),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_95),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_62),
.C(n_69),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_10),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_81),
.B(n_14),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_98),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_103),
.C(n_105),
.Y(n_113)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_86),
.Y(n_104)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_105),
.A2(n_88),
.B1(n_94),
.B2(n_45),
.Y(n_108)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_107),
.Y(n_111)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_104),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_113),
.Y(n_116)
);

OA21x2_ASAP7_75t_SL g114 ( 
.A1(n_113),
.A2(n_99),
.B(n_109),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_111),
.Y(n_118)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_116),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_117),
.A2(n_110),
.B(n_106),
.C(n_100),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_118),
.A2(n_115),
.B(n_110),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_120),
.C(n_109),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_114),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_115),
.B(n_103),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_108),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_102),
.Y(n_125)
);


endmodule