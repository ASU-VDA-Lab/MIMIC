module fake_jpeg_1849_n_427 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_427);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_427;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_292;
wire n_213;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_352;
wire n_350;
wire n_150;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx4f_ASAP7_75t_SL g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_4),
.B(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_46),
.Y(n_128)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_48),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_8),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_49),
.B(n_62),
.Y(n_142)
);

INVx11_ASAP7_75t_SL g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_43),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_51),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_8),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_52),
.B(n_53),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_30),
.B(n_8),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_30),
.B(n_8),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_57),
.B(n_63),
.Y(n_120)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_58),
.Y(n_132)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_59),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_39),
.B(n_2),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_2),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_19),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_64),
.B(n_69),
.Y(n_130)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_43),
.B(n_24),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_67),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx3_ASAP7_75t_SL g109 ( 
.A(n_68),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_40),
.B(n_6),
.Y(n_69)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_70),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_19),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_71),
.B(n_74),
.Y(n_133)
);

BUFx24_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_72),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_73),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_41),
.B(n_6),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_80),
.Y(n_144)
);

BUFx24_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_20),
.B(n_6),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_97),
.Y(n_99)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_19),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_84),
.B(n_85),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_41),
.B(n_7),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_86),
.Y(n_152)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_87),
.B(n_95),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_14),
.Y(n_92)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_28),
.Y(n_93)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_14),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_96),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_14),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_44),
.B(n_7),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_98),
.A2(n_27),
.B1(n_26),
.B2(n_22),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_54),
.A2(n_32),
.B1(n_20),
.B2(n_36),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_100),
.A2(n_117),
.B1(n_125),
.B2(n_126),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_52),
.A2(n_35),
.B1(n_36),
.B2(n_16),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_110),
.A2(n_137),
.B1(n_72),
.B2(n_97),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_111),
.B(n_45),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_50),
.A2(n_32),
.B1(n_36),
.B2(n_27),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_51),
.A2(n_32),
.B1(n_26),
.B2(n_22),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_76),
.A2(n_32),
.B1(n_90),
.B2(n_47),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_83),
.A2(n_17),
.B1(n_16),
.B2(n_15),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_127),
.A2(n_149),
.B1(n_151),
.B2(n_34),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_63),
.A2(n_35),
.B1(n_15),
.B2(n_17),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_92),
.A2(n_28),
.B1(n_35),
.B2(n_31),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_147),
.A2(n_91),
.B1(n_88),
.B2(n_96),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_70),
.A2(n_45),
.B1(n_31),
.B2(n_29),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_72),
.A2(n_45),
.B1(n_42),
.B2(n_34),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_103),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_155),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_156),
.B(n_170),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_124),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_157),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_99),
.B(n_67),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_158),
.B(n_160),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_94),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_165),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_99),
.B(n_67),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_103),
.Y(n_161)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_161),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_162),
.A2(n_163),
.B1(n_112),
.B2(n_109),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_111),
.A2(n_56),
.B1(n_55),
.B2(n_60),
.Y(n_163)
);

BUFx24_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_164),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_95),
.Y(n_165)
);

OR2x2_ASAP7_75t_SL g166 ( 
.A(n_148),
.B(n_81),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_166),
.Y(n_206)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_168),
.Y(n_197)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_144),
.Y(n_169)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_169),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_128),
.B(n_89),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_130),
.B(n_0),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_171),
.B(n_190),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_131),
.B(n_73),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_172),
.B(n_177),
.Y(n_220)
);

AND2x4_ASAP7_75t_L g173 ( 
.A(n_105),
.B(n_81),
.Y(n_173)
);

NOR2x1_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_187),
.Y(n_198)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_145),
.Y(n_174)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_174),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_105),
.B(n_73),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_175),
.B(n_179),
.Y(n_226)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_176),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_142),
.B(n_80),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_178),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_113),
.B(n_0),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_132),
.B(n_78),
.C(n_77),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_194),
.C(n_195),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_114),
.Y(n_181)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_144),
.Y(n_182)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_122),
.Y(n_183)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_183),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_184),
.B(n_186),
.Y(n_224)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_122),
.Y(n_185)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_185),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_133),
.Y(n_186)
);

NAND3xp33_ASAP7_75t_L g187 ( 
.A(n_102),
.B(n_13),
.C(n_7),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_119),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_188),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_119),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_189),
.Y(n_221)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_116),
.Y(n_190)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_143),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_191),
.B(n_193),
.Y(n_211)
);

AO21x2_ASAP7_75t_L g214 ( 
.A1(n_192),
.A2(n_134),
.B(n_118),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_112),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_136),
.B(n_0),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_138),
.B(n_68),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_158),
.A2(n_134),
.B1(n_108),
.B2(n_106),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_209),
.A2(n_214),
.B1(n_217),
.B2(n_222),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_212),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_160),
.A2(n_106),
.B1(n_108),
.B2(n_123),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_184),
.A2(n_113),
.B1(n_123),
.B2(n_121),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_223),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_228),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_219),
.Y(n_229)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_229),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_211),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_230),
.B(n_231),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_202),
.B(n_171),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_196),
.B(n_166),
.C(n_180),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_240),
.C(n_173),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_211),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_233),
.B(n_237),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_194),
.Y(n_234)
);

A2O1A1O1Ixp25_ASAP7_75t_L g267 ( 
.A1(n_234),
.A2(n_236),
.B(n_248),
.C(n_250),
.D(n_251),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_226),
.Y(n_235)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_235),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_195),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_178),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_216),
.A2(n_154),
.B1(n_179),
.B2(n_121),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_238),
.A2(n_241),
.B1(n_206),
.B2(n_209),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_207),
.B(n_183),
.Y(n_239)
);

OAI21xp33_ASAP7_75t_SL g257 ( 
.A1(n_239),
.A2(n_242),
.B(n_173),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_201),
.B(n_185),
.C(n_135),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_214),
.A2(n_220),
.B1(n_200),
.B2(n_206),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_189),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_218),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_243),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_218),
.Y(n_245)
);

NAND2xp33_ASAP7_75t_SL g263 ( 
.A(n_245),
.B(n_247),
.Y(n_263)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_227),
.Y(n_246)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_246),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_215),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_200),
.B(n_179),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_203),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_249),
.A2(n_253),
.B(n_197),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_190),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_173),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_224),
.B(n_152),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_199),
.Y(n_254)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_254),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_255),
.A2(n_258),
.B1(n_259),
.B2(n_261),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_264),
.C(n_268),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_257),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_241),
.A2(n_214),
.B1(n_217),
.B2(n_222),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_252),
.A2(n_238),
.B1(n_230),
.B2(n_233),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_252),
.A2(n_214),
.B1(n_227),
.B2(n_210),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_210),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_262),
.B(n_248),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_135),
.C(n_204),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_243),
.A2(n_214),
.B(n_245),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_266),
.A2(n_197),
.B(n_221),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_240),
.B(n_198),
.Y(n_268)
);

OAI32xp33_ASAP7_75t_L g270 ( 
.A1(n_234),
.A2(n_204),
.A3(n_199),
.B1(n_205),
.B2(n_169),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_270),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_252),
.A2(n_214),
.B1(n_208),
.B2(n_155),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_273),
.A2(n_249),
.B1(n_254),
.B2(n_203),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_276),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_232),
.B(n_198),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_279),
.C(n_232),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_235),
.B(n_175),
.C(n_139),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_274),
.Y(n_281)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_281),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_276),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_282),
.B(n_297),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g283 ( 
.A1(n_278),
.A2(n_244),
.B1(n_247),
.B2(n_237),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_283),
.A2(n_298),
.B1(n_300),
.B2(n_301),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_284),
.B(n_285),
.C(n_293),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_256),
.B(n_277),
.C(n_268),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_286),
.B(n_272),
.Y(n_307)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_287),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_266),
.A2(n_251),
.B(n_239),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_288),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_271),
.B(n_231),
.Y(n_291)
);

INVxp33_ASAP7_75t_L g304 ( 
.A(n_291),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_253),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_292),
.B(n_272),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_262),
.B(n_250),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_246),
.Y(n_295)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_295),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_264),
.B(n_242),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_296),
.B(n_285),
.C(n_280),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_273),
.A2(n_228),
.B1(n_203),
.B2(n_223),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_259),
.A2(n_228),
.B1(n_229),
.B2(n_225),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_275),
.Y(n_302)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_302),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_263),
.A2(n_198),
.B(n_219),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_303),
.Y(n_316)
);

CKINVDCx14_ASAP7_75t_R g342 ( 
.A(n_306),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_307),
.B(n_175),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_279),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_308),
.B(n_289),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_290),
.A2(n_261),
.B1(n_258),
.B2(n_255),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_309),
.B(n_295),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_291),
.B(n_229),
.Y(n_312)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_312),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_290),
.A2(n_267),
.B1(n_269),
.B2(n_260),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_315),
.A2(n_322),
.B1(n_325),
.B2(n_301),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_280),
.B(n_260),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_317),
.B(n_318),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_288),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_299),
.A2(n_269),
.B1(n_267),
.B2(n_228),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_310),
.C(n_308),
.Y(n_331)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_281),
.Y(n_324)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_324),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_299),
.A2(n_225),
.B1(n_221),
.B2(n_161),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_293),
.B(n_205),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_326),
.B(n_302),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_327),
.A2(n_329),
.B1(n_340),
.B2(n_182),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_313),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_328),
.B(n_335),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_307),
.B(n_284),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_330),
.B(n_337),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_331),
.B(n_336),
.C(n_339),
.Y(n_354)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_305),
.Y(n_332)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_332),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_314),
.A2(n_313),
.B(n_316),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_333),
.A2(n_316),
.B(n_325),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_314),
.Y(n_335)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_335),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_323),
.B(n_286),
.C(n_294),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_310),
.B(n_303),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_315),
.B(n_294),
.C(n_287),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_320),
.A2(n_282),
.B1(n_298),
.B2(n_297),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_341),
.B(n_115),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_304),
.B(n_300),
.Y(n_343)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_343),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_344),
.B(n_347),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_320),
.B(n_289),
.Y(n_345)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_345),
.Y(n_364)
);

NOR2x1_ASAP7_75t_L g348 ( 
.A(n_333),
.B(n_345),
.Y(n_348)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_348),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_350),
.A2(n_356),
.B(n_362),
.Y(n_375)
);

AOI322xp5_ASAP7_75t_L g351 ( 
.A1(n_327),
.A2(n_309),
.A3(n_305),
.B1(n_319),
.B2(n_324),
.C1(n_311),
.C2(n_321),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_351),
.B(n_353),
.Y(n_367)
);

AOI322xp5_ASAP7_75t_L g353 ( 
.A1(n_343),
.A2(n_319),
.A3(n_321),
.B1(n_168),
.B2(n_167),
.C1(n_174),
.C2(n_118),
.Y(n_353)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_355),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_339),
.A2(n_191),
.B(n_104),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_334),
.B(n_213),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_357),
.B(n_360),
.Y(n_369)
);

FAx1_ASAP7_75t_SL g360 ( 
.A(n_336),
.B(n_340),
.CI(n_337),
.CON(n_360),
.SN(n_360)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_342),
.B(n_213),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_363),
.A2(n_109),
.B1(n_101),
.B2(n_129),
.Y(n_379)
);

OAI221xp5_ASAP7_75t_L g377 ( 
.A1(n_365),
.A2(n_115),
.B1(n_129),
.B2(n_107),
.C(n_176),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_349),
.B(n_344),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_366),
.B(n_370),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_354),
.B(n_331),
.C(n_330),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_368),
.B(n_372),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_349),
.B(n_338),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_352),
.B(n_347),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_371),
.B(n_380),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_354),
.B(n_346),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_356),
.B(n_332),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_374),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_348),
.A2(n_139),
.B(n_104),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_376),
.A2(n_358),
.B(n_362),
.Y(n_382)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_377),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_359),
.A2(n_181),
.B1(n_101),
.B2(n_146),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_378),
.A2(n_357),
.B1(n_364),
.B2(n_146),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_379),
.A2(n_358),
.B1(n_361),
.B2(n_359),
.Y(n_388)
);

XNOR2x1_ASAP7_75t_L g380 ( 
.A(n_348),
.B(n_143),
.Y(n_380)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_382),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_368),
.B(n_352),
.C(n_361),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_384),
.B(n_390),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_370),
.Y(n_386)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_386),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_388),
.B(n_394),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_369),
.B(n_350),
.C(n_363),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_367),
.A2(n_355),
.B(n_360),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_391),
.A2(n_392),
.B(n_366),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_381),
.B(n_364),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_393),
.B(n_380),
.Y(n_404)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_373),
.Y(n_394)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_396),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_385),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_399),
.B(n_400),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_384),
.B(n_374),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_390),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_402),
.B(n_404),
.Y(n_412)
);

MAJx2_ASAP7_75t_L g403 ( 
.A(n_383),
.B(n_360),
.C(n_371),
.Y(n_403)
);

AOI21x1_ASAP7_75t_L g409 ( 
.A1(n_403),
.A2(n_375),
.B(n_383),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_395),
.B(n_365),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_405),
.B(n_150),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_398),
.A2(n_387),
.B(n_389),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_408),
.A2(n_399),
.B(n_406),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_409),
.A2(n_414),
.B(n_164),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_402),
.A2(n_388),
.B1(n_378),
.B2(n_389),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_410),
.B(n_413),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_401),
.A2(n_107),
.B1(n_150),
.B2(n_164),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_415),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_411),
.B(n_397),
.C(n_403),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_417),
.B(n_418),
.C(n_419),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_408),
.A2(n_42),
.B(n_34),
.Y(n_419)
);

A2O1A1Ixp33_ASAP7_75t_SL g420 ( 
.A1(n_416),
.A2(n_412),
.B(n_410),
.C(n_407),
.Y(n_420)
);

OAI211xp5_ASAP7_75t_L g423 ( 
.A1(n_420),
.A2(n_42),
.B(n_11),
.C(n_13),
.Y(n_423)
);

NOR3xp33_ASAP7_75t_L g425 ( 
.A(n_423),
.B(n_424),
.C(n_422),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_421),
.B(n_10),
.C(n_11),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_425),
.B(n_13),
.C(n_10),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_426),
.A2(n_11),
.B(n_13),
.Y(n_427)
);


endmodule