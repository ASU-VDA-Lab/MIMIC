module fake_jpeg_552_n_191 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_191);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_191;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

INVx8_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_49),
.Y(n_59)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx8_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_45),
.B(n_46),
.Y(n_56)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

HAxp5_ASAP7_75t_SL g48 ( 
.A(n_17),
.B(n_0),
.CON(n_48),
.SN(n_48)
);

AOI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_48),
.A2(n_30),
.B(n_29),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_17),
.B(n_0),
.Y(n_49)
);

CKINVDCx12_ASAP7_75t_R g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_52),
.Y(n_62)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_29),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_53),
.A2(n_23),
.B1(n_21),
.B2(n_26),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_4),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_40),
.A2(n_27),
.B1(n_22),
.B2(n_24),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_61),
.A2(n_63),
.B1(n_5),
.B2(n_6),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_35),
.A2(n_27),
.B1(n_22),
.B2(n_24),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_34),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_64),
.B(n_65),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_34),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_33),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_67),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_33),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_70),
.A2(n_73),
.B1(n_23),
.B2(n_20),
.Y(n_81)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_41),
.A2(n_30),
.B1(n_26),
.B2(n_23),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_32),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_74),
.B(n_76),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_16),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_23),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_77),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_90),
.Y(n_113)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_56),
.A2(n_48),
.B(n_3),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_2),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_91),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_2),
.C(n_4),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_97),
.C(n_103),
.Y(n_117)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_88),
.B(n_57),
.Y(n_107)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_62),
.A2(n_5),
.B(n_7),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_5),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_99),
.Y(n_121)
);

INVx5_ASAP7_75t_SL g93 ( 
.A(n_80),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_95),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_60),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_94),
.A2(n_55),
.B1(n_69),
.B2(n_72),
.Y(n_110)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_9),
.C(n_10),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_80),
.A2(n_9),
.B1(n_11),
.B2(n_15),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_55),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_58),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_101),
.B(n_106),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_80),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_57),
.A2(n_54),
.B(n_71),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_54),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_79),
.Y(n_106)
);

OAI21x1_ASAP7_75t_L g137 ( 
.A1(n_107),
.A2(n_123),
.B(n_124),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_110),
.A2(n_94),
.B1(n_96),
.B2(n_103),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_104),
.B(n_99),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_112),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_100),
.B(n_57),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_85),
.B(n_54),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_122),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_88),
.B(n_55),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_84),
.B(n_54),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_93),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_69),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_103),
.C(n_87),
.Y(n_131)
);

BUFx6f_ASAP7_75t_SL g127 ( 
.A(n_109),
.Y(n_127)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_108),
.A2(n_83),
.B(n_88),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_131),
.C(n_140),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_124),
.A2(n_105),
.B(n_106),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_130),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_91),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_134),
.Y(n_146)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_107),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_116),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_139),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_102),
.B(n_89),
.Y(n_138)
);

NAND3xp33_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_143),
.C(n_113),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_114),
.A2(n_101),
.B(n_95),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_86),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_141),
.B(n_142),
.Y(n_144)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_113),
.A2(n_82),
.B(n_90),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_145),
.B(n_148),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_128),
.B(n_121),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_128),
.B(n_121),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_155),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_117),
.C(n_118),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_154),
.C(n_135),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_141),
.B(n_117),
.C(n_113),
.Y(n_154)
);

BUFx24_ASAP7_75t_SL g155 ( 
.A(n_138),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_129),
.B(n_122),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_157),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_151),
.A2(n_143),
.B1(n_137),
.B2(n_130),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_158),
.A2(n_149),
.B1(n_147),
.B2(n_139),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_159),
.Y(n_172)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

AOI31xp33_ASAP7_75t_L g161 ( 
.A1(n_154),
.A2(n_137),
.A3(n_132),
.B(n_133),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_136),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_132),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_165),
.C(n_167),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_140),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_169),
.B(n_174),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_147),
.C(n_149),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_162),
.C(n_165),
.Y(n_177)
);

NOR3xp33_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_163),
.C(n_164),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_166),
.A2(n_127),
.B(n_134),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_173),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_178),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_168),
.C(n_142),
.Y(n_184)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_172),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_180),
.Y(n_183)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_172),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_175),
.A2(n_158),
.B1(n_170),
.B2(n_168),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_184),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_181),
.A2(n_178),
.B(n_159),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_185),
.A2(n_186),
.B(n_183),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_182),
.A2(n_119),
.B(n_97),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_187),
.Y(n_188)
);

OAI32xp33_ASAP7_75t_SL g190 ( 
.A1(n_188),
.A2(n_189),
.A3(n_119),
.B1(n_96),
.B2(n_110),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_96),
.Y(n_191)
);


endmodule