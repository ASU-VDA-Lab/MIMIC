module fake_jpeg_12499_n_88 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_88);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_88;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_6),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_0),
.B(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_12),
.B(n_8),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_25),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_23),
.A2(n_13),
.B1(n_19),
.B2(n_11),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_12),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_24)
);

NOR2x1_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_13),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_17),
.B(n_2),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

NAND2xp33_ASAP7_75t_SL g31 ( 
.A(n_26),
.B(n_27),
.Y(n_31)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_28),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_10),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_14),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_19),
.B1(n_15),
.B2(n_18),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_35),
.B(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_29),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g37 ( 
.A1(n_26),
.A2(n_16),
.B1(n_14),
.B2(n_21),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_25),
.C(n_23),
.Y(n_43)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx2_ASAP7_75t_SL g47 ( 
.A(n_39),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_24),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_40),
.B(n_43),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_24),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_45),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_18),
.B(n_21),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_46),
.A2(n_34),
.B1(n_49),
.B2(n_43),
.Y(n_60)
);

AND2x2_ASAP7_75t_SL g48 ( 
.A(n_37),
.B(n_38),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_31),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_50),
.B(n_20),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_57),
.Y(n_61)
);

NOR3xp33_ASAP7_75t_SL g54 ( 
.A(n_42),
.B(n_35),
.C(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_54),
.B(n_55),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_45),
.B(n_15),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_37),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_48),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_59),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_65),
.B(n_30),
.Y(n_74)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_67),
.Y(n_70)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_58),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_51),
.B(n_64),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_73),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_53),
.C(n_51),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_31),
.C(n_63),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_68),
.A2(n_44),
.B(n_54),
.C(n_62),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_74),
.A2(n_48),
.B1(n_47),
.B2(n_46),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_70),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_71),
.C(n_63),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_79),
.A2(n_77),
.B1(n_78),
.B2(n_9),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_39),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_39),
.C(n_8),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_81),
.B(n_9),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_84),
.Y(n_85)
);

OAI21x1_ASAP7_75t_SL g87 ( 
.A1(n_86),
.A2(n_83),
.B(n_39),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_85),
.Y(n_88)
);


endmodule