module fake_jpeg_16981_n_353 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_353);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_353;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_39),
.B(n_43),
.Y(n_76)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_46),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_49),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_56),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_32),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_59),
.Y(n_83)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_61),
.Y(n_86)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_19),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_67),
.Y(n_96)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_65),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_19),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_29),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_79),
.A2(n_90),
.B1(n_104),
.B2(n_30),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_82),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_49),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_84),
.B(n_77),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_22),
.B1(n_33),
.B2(n_31),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_89),
.A2(n_75),
.B1(n_46),
.B2(n_65),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_58),
.A2(n_33),
.B1(n_31),
.B2(n_48),
.Y(n_90)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_59),
.B(n_40),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_49),
.C(n_77),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_68),
.A2(n_33),
.B1(n_31),
.B2(n_48),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_L g115 ( 
.A1(n_92),
.A2(n_48),
.B1(n_71),
.B2(n_72),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_53),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_93),
.B(n_30),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_73),
.B(n_26),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_97),
.B(n_98),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_69),
.B(n_24),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_74),
.Y(n_101)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_64),
.B(n_29),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_61),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_74),
.Y(n_106)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_103),
.Y(n_107)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_107),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_40),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_109),
.B(n_126),
.C(n_129),
.Y(n_149)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_111),
.Y(n_140)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

INVxp33_ASAP7_75t_L g163 ( 
.A(n_112),
.Y(n_163)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_115),
.A2(n_119),
.B1(n_131),
.B2(n_101),
.Y(n_143)
);

OAI32xp33_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_25),
.A3(n_21),
.B1(n_20),
.B2(n_24),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_118),
.A2(n_79),
.B1(n_104),
.B2(n_21),
.Y(n_139)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_82),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_121),
.B(n_125),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_25),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_123),
.B(n_124),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_20),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_82),
.Y(n_125)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

INVx11_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_134),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_91),
.B(n_41),
.C(n_37),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

INVx5_ASAP7_75t_SL g160 ( 
.A(n_130),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_132),
.B(n_26),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_91),
.B(n_88),
.C(n_86),
.Y(n_133)
);

FAx1_ASAP7_75t_SL g151 ( 
.A(n_133),
.B(n_88),
.CI(n_35),
.CON(n_151),
.SN(n_151)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_128),
.A2(n_66),
.B1(n_102),
.B2(n_87),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_137),
.A2(n_139),
.B1(n_142),
.B2(n_143),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_129),
.A2(n_79),
.B1(n_104),
.B2(n_92),
.Y(n_142)
);

AO22x1_ASAP7_75t_SL g144 ( 
.A1(n_109),
.A2(n_102),
.B1(n_37),
.B2(n_38),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_144),
.A2(n_147),
.B1(n_94),
.B2(n_113),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_146),
.B(n_155),
.Y(n_164)
);

OA22x2_ASAP7_75t_L g147 ( 
.A1(n_127),
.A2(n_130),
.B1(n_101),
.B2(n_102),
.Y(n_147)
);

AND2x2_ASAP7_75t_SL g148 ( 
.A(n_126),
.B(n_133),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_148),
.A2(n_154),
.B(n_135),
.Y(n_167)
);

XOR2x1_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_34),
.Y(n_181)
);

AO21x2_ASAP7_75t_L g153 ( 
.A1(n_115),
.A2(n_42),
.B(n_99),
.Y(n_153)
);

AO21x2_ASAP7_75t_L g188 ( 
.A1(n_153),
.A2(n_117),
.B(n_99),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_134),
.A2(n_95),
.B(n_78),
.Y(n_154)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_136),
.B(n_16),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_157),
.B(n_158),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_35),
.Y(n_158)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

INVxp33_ASAP7_75t_SL g178 ( 
.A(n_159),
.Y(n_178)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_108),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_161),
.Y(n_179)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_SL g210 ( 
.A(n_167),
.B(n_170),
.C(n_177),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_148),
.A2(n_131),
.B(n_135),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_168),
.A2(n_174),
.B(n_183),
.Y(n_205)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

NAND3xp33_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_35),
.C(n_34),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_162),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_171),
.B(n_152),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_153),
.A2(n_122),
.B1(n_94),
.B2(n_78),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_173),
.A2(n_188),
.B1(n_160),
.B2(n_116),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_122),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_175),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_107),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_185),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_149),
.A2(n_114),
.B(n_95),
.Y(n_177)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_180),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_181),
.A2(n_160),
.B1(n_155),
.B2(n_150),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_182),
.A2(n_184),
.B1(n_186),
.B2(n_153),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_148),
.A2(n_81),
.B(n_34),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_154),
.A2(n_81),
.B(n_34),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_34),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_153),
.A2(n_116),
.B1(n_46),
.B2(n_47),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_149),
.B(n_35),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_137),
.Y(n_211)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_150),
.Y(n_189)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_189),
.Y(n_212)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_190),
.Y(n_233)
);

NOR2xp67_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_139),
.Y(n_191)
);

NOR3xp33_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_184),
.C(n_166),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_178),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_198),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_189),
.B(n_163),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_193),
.B(n_202),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_151),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_211),
.C(n_215),
.Y(n_217)
);

AND2x6_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_151),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_199),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_175),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_188),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_200),
.B(n_203),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_201),
.A2(n_188),
.B1(n_174),
.B2(n_172),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_164),
.B(n_163),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_179),
.B(n_138),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_153),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_204),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_205),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_147),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_209),
.A2(n_152),
.B(n_161),
.Y(n_227)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_186),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_213),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_214),
.A2(n_188),
.B1(n_185),
.B2(n_147),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_147),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_218),
.A2(n_221),
.B1(n_223),
.B2(n_228),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_187),
.C(n_183),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_224),
.C(n_229),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_168),
.C(n_188),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_197),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_225),
.B(n_232),
.Y(n_259)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_227),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_209),
.A2(n_159),
.B1(n_46),
.B2(n_45),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_211),
.C(n_208),
.Y(n_229)
);

MAJx2_ASAP7_75t_L g230 ( 
.A(n_196),
.B(n_81),
.C(n_27),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_230),
.B(n_27),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_206),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_239),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_212),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_236),
.B(n_85),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_199),
.Y(n_237)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_237),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_209),
.A2(n_45),
.B1(n_38),
.B2(n_41),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_238),
.A2(n_204),
.B1(n_85),
.B2(n_54),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_35),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_27),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_235),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_208),
.A2(n_200),
.B(n_192),
.Y(n_242)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_242),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_207),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_243),
.B(n_257),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_219),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_252),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_216),
.C(n_195),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_258),
.C(n_263),
.Y(n_266)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_251),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_233),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_222),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_253),
.B(n_264),
.Y(n_271)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_242),
.Y(n_254)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_254),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_255),
.A2(n_256),
.B1(n_228),
.B2(n_238),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_231),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_220),
.B(n_54),
.C(n_51),
.Y(n_258)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_261),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_262),
.B(n_265),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_28),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_224),
.B(n_51),
.C(n_47),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_28),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_250),
.A2(n_234),
.B(n_227),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_267),
.A2(n_280),
.B(n_5),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_246),
.A2(n_218),
.B1(n_230),
.B2(n_241),
.Y(n_268)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_268),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_226),
.Y(n_272)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_273),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_264),
.A2(n_223),
.B1(n_240),
.B2(n_4),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_284),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_259),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_283),
.Y(n_293)
);

FAx1_ASAP7_75t_SL g278 ( 
.A(n_257),
.B(n_28),
.CI(n_23),
.CON(n_278),
.SN(n_278)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_278),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_260),
.A2(n_2),
.B(n_3),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_262),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_282),
.Y(n_290)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_258),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_245),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_265),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_285),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_263),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_292),
.C(n_294),
.Y(n_306)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_289),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_248),
.C(n_245),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_243),
.C(n_244),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_244),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_297),
.C(n_47),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_6),
.Y(n_296)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_296),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_6),
.Y(n_297)
);

INVx13_ASAP7_75t_L g298 ( 
.A(n_271),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_291),
.Y(n_305)
);

OA21x2_ASAP7_75t_SL g301 ( 
.A1(n_269),
.A2(n_7),
.B(n_8),
.Y(n_301)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_301),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_293),
.A2(n_279),
.B(n_284),
.Y(n_303)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_303),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_281),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_304),
.B(n_308),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_305),
.B(n_307),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_290),
.A2(n_277),
.B(n_267),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_299),
.B(n_268),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_287),
.B(n_280),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_309),
.B(n_297),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_300),
.A2(n_274),
.B1(n_278),
.B2(n_270),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_311),
.C(n_312),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_286),
.B(n_270),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_7),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_47),
.C(n_45),
.Y(n_325)
);

BUFx24_ASAP7_75t_SL g315 ( 
.A(n_288),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_298),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_318),
.B(n_324),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_294),
.C(n_295),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_325),
.C(n_45),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_289),
.Y(n_321)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_321),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_322),
.B(n_327),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_312),
.A2(n_302),
.B(n_8),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_316),
.B(n_7),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_313),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_328),
.Y(n_334)
);

OAI21x1_ASAP7_75t_L g330 ( 
.A1(n_319),
.A2(n_306),
.B(n_314),
.Y(n_330)
);

AOI322xp5_ASAP7_75t_L g340 ( 
.A1(n_330),
.A2(n_332),
.A3(n_333),
.B1(n_10),
.B2(n_11),
.C1(n_12),
.C2(n_13),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_331),
.B(n_335),
.Y(n_342)
);

OA21x2_ASAP7_75t_SL g332 ( 
.A1(n_326),
.A2(n_9),
.B(n_10),
.Y(n_332)
);

AOI31xp67_ASAP7_75t_L g333 ( 
.A1(n_329),
.A2(n_9),
.A3(n_10),
.B(n_11),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_320),
.B(n_41),
.C(n_38),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_328),
.B(n_323),
.Y(n_339)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_339),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_340),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_336),
.B(n_337),
.Y(n_341)
);

AO21x1_ASAP7_75t_L g346 ( 
.A1(n_341),
.A2(n_343),
.B(n_344),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_334),
.B(n_12),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_336),
.B(n_37),
.Y(n_344)
);

OA21x2_ASAP7_75t_L g348 ( 
.A1(n_346),
.A2(n_342),
.B(n_37),
.Y(n_348)
);

BUFx24_ASAP7_75t_SL g349 ( 
.A(n_348),
.Y(n_349)
);

O2A1O1Ixp33_ASAP7_75t_SL g350 ( 
.A1(n_349),
.A2(n_347),
.B(n_345),
.C(n_38),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_350),
.A2(n_12),
.B(n_13),
.Y(n_351)
);

BUFx24_ASAP7_75t_SL g352 ( 
.A(n_351),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_352),
.B(n_41),
.C(n_15),
.Y(n_353)
);


endmodule