module fake_netlist_6_221_n_1786 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_507, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_396, n_495, n_350, n_78, n_84, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_542, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_338, n_522, n_466, n_506, n_56, n_360, n_119, n_235, n_536, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_516, n_153, n_525, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_472, n_270, n_239, n_126, n_414, n_97, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_552, n_216, n_455, n_83, n_521, n_363, n_395, n_323, n_393, n_411, n_503, n_152, n_92, n_513, n_321, n_331, n_105, n_227, n_132, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_481, n_325, n_329, n_464, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_546, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_514, n_528, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1786);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_507;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_542;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_119;
input n_235;
input n_536;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_552;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_481;
input n_325;
input n_329;
input n_464;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_546;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_514;
input n_528;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1786;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_1380;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_830;
wire n_873;
wire n_1285;
wire n_1371;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_699;
wire n_564;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_572;
wire n_813;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_608;
wire n_630;
wire n_792;
wire n_1328;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_1762;
wire n_1075;
wire n_932;
wire n_1697;
wire n_979;
wire n_905;
wire n_1680;
wire n_993;
wire n_689;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1563;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_1165;
wire n_702;
wire n_1175;
wire n_1386;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_593;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_1709;
wire n_1757;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_996;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_791;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_929;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_1358;
wire n_1388;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_811;
wire n_683;
wire n_1207;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1372;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1427;
wire n_1466;
wire n_1080;
wire n_723;
wire n_596;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_1060;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_1745;
wire n_914;
wire n_759;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_1617;
wire n_1470;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_1520;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_1731;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_607;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1095;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_923;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_1694;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_782;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_1361;
wire n_1491;
wire n_662;
wire n_1152;
wire n_1705;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_1222;
wire n_599;
wire n_776;
wire n_1720;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1341;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1640;
wire n_804;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_1522;
wire n_1782;
wire n_1676;
wire n_833;
wire n_1567;
wire n_1319;
wire n_707;
wire n_799;
wire n_1548;
wire n_1155;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_1047;
wire n_1385;
wire n_1269;
wire n_672;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1727;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_853;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1737;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_576;
wire n_1028;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_1276;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_1584;
wire n_924;
wire n_1582;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1525;
wire n_1585;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_570;
wire n_735;
wire n_1770;
wire n_878;
wire n_620;
wire n_1218;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_985;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_849;
wire n_753;
wire n_1753;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_1578;
wire n_1006;
wire n_1632;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_784;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_1423;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_1025;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_364),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_159),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_290),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_80),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_522),
.Y(n_558)
);

BUFx2_ASAP7_75t_L g559 ( 
.A(n_190),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_280),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_66),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_473),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_452),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_189),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_392),
.Y(n_565)
);

INVxp67_ASAP7_75t_L g566 ( 
.A(n_222),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_203),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_178),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_299),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_457),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_511),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_336),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_56),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_156),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_416),
.Y(n_575)
);

INVx1_ASAP7_75t_SL g576 ( 
.A(n_256),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_513),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_168),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_466),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_484),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_239),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_434),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_498),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_505),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_518),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_162),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_271),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_177),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_366),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_464),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_501),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_365),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_482),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_395),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_527),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_340),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_421),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_479),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_460),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_507),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_123),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_490),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_156),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_480),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_437),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_386),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_497),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_347),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_152),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_132),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_458),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_257),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_294),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_524),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_528),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g616 ( 
.A(n_519),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_220),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_523),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_38),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_459),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_521),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_94),
.Y(n_622)
);

BUFx2_ASAP7_75t_L g623 ( 
.A(n_305),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_491),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_422),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_176),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_432),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_60),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_462),
.Y(n_629)
);

BUFx2_ASAP7_75t_SL g630 ( 
.A(n_335),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_18),
.Y(n_631)
);

BUFx5_ASAP7_75t_L g632 ( 
.A(n_525),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_351),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_487),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_495),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_504),
.Y(n_636)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_515),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_526),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_461),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_485),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_81),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_536),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_446),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_488),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_163),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_481),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_492),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_475),
.Y(n_648)
);

CKINVDCx16_ASAP7_75t_R g649 ( 
.A(n_163),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_499),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_106),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_300),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_517),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_508),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_553),
.Y(n_655)
);

CKINVDCx20_ASAP7_75t_R g656 ( 
.A(n_201),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_407),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_181),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_357),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_516),
.Y(n_660)
);

INVx1_ASAP7_75t_SL g661 ( 
.A(n_334),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_467),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_250),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_136),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_530),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_502),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_368),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_39),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_496),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_209),
.Y(n_670)
);

CKINVDCx11_ASAP7_75t_R g671 ( 
.A(n_131),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_79),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_370),
.Y(n_673)
);

BUFx5_ASAP7_75t_L g674 ( 
.A(n_98),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_182),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_450),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_472),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_469),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_449),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_220),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_221),
.Y(n_681)
);

CKINVDCx14_ASAP7_75t_R g682 ( 
.A(n_90),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_213),
.Y(n_683)
);

INVx1_ASAP7_75t_SL g684 ( 
.A(n_73),
.Y(n_684)
);

BUFx10_ASAP7_75t_L g685 ( 
.A(n_39),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_483),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_486),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_403),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_387),
.Y(n_689)
);

INVx1_ASAP7_75t_SL g690 ( 
.A(n_242),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_444),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_198),
.Y(n_692)
);

BUFx2_ASAP7_75t_L g693 ( 
.A(n_188),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_388),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_344),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_232),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_330),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_493),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_11),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_128),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_248),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_234),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_509),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_552),
.Y(n_704)
);

HB1xp67_ASAP7_75t_L g705 ( 
.A(n_476),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_514),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_329),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_535),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_125),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_532),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_129),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_549),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_423),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_183),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_506),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_510),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_398),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_430),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_355),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_451),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_465),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_345),
.Y(n_722)
);

CKINVDCx14_ASAP7_75t_R g723 ( 
.A(n_477),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_207),
.Y(n_724)
);

CKINVDCx20_ASAP7_75t_R g725 ( 
.A(n_474),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_534),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_317),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_211),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_494),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_186),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_309),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_112),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_545),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_438),
.Y(n_734)
);

INVx1_ASAP7_75t_SL g735 ( 
.A(n_339),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_219),
.Y(n_736)
);

CKINVDCx20_ASAP7_75t_R g737 ( 
.A(n_203),
.Y(n_737)
);

INVxp67_ASAP7_75t_SL g738 ( 
.A(n_376),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_78),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_448),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_489),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_463),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_16),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_374),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_96),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_456),
.Y(n_746)
);

INVx1_ASAP7_75t_SL g747 ( 
.A(n_349),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_331),
.Y(n_748)
);

CKINVDCx20_ASAP7_75t_R g749 ( 
.A(n_93),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_533),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_236),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_324),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_417),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_144),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_216),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_89),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_426),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_503),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_128),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_167),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_478),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_249),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_5),
.Y(n_763)
);

CKINVDCx14_ASAP7_75t_R g764 ( 
.A(n_191),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_73),
.Y(n_765)
);

BUFx5_ASAP7_75t_L g766 ( 
.A(n_531),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_384),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_471),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_31),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_520),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_134),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_22),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_1),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_26),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_470),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_241),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_529),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_310),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_350),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_447),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_500),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_468),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_512),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_40),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_674),
.Y(n_785)
);

CKINVDCx16_ASAP7_75t_R g786 ( 
.A(n_649),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_674),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_591),
.B(n_1),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_671),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_559),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_623),
.B(n_2),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_674),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_554),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_674),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_556),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_674),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_711),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_572),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_711),
.Y(n_799)
);

CKINVDCx20_ASAP7_75t_R g800 ( 
.A(n_616),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_558),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_631),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_681),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_555),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_564),
.Y(n_805)
);

CKINVDCx20_ASAP7_75t_R g806 ( 
.A(n_620),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_610),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_622),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_621),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_628),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_797),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_799),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_785),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_792),
.Y(n_814)
);

OAI22xp5_ASAP7_75t_L g815 ( 
.A1(n_790),
.A2(n_764),
.B1(n_682),
.B2(n_723),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_787),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_794),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_796),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_802),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_804),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_805),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_807),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_793),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_808),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_810),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_803),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_786),
.B(n_638),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_795),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_801),
.B(n_624),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_788),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_789),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_791),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_798),
.Y(n_833)
);

BUFx8_ASAP7_75t_L g834 ( 
.A(n_800),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_806),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_809),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_823),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_830),
.B(n_641),
.Y(n_838)
);

BUFx3_ASAP7_75t_L g839 ( 
.A(n_833),
.Y(n_839)
);

BUFx4f_ASAP7_75t_L g840 ( 
.A(n_833),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_820),
.Y(n_841)
);

OAI22xp33_ASAP7_75t_L g842 ( 
.A1(n_832),
.A2(n_693),
.B1(n_684),
.B2(n_690),
.Y(n_842)
);

AOI22xp5_ASAP7_75t_L g843 ( 
.A1(n_815),
.A2(n_697),
.B1(n_725),
.B2(n_666),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_814),
.Y(n_844)
);

NAND3xp33_ASAP7_75t_L g845 ( 
.A(n_826),
.B(n_705),
.C(n_597),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_821),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_813),
.B(n_650),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_824),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_828),
.B(n_637),
.Y(n_849)
);

INVx4_ASAP7_75t_L g850 ( 
.A(n_831),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_825),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_827),
.B(n_661),
.Y(n_852)
);

AO22x2_ASAP7_75t_L g853 ( 
.A1(n_836),
.A2(n_576),
.B1(n_573),
.B2(n_668),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_817),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_818),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_816),
.B(n_673),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_822),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_834),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_811),
.Y(n_859)
);

AND2x6_ASAP7_75t_L g860 ( 
.A(n_819),
.B(n_607),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_812),
.B(n_735),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_812),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_835),
.Y(n_863)
);

OR2x2_ASAP7_75t_L g864 ( 
.A(n_834),
.B(n_566),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_820),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_814),
.Y(n_866)
);

INVx5_ASAP7_75t_L g867 ( 
.A(n_822),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_829),
.B(n_747),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_829),
.Y(n_869)
);

OR2x6_ASAP7_75t_L g870 ( 
.A(n_833),
.B(n_675),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_820),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_822),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_844),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_841),
.Y(n_874)
);

AO22x2_ASAP7_75t_L g875 ( 
.A1(n_845),
.A2(n_692),
.B1(n_699),
.B2(n_683),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_846),
.Y(n_876)
);

OAI221xp5_ASAP7_75t_L g877 ( 
.A1(n_852),
.A2(n_728),
.B1(n_771),
.B2(n_762),
.C(n_739),
.Y(n_877)
);

NAND2x1p5_ASAP7_75t_L g878 ( 
.A(n_850),
.B(n_677),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_848),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_851),
.Y(n_880)
);

BUFx8_ASAP7_75t_L g881 ( 
.A(n_839),
.Y(n_881)
);

AO22x2_ASAP7_75t_L g882 ( 
.A1(n_863),
.A2(n_776),
.B1(n_672),
.B2(n_680),
.Y(n_882)
);

NAND2xp33_ASAP7_75t_L g883 ( 
.A(n_869),
.B(n_562),
.Y(n_883)
);

INVxp67_ASAP7_75t_L g884 ( 
.A(n_849),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_865),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_868),
.B(n_738),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_857),
.B(n_740),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_871),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_854),
.B(n_563),
.Y(n_889)
);

NOR2xp67_ASAP7_75t_L g890 ( 
.A(n_837),
.B(n_843),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_859),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_840),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_862),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_855),
.Y(n_894)
);

OR2x6_ASAP7_75t_L g895 ( 
.A(n_870),
.B(n_864),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_866),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_872),
.B(n_565),
.Y(n_897)
);

AO22x2_ASAP7_75t_L g898 ( 
.A1(n_842),
.A2(n_571),
.B1(n_579),
.B2(n_577),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_872),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_861),
.Y(n_900)
);

INVxp67_ASAP7_75t_L g901 ( 
.A(n_853),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_856),
.Y(n_902)
);

AO22x2_ASAP7_75t_L g903 ( 
.A1(n_847),
.A2(n_595),
.B1(n_596),
.B2(n_590),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_867),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_860),
.Y(n_905)
);

INVxp67_ASAP7_75t_L g906 ( 
.A(n_860),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_841),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_868),
.B(n_557),
.Y(n_908)
);

AO22x2_ASAP7_75t_L g909 ( 
.A1(n_845),
.A2(n_602),
.B1(n_605),
.B2(n_598),
.Y(n_909)
);

CKINVDCx14_ASAP7_75t_R g910 ( 
.A(n_858),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_839),
.B(n_719),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_844),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_839),
.B(n_729),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_841),
.Y(n_914)
);

AO22x2_ASAP7_75t_L g915 ( 
.A1(n_845),
.A2(n_613),
.B1(n_615),
.B2(n_611),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_841),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_841),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_869),
.B(n_775),
.Y(n_918)
);

AO22x2_ASAP7_75t_L g919 ( 
.A1(n_845),
.A2(n_625),
.B1(n_627),
.B2(n_618),
.Y(n_919)
);

OAI221xp5_ASAP7_75t_L g920 ( 
.A1(n_852),
.A2(n_629),
.B1(n_691),
.B2(n_660),
.C(n_646),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_841),
.Y(n_921)
);

NAND3xp33_ASAP7_75t_L g922 ( 
.A(n_852),
.B(n_567),
.C(n_561),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_838),
.B(n_685),
.Y(n_923)
);

BUFx8_ASAP7_75t_L g924 ( 
.A(n_839),
.Y(n_924)
);

AOI22x1_ASAP7_75t_L g925 ( 
.A1(n_841),
.A2(n_582),
.B1(n_589),
.B2(n_560),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_841),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_839),
.B(n_634),
.Y(n_927)
);

INVx2_ASAP7_75t_SL g928 ( 
.A(n_870),
.Y(n_928)
);

OR2x2_ASAP7_75t_SL g929 ( 
.A(n_845),
.B(n_656),
.Y(n_929)
);

INVxp67_ASAP7_75t_L g930 ( 
.A(n_852),
.Y(n_930)
);

OAI221xp5_ASAP7_75t_L g931 ( 
.A1(n_852),
.A2(n_722),
.B1(n_734),
.B2(n_698),
.C(n_679),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_837),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_841),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_841),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_841),
.Y(n_935)
);

AO22x2_ASAP7_75t_L g936 ( 
.A1(n_845),
.A2(n_635),
.B1(n_639),
.B2(n_636),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_868),
.B(n_644),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_839),
.B(n_647),
.Y(n_938)
);

AO22x2_ASAP7_75t_L g939 ( 
.A1(n_845),
.A2(n_652),
.B1(n_665),
.B2(n_659),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_872),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_841),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_868),
.B(n_703),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_841),
.Y(n_943)
);

INVxp67_ASAP7_75t_L g944 ( 
.A(n_852),
.Y(n_944)
);

BUFx8_ASAP7_75t_L g945 ( 
.A(n_839),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_841),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_841),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_884),
.B(n_706),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_930),
.B(n_569),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_900),
.B(n_715),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_944),
.B(n_570),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_908),
.B(n_575),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_886),
.B(n_580),
.Y(n_953)
);

NAND2xp33_ASAP7_75t_L g954 ( 
.A(n_937),
.B(n_632),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_942),
.B(n_583),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_890),
.B(n_584),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_902),
.B(n_585),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_892),
.B(n_587),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_876),
.B(n_592),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_879),
.B(n_718),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_880),
.B(n_885),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_888),
.B(n_726),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_891),
.B(n_593),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_923),
.B(n_568),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_894),
.B(n_594),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_907),
.B(n_599),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_914),
.B(n_727),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_916),
.B(n_731),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_917),
.B(n_600),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_921),
.B(n_604),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_926),
.B(n_741),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_933),
.B(n_606),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_934),
.B(n_608),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_935),
.B(n_753),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_941),
.B(n_614),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_943),
.B(n_758),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_946),
.B(n_640),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_947),
.B(n_642),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_922),
.B(n_643),
.Y(n_979)
);

NAND2xp33_ASAP7_75t_SL g980 ( 
.A(n_932),
.B(n_663),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_928),
.B(n_648),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_893),
.B(n_761),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_873),
.B(n_767),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_896),
.B(n_653),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_912),
.B(n_654),
.Y(n_985)
);

NAND2xp33_ASAP7_75t_SL g986 ( 
.A(n_918),
.B(n_737),
.Y(n_986)
);

NAND2xp33_ASAP7_75t_SL g987 ( 
.A(n_905),
.B(n_749),
.Y(n_987)
);

NAND2xp33_ASAP7_75t_SL g988 ( 
.A(n_904),
.B(n_897),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_927),
.B(n_938),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_889),
.B(n_778),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_883),
.B(n_782),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_887),
.B(n_574),
.Y(n_992)
);

NAND2xp33_ASAP7_75t_SL g993 ( 
.A(n_940),
.B(n_667),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_911),
.B(n_669),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_899),
.B(n_657),
.Y(n_995)
);

NAND2xp33_ASAP7_75t_SL g996 ( 
.A(n_913),
.B(n_676),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_878),
.B(n_678),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_906),
.B(n_686),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_901),
.B(n_687),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_895),
.B(n_270),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_898),
.B(n_882),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_895),
.B(n_272),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_881),
.B(n_688),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_924),
.B(n_689),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_945),
.B(n_694),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_925),
.B(n_695),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_909),
.B(n_273),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_929),
.B(n_704),
.Y(n_1008)
);

NAND2xp33_ASAP7_75t_SL g1009 ( 
.A(n_915),
.B(n_707),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_920),
.B(n_708),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_919),
.B(n_710),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_931),
.B(n_712),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_936),
.B(n_713),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_939),
.B(n_716),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_903),
.B(n_717),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_877),
.B(n_720),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_875),
.B(n_721),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_910),
.B(n_733),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_930),
.B(n_742),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_930),
.B(n_744),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_884),
.B(n_746),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_930),
.B(n_748),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_930),
.B(n_750),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_930),
.B(n_752),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_884),
.B(n_578),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_930),
.B(n_768),
.Y(n_1026)
);

NAND2xp33_ASAP7_75t_SL g1027 ( 
.A(n_892),
.B(n_777),
.Y(n_1027)
);

AND2x4_ASAP7_75t_L g1028 ( 
.A(n_874),
.B(n_274),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_930),
.B(n_779),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_930),
.B(n_780),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_930),
.B(n_781),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_930),
.B(n_783),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_930),
.B(n_607),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_884),
.B(n_630),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_930),
.B(n_757),
.Y(n_1035)
);

AND2x4_ASAP7_75t_L g1036 ( 
.A(n_874),
.B(n_275),
.Y(n_1036)
);

NAND2xp33_ASAP7_75t_SL g1037 ( 
.A(n_892),
.B(n_581),
.Y(n_1037)
);

NAND2xp33_ASAP7_75t_SL g1038 ( 
.A(n_892),
.B(n_586),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_930),
.B(n_633),
.Y(n_1039)
);

NAND2xp33_ASAP7_75t_SL g1040 ( 
.A(n_892),
.B(n_588),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_930),
.B(n_633),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_884),
.B(n_601),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_930),
.B(n_633),
.Y(n_1043)
);

NAND2xp33_ASAP7_75t_SL g1044 ( 
.A(n_892),
.B(n_603),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_930),
.B(n_655),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_884),
.B(n_632),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_930),
.B(n_655),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_884),
.B(n_632),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_884),
.B(n_766),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_930),
.B(n_655),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_930),
.B(n_662),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_930),
.B(n_662),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_884),
.B(n_766),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_930),
.B(n_662),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_884),
.B(n_766),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_884),
.B(n_609),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_930),
.B(n_757),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_930),
.B(n_770),
.Y(n_1058)
);

NAND2xp33_ASAP7_75t_SL g1059 ( 
.A(n_892),
.B(n_612),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_930),
.B(n_770),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_930),
.B(n_770),
.Y(n_1061)
);

NAND2xp33_ASAP7_75t_SL g1062 ( 
.A(n_892),
.B(n_617),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_884),
.B(n_766),
.Y(n_1063)
);

NAND2xp33_ASAP7_75t_SL g1064 ( 
.A(n_892),
.B(n_619),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_930),
.B(n_766),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_884),
.B(n_626),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_961),
.Y(n_1067)
);

INVx2_ASAP7_75t_SL g1068 ( 
.A(n_995),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_986),
.A2(n_651),
.B(n_658),
.C(n_645),
.Y(n_1069)
);

AOI21x1_ASAP7_75t_L g1070 ( 
.A1(n_1065),
.A2(n_277),
.B(n_276),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_983),
.Y(n_1071)
);

OAI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_950),
.A2(n_670),
.B(n_664),
.Y(n_1072)
);

AND2x6_ASAP7_75t_L g1073 ( 
.A(n_1007),
.B(n_278),
.Y(n_1073)
);

INVx3_ASAP7_75t_L g1074 ( 
.A(n_995),
.Y(n_1074)
);

AND2x4_ASAP7_75t_L g1075 ( 
.A(n_989),
.B(n_279),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_1034),
.B(n_696),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_1000),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_982),
.A2(n_282),
.B(n_281),
.Y(n_1078)
);

OAI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_1046),
.A2(n_701),
.B(n_700),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_948),
.B(n_702),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_1048),
.A2(n_714),
.B(n_709),
.Y(n_1081)
);

AO31x2_ASAP7_75t_L g1082 ( 
.A1(n_991),
.A2(n_284),
.A3(n_285),
.B(n_283),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_962),
.Y(n_1083)
);

AO31x2_ASAP7_75t_L g1084 ( 
.A1(n_1049),
.A2(n_287),
.A3(n_288),
.B(n_286),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1025),
.B(n_724),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1042),
.B(n_730),
.Y(n_1086)
);

OAI21x1_ASAP7_75t_L g1087 ( 
.A1(n_967),
.A2(n_291),
.B(n_289),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_968),
.A2(n_293),
.B(n_292),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_960),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_1021),
.B(n_732),
.Y(n_1090)
);

INVx2_ASAP7_75t_SL g1091 ( 
.A(n_992),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_1028),
.Y(n_1092)
);

AO32x2_ASAP7_75t_L g1093 ( 
.A1(n_1001),
.A2(n_3),
.A3(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_1093)
);

O2A1O1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_1066),
.A2(n_743),
.B(n_745),
.C(n_736),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_1000),
.Y(n_1095)
);

AOI21xp33_ASAP7_75t_L g1096 ( 
.A1(n_952),
.A2(n_754),
.B(n_751),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_971),
.A2(n_296),
.B(n_295),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1056),
.B(n_755),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_957),
.A2(n_298),
.B(n_297),
.Y(n_1099)
);

AO31x2_ASAP7_75t_L g1100 ( 
.A1(n_1053),
.A2(n_550),
.A3(n_551),
.B(n_548),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_974),
.Y(n_1101)
);

INVx1_ASAP7_75t_SL g1102 ( 
.A(n_980),
.Y(n_1102)
);

AO21x2_ASAP7_75t_L g1103 ( 
.A1(n_1055),
.A2(n_302),
.B(n_301),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_960),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_1006),
.A2(n_304),
.B(n_303),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_1036),
.A2(n_759),
.B1(n_760),
.B2(n_756),
.Y(n_1106)
);

INVx2_ASAP7_75t_SL g1107 ( 
.A(n_1002),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_949),
.B(n_763),
.Y(n_1108)
);

AO31x2_ASAP7_75t_L g1109 ( 
.A1(n_1063),
.A2(n_307),
.A3(n_308),
.B(n_306),
.Y(n_1109)
);

AOI21x1_ASAP7_75t_L g1110 ( 
.A1(n_990),
.A2(n_312),
.B(n_311),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_964),
.B(n_765),
.Y(n_1111)
);

INVxp67_ASAP7_75t_L g1112 ( 
.A(n_999),
.Y(n_1112)
);

AO31x2_ASAP7_75t_L g1113 ( 
.A1(n_1011),
.A2(n_546),
.A3(n_547),
.B(n_544),
.Y(n_1113)
);

AOI21x1_ASAP7_75t_L g1114 ( 
.A1(n_979),
.A2(n_314),
.B(n_313),
.Y(n_1114)
);

AOI21xp33_ASAP7_75t_L g1115 ( 
.A1(n_953),
.A2(n_772),
.B(n_769),
.Y(n_1115)
);

INVx3_ASAP7_75t_L g1116 ( 
.A(n_1036),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_976),
.Y(n_1117)
);

AOI211x1_ASAP7_75t_L g1118 ( 
.A1(n_1015),
.A2(n_774),
.B(n_784),
.C(n_773),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_976),
.B(n_0),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_1002),
.Y(n_1120)
);

AOI21xp33_ASAP7_75t_L g1121 ( 
.A1(n_1017),
.A2(n_4),
.B(n_5),
.Y(n_1121)
);

OAI22x1_ASAP7_75t_L g1122 ( 
.A1(n_1007),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_955),
.B(n_6),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_984),
.A2(n_316),
.B(n_315),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_998),
.A2(n_319),
.B1(n_320),
.B2(n_318),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_959),
.A2(n_322),
.B(n_321),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_985),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_987),
.B(n_323),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_951),
.B(n_9),
.Y(n_1129)
);

INVxp67_ASAP7_75t_L g1130 ( 
.A(n_1037),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_SL g1131 ( 
.A1(n_997),
.A2(n_326),
.B(n_325),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_981),
.B(n_327),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1019),
.B(n_9),
.Y(n_1133)
);

A2O1A1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_1009),
.A2(n_12),
.B(n_10),
.C(n_11),
.Y(n_1134)
);

BUFx3_ASAP7_75t_L g1135 ( 
.A(n_1038),
.Y(n_1135)
);

O2A1O1Ixp5_ASAP7_75t_L g1136 ( 
.A1(n_1033),
.A2(n_540),
.B(n_541),
.C(n_539),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_1008),
.A2(n_13),
.B(n_10),
.C(n_12),
.Y(n_1137)
);

HB1xp67_ASAP7_75t_L g1138 ( 
.A(n_1013),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_963),
.A2(n_332),
.B(n_328),
.Y(n_1139)
);

BUFx2_ASAP7_75t_L g1140 ( 
.A(n_1040),
.Y(n_1140)
);

AND3x2_ASAP7_75t_L g1141 ( 
.A(n_1044),
.B(n_14),
.C(n_15),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1020),
.B(n_15),
.Y(n_1142)
);

NOR2xp67_ASAP7_75t_L g1143 ( 
.A(n_956),
.B(n_333),
.Y(n_1143)
);

BUFx12f_ASAP7_75t_L g1144 ( 
.A(n_1059),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_1022),
.B(n_16),
.Y(n_1145)
);

INVx4_ASAP7_75t_L g1146 ( 
.A(n_988),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1023),
.B(n_17),
.Y(n_1147)
);

A2O1A1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_965),
.A2(n_966),
.B(n_970),
.C(n_969),
.Y(n_1148)
);

OA21x2_ASAP7_75t_L g1149 ( 
.A1(n_972),
.A2(n_338),
.B(n_337),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_954),
.Y(n_1150)
);

O2A1O1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1014),
.A2(n_20),
.B(n_18),
.C(n_19),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_973),
.A2(n_342),
.B(n_341),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1035),
.Y(n_1153)
);

AO21x2_ASAP7_75t_L g1154 ( 
.A1(n_975),
.A2(n_346),
.B(n_343),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_1024),
.B(n_348),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1039),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1026),
.B(n_20),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1029),
.B(n_21),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_994),
.B(n_352),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1067),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_1112),
.B(n_1030),
.Y(n_1161)
);

OA21x2_ASAP7_75t_L g1162 ( 
.A1(n_1150),
.A2(n_1043),
.B(n_1041),
.Y(n_1162)
);

OR2x6_ASAP7_75t_L g1163 ( 
.A(n_1077),
.B(n_1003),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_L g1164 ( 
.A1(n_1145),
.A2(n_1016),
.B1(n_1012),
.B2(n_1010),
.Y(n_1164)
);

AO32x2_ASAP7_75t_L g1165 ( 
.A1(n_1146),
.A2(n_1047),
.A3(n_1051),
.B1(n_1050),
.B2(n_1045),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1105),
.A2(n_978),
.B(n_977),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_1083),
.B(n_1031),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_L g1168 ( 
.A1(n_1108),
.A2(n_1032),
.B1(n_958),
.B2(n_996),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_1124),
.A2(n_1054),
.B(n_1052),
.Y(n_1169)
);

AO32x2_ASAP7_75t_L g1170 ( 
.A1(n_1106),
.A2(n_1060),
.A3(n_1061),
.B1(n_1058),
.B2(n_1057),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1101),
.Y(n_1171)
);

INVxp67_ASAP7_75t_SL g1172 ( 
.A(n_1092),
.Y(n_1172)
);

OR2x2_ASAP7_75t_L g1173 ( 
.A(n_1085),
.B(n_1018),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1089),
.Y(n_1174)
);

INVx3_ASAP7_75t_L g1175 ( 
.A(n_1077),
.Y(n_1175)
);

OR2x6_ASAP7_75t_L g1176 ( 
.A(n_1095),
.B(n_1004),
.Y(n_1176)
);

AO31x2_ASAP7_75t_L g1177 ( 
.A1(n_1134),
.A2(n_993),
.A3(n_1027),
.B(n_1062),
.Y(n_1177)
);

OAI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_1116),
.A2(n_1005),
.B1(n_1064),
.B2(n_23),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_1095),
.Y(n_1179)
);

OAI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1071),
.A2(n_354),
.B(n_353),
.Y(n_1180)
);

OAI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1148),
.A2(n_358),
.B(n_356),
.Y(n_1181)
);

INVx1_ASAP7_75t_SL g1182 ( 
.A(n_1138),
.Y(n_1182)
);

INVx1_ASAP7_75t_SL g1183 ( 
.A(n_1120),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1104),
.Y(n_1184)
);

OR2x2_ASAP7_75t_L g1185 ( 
.A(n_1086),
.B(n_21),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1117),
.Y(n_1186)
);

NAND2x1p5_ASAP7_75t_L g1187 ( 
.A(n_1120),
.B(n_363),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1107),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_1102),
.B(n_24),
.Y(n_1189)
);

AOI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1114),
.A2(n_360),
.B(n_359),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1127),
.Y(n_1191)
);

AOI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1110),
.A2(n_362),
.B(n_361),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1119),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_1068),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1153),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1070),
.Y(n_1196)
);

BUFx4_ASAP7_75t_R g1197 ( 
.A(n_1135),
.Y(n_1197)
);

OA21x2_ASAP7_75t_L g1198 ( 
.A1(n_1078),
.A2(n_1088),
.B(n_1087),
.Y(n_1198)
);

HB1xp67_ASAP7_75t_L g1199 ( 
.A(n_1074),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_1144),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1156),
.Y(n_1201)
);

OAI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1080),
.A2(n_369),
.B(n_367),
.Y(n_1202)
);

AOI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1073),
.A2(n_1130),
.B1(n_1075),
.B2(n_1159),
.Y(n_1203)
);

AOI222xp33_ASAP7_75t_L g1204 ( 
.A1(n_1122),
.A2(n_27),
.B1(n_29),
.B2(n_25),
.C1(n_26),
.C2(n_28),
.Y(n_1204)
);

OR2x6_ASAP7_75t_L g1205 ( 
.A(n_1140),
.B(n_371),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1098),
.B(n_25),
.Y(n_1206)
);

OA21x2_ASAP7_75t_L g1207 ( 
.A1(n_1097),
.A2(n_373),
.B(n_372),
.Y(n_1207)
);

BUFx2_ASAP7_75t_L g1208 ( 
.A(n_1073),
.Y(n_1208)
);

BUFx2_ASAP7_75t_L g1209 ( 
.A(n_1073),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1149),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1103),
.Y(n_1211)
);

HB1xp67_ASAP7_75t_L g1212 ( 
.A(n_1129),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1133),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1111),
.B(n_30),
.Y(n_1214)
);

AOI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1128),
.A2(n_377),
.B(n_375),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1076),
.A2(n_379),
.B(n_378),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_1132),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1142),
.Y(n_1218)
);

OAI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1090),
.A2(n_381),
.B(n_380),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1154),
.Y(n_1220)
);

AO31x2_ASAP7_75t_L g1221 ( 
.A1(n_1125),
.A2(n_383),
.A3(n_385),
.B(n_382),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1118),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_1222)
);

OA21x2_ASAP7_75t_L g1223 ( 
.A1(n_1136),
.A2(n_390),
.B(n_389),
.Y(n_1223)
);

A2O1A1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1094),
.A2(n_34),
.B(n_32),
.C(n_33),
.Y(n_1224)
);

AO21x2_ASAP7_75t_L g1225 ( 
.A1(n_1155),
.A2(n_393),
.B(n_391),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1072),
.B(n_33),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1099),
.A2(n_1139),
.B(n_1126),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1079),
.B(n_34),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1152),
.A2(n_396),
.B(n_394),
.Y(n_1229)
);

AO31x2_ASAP7_75t_L g1230 ( 
.A1(n_1069),
.A2(n_399),
.A3(n_400),
.B(n_397),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1147),
.Y(n_1231)
);

CKINVDCx8_ASAP7_75t_R g1232 ( 
.A(n_1141),
.Y(n_1232)
);

OA21x2_ASAP7_75t_L g1233 ( 
.A1(n_1123),
.A2(n_402),
.B(n_401),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1131),
.A2(n_405),
.B(n_404),
.Y(n_1234)
);

AO31x2_ASAP7_75t_L g1235 ( 
.A1(n_1157),
.A2(n_408),
.A3(n_409),
.B(n_406),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_1096),
.B(n_1158),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1151),
.A2(n_411),
.B(n_410),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1081),
.B(n_35),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1137),
.A2(n_413),
.B(n_412),
.Y(n_1239)
);

INVx4_ASAP7_75t_L g1240 ( 
.A(n_1143),
.Y(n_1240)
);

OA21x2_ASAP7_75t_L g1241 ( 
.A1(n_1121),
.A2(n_415),
.B(n_414),
.Y(n_1241)
);

CKINVDCx11_ASAP7_75t_R g1242 ( 
.A(n_1113),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_SL g1243 ( 
.A1(n_1093),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_1243)
);

OAI33xp33_ASAP7_75t_L g1244 ( 
.A1(n_1115),
.A2(n_38),
.A3(n_41),
.B1(n_36),
.B2(n_37),
.B3(n_40),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1113),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1084),
.Y(n_1246)
);

OAI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1084),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_1247)
);

OR2x6_ASAP7_75t_L g1248 ( 
.A(n_1100),
.B(n_418),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1082),
.A2(n_420),
.B(n_419),
.Y(n_1249)
);

BUFx10_ASAP7_75t_L g1250 ( 
.A(n_1109),
.Y(n_1250)
);

BUFx3_ASAP7_75t_L g1251 ( 
.A(n_1091),
.Y(n_1251)
);

OAI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1083),
.A2(n_425),
.B(n_424),
.Y(n_1252)
);

NAND2x1p5_ASAP7_75t_L g1253 ( 
.A(n_1077),
.B(n_427),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1077),
.Y(n_1254)
);

BUFx2_ASAP7_75t_L g1255 ( 
.A(n_1251),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1171),
.Y(n_1256)
);

CKINVDCx11_ASAP7_75t_R g1257 ( 
.A(n_1200),
.Y(n_1257)
);

INVx1_ASAP7_75t_SL g1258 ( 
.A(n_1197),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1160),
.Y(n_1259)
);

BUFx2_ASAP7_75t_L g1260 ( 
.A(n_1217),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1203),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1191),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1195),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1201),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1212),
.B(n_45),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1227),
.A2(n_429),
.B(n_428),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1193),
.B(n_47),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1214),
.B(n_47),
.Y(n_1268)
);

OR2x2_ASAP7_75t_L g1269 ( 
.A(n_1213),
.B(n_48),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1174),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_1194),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1182),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1184),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1186),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1181),
.A2(n_543),
.B(n_542),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1218),
.Y(n_1276)
);

OR2x2_ASAP7_75t_L g1277 ( 
.A(n_1231),
.B(n_48),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1206),
.Y(n_1278)
);

BUFx2_ASAP7_75t_L g1279 ( 
.A(n_1179),
.Y(n_1279)
);

OR2x2_ASAP7_75t_L g1280 ( 
.A(n_1185),
.B(n_49),
.Y(n_1280)
);

INVx3_ASAP7_75t_L g1281 ( 
.A(n_1254),
.Y(n_1281)
);

AND2x4_ASAP7_75t_L g1282 ( 
.A(n_1175),
.B(n_431),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1199),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1254),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1226),
.Y(n_1285)
);

INVx3_ASAP7_75t_L g1286 ( 
.A(n_1240),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_SL g1287 ( 
.A1(n_1236),
.A2(n_57),
.B1(n_65),
.B2(n_49),
.Y(n_1287)
);

AND2x4_ASAP7_75t_L g1288 ( 
.A(n_1183),
.B(n_433),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1167),
.B(n_50),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1162),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1246),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1205),
.B(n_50),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1228),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1238),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1196),
.Y(n_1295)
);

OAI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1164),
.A2(n_51),
.B(n_52),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1172),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1235),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1235),
.Y(n_1299)
);

OAI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1205),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_1300)
);

HB1xp67_ASAP7_75t_L g1301 ( 
.A(n_1163),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1190),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1165),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1189),
.B(n_53),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1208),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1161),
.B(n_54),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1209),
.Y(n_1307)
);

INVx3_ASAP7_75t_L g1308 ( 
.A(n_1187),
.Y(n_1308)
);

NOR2x1_ASAP7_75t_R g1309 ( 
.A(n_1200),
.B(n_435),
.Y(n_1309)
);

HB1xp67_ASAP7_75t_L g1310 ( 
.A(n_1163),
.Y(n_1310)
);

INVx2_ASAP7_75t_SL g1311 ( 
.A(n_1176),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1173),
.B(n_1232),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1233),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1166),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1202),
.A2(n_538),
.B(n_537),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1250),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1263),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1264),
.Y(n_1318)
);

OR2x6_ASAP7_75t_L g1319 ( 
.A(n_1311),
.B(n_1253),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_R g1320 ( 
.A(n_1257),
.B(n_1242),
.Y(n_1320)
);

BUFx8_ASAP7_75t_SL g1321 ( 
.A(n_1279),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1289),
.B(n_1224),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_R g1323 ( 
.A(n_1308),
.B(n_1215),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_R g1324 ( 
.A(n_1308),
.B(n_1168),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1285),
.B(n_1204),
.Y(n_1325)
);

NAND2xp33_ASAP7_75t_R g1326 ( 
.A(n_1255),
.B(n_1241),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1258),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1293),
.B(n_1243),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1270),
.Y(n_1329)
);

AND2x4_ASAP7_75t_L g1330 ( 
.A(n_1260),
.B(n_1177),
.Y(n_1330)
);

XNOR2xp5_ASAP7_75t_L g1331 ( 
.A(n_1301),
.B(n_1310),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1262),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1284),
.B(n_1177),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1294),
.B(n_1222),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_1278),
.B(n_1178),
.Y(n_1335)
);

NAND2xp33_ASAP7_75t_R g1336 ( 
.A(n_1312),
.B(n_1207),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1272),
.B(n_1234),
.Y(n_1337)
);

INVxp67_ASAP7_75t_L g1338 ( 
.A(n_1271),
.Y(n_1338)
);

BUFx3_ASAP7_75t_L g1339 ( 
.A(n_1281),
.Y(n_1339)
);

AND2x4_ASAP7_75t_L g1340 ( 
.A(n_1281),
.B(n_1225),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1273),
.Y(n_1341)
);

BUFx3_ASAP7_75t_L g1342 ( 
.A(n_1283),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_R g1343 ( 
.A(n_1286),
.B(n_1192),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1306),
.B(n_1170),
.Y(n_1344)
);

NAND2xp33_ASAP7_75t_R g1345 ( 
.A(n_1288),
.B(n_1248),
.Y(n_1345)
);

NAND2xp33_ASAP7_75t_R g1346 ( 
.A(n_1288),
.B(n_1248),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1305),
.B(n_1230),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1259),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1256),
.Y(n_1349)
);

AND2x4_ASAP7_75t_L g1350 ( 
.A(n_1307),
.B(n_1230),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1268),
.B(n_1244),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1292),
.B(n_1188),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1282),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1267),
.B(n_1170),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_SL g1355 ( 
.A1(n_1335),
.A2(n_1296),
.B(n_1275),
.Y(n_1355)
);

OAI222xp33_ASAP7_75t_L g1356 ( 
.A1(n_1325),
.A2(n_1287),
.B1(n_1261),
.B2(n_1300),
.C1(n_1322),
.C2(n_1328),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1348),
.Y(n_1357)
);

BUFx2_ASAP7_75t_L g1358 ( 
.A(n_1321),
.Y(n_1358)
);

BUFx2_ASAP7_75t_L g1359 ( 
.A(n_1342),
.Y(n_1359)
);

INVx3_ASAP7_75t_L g1360 ( 
.A(n_1333),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1349),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1344),
.B(n_1265),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1354),
.B(n_1276),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1338),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_SL g1365 ( 
.A(n_1324),
.B(n_1297),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1317),
.Y(n_1366)
);

INVxp67_ASAP7_75t_L g1367 ( 
.A(n_1339),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1318),
.B(n_1304),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1329),
.Y(n_1369)
);

AOI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1345),
.A2(n_1315),
.B1(n_1219),
.B2(n_1282),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1320),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1341),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1332),
.B(n_1303),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1347),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1351),
.B(n_1274),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1350),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1330),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1331),
.Y(n_1378)
);

AND2x4_ASAP7_75t_L g1379 ( 
.A(n_1337),
.B(n_1316),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1326),
.Y(n_1380)
);

AOI221xp5_ASAP7_75t_L g1381 ( 
.A1(n_1352),
.A2(n_1247),
.B1(n_1245),
.B2(n_1280),
.C(n_1277),
.Y(n_1381)
);

OR2x2_ASAP7_75t_SL g1382 ( 
.A(n_1334),
.B(n_1269),
.Y(n_1382)
);

BUFx3_ASAP7_75t_L g1383 ( 
.A(n_1327),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1340),
.Y(n_1384)
);

OAI221xp5_ASAP7_75t_L g1385 ( 
.A1(n_1346),
.A2(n_1216),
.B1(n_1252),
.B2(n_1180),
.C(n_1249),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1353),
.B(n_1298),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1343),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1323),
.Y(n_1388)
);

HB1xp67_ASAP7_75t_L g1389 ( 
.A(n_1336),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1319),
.B(n_1295),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1319),
.B(n_1291),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1359),
.B(n_1299),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1372),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1372),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1366),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1362),
.B(n_1290),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1357),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1383),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1364),
.B(n_1291),
.Y(n_1399)
);

INVx2_ASAP7_75t_SL g1400 ( 
.A(n_1358),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1361),
.Y(n_1401)
);

BUFx2_ASAP7_75t_L g1402 ( 
.A(n_1380),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1369),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1373),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1391),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1363),
.B(n_1314),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1389),
.B(n_1313),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1374),
.Y(n_1408)
);

BUFx2_ASAP7_75t_L g1409 ( 
.A(n_1379),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1376),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1384),
.B(n_1302),
.Y(n_1411)
);

NAND2xp33_ASAP7_75t_SL g1412 ( 
.A(n_1371),
.B(n_1365),
.Y(n_1412)
);

OR2x2_ASAP7_75t_L g1413 ( 
.A(n_1382),
.B(n_1211),
.Y(n_1413)
);

OAI221xp5_ASAP7_75t_SL g1414 ( 
.A1(n_1355),
.A2(n_1309),
.B1(n_1220),
.B2(n_57),
.C(n_59),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1390),
.Y(n_1415)
);

INVx1_ASAP7_75t_SL g1416 ( 
.A(n_1378),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1377),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_SL g1418 ( 
.A(n_1356),
.B(n_1210),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_1367),
.Y(n_1419)
);

OAI21xp33_ASAP7_75t_L g1420 ( 
.A1(n_1381),
.A2(n_1239),
.B(n_1237),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1386),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1387),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1360),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1387),
.Y(n_1424)
);

BUFx2_ASAP7_75t_L g1425 ( 
.A(n_1360),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1388),
.Y(n_1426)
);

INVxp67_ASAP7_75t_L g1427 ( 
.A(n_1375),
.Y(n_1427)
);

BUFx2_ASAP7_75t_L g1428 ( 
.A(n_1368),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1370),
.B(n_1221),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1385),
.Y(n_1430)
);

INVx2_ASAP7_75t_SL g1431 ( 
.A(n_1359),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1380),
.B(n_1266),
.Y(n_1432)
);

AND2x2_ASAP7_75t_SL g1433 ( 
.A(n_1389),
.B(n_1198),
.Y(n_1433)
);

BUFx2_ASAP7_75t_L g1434 ( 
.A(n_1379),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1372),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1385),
.A2(n_1229),
.B1(n_1169),
.B2(n_1223),
.Y(n_1436)
);

INVx3_ASAP7_75t_L g1437 ( 
.A(n_1398),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1427),
.B(n_55),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1422),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1415),
.B(n_58),
.Y(n_1440)
);

INVxp67_ASAP7_75t_SL g1441 ( 
.A(n_1424),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1394),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1426),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1402),
.B(n_61),
.Y(n_1444)
);

NAND3xp33_ASAP7_75t_L g1445 ( 
.A(n_1430),
.B(n_61),
.C(n_62),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1405),
.B(n_62),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1435),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1402),
.B(n_63),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1395),
.Y(n_1449)
);

INVx1_ASAP7_75t_SL g1450 ( 
.A(n_1416),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1434),
.B(n_64),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1403),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1428),
.B(n_65),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1408),
.B(n_67),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1423),
.B(n_1425),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1421),
.B(n_68),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1397),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1431),
.B(n_69),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1401),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1410),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_SL g1461 ( 
.A(n_1412),
.B(n_69),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1425),
.B(n_1417),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1407),
.B(n_70),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1396),
.B(n_1392),
.Y(n_1464)
);

INVx3_ASAP7_75t_L g1465 ( 
.A(n_1400),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1399),
.B(n_71),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1406),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1413),
.B(n_72),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1433),
.B(n_74),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1411),
.B(n_75),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1429),
.B(n_76),
.Y(n_1471)
);

NOR3x1_ASAP7_75t_L g1472 ( 
.A(n_1432),
.B(n_77),
.C(n_78),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1419),
.B(n_77),
.Y(n_1473)
);

INVx3_ASAP7_75t_L g1474 ( 
.A(n_1418),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1420),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1436),
.Y(n_1476)
);

NOR2x1_ASAP7_75t_L g1477 ( 
.A(n_1414),
.B(n_79),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1393),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1404),
.B(n_81),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1404),
.B(n_82),
.Y(n_1480)
);

INVx3_ASAP7_75t_L g1481 ( 
.A(n_1398),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1427),
.B(n_83),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1422),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1393),
.Y(n_1484)
);

INVx3_ASAP7_75t_L g1485 ( 
.A(n_1398),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1409),
.B(n_84),
.Y(n_1486)
);

AOI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1477),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1475),
.B(n_88),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1478),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1476),
.B(n_88),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_L g1491 ( 
.A(n_1450),
.B(n_91),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1441),
.B(n_92),
.Y(n_1492)
);

OAI221xp5_ASAP7_75t_L g1493 ( 
.A1(n_1471),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.C(n_95),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1443),
.B(n_95),
.Y(n_1494)
);

NAND2xp33_ASAP7_75t_SL g1495 ( 
.A(n_1444),
.B(n_96),
.Y(n_1495)
);

AO221x2_ASAP7_75t_L g1496 ( 
.A1(n_1445),
.A2(n_99),
.B1(n_97),
.B2(n_98),
.C(n_100),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1455),
.Y(n_1497)
);

AO221x2_ASAP7_75t_L g1498 ( 
.A1(n_1448),
.A2(n_100),
.B1(n_97),
.B2(n_99),
.C(n_101),
.Y(n_1498)
);

AO221x2_ASAP7_75t_L g1499 ( 
.A1(n_1438),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.C(n_105),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1478),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1464),
.B(n_1449),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1452),
.B(n_1457),
.Y(n_1502)
);

OAI22xp33_ASAP7_75t_L g1503 ( 
.A1(n_1474),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1439),
.B(n_110),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1483),
.B(n_111),
.Y(n_1505)
);

OAI221xp5_ASAP7_75t_L g1506 ( 
.A1(n_1468),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.C(n_116),
.Y(n_1506)
);

BUFx2_ASAP7_75t_L g1507 ( 
.A(n_1455),
.Y(n_1507)
);

AO221x2_ASAP7_75t_L g1508 ( 
.A1(n_1482),
.A2(n_117),
.B1(n_119),
.B2(n_116),
.C(n_118),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1462),
.Y(n_1509)
);

AO221x2_ASAP7_75t_L g1510 ( 
.A1(n_1440),
.A2(n_118),
.B1(n_120),
.B2(n_117),
.C(n_119),
.Y(n_1510)
);

NAND2xp33_ASAP7_75t_SL g1511 ( 
.A(n_1469),
.B(n_115),
.Y(n_1511)
);

NAND2xp33_ASAP7_75t_SL g1512 ( 
.A(n_1453),
.B(n_120),
.Y(n_1512)
);

BUFx3_ASAP7_75t_L g1513 ( 
.A(n_1437),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1459),
.B(n_121),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1460),
.B(n_121),
.Y(n_1515)
);

BUFx3_ASAP7_75t_L g1516 ( 
.A(n_1481),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1442),
.B(n_122),
.Y(n_1517)
);

NOR2x1_ASAP7_75t_L g1518 ( 
.A(n_1485),
.B(n_124),
.Y(n_1518)
);

INVxp67_ASAP7_75t_L g1519 ( 
.A(n_1470),
.Y(n_1519)
);

INVx3_ASAP7_75t_L g1520 ( 
.A(n_1465),
.Y(n_1520)
);

AO221x2_ASAP7_75t_L g1521 ( 
.A1(n_1463),
.A2(n_129),
.B1(n_126),
.B2(n_127),
.C(n_130),
.Y(n_1521)
);

XOR2xp5_ASAP7_75t_L g1522 ( 
.A(n_1473),
.B(n_126),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1447),
.B(n_127),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1484),
.B(n_133),
.Y(n_1524)
);

AO221x2_ASAP7_75t_L g1525 ( 
.A1(n_1466),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.C(n_138),
.Y(n_1525)
);

NAND2xp33_ASAP7_75t_SL g1526 ( 
.A(n_1451),
.B(n_137),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1454),
.B(n_139),
.Y(n_1527)
);

AO221x2_ASAP7_75t_L g1528 ( 
.A1(n_1446),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.C(n_143),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_1458),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1479),
.B(n_141),
.Y(n_1530)
);

NAND2xp33_ASAP7_75t_SL g1531 ( 
.A(n_1486),
.B(n_143),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1480),
.B(n_144),
.Y(n_1532)
);

AO221x2_ASAP7_75t_L g1533 ( 
.A1(n_1472),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.C(n_148),
.Y(n_1533)
);

NAND3x1_ASAP7_75t_SL g1534 ( 
.A(n_1456),
.B(n_149),
.C(n_150),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_L g1535 ( 
.A(n_1450),
.B(n_150),
.Y(n_1535)
);

INVx4_ASAP7_75t_L g1536 ( 
.A(n_1437),
.Y(n_1536)
);

NAND2xp33_ASAP7_75t_SL g1537 ( 
.A(n_1461),
.B(n_151),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1478),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1467),
.B(n_153),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1467),
.B(n_154),
.Y(n_1540)
);

AO221x2_ASAP7_75t_L g1541 ( 
.A1(n_1445),
.A2(n_157),
.B1(n_154),
.B2(n_155),
.C(n_158),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_1450),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_SL g1543 ( 
.A(n_1474),
.B(n_159),
.Y(n_1543)
);

NOR2x1_ASAP7_75t_L g1544 ( 
.A(n_1437),
.B(n_160),
.Y(n_1544)
);

AO221x2_ASAP7_75t_L g1545 ( 
.A1(n_1448),
.A2(n_164),
.B1(n_161),
.B2(n_162),
.C(n_165),
.Y(n_1545)
);

NAND2xp33_ASAP7_75t_SL g1546 ( 
.A(n_1461),
.B(n_164),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1519),
.B(n_166),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1489),
.Y(n_1548)
);

A2O1A1Ixp33_ASAP7_75t_SL g1549 ( 
.A1(n_1493),
.A2(n_168),
.B(n_166),
.C(n_167),
.Y(n_1549)
);

AND2x4_ASAP7_75t_SL g1550 ( 
.A(n_1536),
.B(n_169),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1501),
.B(n_170),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1507),
.B(n_170),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1509),
.B(n_171),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1488),
.B(n_171),
.Y(n_1554)
);

NOR2x1_ASAP7_75t_L g1555 ( 
.A(n_1518),
.B(n_172),
.Y(n_1555)
);

INVx1_ASAP7_75t_SL g1556 ( 
.A(n_1513),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1500),
.Y(n_1557)
);

INVx1_ASAP7_75t_SL g1558 ( 
.A(n_1516),
.Y(n_1558)
);

NAND4xp25_ASAP7_75t_L g1559 ( 
.A(n_1487),
.B(n_174),
.C(n_172),
.D(n_173),
.Y(n_1559)
);

NAND2x1p5_ASAP7_75t_L g1560 ( 
.A(n_1520),
.B(n_173),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1538),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1502),
.B(n_175),
.Y(n_1562)
);

AND3x2_ASAP7_75t_L g1563 ( 
.A(n_1491),
.B(n_176),
.C(n_177),
.Y(n_1563)
);

INVx1_ASAP7_75t_SL g1564 ( 
.A(n_1526),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1515),
.B(n_178),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1529),
.B(n_179),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1514),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1504),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1505),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1494),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1492),
.B(n_179),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1532),
.B(n_180),
.Y(n_1572)
);

AOI22x1_ASAP7_75t_L g1573 ( 
.A1(n_1522),
.A2(n_183),
.B1(n_181),
.B2(n_182),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1517),
.Y(n_1574)
);

NAND3xp33_ASAP7_75t_L g1575 ( 
.A(n_1506),
.B(n_184),
.C(n_185),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1544),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1523),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1524),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1539),
.B(n_186),
.Y(n_1579)
);

INVx1_ASAP7_75t_SL g1580 ( 
.A(n_1531),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1540),
.B(n_187),
.Y(n_1581)
);

INVxp67_ASAP7_75t_L g1582 ( 
.A(n_1495),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1490),
.Y(n_1583)
);

BUFx2_ASAP7_75t_L g1584 ( 
.A(n_1511),
.Y(n_1584)
);

INVx2_ASAP7_75t_SL g1585 ( 
.A(n_1533),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1530),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1535),
.B(n_192),
.Y(n_1587)
);

AO21x2_ASAP7_75t_L g1588 ( 
.A1(n_1527),
.A2(n_193),
.B(n_194),
.Y(n_1588)
);

INVxp67_ASAP7_75t_L g1589 ( 
.A(n_1512),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1543),
.B(n_194),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1498),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1499),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_SL g1593 ( 
.A(n_1537),
.B(n_195),
.Y(n_1593)
);

CKINVDCx16_ASAP7_75t_R g1594 ( 
.A(n_1546),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1545),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1521),
.B(n_196),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1510),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1508),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1528),
.B(n_197),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1525),
.Y(n_1600)
);

NAND2xp33_ASAP7_75t_R g1601 ( 
.A(n_1534),
.B(n_198),
.Y(n_1601)
);

INVx3_ASAP7_75t_L g1602 ( 
.A(n_1496),
.Y(n_1602)
);

NAND3xp33_ASAP7_75t_L g1603 ( 
.A(n_1541),
.B(n_199),
.C(n_200),
.Y(n_1603)
);

BUFx2_ASAP7_75t_L g1604 ( 
.A(n_1503),
.Y(n_1604)
);

AND2x4_ASAP7_75t_L g1605 ( 
.A(n_1536),
.B(n_202),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1519),
.B(n_204),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1497),
.B(n_205),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1489),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_1542),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1519),
.B(n_206),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1497),
.B(n_208),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1497),
.B(n_208),
.Y(n_1612)
);

INVx1_ASAP7_75t_SL g1613 ( 
.A(n_1542),
.Y(n_1613)
);

CKINVDCx16_ASAP7_75t_R g1614 ( 
.A(n_1511),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1519),
.B(n_209),
.Y(n_1615)
);

BUFx2_ASAP7_75t_L g1616 ( 
.A(n_1507),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1489),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1489),
.Y(n_1618)
);

OAI21x1_ASAP7_75t_L g1619 ( 
.A1(n_1489),
.A2(n_210),
.B(n_211),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1489),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1519),
.B(n_212),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_L g1622 ( 
.A(n_1519),
.B(n_214),
.Y(n_1622)
);

NAND2x1p5_ASAP7_75t_L g1623 ( 
.A(n_1536),
.B(n_214),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1536),
.B(n_215),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1497),
.B(n_215),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1497),
.B(n_216),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1519),
.B(n_217),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1519),
.B(n_218),
.Y(n_1628)
);

HB1xp67_ASAP7_75t_L g1629 ( 
.A(n_1489),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1489),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1501),
.B(n_223),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1497),
.B(n_224),
.Y(n_1632)
);

OAI322xp33_ASAP7_75t_L g1633 ( 
.A1(n_1591),
.A2(n_230),
.A3(n_229),
.B1(n_227),
.B2(n_225),
.C1(n_226),
.C2(n_228),
.Y(n_1633)
);

OAI31xp33_ASAP7_75t_L g1634 ( 
.A1(n_1584),
.A2(n_230),
.A3(n_228),
.B(n_229),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1629),
.Y(n_1635)
);

AOI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1614),
.A2(n_233),
.B1(n_231),
.B2(n_232),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1548),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_SL g1638 ( 
.A(n_1594),
.B(n_235),
.Y(n_1638)
);

OAI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1595),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1557),
.Y(n_1640)
);

OAI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1592),
.A2(n_239),
.B1(n_237),
.B2(n_238),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1561),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1602),
.B(n_240),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1583),
.B(n_1586),
.Y(n_1644)
);

AOI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1549),
.A2(n_241),
.B(n_242),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1608),
.Y(n_1646)
);

AOI32xp33_ASAP7_75t_L g1647 ( 
.A1(n_1604),
.A2(n_245),
.A3(n_243),
.B1(n_244),
.B2(n_246),
.Y(n_1647)
);

AND2x4_ASAP7_75t_L g1648 ( 
.A(n_1616),
.B(n_243),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1617),
.Y(n_1649)
);

XNOR2x1_ASAP7_75t_L g1650 ( 
.A(n_1596),
.B(n_244),
.Y(n_1650)
);

AOI21xp33_ASAP7_75t_SL g1651 ( 
.A1(n_1601),
.A2(n_245),
.B(n_246),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1618),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1616),
.B(n_247),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1620),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1569),
.B(n_247),
.Y(n_1655)
);

AOI22xp5_ASAP7_75t_L g1656 ( 
.A1(n_1575),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1630),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_SL g1658 ( 
.A(n_1576),
.B(n_251),
.Y(n_1658)
);

AOI211x1_ASAP7_75t_L g1659 ( 
.A1(n_1603),
.A2(n_254),
.B(n_252),
.C(n_253),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1585),
.B(n_254),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1567),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1568),
.Y(n_1662)
);

NAND2x1p5_ASAP7_75t_L g1663 ( 
.A(n_1555),
.B(n_255),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1556),
.B(n_258),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1570),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1574),
.Y(n_1666)
);

NAND2x1_ASAP7_75t_SL g1667 ( 
.A(n_1598),
.B(n_259),
.Y(n_1667)
);

AOI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1597),
.A2(n_262),
.B1(n_260),
.B2(n_261),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1577),
.B(n_262),
.Y(n_1669)
);

OAI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1582),
.A2(n_1589),
.B(n_1593),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1578),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1547),
.Y(n_1672)
);

INVx1_ASAP7_75t_SL g1673 ( 
.A(n_1609),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1551),
.B(n_263),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1588),
.B(n_263),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1562),
.B(n_264),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1558),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1552),
.B(n_265),
.Y(n_1678)
);

INVx1_ASAP7_75t_SL g1679 ( 
.A(n_1613),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1606),
.Y(n_1680)
);

OAI322xp33_ASAP7_75t_L g1681 ( 
.A1(n_1599),
.A2(n_266),
.A3(n_267),
.B1(n_268),
.B2(n_269),
.C1(n_436),
.C2(n_439),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1605),
.Y(n_1682)
);

A2O1A1Ixp33_ASAP7_75t_L g1683 ( 
.A1(n_1600),
.A2(n_269),
.B(n_267),
.C(n_268),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1564),
.B(n_440),
.Y(n_1684)
);

AOI211xp5_ASAP7_75t_L g1685 ( 
.A1(n_1559),
.A2(n_443),
.B(n_441),
.C(n_442),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1615),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1621),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1627),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1628),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1580),
.B(n_445),
.Y(n_1690)
);

INVx2_ASAP7_75t_SL g1691 ( 
.A(n_1624),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1619),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1553),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1607),
.Y(n_1694)
);

INVx2_ASAP7_75t_SL g1695 ( 
.A(n_1667),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1637),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1640),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1642),
.Y(n_1698)
);

AND2x4_ASAP7_75t_L g1699 ( 
.A(n_1677),
.B(n_1550),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1646),
.Y(n_1700)
);

OAI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1636),
.A2(n_1631),
.B1(n_1623),
.B2(n_1560),
.Y(n_1701)
);

OAI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1659),
.A2(n_1573),
.B1(n_1622),
.B2(n_1610),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1649),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1694),
.B(n_1563),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1693),
.B(n_1579),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1652),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1692),
.B(n_1581),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1654),
.Y(n_1708)
);

HB1xp67_ASAP7_75t_L g1709 ( 
.A(n_1648),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_L g1710 ( 
.A(n_1673),
.B(n_1565),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1691),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1679),
.B(n_1571),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1650),
.A2(n_1587),
.B1(n_1572),
.B2(n_1590),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1657),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1653),
.B(n_1611),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1647),
.B(n_1672),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1680),
.B(n_1612),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_L g1718 ( 
.A(n_1682),
.B(n_1554),
.Y(n_1718)
);

INVxp67_ASAP7_75t_L g1719 ( 
.A(n_1638),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1670),
.B(n_1625),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1686),
.B(n_1687),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1688),
.B(n_1632),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1689),
.B(n_1626),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_SL g1724 ( 
.A(n_1634),
.B(n_1566),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1651),
.B(n_453),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1664),
.B(n_454),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1635),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1666),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1671),
.B(n_455),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1661),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1662),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1709),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1699),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1721),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1696),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1697),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1698),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1700),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1703),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1706),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1708),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1714),
.Y(n_1742)
);

INVx3_ASAP7_75t_L g1743 ( 
.A(n_1699),
.Y(n_1743)
);

AND2x4_ASAP7_75t_L g1744 ( 
.A(n_1695),
.B(n_1665),
.Y(n_1744)
);

INVx1_ASAP7_75t_SL g1745 ( 
.A(n_1712),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1727),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1728),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1730),
.Y(n_1748)
);

INVxp33_ASAP7_75t_SL g1749 ( 
.A(n_1710),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1731),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1705),
.Y(n_1751)
);

XNOR2xp5_ASAP7_75t_L g1752 ( 
.A(n_1702),
.B(n_1685),
.Y(n_1752)
);

XNOR2x1_ASAP7_75t_L g1753 ( 
.A(n_1716),
.B(n_1656),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1722),
.Y(n_1754)
);

NAND3xp33_ASAP7_75t_SL g1755 ( 
.A(n_1745),
.B(n_1724),
.C(n_1645),
.Y(n_1755)
);

OAI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1753),
.A2(n_1719),
.B1(n_1668),
.B2(n_1683),
.Y(n_1756)
);

INVx2_ASAP7_75t_SL g1757 ( 
.A(n_1743),
.Y(n_1757)
);

NAND4xp25_ASAP7_75t_L g1758 ( 
.A(n_1749),
.B(n_1711),
.C(n_1704),
.D(n_1707),
.Y(n_1758)
);

NAND4xp25_ASAP7_75t_L g1759 ( 
.A(n_1733),
.B(n_1718),
.C(n_1713),
.D(n_1720),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1744),
.B(n_1723),
.Y(n_1760)
);

NOR2x1_ASAP7_75t_L g1761 ( 
.A(n_1732),
.B(n_1643),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1754),
.B(n_1734),
.Y(n_1762)
);

NOR3x1_ASAP7_75t_L g1763 ( 
.A(n_1751),
.B(n_1644),
.C(n_1717),
.Y(n_1763)
);

AOI211xp5_ASAP7_75t_L g1764 ( 
.A1(n_1752),
.A2(n_1633),
.B(n_1639),
.C(n_1681),
.Y(n_1764)
);

AOI221xp5_ASAP7_75t_L g1765 ( 
.A1(n_1755),
.A2(n_1746),
.B1(n_1737),
.B2(n_1738),
.C(n_1736),
.Y(n_1765)
);

OAI31xp33_ASAP7_75t_L g1766 ( 
.A1(n_1756),
.A2(n_1663),
.A3(n_1701),
.B(n_1641),
.Y(n_1766)
);

NOR4xp25_ASAP7_75t_L g1767 ( 
.A(n_1758),
.B(n_1735),
.C(n_1740),
.D(n_1739),
.Y(n_1767)
);

O2A1O1Ixp33_ASAP7_75t_L g1768 ( 
.A1(n_1764),
.A2(n_1675),
.B(n_1660),
.C(n_1658),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1757),
.B(n_1715),
.Y(n_1769)
);

XNOR2xp5_ASAP7_75t_L g1770 ( 
.A(n_1769),
.B(n_1759),
.Y(n_1770)
);

NAND4xp75_ASAP7_75t_L g1771 ( 
.A(n_1765),
.B(n_1761),
.C(n_1763),
.D(n_1762),
.Y(n_1771)
);

OR2x2_ASAP7_75t_L g1772 ( 
.A(n_1767),
.B(n_1760),
.Y(n_1772)
);

NOR2xp67_ASAP7_75t_L g1773 ( 
.A(n_1766),
.B(n_1741),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1768),
.B(n_1742),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_R g1775 ( 
.A(n_1770),
.B(n_1772),
.Y(n_1775)
);

NAND2xp33_ASAP7_75t_SL g1776 ( 
.A(n_1774),
.B(n_1669),
.Y(n_1776)
);

NAND2xp33_ASAP7_75t_SL g1777 ( 
.A(n_1771),
.B(n_1655),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1776),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1778),
.Y(n_1779)
);

AOI22xp33_ASAP7_75t_L g1780 ( 
.A1(n_1779),
.A2(n_1777),
.B1(n_1775),
.B2(n_1773),
.Y(n_1780)
);

AOI22xp33_ASAP7_75t_L g1781 ( 
.A1(n_1780),
.A2(n_1748),
.B1(n_1750),
.B2(n_1747),
.Y(n_1781)
);

XNOR2x1_ASAP7_75t_L g1782 ( 
.A(n_1781),
.B(n_1726),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1782),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1783),
.Y(n_1784)
);

OAI221xp5_ASAP7_75t_R g1785 ( 
.A1(n_1784),
.A2(n_1674),
.B1(n_1678),
.B2(n_1676),
.C(n_1729),
.Y(n_1785)
);

AOI211xp5_ASAP7_75t_L g1786 ( 
.A1(n_1785),
.A2(n_1690),
.B(n_1684),
.C(n_1725),
.Y(n_1786)
);


endmodule