module real_jpeg_32333_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_288;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_249;
wire n_286;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_11;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_110;
wire n_195;
wire n_205;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_127;
wire n_53;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_0),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g189 ( 
.A(n_0),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_1),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_2),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_3),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_3),
.Y(n_142)
);

OAI32xp33_ASAP7_75t_L g17 ( 
.A1(n_4),
.A2(n_18),
.A3(n_21),
.B1(n_25),
.B2(n_36),
.Y(n_17)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_4),
.A2(n_42),
.B1(n_45),
.B2(n_48),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_4),
.A2(n_42),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

AO22x1_ASAP7_75t_SL g126 ( 
.A1(n_4),
.A2(n_42),
.B1(n_116),
.B2(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_4),
.B(n_98),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_4),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_4),
.B(n_133),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_4),
.B(n_210),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_5),
.Y(n_87)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_6),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_6),
.Y(n_265)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_7),
.Y(n_71)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_7),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_8),
.Y(n_117)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_8),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_9),
.A2(n_90),
.B1(n_93),
.B2(n_94),
.Y(n_89)
);

INVx2_ASAP7_75t_R g93 ( 
.A(n_9),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_9),
.A2(n_93),
.B1(n_140),
.B2(n_143),
.Y(n_139)
);

AOI22x1_ASAP7_75t_L g246 ( 
.A1(n_9),
.A2(n_93),
.B1(n_247),
.B2(n_250),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_231),
.Y(n_10)
);

HB1xp67_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

AOI21x1_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_202),
.B(n_230),
.Y(n_12)
);

OAI21x1_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_150),
.B(n_201),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_130),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_15),
.B(n_130),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_62),
.Y(n_15)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_16),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_43),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_17),
.B(n_43),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_19),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx8_ASAP7_75t_L g275 ( 
.A(n_20),
.Y(n_275)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_24),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_27),
.Y(n_284)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_28),
.Y(n_112)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_28),
.Y(n_125)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_29),
.Y(n_127)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_34),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_35),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_42),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_42),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_42),
.B(n_176),
.Y(n_175)
);

OAI21x1_ASAP7_75t_SL g255 ( 
.A1(n_42),
.A2(n_256),
.B(n_258),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_42),
.B(n_259),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_51),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_44),
.A2(n_53),
.B1(n_139),
.B2(n_146),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_44),
.B(n_53),
.Y(n_159)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_47),
.Y(n_182)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_59),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_58),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_57),
.Y(n_148)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_96),
.B1(n_128),
.B2(n_129),
.Y(n_62)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_63),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_63),
.B(n_161),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_88),
.Y(n_63)
);

NOR2x1_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_82),
.Y(n_64)
);

INVxp67_ASAP7_75t_SL g136 ( 
.A(n_65),
.Y(n_136)
);

NAND2x1p5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_75),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_66),
.B(n_75),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_69),
.B1(n_72),
.B2(n_74),
.Y(n_66)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_68),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_68),
.Y(n_179)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_71),
.Y(n_174)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_75),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_75),
.B(n_239),
.Y(n_238)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_79),
.B2(n_81),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_80),
.Y(n_145)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

INVxp33_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_111),
.B(n_113),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_96),
.A2(n_129),
.B1(n_237),
.B2(n_240),
.Y(n_236)
);

AND2x4_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_118),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_110),
.Y(n_97)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_98),
.Y(n_220)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_120),
.Y(n_119)
);

AOI22x1_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_102),
.B1(n_104),
.B2(n_108),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp33_ASAP7_75t_SL g221 ( 
.A(n_110),
.B(n_119),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_117),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_126),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_126),
.Y(n_219)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_128),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_129),
.B(n_199),
.C(n_229),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_137),
.C(n_149),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_131),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_131),
.Y(n_288)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_132),
.B(n_149),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_132),
.Y(n_225)
);

AO22x2_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_134),
.B(n_238),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_138),
.B(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_138),
.B(n_191),
.Y(n_192)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_138),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_138),
.A2(n_196),
.B1(n_271),
.B2(n_285),
.Y(n_270)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx4f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_SL g146 ( 
.A(n_147),
.Y(n_146)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_194),
.B(n_200),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_183),
.B(n_193),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_160),
.Y(n_152)
);

NAND2xp33_ASAP7_75t_SL g193 ( 
.A(n_153),
.B(n_160),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_153),
.A2(n_154),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_153),
.B(n_208),
.C(n_222),
.Y(n_286)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_185),
.Y(n_184)
);

OA21x2_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_158),
.B(n_159),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_167),
.B1(n_175),
.B2(n_180),
.Y(n_161)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_180),
.B(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_190),
.B(n_192),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx4_ASAP7_75t_SL g188 ( 
.A(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_198),
.Y(n_194)
);

NOR2xp67_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_198),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_228),
.Y(n_202)
);

NOR2xp67_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_228),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_223),
.B2(n_227),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_204),
.B(n_224),
.C(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_218),
.B2(n_222),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_211),
.Y(n_245)
);

NOR2x1_ASAP7_75t_L g260 ( 
.A(n_211),
.B(n_261),
.Y(n_260)
);

AO22x1_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_214),
.B1(n_215),
.B2(n_217),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_216),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_218),
.Y(n_222)
);

OA21x2_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B(n_221),
.Y(n_218)
);

INVxp67_ASAP7_75t_SL g227 ( 
.A(n_223),
.Y(n_227)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_224),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_289),
.Y(n_231)
);

INVxp33_ASAP7_75t_SL g232 ( 
.A(n_233),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_287),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_234),
.B(n_287),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_269),
.Y(n_234)
);

XNOR2x1_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_241),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_237),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_246),
.B(n_254),
.Y(n_244)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_249),
.Y(n_253)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_249),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_249),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_253),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_260),
.Y(n_254)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

OAI32xp33_ASAP7_75t_L g271 ( 
.A1(n_258),
.A2(n_272),
.A3(n_276),
.B1(n_279),
.B2(n_281),
.Y(n_271)
);

AOI22x1_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_266),
.B2(n_267),
.Y(n_261)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_265),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

INVx3_ASAP7_75t_SL g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g280 ( 
.A(n_268),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_286),
.Y(n_269)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_271),
.Y(n_285)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx3_ASAP7_75t_SL g273 ( 
.A(n_274),
.Y(n_273)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx11_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_284),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);


endmodule