module real_jpeg_25521_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_356, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_356;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_286;
wire n_176;
wire n_215;
wire n_166;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_1),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_2),
.A2(n_49),
.B1(n_50),
.B2(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_2),
.A2(n_62),
.B1(n_66),
.B2(n_69),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_62),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_2),
.A2(n_62),
.B1(n_81),
.B2(n_84),
.Y(n_258)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx8_ASAP7_75t_SL g88 ( 
.A(n_4),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_5),
.A2(n_66),
.B1(n_69),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_5),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_5),
.A2(n_30),
.B1(n_31),
.B2(n_77),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_5),
.A2(n_49),
.B1(n_50),
.B2(n_77),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_5),
.A2(n_77),
.B1(n_81),
.B2(n_84),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_6),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_48)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_6),
.A2(n_30),
.B1(n_31),
.B2(n_52),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_6),
.A2(n_52),
.B1(n_66),
.B2(n_69),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_6),
.A2(n_52),
.B1(n_81),
.B2(n_84),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_7),
.A2(n_66),
.B1(n_68),
.B2(n_69),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_7),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_7),
.A2(n_68),
.B1(n_81),
.B2(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_7),
.A2(n_49),
.B1(n_50),
.B2(n_68),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_7),
.A2(n_30),
.B1(n_31),
.B2(n_68),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_8),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_8),
.B(n_92),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_8),
.B(n_31),
.C(n_47),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_8),
.A2(n_49),
.B1(n_50),
.B2(n_82),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_8),
.B(n_75),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_8),
.A2(n_28),
.B1(n_171),
.B2(n_174),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_9),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_10),
.A2(n_84),
.B1(n_91),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_10),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_10),
.A2(n_66),
.B1(n_69),
.B2(n_95),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_10),
.A2(n_49),
.B1(n_50),
.B2(n_95),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_95),
.Y(n_171)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_11),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_12),
.A2(n_30),
.B1(n_31),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_12),
.A2(n_36),
.B1(n_49),
.B2(n_50),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_12),
.A2(n_36),
.B1(n_66),
.B2(n_69),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_12),
.A2(n_36),
.B1(n_323),
.B2(n_325),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_14),
.A2(n_39),
.B1(n_49),
.B2(n_50),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_14),
.A2(n_39),
.B1(n_66),
.B2(n_69),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_14),
.A2(n_39),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_15),
.Y(n_247)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_349),
.C(n_354),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_347),
.B(n_352),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_334),
.B(n_346),
.Y(n_18)
);

OAI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_297),
.A3(n_327),
.B1(n_332),
.B2(n_333),
.C(n_356),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_269),
.B(n_296),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_240),
.B(n_268),
.Y(n_21)
);

O2A1O1Ixp33_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_133),
.B(n_219),
.C(n_239),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_117),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_24),
.B(n_117),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_96),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_59),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_26),
.B(n_59),
.C(n_96),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_44),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_27),
.B(n_44),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_34),
.B(n_37),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_28),
.A2(n_149),
.B(n_150),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_28),
.A2(n_41),
.B1(n_164),
.B2(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_28),
.A2(n_37),
.B(n_153),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_28),
.A2(n_153),
.B(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_29),
.A2(n_35),
.B1(n_40),
.B2(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_29),
.B(n_38),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_29),
.A2(n_151),
.B1(n_163),
.B2(n_165),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_30),
.A2(n_31),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_30),
.B(n_176),
.Y(n_175)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_32),
.Y(n_174)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_33),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_33),
.B(n_82),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_40),
.Y(n_37)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g151 ( 
.A(n_43),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_48),
.B(n_53),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_58),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_45),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_45),
.A2(n_55),
.B1(n_146),
.B2(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_45),
.B(n_82),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_45),
.A2(n_55),
.B(n_308),
.Y(n_307)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_46),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_48),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_50),
.B1(n_72),
.B2(n_73),
.Y(n_74)
);

O2A1O1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_49),
.A2(n_73),
.B(n_185),
.C(n_187),
.Y(n_184)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_50),
.B(n_141),
.Y(n_140)
);

NOR3xp33_ASAP7_75t_L g187 ( 
.A(n_50),
.B(n_69),
.C(n_72),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_53),
.B(n_209),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_54),
.A2(n_61),
.B(n_63),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_54),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_54),
.A2(n_144),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_54),
.A2(n_144),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_55),
.A2(n_208),
.B(n_209),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_55),
.A2(n_249),
.B(n_250),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_64),
.C(n_78),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_60),
.B(n_64),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_61),
.B(n_144),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_61),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_63),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_70),
.B1(n_75),
.B2(n_76),
.Y(n_64)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_69),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_69),
.B1(n_87),
.B2(n_89),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_66),
.A2(n_83),
.B(n_87),
.C(n_115),
.Y(n_114)
);

HAxp5_ASAP7_75t_SL g186 ( 
.A(n_66),
.B(n_82),
.CON(n_186),
.SN(n_186)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND3xp33_ASAP7_75t_L g115 ( 
.A(n_69),
.B(n_84),
.C(n_89),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_70),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_70),
.A2(n_75),
.B1(n_131),
.B2(n_186),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_70),
.A2(n_108),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_70),
.B(n_263),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_70),
.A2(n_75),
.B1(n_275),
.B2(n_276),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_70),
.A2(n_236),
.B(n_276),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_70),
.A2(n_75),
.B(n_108),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_74),
.A2(n_106),
.B1(n_130),
.B2(n_132),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_74),
.B(n_237),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_74),
.A2(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_75),
.B(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_76),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_78),
.B(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_85),
.B1(n_92),
.B2(n_93),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_82),
.B(n_83),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_87),
.B1(n_89),
.B2(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_80),
.Y(n_289)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

INVx8_ASAP7_75t_L g288 ( 
.A(n_81),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_82),
.B(n_84),
.Y(n_83)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_85),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_85),
.A2(n_92),
.B1(n_102),
.B2(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_85),
.B(n_287),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_85),
.A2(n_92),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_85),
.A2(n_322),
.B(n_341),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_85),
.A2(n_92),
.B(n_258),
.Y(n_354)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_90),
.Y(n_85)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_86),
.A2(n_94),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_86),
.A2(n_302),
.B(n_303),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g89 ( 
.A(n_87),
.Y(n_89)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_92),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_92),
.B(n_287),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_109),
.B2(n_116),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_104),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_99),
.B(n_104),
.C(n_116),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_100),
.A2(n_256),
.B(n_257),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_100),
.A2(n_285),
.B(n_286),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

INVx8_ASAP7_75t_L g324 ( 
.A(n_103),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B(n_107),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_107),
.B(n_262),
.Y(n_319)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_110),
.A2(n_111),
.B1(n_114),
.B2(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_113),
.A2(n_124),
.B(n_126),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_114),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_120),
.C(n_122),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_118),
.B(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_120),
.B(n_122),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_127),
.C(n_129),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_123),
.A2(n_127),
.B1(n_128),
.B2(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_123),
.Y(n_203)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_126),
.B(n_150),
.Y(n_225)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_129),
.B(n_202),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_218),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_213),
.B(n_217),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_197),
.B(n_212),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_180),
.B(n_196),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_160),
.B(n_179),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_147),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_147),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_142),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_154),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_148),
.B(n_155),
.C(n_158),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_149),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_159),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_167),
.B(n_178),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_166),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_166),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_172),
.B(n_177),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_170),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_175),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_195),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_195),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_190),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_191),
.C(n_192),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_188),
.B2(n_189),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_189),
.Y(n_206)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_194),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_199),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_204),
.B2(n_205),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_207),
.C(n_210),
.Y(n_216)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_210),
.B2(n_211),
.Y(n_205)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_216),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_216),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_221),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_238),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_230),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_230),
.C(n_238),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_229),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_229),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_226),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_228),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_231),
.B(n_233),
.C(n_235),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_234),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_241),
.B(n_242),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_267),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_252),
.B1(n_265),
.B2(n_266),
.Y(n_243)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_244),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_266),
.C(n_267),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_248),
.B2(n_251),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_245),
.A2(n_246),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_245),
.A2(n_280),
.B(n_284),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_246),
.B(n_248),
.Y(n_281)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_248),
.Y(n_251)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_252),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_253),
.B(n_259),
.C(n_264),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_259),
.B1(n_260),
.B2(n_264),
.Y(n_254)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_255),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_257),
.B(n_303),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_258),
.Y(n_285)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_261),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_270),
.B(n_271),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_271)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_279),
.B1(n_291),
.B2(n_292),
.Y(n_272)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_273),
.Y(n_291)
);

OAI21xp33_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_277),
.B(n_278),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_274),
.B(n_277),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_278),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_278),
.A2(n_299),
.B1(n_311),
.B2(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_279),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_279),
.B(n_291),
.C(n_295),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_282),
.B2(n_290),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_282),
.Y(n_290)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_286),
.Y(n_341)
);

INVx11_ASAP7_75t_L g325 ( 
.A(n_288),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_293),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_313),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_298),
.B(n_313),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_311),
.C(n_312),
.Y(n_298)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_299),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_304),
.B2(n_305),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_300),
.A2(n_301),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_301),
.B(n_306),
.C(n_310),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_301),
.B(n_316),
.C(n_326),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_302),
.Y(n_321)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_309),
.B2(n_310),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_306),
.A2(n_307),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_307),
.B(n_318),
.C(n_320),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_310),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_312),
.B(n_330),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_326),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_320),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_319),
.Y(n_318)
);

INVx8_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_328),
.B(n_329),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_335),
.B(n_336),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_338),
.B1(n_344),
.B2(n_345),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_340),
.B1(n_342),
.B2(n_343),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_339),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_340),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_340),
.B(n_342),
.C(n_344),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_345),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_349),
.Y(n_353)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_351),
.B(n_353),
.Y(n_352)
);


endmodule