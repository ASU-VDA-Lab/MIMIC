module fake_netlist_1_6731_n_13 (n_1, n_2, n_0, n_13);
input n_1;
input n_2;
input n_0;
output n_13;
wire n_11;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx1_ASAP7_75t_L g3 ( .A(n_1), .Y(n_3) );
NAND2xp33_ASAP7_75t_L g4 ( .A(n_2), .B(n_0), .Y(n_4) );
OAI21x1_ASAP7_75t_L g5 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_5) );
HB1xp67_ASAP7_75t_L g6 ( .A(n_3), .Y(n_6) );
NAND3xp33_ASAP7_75t_L g7 ( .A(n_6), .B(n_4), .C(n_1), .Y(n_7) );
BUFx2_ASAP7_75t_L g8 ( .A(n_5), .Y(n_8) );
NAND3xp33_ASAP7_75t_SL g9 ( .A(n_7), .B(n_4), .C(n_1), .Y(n_9) );
AOI21xp33_ASAP7_75t_L g10 ( .A1(n_8), .A2(n_5), .B(n_0), .Y(n_10) );
AOI21xp5_ASAP7_75t_L g11 ( .A1(n_10), .A2(n_0), .B(n_2), .Y(n_11) );
NAND2xp5_ASAP7_75t_L g12 ( .A(n_11), .B(n_9), .Y(n_12) );
NOR3xp33_ASAP7_75t_L g13 ( .A(n_12), .B(n_2), .C(n_9), .Y(n_13) );
endmodule