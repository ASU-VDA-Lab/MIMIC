module fake_jpeg_5599_n_131 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_131);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx4f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx2_ASAP7_75t_R g24 ( 
.A(n_18),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_24),
.Y(n_49)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_20),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_28),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_20),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_29),
.B(n_19),
.Y(n_34)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_32),
.A2(n_13),
.B1(n_17),
.B2(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx9p33_ASAP7_75t_R g41 ( 
.A(n_24),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_28),
.B(n_14),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_47),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_13),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_28),
.B(n_14),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_29),
.B(n_14),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_19),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_35),
.A2(n_13),
.B1(n_30),
.B2(n_32),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_52),
.A2(n_60),
.B1(n_40),
.B2(n_25),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_21),
.Y(n_57)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_32),
.B1(n_25),
.B2(n_17),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_21),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_61),
.B(n_35),
.Y(n_69)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_29),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_33),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_65),
.Y(n_80)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

AND2x4_ASAP7_75t_SL g67 ( 
.A(n_37),
.B(n_27),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_41),
.B(n_37),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_69),
.B(n_77),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_73),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_34),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_84),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_52),
.A2(n_25),
.B1(n_32),
.B2(n_39),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_74),
.A2(n_75),
.B1(n_65),
.B2(n_62),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_66),
.A2(n_39),
.B1(n_49),
.B2(n_31),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_SL g88 ( 
.A(n_78),
.B(n_81),
.C(n_67),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_37),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_21),
.Y(n_82)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_45),
.Y(n_83)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_47),
.Y(n_84)
);

AO21x2_ASAP7_75t_L g85 ( 
.A1(n_74),
.A2(n_67),
.B(n_56),
.Y(n_85)
);

AOI21x1_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_89),
.B(n_68),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_63),
.B(n_55),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_55),
.C(n_56),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_92),
.C(n_79),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_56),
.C(n_37),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_94),
.A2(n_70),
.B1(n_75),
.B2(n_77),
.Y(n_101)
);

AND2x6_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_54),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_99),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_77),
.B(n_79),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_98),
.Y(n_100)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_90),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_54),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_105),
.A2(n_85),
.B(n_95),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_31),
.B1(n_45),
.B2(n_26),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_109),
.A2(n_102),
.B1(n_106),
.B2(n_105),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_110),
.A2(n_112),
.B(n_113),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_104),
.A2(n_103),
.B(n_100),
.C(n_101),
.Y(n_111)
);

OAI21xp33_ASAP7_75t_L g112 ( 
.A1(n_108),
.A2(n_88),
.B(n_93),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_107),
.A2(n_92),
.B(n_89),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_97),
.B(n_87),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_114),
.Y(n_116)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_116),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_26),
.C(n_76),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_16),
.C(n_22),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_117),
.B(n_111),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_122),
.B(n_121),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_22),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_123),
.Y(n_125)
);

INVxp33_ASAP7_75t_L g126 ( 
.A(n_124),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_127),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_125),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_8),
.C(n_9),
.Y(n_129)
);

XNOR2x2_ASAP7_75t_SL g130 ( 
.A(n_129),
.B(n_18),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_18),
.Y(n_131)
);


endmodule