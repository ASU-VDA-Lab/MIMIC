module fake_jpeg_18412_n_314 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_314);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_314;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_SL g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_25),
.Y(n_43)
);

AND2x4_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_44),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_25),
.B(n_0),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_22),
.B1(n_21),
.B2(n_30),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_47),
.A2(n_56),
.B1(n_39),
.B2(n_38),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_42),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_48),
.B(n_55),
.Y(n_68)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_36),
.A2(n_22),
.B1(n_21),
.B2(n_30),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_30),
.B1(n_17),
.B2(n_18),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_57),
.A2(n_9),
.B1(n_11),
.B2(n_14),
.Y(n_106)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_65),
.B(n_42),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_52),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_66),
.B(n_85),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_44),
.B1(n_38),
.B2(n_40),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_70),
.A2(n_78),
.B1(n_95),
.B2(n_96),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_43),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_74),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_40),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

OAI21xp33_ASAP7_75t_L g77 ( 
.A1(n_50),
.A2(n_39),
.B(n_20),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_77),
.A2(n_83),
.B(n_90),
.Y(n_136)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_42),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_24),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_87),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_49),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_86),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_24),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_53),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_94),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_62),
.A2(n_20),
.B1(n_33),
.B2(n_34),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_53),
.A2(n_39),
.B1(n_38),
.B2(n_18),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_93),
.A2(n_102),
.B1(n_41),
.B2(n_42),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_51),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_63),
.A2(n_16),
.B1(n_17),
.B2(n_23),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_46),
.A2(n_31),
.B1(n_23),
.B2(n_26),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_65),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_101),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_46),
.A2(n_31),
.B1(n_26),
.B2(n_16),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_99),
.B1(n_105),
.B2(n_45),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_46),
.A2(n_32),
.B1(n_27),
.B2(n_34),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_106),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_61),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_64),
.A2(n_32),
.B1(n_33),
.B2(n_27),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_60),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_104),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_60),
.A2(n_24),
.B1(n_28),
.B2(n_25),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_35),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_109),
.B(n_114),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_84),
.C(n_83),
.Y(n_114)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_132),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_68),
.A2(n_45),
.B1(n_64),
.B2(n_48),
.Y(n_120)
);

AO21x2_ASAP7_75t_L g137 ( 
.A1(n_120),
.A2(n_135),
.B(n_105),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_122),
.A2(n_129),
.B1(n_86),
.B2(n_100),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_42),
.C(n_61),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_124),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_29),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_41),
.B1(n_28),
.B2(n_42),
.Y(n_129)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_66),
.B(n_35),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_134),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_95),
.A2(n_28),
.B1(n_35),
.B2(n_29),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_137),
.A2(n_117),
.B1(n_75),
.B2(n_91),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_115),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_140),
.B(n_142),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_71),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_141),
.B(n_159),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_116),
.Y(n_142)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

NOR2x1_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_90),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_147),
.B(n_154),
.Y(n_193)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_162),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_125),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_149),
.B(n_160),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_136),
.A2(n_71),
.B(n_72),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_150),
.A2(n_124),
.B(n_133),
.Y(n_175)
);

AND2x2_ASAP7_75t_SL g151 ( 
.A(n_121),
.B(n_72),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_151),
.A2(n_156),
.B(n_141),
.Y(n_171)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_113),
.Y(n_152)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_153),
.Y(n_194)
);

NOR2x1_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_98),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_155),
.Y(n_178)
);

AND2x2_ASAP7_75t_SL g156 ( 
.A(n_121),
.B(n_79),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_128),
.A2(n_75),
.B1(n_85),
.B2(n_103),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_157),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_108),
.B(n_92),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_110),
.B(n_67),
.Y(n_160)
);

BUFx24_ASAP7_75t_SL g162 ( 
.A(n_109),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_114),
.B(n_80),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_166),
.Y(n_187)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_165),
.Y(n_195)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_167),
.B(n_0),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_129),
.B1(n_131),
.B2(n_107),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_169),
.A2(n_177),
.B1(n_152),
.B2(n_146),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_158),
.A2(n_131),
.B(n_133),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_170),
.A2(n_198),
.B(n_199),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_171),
.B(n_183),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_123),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_192),
.Y(n_205)
);

AND2x6_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_107),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_173),
.B(n_191),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_175),
.A2(n_196),
.B(n_149),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_132),
.C(n_118),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_139),
.C(n_156),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_167),
.A2(n_88),
.B1(n_126),
.B2(n_112),
.Y(n_177)
);

AO22x1_ASAP7_75t_L g183 ( 
.A1(n_159),
.A2(n_88),
.B1(n_42),
.B2(n_91),
.Y(n_183)
);

OA21x2_ASAP7_75t_L g184 ( 
.A1(n_154),
.A2(n_117),
.B(n_69),
.Y(n_184)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_184),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_188),
.A2(n_137),
.B1(n_3),
.B2(n_4),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_76),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_190),
.B(n_197),
.Y(n_204)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_153),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_29),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_150),
.A2(n_0),
.B(n_1),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_6),
.Y(n_197)
);

A2O1A1Ixp33_ASAP7_75t_SL g199 ( 
.A1(n_158),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_179),
.Y(n_200)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_200),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_174),
.B(n_166),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_202),
.B(n_216),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_210),
.C(n_211),
.Y(n_228)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_206),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_155),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_207),
.A2(n_219),
.B(n_182),
.Y(n_241)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_181),
.Y(n_208)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_208),
.Y(n_244)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_181),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_226),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_172),
.B(n_176),
.C(n_139),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_156),
.C(n_151),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_213),
.A2(n_169),
.B1(n_182),
.B2(n_137),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_196),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_151),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_185),
.Y(n_233)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_186),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_187),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_218),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_173),
.A2(n_137),
.B1(n_168),
.B2(n_145),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_189),
.B(n_144),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_222),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_194),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_171),
.B(n_144),
.C(n_143),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_170),
.C(n_184),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_185),
.B(n_143),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_178),
.Y(n_231)
);

AOI322xp5_ASAP7_75t_L g225 ( 
.A1(n_180),
.A2(n_137),
.A3(n_138),
.B1(n_148),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_225)
);

NAND3xp33_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_199),
.C(n_191),
.Y(n_234)
);

MAJx2_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_210),
.C(n_175),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_241),
.Y(n_249)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_231),
.Y(n_255)
);

OAI21xp33_ASAP7_75t_L g232 ( 
.A1(n_212),
.A2(n_193),
.B(n_184),
.Y(n_232)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_232),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_211),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_234),
.A2(n_242),
.B1(n_209),
.B2(n_206),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_183),
.Y(n_235)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_235),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_247),
.C(n_205),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_207),
.B(n_183),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_246),
.Y(n_253)
);

FAx1_ASAP7_75t_SL g261 ( 
.A(n_240),
.B(n_207),
.CI(n_220),
.CON(n_261),
.SN(n_261)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_204),
.B(n_194),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_203),
.B(n_177),
.C(n_199),
.Y(n_247)
);

XOR2x2_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_223),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_248),
.B(n_252),
.Y(n_270)
);

NAND2x1_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_220),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_250),
.A2(n_239),
.B(n_243),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_230),
.A2(n_226),
.B1(n_217),
.B2(n_201),
.Y(n_251)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_251),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_247),
.Y(n_254)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_257),
.C(n_260),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_212),
.C(n_214),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_227),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_262),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_228),
.B(n_238),
.C(n_233),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_261),
.B(n_243),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_219),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_201),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_266),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_265),
.A2(n_213),
.B1(n_236),
.B2(n_199),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_245),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_250),
.A2(n_230),
.B1(n_242),
.B2(n_257),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_2),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_269),
.A2(n_272),
.B(n_13),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_237),
.C(n_244),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_276),
.C(n_280),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_274),
.A2(n_264),
.B1(n_261),
.B2(n_263),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_8),
.C(n_12),
.Y(n_276)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_253),
.Y(n_279)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_279),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_9),
.C(n_12),
.Y(n_280)
);

A2O1A1O1Ixp25_ASAP7_75t_L g281 ( 
.A1(n_269),
.A2(n_248),
.B(n_261),
.C(n_258),
.D(n_262),
.Y(n_281)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_281),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_255),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_277),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_283),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_249),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_286),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_249),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_289),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_278),
.Y(n_290)
);

INVx11_ASAP7_75t_L g299 ( 
.A(n_290),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_7),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_291),
.B(n_280),
.Y(n_293)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_293),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_294),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_268),
.C(n_267),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_268),
.C(n_285),
.Y(n_305)
);

AOI322xp5_ASAP7_75t_L g300 ( 
.A1(n_295),
.A2(n_288),
.A3(n_275),
.B1(n_284),
.B2(n_281),
.C1(n_271),
.C2(n_286),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_300),
.A2(n_299),
.B1(n_11),
.B2(n_7),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_274),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_303),
.C(n_305),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_292),
.A2(n_297),
.B(n_295),
.Y(n_303)
);

AOI31xp67_ASAP7_75t_L g306 ( 
.A1(n_304),
.A2(n_299),
.A3(n_296),
.B(n_298),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_306),
.A2(n_301),
.B(n_305),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_307),
.B(n_13),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_309),
.B(n_310),
.Y(n_311)
);

AOI322xp5_ASAP7_75t_L g312 ( 
.A1(n_311),
.A2(n_3),
.A3(n_4),
.B1(n_9),
.B2(n_12),
.C1(n_308),
.C2(n_306),
.Y(n_312)
);

NAND2xp33_ASAP7_75t_R g313 ( 
.A(n_312),
.B(n_3),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_3),
.Y(n_314)
);


endmodule