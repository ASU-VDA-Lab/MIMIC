module fake_jpeg_17632_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_11),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_34),
.Y(n_57)
);

INVxp67_ASAP7_75t_SL g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_21),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_43),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_39),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_44),
.B(n_50),
.Y(n_77)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_58),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_39),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_34),
.Y(n_69)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx4_ASAP7_75t_SL g53 ( 
.A(n_35),
.Y(n_53)
);

CKINVDCx6p67_ASAP7_75t_R g83 ( 
.A(n_53),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_19),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_25),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_37),
.Y(n_84)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

AO22x2_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_35),
.B1(n_34),
.B2(n_36),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_67),
.A2(n_34),
.B1(n_59),
.B2(n_54),
.Y(n_92)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_29),
.Y(n_70)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_21),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_74),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_29),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_25),
.Y(n_94)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_81),
.Y(n_105)
);

HAxp5_ASAP7_75t_SL g80 ( 
.A(n_58),
.B(n_21),
.CON(n_80),
.SN(n_80)
);

MAJx2_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_34),
.C(n_53),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_54),
.Y(n_81)
);

BUFx6f_ASAP7_75t_SL g82 ( 
.A(n_60),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_38),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

BUFx4f_ASAP7_75t_SL g108 ( 
.A(n_88),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

O2A1O1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_92),
.A2(n_117),
.B(n_97),
.C(n_79),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_94),
.B(n_107),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_16),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_95),
.B(n_103),
.Y(n_119)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_104),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_67),
.A2(n_17),
.B1(n_32),
.B2(n_36),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_98),
.A2(n_115),
.B1(n_117),
.B2(n_33),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_38),
.Y(n_121)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_42),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_87),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_68),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_68),
.B(n_24),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_111),
.Y(n_128)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_80),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_113),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_67),
.B(n_16),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_67),
.A2(n_65),
.B1(n_45),
.B2(n_52),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_121),
.B(n_83),
.Y(n_165)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_20),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_125),
.A2(n_130),
.B1(n_133),
.B2(n_141),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_129),
.Y(n_153)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_98),
.A2(n_48),
.B1(n_90),
.B2(n_71),
.Y(n_130)
);

OR2x2_ASAP7_75t_SL g132 ( 
.A(n_100),
.B(n_26),
.Y(n_132)
);

MAJx2_ASAP7_75t_L g174 ( 
.A(n_132),
.B(n_83),
.C(n_33),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_111),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_134),
.B(n_140),
.Y(n_149)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_136),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_106),
.A2(n_78),
.B1(n_71),
.B2(n_17),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_99),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_138),
.Y(n_154)
);

INVxp33_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_92),
.A2(n_17),
.B1(n_32),
.B2(n_78),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_143),
.A2(n_64),
.B1(n_46),
.B2(n_114),
.Y(n_147)
);

NOR2x1_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_83),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_145),
.B(n_22),
.Y(n_157)
);

OAI21xp33_ASAP7_75t_SL g188 ( 
.A1(n_147),
.A2(n_171),
.B(n_174),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_93),
.B1(n_101),
.B2(n_72),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_148),
.A2(n_172),
.B1(n_140),
.B2(n_126),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_135),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_161),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_72),
.Y(n_155)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_156),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_145),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_122),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_119),
.B(n_134),
.Y(n_162)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_162),
.Y(n_185)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_163),
.Y(n_190)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_120),
.Y(n_164)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_165),
.B(n_170),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_142),
.B(n_24),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_167),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_128),
.B(n_26),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_168),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_128),
.B(n_31),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_173),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_43),
.C(n_57),
.Y(n_170)
);

OAI32xp33_ASAP7_75t_L g171 ( 
.A1(n_132),
.A2(n_83),
.A3(n_28),
.B1(n_22),
.B2(n_16),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_125),
.A2(n_101),
.B1(n_42),
.B2(n_82),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_125),
.B(n_43),
.C(n_57),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_160),
.A2(n_139),
.B1(n_143),
.B2(n_130),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_175),
.A2(n_179),
.B1(n_184),
.B2(n_196),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_177),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_149),
.Y(n_178)
);

O2A1O1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_178),
.A2(n_28),
.B(n_20),
.C(n_23),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_152),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_191),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_158),
.A2(n_136),
.B(n_122),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_182),
.A2(n_22),
.B(n_28),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_146),
.A2(n_85),
.B1(n_123),
.B2(n_129),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_186),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_152),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_151),
.Y(n_192)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_192),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_151),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_200),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_158),
.A2(n_138),
.B1(n_123),
.B2(n_144),
.Y(n_196)
);

AND2x6_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_1),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_SL g204 ( 
.A(n_197),
.B(n_171),
.C(n_174),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_144),
.Y(n_198)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_163),
.Y(n_199)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_199),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_160),
.B(n_113),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_204),
.A2(n_209),
.B1(n_210),
.B2(n_181),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_183),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_214),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_155),
.C(n_173),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_208),
.B(n_212),
.C(n_216),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_188),
.A2(n_146),
.B1(n_162),
.B2(n_170),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_178),
.A2(n_147),
.B1(n_148),
.B2(n_172),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_154),
.Y(n_211)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_42),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_186),
.Y(n_213)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_213),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_194),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_154),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_179),
.B(n_43),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_218),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_108),
.C(n_43),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_177),
.B(n_18),
.Y(n_219)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_220),
.A2(n_185),
.B(n_196),
.Y(n_233)
);

INVxp33_ASAP7_75t_SL g223 ( 
.A(n_190),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_223),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_187),
.B(n_31),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_224),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_57),
.Y(n_245)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_228),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_222),
.B(n_176),
.Y(n_229)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

XOR2x1_ASAP7_75t_SL g232 ( 
.A(n_223),
.B(n_209),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_23),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_233),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_182),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_237),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_185),
.Y(n_236)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_184),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_203),
.B(n_201),
.Y(n_240)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_220),
.A2(n_199),
.B(n_192),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_241),
.A2(n_4),
.B(n_5),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_190),
.Y(n_243)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_243),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_245),
.A2(n_227),
.B1(n_213),
.B2(n_85),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_216),
.B(n_197),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_247),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_27),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_232),
.A2(n_205),
.B1(n_225),
.B2(n_215),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_249),
.A2(n_261),
.B1(n_262),
.B2(n_264),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_218),
.C(n_226),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_265),
.C(n_238),
.Y(n_270)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_254),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_226),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_255),
.B(n_247),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_256),
.A2(n_5),
.B(n_6),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_233),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_257),
.A2(n_245),
.B1(n_241),
.B2(n_242),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_231),
.A2(n_91),
.B1(n_88),
.B2(n_86),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_91),
.C(n_21),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_250),
.A2(n_237),
.B1(n_230),
.B2(n_235),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_266),
.A2(n_274),
.B1(n_278),
.B2(n_18),
.Y(n_289)
);

NAND4xp25_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_234),
.C(n_246),
.D(n_252),
.Y(n_267)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_267),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_268),
.B(n_271),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_273),
.C(n_275),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_239),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_261),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_238),
.C(n_21),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_258),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_27),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_249),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_276),
.A2(n_277),
.B1(n_279),
.B2(n_27),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_253),
.A2(n_256),
.B1(n_265),
.B2(n_263),
.Y(n_278)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_280),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_263),
.C(n_262),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_287),
.C(n_30),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_276),
.A2(n_7),
.B(n_8),
.Y(n_283)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_283),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_285),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_19),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_290),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_18),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_273),
.A2(n_8),
.B(n_9),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_288),
.A2(n_292),
.B(n_10),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_30),
.Y(n_296)
);

INVx6_ASAP7_75t_L g290 ( 
.A(n_269),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_9),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_275),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_10),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_274),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_295),
.B(n_301),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_298),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_292),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_291),
.B(n_10),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_294),
.A2(n_284),
.B1(n_285),
.B2(n_290),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_304),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_308),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_30),
.C(n_11),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_307),
.A2(n_302),
.B(n_294),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_11),
.Y(n_309)
);

AOI322xp5_ASAP7_75t_L g311 ( 
.A1(n_309),
.A2(n_12),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.C1(n_300),
.C2(n_303),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_310),
.A2(n_311),
.B(n_312),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_313),
.C(n_308),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_307),
.C(n_305),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_316),
.B(n_12),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_13),
.C(n_15),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_13),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_319),
.Y(n_320)
);


endmodule