module fake_netlist_1_12256_n_558 (n_117, n_44, n_133, n_149, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_125, n_9, n_161, n_10, n_130, n_103, n_19, n_87, n_137, n_104, n_160, n_98, n_74, n_154, n_7, n_29, n_165, n_146, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_169, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_24, n_78, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_38, n_64, n_142, n_46, n_31, n_58, n_122, n_138, n_126, n_118, n_32, n_0, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_166, n_162, n_75, n_163, n_105, n_159, n_72, n_136, n_43, n_76, n_89, n_68, n_144, n_27, n_53, n_67, n_77, n_20, n_2, n_147, n_54, n_148, n_123, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_15, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_558);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_125;
input n_9;
input n_161;
input n_10;
input n_130;
input n_103;
input n_19;
input n_87;
input n_137;
input n_104;
input n_160;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_165;
input n_146;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_169;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_38;
input n_64;
input n_142;
input n_46;
input n_31;
input n_58;
input n_122;
input n_138;
input n_126;
input n_118;
input n_32;
input n_0;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_166;
input n_162;
input n_75;
input n_163;
input n_105;
input n_159;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_68;
input n_144;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_54;
input n_148;
input n_123;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_15;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_558;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_431;
wire n_484;
wire n_496;
wire n_177;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_202;
wire n_386;
wire n_432;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_205;
wire n_330;
wire n_387;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_517;
wire n_479;
wire n_554;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_207;
wire n_224;
wire n_219;
wire n_475;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_450;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_379;
wire n_527;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_514;
wire n_486;
wire n_357;
wire n_245;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_178;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_295;
wire n_263;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_552;
wire n_344;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_300;
wire n_524;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_198;
wire n_424;
wire n_297;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_291;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_187;
wire n_375;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_421;
wire n_175;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g171 ( .A(n_45), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_126), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_69), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_116), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_51), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_146), .Y(n_176) );
BUFx5_ASAP7_75t_L g177 ( .A(n_82), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_81), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_80), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_48), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_164), .Y(n_181) );
INVxp67_ASAP7_75t_SL g182 ( .A(n_26), .Y(n_182) );
HB1xp67_ASAP7_75t_L g183 ( .A(n_40), .Y(n_183) );
CKINVDCx16_ASAP7_75t_R g184 ( .A(n_168), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_169), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_160), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_153), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_83), .Y(n_188) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_97), .Y(n_189) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_73), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_1), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_162), .Y(n_192) );
INVxp67_ASAP7_75t_L g193 ( .A(n_46), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_120), .Y(n_194) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_15), .Y(n_195) );
BUFx3_ASAP7_75t_L g196 ( .A(n_148), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_133), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_67), .Y(n_198) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_135), .Y(n_199) );
BUFx8_ASAP7_75t_SL g200 ( .A(n_150), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_100), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_54), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_159), .Y(n_203) );
INVx1_ASAP7_75t_SL g204 ( .A(n_99), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_147), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_50), .Y(n_206) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_107), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_104), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_149), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_66), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_165), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_108), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_77), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_42), .Y(n_214) );
HB1xp67_ASAP7_75t_L g215 ( .A(n_25), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_30), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_145), .Y(n_217) );
INVxp67_ASAP7_75t_L g218 ( .A(n_111), .Y(n_218) );
INVx1_ASAP7_75t_SL g219 ( .A(n_161), .Y(n_219) );
CKINVDCx5p33_ASAP7_75t_R g220 ( .A(n_109), .Y(n_220) );
INVxp67_ASAP7_75t_L g221 ( .A(n_13), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_62), .Y(n_222) );
INVx1_ASAP7_75t_SL g223 ( .A(n_75), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_79), .Y(n_224) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_114), .Y(n_225) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_170), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_37), .Y(n_227) );
INVxp67_ASAP7_75t_L g228 ( .A(n_130), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_39), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_31), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_64), .Y(n_231) );
BUFx3_ASAP7_75t_L g232 ( .A(n_72), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_124), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_26), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_89), .Y(n_235) );
BUFx5_ASAP7_75t_L g236 ( .A(n_88), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_136), .Y(n_237) );
INVx3_ASAP7_75t_L g238 ( .A(n_121), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_141), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_163), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_84), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_112), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_119), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_59), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_95), .Y(n_245) );
CKINVDCx5p33_ASAP7_75t_R g246 ( .A(n_118), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_138), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_139), .Y(n_248) );
BUFx10_ASAP7_75t_L g249 ( .A(n_7), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_74), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_19), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_76), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_166), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_144), .Y(n_254) );
INVxp67_ASAP7_75t_L g255 ( .A(n_70), .Y(n_255) );
INVx1_ASAP7_75t_SL g256 ( .A(n_105), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_29), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_85), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_142), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_63), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_106), .Y(n_261) );
BUFx3_ASAP7_75t_L g262 ( .A(n_55), .Y(n_262) );
CKINVDCx16_ASAP7_75t_R g263 ( .A(n_86), .Y(n_263) );
INVx3_ASAP7_75t_L g264 ( .A(n_41), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_102), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_184), .A2(n_3), .B1(n_0), .B2(n_2), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g267 ( .A(n_263), .Y(n_267) );
INVx2_ASAP7_75t_SL g268 ( .A(n_249), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_238), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_183), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_200), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_215), .B(n_0), .Y(n_272) );
BUFx6f_ASAP7_75t_L g273 ( .A(n_190), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_238), .Y(n_274) );
BUFx6f_ASAP7_75t_L g275 ( .A(n_190), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_264), .Y(n_276) );
OAI21x1_ASAP7_75t_L g277 ( .A1(n_264), .A2(n_34), .B(n_33), .Y(n_277) );
INVx5_ASAP7_75t_L g278 ( .A(n_190), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_177), .Y(n_279) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_171), .Y(n_280) );
AOI22xp5_ASAP7_75t_SL g281 ( .A1(n_182), .A2(n_6), .B1(n_4), .B2(n_5), .Y(n_281) );
OAI21x1_ASAP7_75t_L g282 ( .A1(n_173), .A2(n_36), .B(n_35), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_230), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_177), .Y(n_284) );
INVx6_ASAP7_75t_L g285 ( .A(n_249), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_279), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_269), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_269), .Y(n_288) );
OAI22xp33_ASAP7_75t_L g289 ( .A1(n_266), .A2(n_182), .B1(n_221), .B2(n_216), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_274), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_270), .B(n_193), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_284), .Y(n_292) );
INVx3_ASAP7_75t_L g293 ( .A(n_276), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_284), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_285), .B(n_218), .Y(n_295) );
NAND3xp33_ASAP7_75t_L g296 ( .A(n_272), .B(n_234), .C(n_195), .Y(n_296) );
OR2x2_ASAP7_75t_L g297 ( .A(n_268), .B(n_191), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_283), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_280), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_271), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_295), .B(n_267), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_291), .B(n_218), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_293), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g304 ( .A1(n_288), .A2(n_280), .B1(n_257), .B2(n_251), .Y(n_304) );
INVxp67_ASAP7_75t_L g305 ( .A(n_290), .Y(n_305) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_299), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_297), .B(n_228), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_298), .B(n_255), .Y(n_308) );
AND2x6_ASAP7_75t_SL g309 ( .A(n_289), .B(n_281), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_292), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_292), .B(n_255), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_294), .B(n_172), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_286), .Y(n_313) );
INVxp67_ASAP7_75t_SL g314 ( .A(n_287), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_295), .B(n_174), .Y(n_315) );
INVx8_ASAP7_75t_L g316 ( .A(n_300), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g317 ( .A(n_296), .B(n_180), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_287), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_287), .Y(n_319) );
OAI21xp5_ASAP7_75t_L g320 ( .A1(n_305), .A2(n_282), .B(n_277), .Y(n_320) );
O2A1O1Ixp33_ASAP7_75t_SL g321 ( .A1(n_317), .A2(n_176), .B(n_178), .C(n_175), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g322 ( .A1(n_312), .A2(n_181), .B(n_179), .Y(n_322) );
NAND3xp33_ASAP7_75t_L g323 ( .A(n_301), .B(n_186), .C(n_185), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_303), .Y(n_324) );
AOI21xp5_ASAP7_75t_L g325 ( .A1(n_310), .A2(n_188), .B(n_187), .Y(n_325) );
INVx4_ASAP7_75t_L g326 ( .A(n_316), .Y(n_326) );
O2A1O1Ixp33_ASAP7_75t_SL g327 ( .A1(n_302), .A2(n_197), .B(n_198), .C(n_194), .Y(n_327) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_319), .Y(n_328) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_307), .A2(n_205), .B(n_203), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_308), .B(n_189), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_313), .A2(n_208), .B(n_206), .Y(n_331) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_318), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g333 ( .A1(n_311), .A2(n_210), .B1(n_213), .B2(n_209), .Y(n_333) );
OAI21xp5_ASAP7_75t_L g334 ( .A1(n_315), .A2(n_217), .B(n_214), .Y(n_334) );
O2A1O1Ixp33_ASAP7_75t_L g335 ( .A1(n_304), .A2(n_227), .B(n_231), .C(n_224), .Y(n_335) );
INVx3_ASAP7_75t_L g336 ( .A(n_309), .Y(n_336) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_304), .B(n_192), .Y(n_337) );
AOI21xp5_ASAP7_75t_L g338 ( .A1(n_306), .A2(n_243), .B(n_242), .Y(n_338) );
INVx3_ASAP7_75t_L g339 ( .A(n_306), .Y(n_339) );
AOI22xp5_ASAP7_75t_L g340 ( .A1(n_306), .A2(n_252), .B1(n_253), .B2(n_247), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_314), .Y(n_341) );
OAI21x1_ASAP7_75t_L g342 ( .A1(n_320), .A2(n_260), .B(n_258), .Y(n_342) );
OA21x2_ASAP7_75t_L g343 ( .A1(n_338), .A2(n_254), .B(n_233), .Y(n_343) );
NOR2x1_ASAP7_75t_L g344 ( .A(n_341), .B(n_196), .Y(n_344) );
OAI21xp5_ASAP7_75t_L g345 ( .A1(n_329), .A2(n_219), .B(n_204), .Y(n_345) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_328), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_328), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_334), .B(n_199), .Y(n_348) );
AO31x2_ASAP7_75t_L g349 ( .A1(n_333), .A2(n_236), .A3(n_177), .B(n_273), .Y(n_349) );
AOI221xp5_ASAP7_75t_L g350 ( .A1(n_336), .A2(n_256), .B1(n_223), .B2(n_202), .C(n_207), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_330), .B(n_201), .Y(n_351) );
INVx5_ASAP7_75t_L g352 ( .A(n_326), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_322), .A2(n_212), .B(n_211), .Y(n_353) );
OAI21x1_ASAP7_75t_L g354 ( .A1(n_339), .A2(n_236), .B(n_177), .Y(n_354) );
AO31x2_ASAP7_75t_L g355 ( .A1(n_325), .A2(n_236), .A3(n_275), .B(n_273), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_328), .Y(n_356) );
INVx1_ASAP7_75t_SL g357 ( .A(n_332), .Y(n_357) );
O2A1O1Ixp33_ASAP7_75t_L g358 ( .A1(n_327), .A2(n_262), .B(n_232), .C(n_10), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_324), .Y(n_359) );
INVx2_ASAP7_75t_SL g360 ( .A(n_323), .Y(n_360) );
A2O1A1Ixp33_ASAP7_75t_L g361 ( .A1(n_331), .A2(n_222), .B(n_225), .C(n_220), .Y(n_361) );
AOI21xp5_ASAP7_75t_L g362 ( .A1(n_337), .A2(n_229), .B(n_226), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_335), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_340), .B(n_8), .Y(n_364) );
INVx2_ASAP7_75t_SL g365 ( .A(n_321), .Y(n_365) );
OAI21x1_ASAP7_75t_L g366 ( .A1(n_354), .A2(n_275), .B(n_273), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_359), .Y(n_367) );
OAI21x1_ASAP7_75t_L g368 ( .A1(n_342), .A2(n_275), .B(n_38), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_364), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_344), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_357), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_344), .Y(n_372) );
AND2x4_ASAP7_75t_L g373 ( .A(n_352), .B(n_9), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_363), .B(n_10), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_363), .B(n_11), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_360), .B(n_11), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_345), .B(n_12), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_346), .Y(n_378) );
INVxp67_ASAP7_75t_SL g379 ( .A(n_346), .Y(n_379) );
OAI21x1_ASAP7_75t_L g380 ( .A1(n_347), .A2(n_44), .B(n_43), .Y(n_380) );
OAI21xp5_ASAP7_75t_L g381 ( .A1(n_358), .A2(n_278), .B(n_237), .Y(n_381) );
AO31x2_ASAP7_75t_L g382 ( .A1(n_356), .A2(n_278), .A3(n_16), .B(n_14), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_352), .Y(n_383) );
AOI21xp5_ASAP7_75t_L g384 ( .A1(n_343), .A2(n_278), .B(n_239), .Y(n_384) );
OAI21xp5_ASAP7_75t_L g385 ( .A1(n_343), .A2(n_278), .B(n_240), .Y(n_385) );
INVx1_ASAP7_75t_SL g386 ( .A(n_365), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_349), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_348), .B(n_17), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_361), .B(n_17), .Y(n_389) );
OA21x2_ASAP7_75t_L g390 ( .A1(n_349), .A2(n_241), .B(n_235), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_351), .B(n_18), .Y(n_391) );
OA21x2_ASAP7_75t_L g392 ( .A1(n_349), .A2(n_245), .B(n_244), .Y(n_392) );
OAI21x1_ASAP7_75t_L g393 ( .A1(n_353), .A2(n_49), .B(n_47), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_355), .Y(n_394) );
AOI22x1_ASAP7_75t_L g395 ( .A1(n_362), .A2(n_248), .B1(n_250), .B2(n_246), .Y(n_395) );
OAI21x1_ASAP7_75t_L g396 ( .A1(n_350), .A2(n_53), .B(n_52), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_369), .B(n_20), .Y(n_397) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_371), .Y(n_398) );
AO21x2_ASAP7_75t_L g399 ( .A1(n_384), .A2(n_20), .B(n_21), .Y(n_399) );
AO21x2_ASAP7_75t_L g400 ( .A1(n_384), .A2(n_21), .B(n_22), .Y(n_400) );
OAI21x1_ASAP7_75t_L g401 ( .A1(n_366), .A2(n_57), .B(n_56), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_374), .B(n_23), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_375), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_375), .B(n_23), .Y(n_404) );
OA21x2_ASAP7_75t_L g405 ( .A1(n_385), .A2(n_261), .B(n_259), .Y(n_405) );
OA21x2_ASAP7_75t_L g406 ( .A1(n_387), .A2(n_265), .B(n_58), .Y(n_406) );
OAI21x1_ASAP7_75t_SL g407 ( .A1(n_377), .A2(n_24), .B(n_25), .Y(n_407) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_383), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_378), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_382), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_382), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_376), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_382), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_394), .Y(n_414) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_379), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_390), .Y(n_416) );
AO21x2_ASAP7_75t_L g417 ( .A1(n_381), .A2(n_27), .B(n_28), .Y(n_417) );
AO21x2_ASAP7_75t_L g418 ( .A1(n_368), .A2(n_30), .B(n_31), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_388), .B(n_32), .Y(n_419) );
BUFx4f_ASAP7_75t_L g420 ( .A(n_370), .Y(n_420) );
OAI21x1_ASAP7_75t_L g421 ( .A1(n_380), .A2(n_61), .B(n_60), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_390), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_372), .B(n_386), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_389), .Y(n_424) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_392), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_391), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_392), .Y(n_427) );
HB1xp67_ASAP7_75t_SL g428 ( .A(n_396), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_393), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_395), .Y(n_430) );
OAI21x1_ASAP7_75t_L g431 ( .A1(n_366), .A2(n_65), .B(n_68), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_367), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_371), .Y(n_433) );
INVx3_ASAP7_75t_L g434 ( .A(n_373), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_432), .Y(n_435) );
INVx3_ASAP7_75t_L g436 ( .A(n_420), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_403), .B(n_71), .Y(n_437) );
INVx3_ASAP7_75t_L g438 ( .A(n_420), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_424), .B(n_78), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_409), .Y(n_440) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_408), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_397), .Y(n_442) );
AND2x4_ASAP7_75t_L g443 ( .A(n_434), .B(n_87), .Y(n_443) );
AO21x2_ASAP7_75t_L g444 ( .A1(n_429), .A2(n_90), .B(n_91), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_415), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_397), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_398), .B(n_92), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_398), .B(n_93), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_426), .B(n_94), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_412), .B(n_96), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_433), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_414), .Y(n_452) );
INVx1_ASAP7_75t_SL g453 ( .A(n_433), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_408), .B(n_98), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_423), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_418), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_402), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_402), .B(n_101), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_404), .B(n_103), .Y(n_459) );
OA21x2_ASAP7_75t_L g460 ( .A1(n_410), .A2(n_413), .B(n_411), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_419), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_407), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_399), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_416), .B(n_110), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_399), .B(n_167), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_400), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_400), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_427), .Y(n_468) );
NOR2x1_ASAP7_75t_SL g469 ( .A(n_417), .B(n_113), .Y(n_469) );
AND2x4_ASAP7_75t_SL g470 ( .A(n_430), .B(n_115), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_422), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_405), .B(n_117), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_425), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_425), .Y(n_474) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_406), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_421), .Y(n_476) );
INVx3_ASAP7_75t_L g477 ( .A(n_401), .Y(n_477) );
INVx3_ASAP7_75t_L g478 ( .A(n_431), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_435), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_461), .B(n_122), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_455), .B(n_457), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_453), .B(n_428), .Y(n_482) );
AND2x4_ASAP7_75t_L g483 ( .A(n_445), .B(n_123), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_451), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_452), .B(n_125), .Y(n_485) );
BUFx2_ASAP7_75t_L g486 ( .A(n_441), .Y(n_486) );
AND2x4_ASAP7_75t_L g487 ( .A(n_473), .B(n_127), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_440), .B(n_128), .Y(n_488) );
AND2x4_ASAP7_75t_L g489 ( .A(n_474), .B(n_129), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_442), .B(n_131), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_468), .Y(n_491) );
INVxp67_ASAP7_75t_L g492 ( .A(n_466), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_446), .B(n_132), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_471), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_447), .B(n_448), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_462), .Y(n_496) );
AND2x4_ASAP7_75t_L g497 ( .A(n_436), .B(n_134), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_463), .B(n_137), .Y(n_498) );
BUFx2_ASAP7_75t_L g499 ( .A(n_438), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_467), .B(n_140), .Y(n_500) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_460), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_437), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_456), .B(n_143), .Y(n_503) );
INVx4_ASAP7_75t_L g504 ( .A(n_443), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_476), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_450), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_454), .B(n_151), .Y(n_507) );
AND2x2_ASAP7_75t_SL g508 ( .A(n_470), .B(n_152), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_443), .B(n_154), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_484), .B(n_464), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_481), .B(n_439), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_494), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_479), .B(n_465), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_495), .B(n_472), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_491), .B(n_449), .Y(n_515) );
AND2x4_ASAP7_75t_L g516 ( .A(n_504), .B(n_478), .Y(n_516) );
INVx2_ASAP7_75t_SL g517 ( .A(n_508), .Y(n_517) );
AND2x4_ASAP7_75t_L g518 ( .A(n_482), .B(n_477), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_499), .B(n_475), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_505), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_505), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_486), .B(n_477), .Y(n_522) );
AND2x4_ASAP7_75t_L g523 ( .A(n_496), .B(n_469), .Y(n_523) );
AND2x4_ASAP7_75t_L g524 ( .A(n_492), .B(n_444), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_501), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_502), .B(n_458), .Y(n_526) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_512), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_514), .B(n_506), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_525), .Y(n_529) );
NAND2x1p5_ASAP7_75t_L g530 ( .A(n_517), .B(n_509), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_520), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_510), .B(n_513), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_528), .B(n_526), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_527), .B(n_511), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_532), .B(n_519), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_531), .Y(n_536) );
INVxp67_ASAP7_75t_SL g537 ( .A(n_529), .Y(n_537) );
AOI31xp33_ASAP7_75t_L g538 ( .A1(n_530), .A2(n_516), .A3(n_524), .B(n_523), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_534), .Y(n_539) );
AOI21xp33_ASAP7_75t_L g540 ( .A1(n_538), .A2(n_518), .B(n_524), .Y(n_540) );
INVx1_ASAP7_75t_SL g541 ( .A(n_535), .Y(n_541) );
AOI21xp5_ASAP7_75t_SL g542 ( .A1(n_537), .A2(n_483), .B(n_497), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_542), .A2(n_533), .B(n_536), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_541), .B(n_522), .Y(n_544) );
INVx1_ASAP7_75t_SL g545 ( .A(n_544), .Y(n_545) );
OAI21xp5_ASAP7_75t_SL g546 ( .A1(n_543), .A2(n_540), .B(n_539), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_545), .Y(n_547) );
NOR3xp33_ASAP7_75t_L g548 ( .A(n_546), .B(n_459), .C(n_493), .Y(n_548) );
INVx2_ASAP7_75t_SL g549 ( .A(n_547), .Y(n_549) );
NAND3xp33_ASAP7_75t_L g550 ( .A(n_548), .B(n_490), .C(n_480), .Y(n_550) );
BUFx3_ASAP7_75t_L g551 ( .A(n_549), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_551), .A2(n_550), .B1(n_515), .B2(n_521), .Y(n_552) );
OAI21xp5_ASAP7_75t_L g553 ( .A1(n_552), .A2(n_489), .B(n_487), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_553), .A2(n_483), .B1(n_485), .B2(n_507), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_554), .A2(n_500), .B1(n_498), .B2(n_503), .Y(n_555) );
OAI21xp5_ASAP7_75t_L g556 ( .A1(n_555), .A2(n_500), .B(n_488), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_556), .B(n_155), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_557), .A2(n_156), .B1(n_157), .B2(n_158), .Y(n_558) );
endmodule