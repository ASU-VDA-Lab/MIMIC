module fake_jpeg_8245_n_206 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_206);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_17),
.Y(n_34)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_37),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_24),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_39),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_1),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

HAxp5_ASAP7_75t_SL g46 ( 
.A(n_43),
.B(n_18),
.CON(n_46),
.SN(n_46)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_30),
.Y(n_47)
);

O2A1O1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_46),
.A2(n_34),
.B(n_36),
.C(n_18),
.Y(n_75)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_30),
.B1(n_22),
.B2(n_26),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_48),
.A2(n_49),
.B1(n_50),
.B2(n_61),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_44),
.B1(n_39),
.B2(n_38),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_25),
.B1(n_26),
.B2(n_31),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_52),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_54),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_25),
.Y(n_55)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_34),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_23),
.Y(n_58)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_23),
.Y(n_60)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_43),
.A2(n_16),
.B1(n_32),
.B2(n_31),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_32),
.B1(n_29),
.B2(n_33),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_63),
.A2(n_62),
.B1(n_56),
.B2(n_53),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_34),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_87),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_67),
.A2(n_20),
.B1(n_27),
.B2(n_19),
.Y(n_95)
);

BUFx8_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_68),
.Y(n_110)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_53),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_80),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_21),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_72),
.B(n_78),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_45),
.B(n_2),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_65),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_21),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_81),
.B(n_90),
.Y(n_108)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_88),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_51),
.A2(n_20),
.B1(n_41),
.B2(n_27),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_85),
.A2(n_41),
.B1(n_19),
.B2(n_54),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_27),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_57),
.B(n_2),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_93),
.Y(n_114)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_27),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_19),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_95),
.A2(n_71),
.B1(n_76),
.B2(n_86),
.Y(n_124)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_109),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_4),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_106),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_4),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_66),
.B(n_19),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_107),
.B(n_112),
.Y(n_127)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_87),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_113),
.B(n_74),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_115),
.A2(n_69),
.B1(n_84),
.B2(n_74),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_93),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_4),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_103),
.C(n_96),
.Y(n_132)
);

NOR2xp67_ASAP7_75t_SL g118 ( 
.A(n_103),
.B(n_75),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_118),
.A2(n_134),
.B(n_105),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_133),
.B1(n_113),
.B2(n_101),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_114),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_122),
.B(n_123),
.Y(n_155)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_111),
.B1(n_86),
.B2(n_76),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_125),
.B(n_128),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_126),
.B(n_136),
.Y(n_141)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_131),
.Y(n_144)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_108),
.Y(n_140)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_135),
.Y(n_139)
);

A2O1A1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_105),
.A2(n_73),
.B(n_77),
.C(n_83),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_71),
.Y(n_137)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_89),
.Y(n_138)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_140),
.B(n_119),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_142),
.B(n_147),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_117),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_145),
.C(n_124),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_102),
.C(n_108),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_136),
.B(n_96),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_149),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_123),
.B(n_102),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_130),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_153),
.A2(n_104),
.B1(n_6),
.B2(n_5),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_134),
.A2(n_111),
.B(n_106),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_154),
.A2(n_125),
.B(n_131),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_154),
.A2(n_121),
.B1(n_119),
.B2(n_127),
.Y(n_157)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_164),
.C(n_165),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_166),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_161),
.A2(n_168),
.B(n_159),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_140),
.B(n_106),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_144),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_135),
.C(n_68),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_109),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_167),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_142),
.A2(n_104),
.B1(n_129),
.B2(n_68),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_169),
.A2(n_146),
.B1(n_148),
.B2(n_139),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_153),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_170),
.A2(n_8),
.B(n_10),
.Y(n_181)
);

AO22x1_ASAP7_75t_L g171 ( 
.A1(n_168),
.A2(n_141),
.B1(n_156),
.B2(n_144),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_171),
.A2(n_174),
.B1(n_180),
.B2(n_181),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_12),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_145),
.C(n_139),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_179),
.C(n_6),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_151),
.C(n_8),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_158),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_183),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_161),
.C(n_162),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_163),
.C(n_151),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_185),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_12),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_186),
.A2(n_173),
.B(n_180),
.Y(n_192)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_188),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_15),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_189),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_193),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_186),
.A2(n_177),
.B(n_172),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_190),
.B(n_174),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_196),
.B(n_198),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_188),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_187),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_199),
.A2(n_15),
.B(n_196),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_194),
.C(n_171),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_201),
.Y(n_204)
);

INVxp33_ASAP7_75t_L g203 ( 
.A(n_202),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_200),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_203),
.Y(n_206)
);


endmodule