module fake_aes_9120_n_760 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_760);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_760;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_751;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_420;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_195;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_733;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_723;
wire n_597;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g83 ( .A(n_68), .Y(n_83) );
CKINVDCx16_ASAP7_75t_R g84 ( .A(n_60), .Y(n_84) );
CKINVDCx20_ASAP7_75t_R g85 ( .A(n_6), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_78), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_31), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_64), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_73), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_82), .Y(n_90) );
BUFx3_ASAP7_75t_L g91 ( .A(n_63), .Y(n_91) );
BUFx3_ASAP7_75t_L g92 ( .A(n_4), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_19), .Y(n_93) );
CKINVDCx16_ASAP7_75t_R g94 ( .A(n_42), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_20), .Y(n_95) );
INVx1_ASAP7_75t_SL g96 ( .A(n_9), .Y(n_96) );
INVxp67_ASAP7_75t_SL g97 ( .A(n_76), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_72), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_59), .Y(n_99) );
BUFx6f_ASAP7_75t_L g100 ( .A(n_74), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_3), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_12), .Y(n_102) );
INVx1_ASAP7_75t_SL g103 ( .A(n_28), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_23), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_24), .Y(n_105) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_32), .Y(n_106) );
BUFx3_ASAP7_75t_L g107 ( .A(n_30), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_77), .Y(n_108) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_17), .Y(n_109) );
BUFx2_ASAP7_75t_L g110 ( .A(n_12), .Y(n_110) );
BUFx10_ASAP7_75t_L g111 ( .A(n_13), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_47), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_44), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_9), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_1), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_40), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_37), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_56), .Y(n_118) );
INVx4_ASAP7_75t_R g119 ( .A(n_35), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_6), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_1), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_81), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_0), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_52), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_25), .Y(n_125) );
INVxp67_ASAP7_75t_SL g126 ( .A(n_80), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_29), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_57), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_71), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_33), .Y(n_130) );
BUFx2_ASAP7_75t_SL g131 ( .A(n_39), .Y(n_131) );
BUFx5_ASAP7_75t_L g132 ( .A(n_70), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_15), .Y(n_133) );
INVxp67_ASAP7_75t_L g134 ( .A(n_110), .Y(n_134) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_115), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_92), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_121), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_109), .B(n_0), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_84), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_132), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_121), .Y(n_141) );
AOI22xp5_ASAP7_75t_L g142 ( .A1(n_94), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_106), .B(n_2), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_132), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_132), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_85), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_100), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_113), .Y(n_148) );
AOI22xp5_ASAP7_75t_L g149 ( .A1(n_115), .A2(n_5), .B1(n_7), .B2(n_8), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_92), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_101), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_114), .Y(n_152) );
CKINVDCx16_ASAP7_75t_R g153 ( .A(n_111), .Y(n_153) );
OA21x2_ASAP7_75t_L g154 ( .A1(n_86), .A2(n_43), .B(n_75), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_132), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_83), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_87), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_132), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_133), .B(n_5), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_91), .B(n_7), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_100), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_132), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_88), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_89), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_133), .B(n_8), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_90), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_123), .B(n_10), .Y(n_167) );
OA21x2_ASAP7_75t_L g168 ( .A1(n_86), .A2(n_45), .B(n_69), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_93), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_132), .Y(n_170) );
CKINVDCx6p67_ASAP7_75t_R g171 ( .A(n_91), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_100), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_95), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_100), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_129), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_129), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_98), .B(n_10), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_113), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_105), .Y(n_179) );
AND2x4_ASAP7_75t_L g180 ( .A(n_160), .B(n_107), .Y(n_180) );
BUFx10_ASAP7_75t_L g181 ( .A(n_139), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_136), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_156), .B(n_112), .Y(n_183) );
BUFx3_ASAP7_75t_L g184 ( .A(n_136), .Y(n_184) );
BUFx2_ASAP7_75t_L g185 ( .A(n_139), .Y(n_185) );
OR2x2_ASAP7_75t_L g186 ( .A(n_134), .B(n_96), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_153), .B(n_111), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_136), .Y(n_188) );
INVx3_ASAP7_75t_L g189 ( .A(n_160), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_150), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_160), .Y(n_191) );
AND2x4_ASAP7_75t_L g192 ( .A(n_156), .B(n_107), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_157), .B(n_124), .Y(n_193) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_147), .Y(n_194) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_147), .Y(n_195) );
BUFx3_ASAP7_75t_L g196 ( .A(n_171), .Y(n_196) );
OR2x2_ASAP7_75t_L g197 ( .A(n_135), .B(n_151), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_157), .B(n_112), .Y(n_198) );
AND2x6_ASAP7_75t_L g199 ( .A(n_143), .B(n_124), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_163), .B(n_127), .Y(n_200) );
XNOR2xp5_ASAP7_75t_L g201 ( .A(n_148), .B(n_85), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_152), .Y(n_202) );
NAND3xp33_ASAP7_75t_SL g203 ( .A(n_142), .B(n_122), .C(n_127), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_163), .B(n_104), .Y(n_204) );
BUFx3_ASAP7_75t_L g205 ( .A(n_171), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_137), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_140), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_140), .Y(n_208) );
INVx4_ASAP7_75t_L g209 ( .A(n_154), .Y(n_209) );
NAND2xp33_ASAP7_75t_L g210 ( .A(n_179), .B(n_129), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_137), .Y(n_211) );
INVx4_ASAP7_75t_L g212 ( .A(n_154), .Y(n_212) );
OR2x6_ASAP7_75t_L g213 ( .A(n_143), .B(n_131), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_144), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_144), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_145), .Y(n_216) );
OR2x2_ASAP7_75t_L g217 ( .A(n_138), .B(n_130), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_141), .Y(n_218) );
AND2x6_ASAP7_75t_L g219 ( .A(n_164), .B(n_118), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_164), .B(n_117), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_166), .B(n_116), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_145), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_155), .Y(n_223) );
BUFx2_ASAP7_75t_L g224 ( .A(n_146), .Y(n_224) );
NOR2x1p5_ASAP7_75t_L g225 ( .A(n_148), .B(n_97), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_166), .B(n_111), .Y(n_226) );
AND2x6_ASAP7_75t_L g227 ( .A(n_169), .B(n_128), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_155), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_169), .B(n_99), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_141), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_173), .B(n_126), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_167), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_173), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_158), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_179), .B(n_125), .Y(n_235) );
HB1xp67_ASAP7_75t_L g236 ( .A(n_159), .Y(n_236) );
AND2x6_ASAP7_75t_L g237 ( .A(n_158), .B(n_108), .Y(n_237) );
INVx4_ASAP7_75t_L g238 ( .A(n_154), .Y(n_238) );
AND2x4_ASAP7_75t_L g239 ( .A(n_177), .B(n_129), .Y(n_239) );
INVx4_ASAP7_75t_L g240 ( .A(n_154), .Y(n_240) );
BUFx10_ASAP7_75t_L g241 ( .A(n_178), .Y(n_241) );
INVx4_ASAP7_75t_SL g242 ( .A(n_147), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_162), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_178), .B(n_120), .Y(n_244) );
AND2x4_ASAP7_75t_L g245 ( .A(n_162), .B(n_103), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_170), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_170), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_165), .B(n_122), .Y(n_248) );
INVx2_ASAP7_75t_SL g249 ( .A(n_226), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_232), .B(n_168), .Y(n_250) );
OAI22xp33_ASAP7_75t_L g251 ( .A1(n_213), .A2(n_149), .B1(n_120), .B2(n_102), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_236), .B(n_168), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_236), .B(n_168), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_207), .Y(n_254) );
OAI21xp5_ASAP7_75t_L g255 ( .A1(n_209), .A2(n_168), .B(n_119), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_226), .B(n_102), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_189), .B(n_176), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_182), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_188), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_207), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_181), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_208), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_206), .Y(n_263) );
NAND2x2_ASAP7_75t_L g264 ( .A(n_225), .B(n_11), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_231), .B(n_11), .Y(n_265) );
INVxp67_ASAP7_75t_SL g266 ( .A(n_189), .Y(n_266) );
INVx4_ASAP7_75t_L g267 ( .A(n_189), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_211), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_217), .B(n_50), .Y(n_269) );
NOR2xp67_ASAP7_75t_L g270 ( .A(n_203), .B(n_13), .Y(n_270) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_197), .A2(n_175), .B1(n_174), .B2(n_172), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_187), .B(n_14), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_191), .B(n_175), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_208), .Y(n_274) );
AND2x6_ASAP7_75t_SL g275 ( .A(n_244), .B(n_14), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_218), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_183), .B(n_176), .Y(n_277) );
BUFx6f_ASAP7_75t_SL g278 ( .A(n_196), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_198), .B(n_53), .Y(n_279) );
NOR2xp33_ASAP7_75t_R g280 ( .A(n_196), .B(n_15), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_209), .A2(n_176), .B(n_175), .Y(n_281) );
INVx3_ASAP7_75t_L g282 ( .A(n_184), .Y(n_282) );
INVx4_ASAP7_75t_L g283 ( .A(n_219), .Y(n_283) );
CKINVDCx20_ASAP7_75t_R g284 ( .A(n_201), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_214), .Y(n_285) );
NOR3xp33_ASAP7_75t_SL g286 ( .A(n_248), .B(n_16), .C(n_17), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_230), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_209), .B(n_175), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_200), .B(n_231), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_202), .B(n_16), .Y(n_290) );
BUFx2_ASAP7_75t_L g291 ( .A(n_187), .Y(n_291) );
BUFx6f_ASAP7_75t_L g292 ( .A(n_212), .Y(n_292) );
AND2x4_ASAP7_75t_L g293 ( .A(n_213), .B(n_176), .Y(n_293) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_212), .B(n_176), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_190), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_204), .B(n_174), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_192), .Y(n_297) );
NOR2xp33_ASAP7_75t_SL g298 ( .A(n_205), .B(n_175), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_229), .B(n_174), .Y(n_299) );
OR2x2_ASAP7_75t_SL g300 ( .A(n_186), .B(n_174), .Y(n_300) );
INVxp33_ASAP7_75t_L g301 ( .A(n_185), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_245), .B(n_174), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_192), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_192), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_181), .B(n_161), .Y(n_305) );
BUFx2_ASAP7_75t_L g306 ( .A(n_205), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_245), .B(n_161), .Y(n_307) );
OAI22xp5_ASAP7_75t_SL g308 ( .A1(n_224), .A2(n_172), .B1(n_161), .B2(n_147), .Y(n_308) );
NAND2xp5_ASAP7_75t_SL g309 ( .A(n_212), .B(n_161), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_214), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_245), .B(n_161), .Y(n_311) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_199), .A2(n_172), .B1(n_147), .B2(n_22), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_233), .B(n_172), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_199), .B(n_172), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_184), .Y(n_315) );
AOI22xp5_ASAP7_75t_L g316 ( .A1(n_199), .A2(n_18), .B1(n_21), .B2(n_26), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_199), .A2(n_27), .B1(n_34), .B2(n_36), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_238), .A2(n_38), .B(n_41), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_199), .B(n_46), .Y(n_319) );
BUFx3_ASAP7_75t_L g320 ( .A(n_219), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_181), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_215), .Y(n_322) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_283), .Y(n_323) );
NOR2x1_ASAP7_75t_L g324 ( .A(n_270), .B(n_213), .Y(n_324) );
O2A1O1Ixp5_ASAP7_75t_L g325 ( .A1(n_288), .A2(n_238), .B(n_240), .C(n_193), .Y(n_325) );
BUFx2_ASAP7_75t_L g326 ( .A(n_280), .Y(n_326) );
INVx2_ASAP7_75t_SL g327 ( .A(n_283), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_301), .B(n_213), .Y(n_328) );
A2O1A1Ixp33_ASAP7_75t_L g329 ( .A1(n_250), .A2(n_221), .B(n_235), .C(n_180), .Y(n_329) );
BUFx2_ASAP7_75t_L g330 ( .A(n_280), .Y(n_330) );
OAI22xp5_ASAP7_75t_L g331 ( .A1(n_283), .A2(n_180), .B1(n_239), .B2(n_221), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_292), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_292), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_297), .Y(n_334) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_320), .Y(n_335) );
INVx3_ASAP7_75t_L g336 ( .A(n_267), .Y(n_336) );
INVx3_ASAP7_75t_L g337 ( .A(n_267), .Y(n_337) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_249), .A2(n_180), .B1(n_239), .B2(n_240), .Y(n_338) );
BUFx3_ASAP7_75t_L g339 ( .A(n_320), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_249), .B(n_219), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_303), .Y(n_341) );
OAI22xp33_ASAP7_75t_L g342 ( .A1(n_301), .A2(n_241), .B1(n_220), .B2(n_240), .Y(n_342) );
O2A1O1Ixp33_ASAP7_75t_L g343 ( .A1(n_289), .A2(n_220), .B(n_193), .C(n_247), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_304), .Y(n_344) );
CKINVDCx8_ASAP7_75t_R g345 ( .A(n_275), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_292), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_265), .B(n_227), .Y(n_347) );
CKINVDCx16_ASAP7_75t_R g348 ( .A(n_278), .Y(n_348) );
INVx2_ASAP7_75t_SL g349 ( .A(n_267), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_291), .B(n_241), .Y(n_350) );
BUFx3_ASAP7_75t_L g351 ( .A(n_282), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_261), .Y(n_352) );
INVx2_ASAP7_75t_SL g353 ( .A(n_293), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_265), .B(n_227), .Y(n_354) );
NAND2xp5_ASAP7_75t_SL g355 ( .A(n_292), .B(n_238), .Y(n_355) );
AOI21xp5_ASAP7_75t_L g356 ( .A1(n_288), .A2(n_246), .B(n_215), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_254), .Y(n_357) );
BUFx2_ASAP7_75t_L g358 ( .A(n_256), .Y(n_358) );
AOI211xp5_ASAP7_75t_L g359 ( .A1(n_251), .A2(n_239), .B(n_241), .C(n_210), .Y(n_359) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_282), .Y(n_360) );
INVxp67_ASAP7_75t_L g361 ( .A(n_306), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_295), .B(n_227), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_290), .Y(n_363) );
BUFx2_ASAP7_75t_L g364 ( .A(n_261), .Y(n_364) );
BUFx3_ASAP7_75t_L g365 ( .A(n_282), .Y(n_365) );
BUFx2_ASAP7_75t_L g366 ( .A(n_321), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_263), .B(n_227), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_254), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_260), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_268), .B(n_227), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_276), .B(n_219), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_290), .B(n_219), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_287), .B(n_266), .Y(n_373) );
AOI21xp5_ASAP7_75t_L g374 ( .A1(n_294), .A2(n_246), .B(n_216), .Y(n_374) );
OR2x6_ASAP7_75t_L g375 ( .A(n_272), .B(n_222), .Y(n_375) );
NOR2xp67_ASAP7_75t_SL g376 ( .A(n_321), .B(n_243), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_258), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_260), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_293), .A2(n_237), .B1(n_222), .B2(n_234), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_259), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_363), .B(n_253), .Y(n_381) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_361), .Y(n_382) );
BUFx3_ASAP7_75t_L g383 ( .A(n_323), .Y(n_383) );
OA21x2_ASAP7_75t_L g384 ( .A1(n_329), .A2(n_255), .B(n_318), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_328), .B(n_278), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_358), .A2(n_293), .B1(n_264), .B2(n_278), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g387 ( .A1(n_375), .A2(n_252), .B1(n_300), .B2(n_269), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_358), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_377), .B(n_274), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_352), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_350), .B(n_284), .Y(n_391) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_364), .Y(n_392) );
INVx1_ASAP7_75t_SL g393 ( .A(n_372), .Y(n_393) );
OA21x2_ASAP7_75t_L g394 ( .A1(n_329), .A2(n_281), .B(n_294), .Y(n_394) );
OA21x2_ASAP7_75t_L g395 ( .A1(n_325), .A2(n_309), .B(n_316), .Y(n_395) );
OAI21x1_ASAP7_75t_L g396 ( .A1(n_355), .A2(n_309), .B(n_319), .Y(n_396) );
O2A1O1Ixp33_ASAP7_75t_L g397 ( .A1(n_338), .A2(n_286), .B(n_307), .C(n_302), .Y(n_397) );
OA21x2_ASAP7_75t_L g398 ( .A1(n_355), .A2(n_296), .B(n_299), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_380), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_364), .B(n_322), .Y(n_400) );
OAI21x1_ASAP7_75t_L g401 ( .A1(n_356), .A2(n_314), .B(n_277), .Y(n_401) );
O2A1O1Ixp33_ASAP7_75t_L g402 ( .A1(n_331), .A2(n_311), .B(n_273), .C(n_271), .Y(n_402) );
OAI22xp5_ASAP7_75t_SL g403 ( .A1(n_345), .A2(n_284), .B1(n_264), .B2(n_308), .Y(n_403) );
AND2x4_ASAP7_75t_SL g404 ( .A(n_375), .B(n_305), .Y(n_404) );
INVxp67_ASAP7_75t_SL g405 ( .A(n_335), .Y(n_405) );
OAI21x1_ASAP7_75t_L g406 ( .A1(n_374), .A2(n_317), .B(n_313), .Y(n_406) );
INVx1_ASAP7_75t_SL g407 ( .A(n_366), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_357), .Y(n_408) );
OR2x6_ASAP7_75t_L g409 ( .A(n_375), .B(n_315), .Y(n_409) );
AND2x2_ASAP7_75t_SL g410 ( .A(n_372), .B(n_298), .Y(n_410) );
NAND2x1_ASAP7_75t_L g411 ( .A(n_357), .B(n_322), .Y(n_411) );
OAI21x1_ASAP7_75t_L g412 ( .A1(n_332), .A2(n_279), .B(n_312), .Y(n_412) );
OAI21x1_ASAP7_75t_L g413 ( .A1(n_332), .A2(n_257), .B(n_273), .Y(n_413) );
OAI21x1_ASAP7_75t_L g414 ( .A1(n_333), .A2(n_257), .B(n_285), .Y(n_414) );
OAI21x1_ASAP7_75t_L g415 ( .A1(n_333), .A2(n_310), .B(n_285), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_375), .A2(n_310), .B1(n_274), .B2(n_262), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_407), .B(n_352), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g418 ( .A1(n_411), .A2(n_347), .B(n_354), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_403), .A2(n_326), .B1(n_330), .B2(n_324), .Y(n_419) );
AOI21xp5_ASAP7_75t_L g420 ( .A1(n_411), .A2(n_416), .B(n_384), .Y(n_420) );
OAI221xp5_ASAP7_75t_L g421 ( .A1(n_386), .A2(n_359), .B1(n_345), .B2(n_330), .C(n_326), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_400), .B(n_334), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_381), .B(n_378), .Y(n_423) );
OAI222xp33_ASAP7_75t_L g424 ( .A1(n_409), .A2(n_376), .B1(n_348), .B2(n_342), .C1(n_344), .C2(n_341), .Y(n_424) );
AND2x4_ASAP7_75t_L g425 ( .A(n_399), .B(n_351), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_381), .B(n_378), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_399), .B(n_369), .Y(n_427) );
OAI221xp5_ASAP7_75t_L g428 ( .A1(n_388), .A2(n_403), .B1(n_391), .B2(n_382), .C(n_392), .Y(n_428) );
OAI221xp5_ASAP7_75t_L g429 ( .A1(n_385), .A2(n_373), .B1(n_379), .B2(n_340), .C(n_362), .Y(n_429) );
INVx3_ASAP7_75t_L g430 ( .A(n_383), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_389), .Y(n_431) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_400), .Y(n_432) );
AOI222xp33_ASAP7_75t_L g433 ( .A1(n_390), .A2(n_353), .B1(n_370), .B2(n_367), .C1(n_371), .C2(n_369), .Y(n_433) );
AOI222xp33_ASAP7_75t_L g434 ( .A1(n_390), .A2(n_353), .B1(n_368), .B2(n_337), .C1(n_336), .C2(n_351), .Y(n_434) );
OAI221xp5_ASAP7_75t_L g435 ( .A1(n_397), .A2(n_343), .B1(n_349), .B2(n_336), .C(n_337), .Y(n_435) );
OAI211xp5_ASAP7_75t_SL g436 ( .A1(n_393), .A2(n_210), .B(n_336), .C(n_337), .Y(n_436) );
BUFx2_ASAP7_75t_L g437 ( .A(n_409), .Y(n_437) );
AO21x2_ASAP7_75t_L g438 ( .A1(n_415), .A2(n_346), .B(n_368), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_408), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_408), .Y(n_440) );
AOI21xp5_ASAP7_75t_L g441 ( .A1(n_384), .A2(n_346), .B(n_349), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_393), .B(n_262), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_414), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_384), .B(n_360), .Y(n_444) );
OAI21x1_ASAP7_75t_L g445 ( .A1(n_415), .A2(n_216), .B(n_223), .Y(n_445) );
AO21x2_ASAP7_75t_L g446 ( .A1(n_412), .A2(n_223), .B(n_228), .Y(n_446) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_383), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_423), .B(n_409), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_440), .Y(n_449) );
NOR2x1_ASAP7_75t_L g450 ( .A(n_437), .B(n_409), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_438), .Y(n_451) );
BUFx2_ASAP7_75t_L g452 ( .A(n_437), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_428), .B(n_409), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_423), .B(n_384), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_440), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_439), .Y(n_456) );
BUFx3_ASAP7_75t_L g457 ( .A(n_447), .Y(n_457) );
OAI21xp5_ASAP7_75t_L g458 ( .A1(n_441), .A2(n_444), .B(n_420), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_438), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_439), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_426), .B(n_394), .Y(n_461) );
INVx2_ASAP7_75t_SL g462 ( .A(n_447), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_426), .B(n_427), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_432), .B(n_387), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_427), .B(n_394), .Y(n_465) );
NOR4xp25_ASAP7_75t_SL g466 ( .A(n_421), .B(n_405), .C(n_410), .D(n_395), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_438), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_431), .B(n_394), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_431), .B(n_394), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_425), .B(n_398), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_422), .B(n_404), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_425), .B(n_398), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_444), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_425), .B(n_398), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_422), .B(n_395), .Y(n_475) );
NOR2x1p5_ASAP7_75t_L g476 ( .A(n_430), .B(n_447), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_443), .Y(n_477) );
BUFx2_ASAP7_75t_L g478 ( .A(n_447), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_425), .B(n_404), .Y(n_479) );
INVxp33_ASAP7_75t_SL g480 ( .A(n_417), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_443), .Y(n_481) );
AND2x4_ASAP7_75t_L g482 ( .A(n_430), .B(n_396), .Y(n_482) );
AND2x4_ASAP7_75t_L g483 ( .A(n_430), .B(n_396), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_442), .Y(n_484) );
OAI21xp5_ASAP7_75t_L g485 ( .A1(n_469), .A2(n_424), .B(n_419), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_481), .Y(n_486) );
INVx3_ASAP7_75t_L g487 ( .A(n_457), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_477), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_471), .A2(n_429), .B1(n_435), .B2(n_442), .Y(n_489) );
AOI211xp5_ASAP7_75t_L g490 ( .A1(n_453), .A2(n_436), .B(n_447), .C(n_402), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_463), .B(n_461), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_448), .A2(n_434), .B1(n_433), .B2(n_410), .Y(n_492) );
BUFx2_ASAP7_75t_L g493 ( .A(n_478), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_463), .B(n_434), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_471), .A2(n_410), .B1(n_418), .B2(n_365), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_477), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_473), .B(n_446), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_468), .Y(n_498) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_456), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_448), .A2(n_433), .B1(n_395), .B2(n_365), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_481), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_461), .B(n_446), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_461), .B(n_446), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_468), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_468), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_481), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_473), .B(n_445), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_469), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_456), .Y(n_509) );
AND2x4_ASAP7_75t_L g510 ( .A(n_470), .B(n_445), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_480), .B(n_360), .Y(n_511) );
INVxp67_ASAP7_75t_L g512 ( .A(n_449), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_454), .B(n_398), .Y(n_513) );
BUFx3_ASAP7_75t_L g514 ( .A(n_478), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_449), .B(n_395), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_455), .Y(n_516) );
NAND3xp33_ASAP7_75t_L g517 ( .A(n_455), .B(n_360), .C(n_194), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_465), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_465), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_484), .B(n_237), .Y(n_520) );
OAI33xp33_ASAP7_75t_L g521 ( .A1(n_464), .A2(n_228), .A3(n_234), .B1(n_237), .B2(n_54), .B3(n_55), .Y(n_521) );
INVxp67_ASAP7_75t_SL g522 ( .A(n_460), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_484), .B(n_237), .Y(n_523) );
AND2x4_ASAP7_75t_L g524 ( .A(n_470), .B(n_414), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_460), .Y(n_525) );
INVx5_ASAP7_75t_SL g526 ( .A(n_483), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_454), .B(n_360), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_465), .B(n_401), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_475), .Y(n_529) );
BUFx2_ASAP7_75t_L g530 ( .A(n_472), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_475), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_451), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_472), .B(n_401), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_451), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_474), .B(n_413), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_451), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_491), .B(n_474), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_491), .B(n_464), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_488), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_518), .B(n_467), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_488), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_498), .B(n_452), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_518), .B(n_519), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_519), .B(n_467), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_498), .B(n_452), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_530), .B(n_459), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_530), .B(n_504), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_504), .B(n_467), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_505), .B(n_459), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_496), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_505), .B(n_450), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_502), .B(n_459), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_502), .B(n_483), .Y(n_553) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_499), .Y(n_554) );
AND2x4_ASAP7_75t_L g555 ( .A(n_510), .B(n_483), .Y(n_555) );
NAND4xp25_ASAP7_75t_L g556 ( .A(n_492), .B(n_450), .C(n_458), .D(n_479), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_503), .B(n_483), .Y(n_557) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_522), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_503), .B(n_482), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_496), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_517), .A2(n_466), .B(n_458), .Y(n_561) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_493), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_516), .Y(n_563) );
NAND3xp33_ASAP7_75t_SL g564 ( .A(n_511), .B(n_466), .C(n_479), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_516), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_533), .B(n_482), .Y(n_566) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_509), .B(n_482), .Y(n_567) );
NAND2xp33_ASAP7_75t_SL g568 ( .A(n_494), .B(n_476), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_533), .B(n_482), .Y(n_569) );
OAI33xp33_ASAP7_75t_L g570 ( .A1(n_512), .A2(n_476), .A3(n_49), .B1(n_51), .B2(n_58), .B3(n_61), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_528), .B(n_462), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_528), .B(n_462), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_513), .B(n_462), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_513), .B(n_457), .Y(n_574) );
AND2x4_ASAP7_75t_L g575 ( .A(n_510), .B(n_457), .Y(n_575) );
INVx3_ASAP7_75t_L g576 ( .A(n_526), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_535), .B(n_406), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_535), .B(n_406), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_529), .B(n_412), .Y(n_579) );
AOI31xp33_ASAP7_75t_L g580 ( .A1(n_500), .A2(n_327), .A3(n_62), .B(n_65), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_534), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_529), .B(n_48), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_531), .B(n_66), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_531), .B(n_67), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_509), .B(n_237), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_525), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_508), .B(n_506), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_534), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_508), .B(n_79), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_506), .B(n_413), .Y(n_590) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_493), .Y(n_591) );
AND2x4_ASAP7_75t_L g592 ( .A(n_510), .B(n_242), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_525), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_497), .B(n_194), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_536), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_486), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_486), .B(n_194), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_501), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_554), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_547), .B(n_497), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_538), .B(n_485), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_537), .B(n_510), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_543), .B(n_501), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_537), .B(n_524), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_543), .B(n_532), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_539), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_539), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_547), .B(n_532), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_541), .Y(n_609) );
NAND2x1p5_ASAP7_75t_L g610 ( .A(n_576), .B(n_514), .Y(n_610) );
NAND2x1p5_ASAP7_75t_L g611 ( .A(n_576), .B(n_514), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_587), .B(n_527), .Y(n_612) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_558), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_556), .A2(n_521), .B1(n_489), .B2(n_524), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_581), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_552), .B(n_524), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_581), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_541), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_588), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_552), .B(n_524), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_546), .B(n_507), .Y(n_621) );
NOR4xp25_ASAP7_75t_L g622 ( .A(n_556), .B(n_495), .C(n_520), .D(n_523), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_553), .B(n_526), .Y(n_623) );
OR2x2_ASAP7_75t_L g624 ( .A(n_546), .B(n_507), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_553), .B(n_526), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_587), .B(n_527), .Y(n_626) );
NOR2x1_ASAP7_75t_L g627 ( .A(n_580), .B(n_517), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_550), .B(n_514), .Y(n_628) );
INVx1_ASAP7_75t_SL g629 ( .A(n_574), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_550), .B(n_536), .Y(n_630) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_562), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_560), .Y(n_632) );
NAND2xp5_ASAP7_75t_SL g633 ( .A(n_568), .B(n_487), .Y(n_633) );
AO21x1_ASAP7_75t_L g634 ( .A1(n_560), .A2(n_490), .B(n_515), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_563), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g636 ( .A(n_576), .B(n_487), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_563), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_557), .B(n_526), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_565), .B(n_490), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_557), .B(n_487), .Y(n_640) );
OR2x2_ASAP7_75t_SL g641 ( .A(n_591), .B(n_323), .Y(n_641) );
BUFx3_ASAP7_75t_L g642 ( .A(n_575), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_565), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_586), .Y(n_644) );
INVxp67_ASAP7_75t_SL g645 ( .A(n_588), .Y(n_645) );
OR2x2_ASAP7_75t_L g646 ( .A(n_549), .B(n_194), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_559), .B(n_195), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_559), .B(n_195), .Y(n_648) );
AO21x1_ASAP7_75t_SL g649 ( .A1(n_586), .A2(n_242), .B(n_323), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_595), .Y(n_650) );
OAI21xp5_ASAP7_75t_L g651 ( .A1(n_582), .A2(n_327), .B(n_339), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_566), .B(n_195), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_566), .B(n_195), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_540), .B(n_242), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_601), .B(n_639), .Y(n_655) );
NOR2x1_ASAP7_75t_L g656 ( .A(n_627), .B(n_564), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_613), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_599), .B(n_544), .Y(n_658) );
OAI21xp33_ASAP7_75t_L g659 ( .A1(n_602), .A2(n_569), .B(n_572), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_631), .B(n_551), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_605), .B(n_544), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_618), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_608), .Y(n_663) );
INVxp67_ASAP7_75t_SL g664 ( .A(n_645), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g665 ( .A1(n_634), .A2(n_572), .B1(n_571), .B2(n_555), .Y(n_665) );
AOI21xp33_ASAP7_75t_L g666 ( .A1(n_634), .A2(n_542), .B(n_545), .Y(n_666) );
INVxp67_ASAP7_75t_L g667 ( .A(n_644), .Y(n_667) );
OAI33xp33_ASAP7_75t_L g668 ( .A1(n_608), .A2(n_567), .A3(n_549), .B1(n_593), .B2(n_585), .B3(n_598), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_618), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_629), .B(n_569), .Y(n_670) );
NOR3xp33_ASAP7_75t_L g671 ( .A(n_652), .B(n_570), .C(n_584), .Y(n_671) );
AOI21x1_ASAP7_75t_L g672 ( .A1(n_633), .A2(n_561), .B(n_589), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_643), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g674 ( .A1(n_614), .A2(n_622), .B1(n_653), .B2(n_652), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_643), .Y(n_675) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_621), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_641), .A2(n_555), .B1(n_575), .B2(n_571), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_606), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_602), .B(n_555), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_612), .B(n_626), .Y(n_680) );
INVx1_ASAP7_75t_SL g681 ( .A(n_641), .Y(n_681) );
NAND3xp33_ASAP7_75t_L g682 ( .A(n_644), .B(n_593), .C(n_579), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_640), .A2(n_555), .B1(n_575), .B2(n_573), .Y(n_683) );
OAI21xp33_ASAP7_75t_L g684 ( .A1(n_604), .A2(n_540), .B(n_573), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_607), .Y(n_685) );
OAI22xp33_ASAP7_75t_L g686 ( .A1(n_610), .A2(n_598), .B1(n_596), .B2(n_583), .Y(n_686) );
OAI21xp5_ASAP7_75t_L g687 ( .A1(n_651), .A2(n_582), .B(n_584), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_604), .B(n_574), .Y(n_688) );
O2A1O1Ixp33_ASAP7_75t_L g689 ( .A1(n_636), .A2(n_583), .B(n_589), .C(n_594), .Y(n_689) );
OAI21xp33_ASAP7_75t_SL g690 ( .A1(n_623), .A2(n_596), .B(n_548), .Y(n_690) );
NAND2xp33_ASAP7_75t_SL g691 ( .A(n_623), .B(n_575), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g692 ( .A1(n_610), .A2(n_592), .B(n_579), .Y(n_692) );
INVxp67_ASAP7_75t_SL g693 ( .A(n_646), .Y(n_693) );
AO22x1_ASAP7_75t_L g694 ( .A1(n_642), .A2(n_592), .B1(n_548), .B2(n_595), .Y(n_694) );
INVxp67_ASAP7_75t_SL g695 ( .A(n_664), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_676), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_664), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_679), .B(n_642), .Y(n_698) );
NAND2xp5_ASAP7_75t_SL g699 ( .A(n_690), .B(n_610), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_667), .Y(n_700) );
INVx1_ASAP7_75t_SL g701 ( .A(n_657), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_667), .Y(n_702) );
AND2x2_ASAP7_75t_L g703 ( .A(n_688), .B(n_620), .Y(n_703) );
XOR2x2_ASAP7_75t_L g704 ( .A(n_656), .B(n_611), .Y(n_704) );
AOI211xp5_ASAP7_75t_L g705 ( .A1(n_666), .A2(n_640), .B(n_625), .C(n_638), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_662), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_669), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_655), .B(n_603), .Y(n_708) );
INVx3_ASAP7_75t_L g709 ( .A(n_681), .Y(n_709) );
NOR2xp67_ASAP7_75t_L g710 ( .A(n_672), .B(n_625), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_673), .Y(n_711) );
NAND2xp5_ASAP7_75t_SL g712 ( .A(n_665), .B(n_611), .Y(n_712) );
O2A1O1Ixp33_ASAP7_75t_SL g713 ( .A1(n_677), .A2(n_600), .B(n_628), .C(n_621), .Y(n_713) );
AO22x1_ASAP7_75t_L g714 ( .A1(n_687), .A2(n_638), .B1(n_616), .B2(n_620), .Y(n_714) );
AOI32xp33_ASAP7_75t_L g715 ( .A1(n_691), .A2(n_616), .A3(n_653), .B1(n_647), .B2(n_648), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_674), .A2(n_600), .B1(n_609), .B2(n_632), .Y(n_716) );
AOI32xp33_ASAP7_75t_L g717 ( .A1(n_670), .A2(n_648), .A3(n_647), .B1(n_624), .B2(n_635), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_663), .B(n_637), .Y(n_718) );
AND2x2_ASAP7_75t_L g719 ( .A(n_683), .B(n_624), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g720 ( .A1(n_710), .A2(n_659), .B1(n_684), .B2(n_680), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_708), .B(n_660), .Y(n_721) );
AOI21xp33_ASAP7_75t_L g722 ( .A1(n_716), .A2(n_693), .B(n_689), .Y(n_722) );
INVx1_ASAP7_75t_SL g723 ( .A(n_701), .Y(n_723) );
OA22x2_ASAP7_75t_L g724 ( .A1(n_699), .A2(n_658), .B1(n_693), .B2(n_694), .Y(n_724) );
OAI22xp33_ASAP7_75t_L g725 ( .A1(n_699), .A2(n_686), .B1(n_611), .B2(n_692), .Y(n_725) );
OAI21xp33_ASAP7_75t_L g726 ( .A1(n_704), .A2(n_661), .B(n_671), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_696), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_706), .Y(n_728) );
AOI21xp33_ASAP7_75t_L g729 ( .A1(n_695), .A2(n_682), .B(n_685), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_707), .Y(n_730) );
AOI332xp33_ASAP7_75t_L g731 ( .A1(n_709), .A2(n_678), .A3(n_675), .B1(n_617), .B2(n_650), .B3(n_619), .C1(n_615), .C2(n_578), .Y(n_731) );
OAI21xp33_ASAP7_75t_SL g732 ( .A1(n_712), .A2(n_668), .B(n_630), .Y(n_732) );
NAND2xp33_ASAP7_75t_R g733 ( .A(n_709), .B(n_592), .Y(n_733) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_719), .B(n_668), .Y(n_734) );
AOI221xp5_ASAP7_75t_L g735 ( .A1(n_732), .A2(n_713), .B1(n_695), .B2(n_712), .C(n_717), .Y(n_735) );
INVxp67_ASAP7_75t_L g736 ( .A(n_723), .Y(n_736) );
NOR2x1_ASAP7_75t_L g737 ( .A(n_725), .B(n_697), .Y(n_737) );
OAI311xp33_ASAP7_75t_L g738 ( .A1(n_726), .A2(n_715), .A3(n_704), .B1(n_702), .C1(n_700), .Y(n_738) );
AOI221x1_ASAP7_75t_L g739 ( .A1(n_720), .A2(n_734), .B1(n_722), .B2(n_729), .C(n_727), .Y(n_739) );
OAI211xp5_ASAP7_75t_SL g740 ( .A1(n_724), .A2(n_705), .B(n_713), .C(n_697), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_724), .A2(n_698), .B1(n_703), .B2(n_718), .Y(n_741) );
AOI21xp5_ASAP7_75t_L g742 ( .A1(n_721), .A2(n_714), .B(n_711), .Y(n_742) );
AOI222xp33_ASAP7_75t_L g743 ( .A1(n_728), .A2(n_578), .B1(n_577), .B2(n_650), .C1(n_615), .C2(n_619), .Y(n_743) );
NOR3xp33_ASAP7_75t_L g744 ( .A(n_740), .B(n_730), .C(n_671), .Y(n_744) );
AND2x4_ASAP7_75t_L g745 ( .A(n_736), .B(n_592), .Y(n_745) );
NOR2xp67_ASAP7_75t_L g746 ( .A(n_741), .B(n_733), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_737), .Y(n_747) );
NAND4xp75_ASAP7_75t_L g748 ( .A(n_739), .B(n_731), .C(n_654), .D(n_577), .Y(n_748) );
NAND3xp33_ASAP7_75t_SL g749 ( .A(n_744), .B(n_735), .C(n_742), .Y(n_749) );
AND2x4_ASAP7_75t_L g750 ( .A(n_745), .B(n_617), .Y(n_750) );
AND2x2_ASAP7_75t_L g751 ( .A(n_746), .B(n_743), .Y(n_751) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_751), .Y(n_752) );
AOI21xp33_ASAP7_75t_SL g753 ( .A1(n_749), .A2(n_747), .B(n_738), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_752), .A2(n_750), .B1(n_748), .B2(n_646), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_753), .Y(n_755) );
BUFx2_ASAP7_75t_SL g756 ( .A(n_755), .Y(n_756) );
AOI22xp33_ASAP7_75t_R g757 ( .A1(n_754), .A2(n_750), .B1(n_649), .B2(n_594), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_756), .Y(n_758) );
AOI322xp5_ASAP7_75t_L g759 ( .A1(n_758), .A2(n_757), .A3(n_597), .B1(n_649), .B2(n_339), .C1(n_335), .C2(n_323), .Y(n_759) );
AOI222xp33_ASAP7_75t_L g760 ( .A1(n_759), .A2(n_335), .B1(n_590), .B2(n_597), .C1(n_749), .C2(n_758), .Y(n_760) );
endmodule