module fake_netlist_6_4642_n_781 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_781);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_781;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_760;
wire n_741;
wire n_680;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_726;
wire n_671;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_685;
wire n_597;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_156;
wire n_491;
wire n_656;
wire n_772;
wire n_666;
wire n_371;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_731;
wire n_570;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_683;
wire n_620;
wire n_420;
wire n_608;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

BUFx10_ASAP7_75t_L g155 ( 
.A(n_22),
.Y(n_155)
);

BUFx10_ASAP7_75t_L g156 ( 
.A(n_35),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_48),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_57),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_112),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_88),
.Y(n_161)
);

BUFx10_ASAP7_75t_L g162 ( 
.A(n_41),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_36),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_100),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_4),
.Y(n_167)
);

BUFx2_ASAP7_75t_SL g168 ( 
.A(n_58),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_101),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_125),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_37),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_109),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_117),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_40),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_91),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_144),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_27),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_114),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_12),
.B(n_93),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_59),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_133),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_84),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_150),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_44),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_46),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_50),
.Y(n_186)
);

BUFx10_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_64),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_45),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_111),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_146),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_6),
.B(n_78),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_147),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_89),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_26),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_39),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_87),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_90),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_65),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_69),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_81),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_21),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_131),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_128),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_3),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_122),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_6),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_134),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_33),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_145),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_148),
.Y(n_211)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_155),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_205),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_206),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_167),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_206),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_171),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_157),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_161),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_164),
.Y(n_221)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_155),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_160),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_160),
.Y(n_224)
);

OAI22x1_ASAP7_75t_R g225 ( 
.A1(n_182),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_156),
.Y(n_226)
);

AND2x4_ASAP7_75t_L g227 ( 
.A(n_175),
.B(n_3),
.Y(n_227)
);

BUFx12f_ASAP7_75t_L g228 ( 
.A(n_156),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_175),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_179),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_230)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_161),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_165),
.Y(n_232)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_162),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_166),
.Y(n_234)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_162),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_179),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_236)
);

AND2x4_ASAP7_75t_L g237 ( 
.A(n_184),
.B(n_18),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_192),
.Y(n_238)
);

OAI22x1_ASAP7_75t_SL g239 ( 
.A1(n_182),
.A2(n_197),
.B1(n_209),
.B2(n_194),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_170),
.Y(n_240)
);

AND2x4_ASAP7_75t_L g241 ( 
.A(n_174),
.B(n_8),
.Y(n_241)
);

AND2x4_ASAP7_75t_L g242 ( 
.A(n_176),
.B(n_9),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_187),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_177),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_178),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_187),
.B(n_9),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_209),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_180),
.Y(n_248)
);

BUFx12f_ASAP7_75t_L g249 ( 
.A(n_158),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_191),
.B(n_10),
.Y(n_250)
);

BUFx8_ASAP7_75t_SL g251 ( 
.A(n_197),
.Y(n_251)
);

INVx5_ASAP7_75t_L g252 ( 
.A(n_168),
.Y(n_252)
);

AND2x4_ASAP7_75t_L g253 ( 
.A(n_185),
.B(n_19),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_159),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_R g255 ( 
.A(n_220),
.B(n_163),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_251),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_229),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_229),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_229),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_251),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_215),
.Y(n_261)
);

NOR2x1p5_ASAP7_75t_L g262 ( 
.A(n_233),
.B(n_228),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_229),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_232),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_214),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_249),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_249),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_220),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_215),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_R g270 ( 
.A(n_247),
.B(n_169),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_R g271 ( 
.A(n_247),
.B(n_172),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_232),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_228),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_214),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_231),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_223),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_231),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_226),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_233),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_226),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_234),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_238),
.B(n_188),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_243),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_238),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_243),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_234),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_225),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_239),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_240),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_212),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_212),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_222),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_222),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_240),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_223),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_222),
.Y(n_296)
);

BUFx16f_ASAP7_75t_R g297 ( 
.A(n_227),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_222),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_224),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_235),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_235),
.Y(n_301)
);

AOI221xp5_ASAP7_75t_L g302 ( 
.A1(n_282),
.A2(n_250),
.B1(n_213),
.B2(n_236),
.C(n_230),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_257),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_263),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_276),
.B(n_253),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_265),
.B(n_235),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_259),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_263),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_276),
.B(n_253),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_275),
.B(n_235),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_279),
.B(n_246),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_277),
.B(n_217),
.Y(n_312)
);

NAND2xp33_ASAP7_75t_L g313 ( 
.A(n_270),
.B(n_173),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_265),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_274),
.B(n_252),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_271),
.B(n_252),
.Y(n_316)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_255),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_278),
.B(n_217),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_258),
.Y(n_319)
);

BUFx5_ASAP7_75t_L g320 ( 
.A(n_295),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_299),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_280),
.B(n_252),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_299),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_264),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_283),
.B(n_250),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_272),
.B(n_253),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_258),
.B(n_237),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_281),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_261),
.B(n_213),
.Y(n_329)
);

BUFx6f_ASAP7_75t_SL g330 ( 
.A(n_297),
.Y(n_330)
);

NAND2xp33_ASAP7_75t_L g331 ( 
.A(n_290),
.B(n_181),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_258),
.B(n_237),
.Y(n_332)
);

NAND2x1_ASAP7_75t_L g333 ( 
.A(n_258),
.B(n_237),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_285),
.B(n_219),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_286),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_291),
.B(n_241),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_289),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_293),
.B(n_227),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_292),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_269),
.B(n_241),
.Y(n_340)
);

AO221x1_ASAP7_75t_L g341 ( 
.A1(n_294),
.A2(n_189),
.B1(n_208),
.B2(n_210),
.C(n_201),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_296),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_300),
.B(n_242),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_301),
.B(n_242),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_298),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_262),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_273),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_266),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_267),
.B(n_224),
.Y(n_349)
);

BUFx6f_ASAP7_75t_SL g350 ( 
.A(n_260),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_268),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_284),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_288),
.B(n_183),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_284),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_287),
.B(n_245),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_287),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_256),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_256),
.B(n_245),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_258),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_276),
.B(n_245),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_257),
.Y(n_361)
);

NOR2xp67_ASAP7_75t_L g362 ( 
.A(n_261),
.B(n_186),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_276),
.B(n_245),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_275),
.B(n_190),
.Y(n_364)
);

OA22x2_ASAP7_75t_L g365 ( 
.A1(n_338),
.A2(n_218),
.B1(n_254),
.B2(n_216),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_324),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_317),
.B(n_193),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_R g368 ( 
.A(n_313),
.B(n_198),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_359),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_329),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_311),
.B(n_195),
.Y(n_371)
);

INVx5_ASAP7_75t_L g372 ( 
.A(n_359),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_321),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_325),
.B(n_199),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_305),
.A2(n_221),
.B(n_244),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_334),
.B(n_248),
.Y(n_376)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_359),
.Y(n_377)
);

BUFx8_ASAP7_75t_L g378 ( 
.A(n_330),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_340),
.B(n_312),
.Y(n_379)
);

NAND2x1p5_ASAP7_75t_L g380 ( 
.A(n_339),
.B(n_196),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_323),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g382 ( 
.A(n_314),
.B(n_200),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_328),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_335),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_337),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_326),
.B(n_204),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_364),
.B(n_202),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_302),
.A2(n_336),
.B1(n_343),
.B2(n_326),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_305),
.B(n_248),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_349),
.B(n_203),
.Y(n_390)
);

AND2x4_ASAP7_75t_L g391 ( 
.A(n_345),
.B(n_211),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_R g392 ( 
.A(n_348),
.B(n_20),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_333),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_362),
.A2(n_318),
.B1(n_344),
.B2(n_309),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_304),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_349),
.B(n_248),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_308),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_309),
.Y(n_398)
);

BUFx12f_ASAP7_75t_L g399 ( 
.A(n_342),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_303),
.Y(n_400)
);

NAND3xp33_ASAP7_75t_L g401 ( 
.A(n_322),
.B(n_248),
.C(n_13),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_327),
.B(n_23),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_316),
.B(n_11),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_307),
.Y(n_404)
);

AND2x4_ASAP7_75t_L g405 ( 
.A(n_306),
.B(n_24),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_332),
.B(n_25),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_360),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g408 ( 
.A(n_352),
.B(n_13),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_360),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_358),
.B(n_14),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_361),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_363),
.Y(n_412)
);

INVx5_ASAP7_75t_L g413 ( 
.A(n_319),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_363),
.Y(n_414)
);

INVx5_ASAP7_75t_L g415 ( 
.A(n_319),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_355),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_358),
.B(n_14),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_320),
.B(n_28),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_350),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_310),
.B(n_15),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_355),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_320),
.B(n_29),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_320),
.B(n_30),
.Y(n_423)
);

BUFx3_ASAP7_75t_L g424 ( 
.A(n_351),
.Y(n_424)
);

INVx5_ASAP7_75t_L g425 ( 
.A(n_341),
.Y(n_425)
);

NAND2xp33_ASAP7_75t_SL g426 ( 
.A(n_346),
.B(n_15),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_320),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_L g428 ( 
.A1(n_320),
.A2(n_16),
.B1(n_17),
.B2(n_31),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_L g429 ( 
.A1(n_315),
.A2(n_16),
.B1(n_17),
.B2(n_32),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_353),
.B(n_34),
.Y(n_430)
);

INVx2_ASAP7_75t_SL g431 ( 
.A(n_354),
.Y(n_431)
);

OR2x2_ASAP7_75t_L g432 ( 
.A(n_356),
.B(n_38),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_331),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_416),
.B(n_421),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_398),
.A2(n_347),
.B(n_357),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_388),
.A2(n_374),
.B1(n_394),
.B2(n_433),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_389),
.A2(n_42),
.B(n_43),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_396),
.B(n_47),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_373),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_376),
.B(n_330),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_366),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_383),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_390),
.B(n_49),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_407),
.A2(n_350),
.B1(n_52),
.B2(n_53),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_409),
.A2(n_51),
.B1(n_54),
.B2(n_55),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_412),
.B(n_56),
.Y(n_446)
);

OAI21x1_ASAP7_75t_L g447 ( 
.A1(n_402),
.A2(n_60),
.B(n_61),
.Y(n_447)
);

BUFx12f_ASAP7_75t_L g448 ( 
.A(n_399),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_419),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_381),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_410),
.B(n_62),
.Y(n_451)
);

O2A1O1Ixp33_ASAP7_75t_L g452 ( 
.A1(n_417),
.A2(n_63),
.B(n_66),
.C(n_67),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_369),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_414),
.A2(n_68),
.B(n_70),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_384),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_386),
.A2(n_71),
.B(n_72),
.Y(n_456)
);

INVx5_ASAP7_75t_L g457 ( 
.A(n_369),
.Y(n_457)
);

OAI22xp33_ASAP7_75t_L g458 ( 
.A1(n_365),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_371),
.B(n_76),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_385),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_406),
.A2(n_77),
.B(n_79),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_379),
.B(n_80),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_387),
.B(n_82),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_395),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_370),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_R g466 ( 
.A(n_431),
.B(n_83),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_372),
.A2(n_427),
.B(n_377),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_397),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_391),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_400),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g471 ( 
.A(n_424),
.B(n_85),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_391),
.B(n_86),
.Y(n_472)
);

A2O1A1Ixp33_ASAP7_75t_L g473 ( 
.A1(n_430),
.A2(n_92),
.B(n_94),
.C(n_95),
.Y(n_473)
);

OR2x6_ASAP7_75t_L g474 ( 
.A(n_432),
.B(n_96),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_408),
.Y(n_475)
);

A2O1A1Ixp33_ASAP7_75t_L g476 ( 
.A1(n_405),
.A2(n_97),
.B(n_98),
.C(n_99),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_367),
.B(n_102),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_375),
.B(n_103),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_378),
.Y(n_479)
);

OAI21xp33_ASAP7_75t_L g480 ( 
.A1(n_429),
.A2(n_104),
.B(n_105),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_393),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_393),
.A2(n_110),
.B1(n_113),
.B2(n_115),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_392),
.B(n_116),
.Y(n_483)
);

A2O1A1Ixp33_ASAP7_75t_L g484 ( 
.A1(n_405),
.A2(n_118),
.B(n_120),
.C(n_121),
.Y(n_484)
);

INVx4_ASAP7_75t_L g485 ( 
.A(n_369),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_393),
.B(n_411),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_404),
.Y(n_487)
);

AO22x1_ASAP7_75t_L g488 ( 
.A1(n_420),
.A2(n_123),
.B1(n_124),
.B2(n_126),
.Y(n_488)
);

NOR2xp67_ASAP7_75t_SL g489 ( 
.A(n_372),
.B(n_127),
.Y(n_489)
);

OAI21x1_ASAP7_75t_L g490 ( 
.A1(n_447),
.A2(n_423),
.B(n_422),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_436),
.A2(n_418),
.B(n_372),
.Y(n_491)
);

INVx5_ASAP7_75t_SL g492 ( 
.A(n_474),
.Y(n_492)
);

AO21x2_ASAP7_75t_L g493 ( 
.A1(n_443),
.A2(n_459),
.B(n_463),
.Y(n_493)
);

CKINVDCx6p67_ASAP7_75t_R g494 ( 
.A(n_448),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_438),
.A2(n_377),
.B(n_428),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_465),
.Y(n_496)
);

OAI21x1_ASAP7_75t_L g497 ( 
.A1(n_467),
.A2(n_380),
.B(n_403),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_441),
.Y(n_498)
);

OAI21x1_ASAP7_75t_L g499 ( 
.A1(n_446),
.A2(n_401),
.B(n_415),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_434),
.B(n_382),
.Y(n_500)
);

OR2x6_ASAP7_75t_L g501 ( 
.A(n_474),
.B(n_382),
.Y(n_501)
);

INVx8_ASAP7_75t_L g502 ( 
.A(n_457),
.Y(n_502)
);

INVx5_ASAP7_75t_L g503 ( 
.A(n_453),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_455),
.B(n_425),
.Y(n_504)
);

BUFx12f_ASAP7_75t_L g505 ( 
.A(n_449),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_453),
.Y(n_506)
);

AO21x2_ASAP7_75t_L g507 ( 
.A1(n_456),
.A2(n_368),
.B(n_425),
.Y(n_507)
);

BUFx2_ASAP7_75t_R g508 ( 
.A(n_479),
.Y(n_508)
);

OAI21x1_ASAP7_75t_L g509 ( 
.A1(n_462),
.A2(n_415),
.B(n_413),
.Y(n_509)
);

OAI21x1_ASAP7_75t_L g510 ( 
.A1(n_486),
.A2(n_413),
.B(n_425),
.Y(n_510)
);

OAI21x1_ASAP7_75t_L g511 ( 
.A1(n_478),
.A2(n_129),
.B(n_130),
.Y(n_511)
);

OAI21x1_ASAP7_75t_L g512 ( 
.A1(n_454),
.A2(n_132),
.B(n_135),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_442),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_460),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_468),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_453),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_466),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_451),
.A2(n_426),
.B(n_137),
.Y(n_518)
);

AO21x1_ASAP7_75t_SL g519 ( 
.A1(n_480),
.A2(n_136),
.B(n_138),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_457),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_457),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_480),
.A2(n_139),
.B(n_141),
.Y(n_522)
);

OAI21x1_ASAP7_75t_L g523 ( 
.A1(n_456),
.A2(n_142),
.B(n_149),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_470),
.Y(n_524)
);

NAND2x1p5_ASAP7_75t_L g525 ( 
.A(n_485),
.B(n_151),
.Y(n_525)
);

INVx1_ASAP7_75t_SL g526 ( 
.A(n_475),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_474),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_475),
.B(n_152),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_435),
.A2(n_154),
.B(n_378),
.Y(n_529)
);

INVx5_ASAP7_75t_L g530 ( 
.A(n_485),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_472),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_487),
.Y(n_532)
);

AO21x2_ASAP7_75t_L g533 ( 
.A1(n_473),
.A2(n_458),
.B(n_476),
.Y(n_533)
);

NAND2x1p5_ASAP7_75t_L g534 ( 
.A(n_487),
.B(n_489),
.Y(n_534)
);

AO21x2_ASAP7_75t_L g535 ( 
.A1(n_484),
.A2(n_437),
.B(n_461),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_471),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_464),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_439),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_522),
.A2(n_477),
.B1(n_469),
.B2(n_440),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_502),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_498),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_513),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_530),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_L g544 ( 
.A1(n_495),
.A2(n_450),
.B(n_452),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_500),
.B(n_444),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_SL g546 ( 
.A1(n_529),
.A2(n_481),
.B(n_482),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_530),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_514),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_515),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_503),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_526),
.B(n_483),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_531),
.B(n_488),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_504),
.A2(n_445),
.B1(n_501),
.B2(n_533),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_L g554 ( 
.A1(n_518),
.A2(n_536),
.B1(n_527),
.B2(n_538),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_537),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_524),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_L g557 ( 
.A1(n_536),
.A2(n_527),
.B1(n_538),
.B2(n_533),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_523),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_510),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_502),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_531),
.B(n_519),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_532),
.Y(n_562)
);

OR2x6_ASAP7_75t_L g563 ( 
.A(n_501),
.B(n_534),
.Y(n_563)
);

OAI21x1_ASAP7_75t_L g564 ( 
.A1(n_509),
.A2(n_490),
.B(n_491),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_532),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_516),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_512),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_516),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_531),
.A2(n_504),
.B1(n_507),
.B2(n_501),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_530),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_496),
.Y(n_571)
);

CKINVDCx6p67_ASAP7_75t_R g572 ( 
.A(n_505),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_511),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_531),
.A2(n_517),
.B1(n_492),
.B2(n_495),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_516),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_520),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_516),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_534),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_504),
.A2(n_507),
.B1(n_528),
.B2(n_492),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_530),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_521),
.Y(n_581)
);

OR2x6_ASAP7_75t_L g582 ( 
.A(n_563),
.B(n_525),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_SL g583 ( 
.A1(n_545),
.A2(n_492),
.B1(n_523),
.B2(n_517),
.Y(n_583)
);

OR2x6_ASAP7_75t_L g584 ( 
.A(n_563),
.B(n_561),
.Y(n_584)
);

INVx4_ASAP7_75t_L g585 ( 
.A(n_540),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_541),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_574),
.B(n_508),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_541),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_548),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_542),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_542),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_539),
.A2(n_503),
.B1(n_525),
.B2(n_520),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_572),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_549),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_571),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_572),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_R g597 ( 
.A(n_540),
.B(n_505),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_545),
.B(n_506),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_540),
.Y(n_599)
);

AO21x2_ASAP7_75t_L g600 ( 
.A1(n_564),
.A2(n_491),
.B(n_490),
.Y(n_600)
);

CKINVDCx12_ASAP7_75t_R g601 ( 
.A(n_563),
.Y(n_601)
);

CKINVDCx16_ASAP7_75t_R g602 ( 
.A(n_560),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_549),
.Y(n_603)
);

CKINVDCx16_ASAP7_75t_R g604 ( 
.A(n_560),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_553),
.B(n_493),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_548),
.A2(n_493),
.B1(n_535),
.B2(n_499),
.Y(n_606)
);

NAND2xp33_ASAP7_75t_SL g607 ( 
.A(n_554),
.B(n_521),
.Y(n_607)
);

NOR2x1_ASAP7_75t_L g608 ( 
.A(n_560),
.B(n_506),
.Y(n_608)
);

OR2x6_ASAP7_75t_L g609 ( 
.A(n_563),
.B(n_502),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_556),
.Y(n_610)
);

OR2x2_ASAP7_75t_L g611 ( 
.A(n_556),
.B(n_497),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_551),
.B(n_521),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_562),
.B(n_521),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_555),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_565),
.Y(n_615)
);

NAND2xp33_ASAP7_75t_R g616 ( 
.A(n_552),
.B(n_561),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_565),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_576),
.Y(n_618)
);

NAND3xp33_ASAP7_75t_L g619 ( 
.A(n_546),
.B(n_503),
.C(n_535),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_543),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_562),
.B(n_503),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_580),
.Y(n_622)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_566),
.B(n_497),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_580),
.Y(n_624)
);

CKINVDCx16_ASAP7_75t_R g625 ( 
.A(n_563),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_566),
.Y(n_626)
);

NAND3xp33_ASAP7_75t_SL g627 ( 
.A(n_557),
.B(n_499),
.C(n_494),
.Y(n_627)
);

BUFx6f_ASAP7_75t_SL g628 ( 
.A(n_568),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_R g629 ( 
.A(n_581),
.B(n_543),
.Y(n_629)
);

OR2x2_ASAP7_75t_L g630 ( 
.A(n_605),
.B(n_558),
.Y(n_630)
);

INVx1_ASAP7_75t_SL g631 ( 
.A(n_618),
.Y(n_631)
);

HB1xp67_ASAP7_75t_L g632 ( 
.A(n_622),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_624),
.Y(n_633)
);

OAI221xp5_ASAP7_75t_L g634 ( 
.A1(n_587),
.A2(n_579),
.B1(n_553),
.B2(n_569),
.C(n_544),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_586),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_588),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_589),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_590),
.Y(n_638)
);

AND2x4_ASAP7_75t_L g639 ( 
.A(n_584),
.B(n_578),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_602),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_595),
.B(n_581),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_584),
.B(n_578),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_598),
.B(n_552),
.Y(n_643)
);

INVx4_ASAP7_75t_R g644 ( 
.A(n_599),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_591),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_604),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_612),
.B(n_568),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_594),
.B(n_558),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_629),
.Y(n_649)
);

NOR2x1_ASAP7_75t_L g650 ( 
.A(n_585),
.B(n_543),
.Y(n_650)
);

BUFx2_ASAP7_75t_L g651 ( 
.A(n_584),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_610),
.B(n_577),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_593),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_603),
.Y(n_654)
);

HB1xp67_ASAP7_75t_L g655 ( 
.A(n_626),
.Y(n_655)
);

NAND3xp33_ASAP7_75t_L g656 ( 
.A(n_583),
.B(n_619),
.C(n_607),
.Y(n_656)
);

BUFx2_ASAP7_75t_L g657 ( 
.A(n_623),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_614),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_611),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_613),
.B(n_615),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_617),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_605),
.B(n_559),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_583),
.B(n_559),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_621),
.B(n_577),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_625),
.B(n_575),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_628),
.Y(n_666)
);

AOI221xp5_ASAP7_75t_L g667 ( 
.A1(n_592),
.A2(n_573),
.B1(n_567),
.B2(n_575),
.C(n_581),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_662),
.B(n_606),
.Y(n_668)
);

AND2x4_ASAP7_75t_SL g669 ( 
.A(n_639),
.B(n_609),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_662),
.B(n_606),
.Y(n_670)
);

NAND2xp67_ASAP7_75t_L g671 ( 
.A(n_665),
.B(n_573),
.Y(n_671)
);

INVx4_ASAP7_75t_L g672 ( 
.A(n_640),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_636),
.Y(n_673)
);

INVx1_ASAP7_75t_SL g674 ( 
.A(n_631),
.Y(n_674)
);

INVxp67_ASAP7_75t_L g675 ( 
.A(n_647),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_663),
.B(n_600),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_663),
.B(n_600),
.Y(n_677)
);

NOR2xp67_ASAP7_75t_L g678 ( 
.A(n_640),
.B(n_619),
.Y(n_678)
);

INVxp67_ASAP7_75t_L g679 ( 
.A(n_660),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_659),
.B(n_582),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_636),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_659),
.B(n_582),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_637),
.B(n_620),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_658),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_648),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_648),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_655),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_635),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_638),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_651),
.B(n_609),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_645),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_654),
.Y(n_692)
);

BUFx2_ASAP7_75t_L g693 ( 
.A(n_651),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_673),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_676),
.B(n_657),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_675),
.B(n_679),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_676),
.B(n_657),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_691),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_691),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_673),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_688),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_689),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_677),
.B(n_668),
.Y(n_703)
);

AOI221xp5_ASAP7_75t_L g704 ( 
.A1(n_684),
.A2(n_656),
.B1(n_634),
.B2(n_643),
.C(n_666),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_678),
.A2(n_674),
.B1(n_646),
.B2(n_627),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_692),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_693),
.B(n_646),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_693),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_687),
.B(n_661),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_677),
.B(n_630),
.Y(n_710)
);

OR2x2_ASAP7_75t_L g711 ( 
.A(n_668),
.B(n_670),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_694),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_696),
.B(n_711),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_694),
.Y(n_714)
);

OA222x2_ASAP7_75t_L g715 ( 
.A1(n_698),
.A2(n_630),
.B1(n_582),
.B2(n_685),
.C1(n_686),
.C2(n_609),
.Y(n_715)
);

OR2x6_ASAP7_75t_L g716 ( 
.A(n_707),
.B(n_672),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_704),
.A2(n_690),
.B1(n_601),
.B2(n_616),
.Y(n_717)
);

AO221x1_ASAP7_75t_L g718 ( 
.A1(n_699),
.A2(n_686),
.B1(n_685),
.B2(n_592),
.C(n_681),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_701),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_702),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_705),
.A2(n_690),
.B1(n_616),
.B2(n_627),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_706),
.Y(n_722)
);

AO22x1_ASAP7_75t_L g723 ( 
.A1(n_719),
.A2(n_708),
.B1(n_596),
.B2(n_672),
.Y(n_723)
);

OAI22xp33_ASAP7_75t_L g724 ( 
.A1(n_721),
.A2(n_672),
.B1(n_708),
.B2(n_690),
.Y(n_724)
);

AOI21xp33_ASAP7_75t_L g725 ( 
.A1(n_717),
.A2(n_705),
.B(n_709),
.Y(n_725)
);

OAI22xp33_ASAP7_75t_L g726 ( 
.A1(n_716),
.A2(n_649),
.B1(n_703),
.B2(n_670),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_720),
.Y(n_727)
);

NAND4xp75_ASAP7_75t_L g728 ( 
.A(n_725),
.B(n_649),
.C(n_715),
.D(n_650),
.Y(n_728)
);

INVx1_ASAP7_75t_SL g729 ( 
.A(n_723),
.Y(n_729)
);

NOR2xp67_ASAP7_75t_L g730 ( 
.A(n_727),
.B(n_722),
.Y(n_730)
);

AOI21xp33_ASAP7_75t_L g731 ( 
.A1(n_724),
.A2(n_713),
.B(n_641),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_729),
.B(n_731),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_730),
.A2(n_726),
.B(n_718),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_728),
.B(n_703),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_730),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_732),
.B(n_710),
.Y(n_736)
);

AOI221xp5_ASAP7_75t_L g737 ( 
.A1(n_734),
.A2(n_714),
.B1(n_712),
.B2(n_695),
.C(n_697),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_L g738 ( 
.A1(n_737),
.A2(n_733),
.B1(n_735),
.B2(n_669),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_736),
.Y(n_739)
);

NOR2x1_ASAP7_75t_L g740 ( 
.A(n_736),
.B(n_653),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_739),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_740),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_738),
.B(n_653),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_740),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_740),
.B(n_716),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_740),
.B(n_710),
.Y(n_746)
);

AND2x2_ASAP7_75t_SL g747 ( 
.A(n_744),
.B(n_597),
.Y(n_747)
);

OAI21xp5_ASAP7_75t_SL g748 ( 
.A1(n_742),
.A2(n_669),
.B(n_665),
.Y(n_748)
);

AOI221xp5_ASAP7_75t_L g749 ( 
.A1(n_741),
.A2(n_745),
.B1(n_743),
.B2(n_746),
.C(n_667),
.Y(n_749)
);

INVx1_ASAP7_75t_SL g750 ( 
.A(n_745),
.Y(n_750)
);

NOR2xp67_ASAP7_75t_L g751 ( 
.A(n_741),
.B(n_585),
.Y(n_751)
);

AOI221xp5_ASAP7_75t_L g752 ( 
.A1(n_743),
.A2(n_628),
.B1(n_683),
.B2(n_664),
.C(n_700),
.Y(n_752)
);

OR2x2_ASAP7_75t_L g753 ( 
.A(n_744),
.B(n_697),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_753),
.Y(n_754)
);

BUFx2_ASAP7_75t_L g755 ( 
.A(n_750),
.Y(n_755)
);

AND2x4_ASAP7_75t_L g756 ( 
.A(n_751),
.B(n_695),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_747),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_748),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_749),
.B(n_700),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_755),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_758),
.A2(n_752),
.B1(n_608),
.B2(n_639),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_757),
.B(n_671),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_756),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_754),
.Y(n_764)
);

NAND2xp33_ASAP7_75t_L g765 ( 
.A(n_756),
.B(n_644),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_759),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_760),
.Y(n_767)
);

AOI31xp33_ASAP7_75t_L g768 ( 
.A1(n_764),
.A2(n_550),
.A3(n_682),
.B(n_680),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_763),
.Y(n_769)
);

AOI31xp33_ASAP7_75t_L g770 ( 
.A1(n_766),
.A2(n_550),
.A3(n_682),
.B(n_680),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_SL g771 ( 
.A(n_762),
.B(n_581),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_769),
.Y(n_772)
);

CKINVDCx20_ASAP7_75t_R g773 ( 
.A(n_767),
.Y(n_773)
);

OAI221xp5_ASAP7_75t_L g774 ( 
.A1(n_771),
.A2(n_765),
.B1(n_761),
.B2(n_652),
.C(n_633),
.Y(n_774)
);

OAI31xp67_ASAP7_75t_SL g775 ( 
.A1(n_773),
.A2(n_770),
.A3(n_768),
.B(n_543),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_772),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_774),
.A2(n_639),
.B1(n_642),
.B2(n_632),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_776),
.B(n_547),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_SL g779 ( 
.A1(n_778),
.A2(n_775),
.B1(n_777),
.B2(n_570),
.Y(n_779)
);

AOI221x1_ASAP7_75t_L g780 ( 
.A1(n_779),
.A2(n_547),
.B1(n_570),
.B2(n_620),
.C(n_642),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_SL g781 ( 
.A1(n_780),
.A2(n_547),
.B1(n_570),
.B2(n_642),
.Y(n_781)
);


endmodule