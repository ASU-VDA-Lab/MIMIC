module fake_netlist_5_630_n_802 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_802);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_802;

wire n_676;
wire n_294;
wire n_431;
wire n_380;
wire n_419;
wire n_318;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_316;
wire n_785;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_523;
wire n_268;
wire n_315;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_525;
wire n_493;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_443;
wire n_372;
wire n_244;
wire n_677;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_433;
wire n_314;
wire n_368;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_779;
wire n_576;
wire n_537;
wire n_587;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_524;
wire n_399;
wire n_579;
wire n_204;
wire n_394;
wire n_250;
wire n_341;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_782;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_234;
wire n_343;
wire n_379;
wire n_428;
wire n_308;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_432;
wire n_395;
wire n_553;
wire n_727;
wire n_311;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_772;
wire n_691;
wire n_717;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_796;
wire n_573;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_477;
wire n_338;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_466;
wire n_239;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_332;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_557;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_707;
wire n_710;
wire n_795;
wire n_695;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_403;
wire n_453;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_794;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_246;
wire n_596;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_565;
wire n_426;
wire n_520;
wire n_566;
wire n_409;
wire n_797;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_334;
wire n_599;
wire n_766;
wire n_541;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_538;
wire n_666;
wire n_262;
wire n_238;
wire n_639;
wire n_799;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_759;
wire n_222;
wire n_438;
wire n_713;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_401;
wire n_348;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;
wire n_784;

INVx1_ASAP7_75t_L g198 ( 
.A(n_10),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_144),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_171),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_154),
.Y(n_201)
);

NOR2xp67_ASAP7_75t_L g202 ( 
.A(n_37),
.B(n_167),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_118),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_91),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_12),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_110),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_113),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_18),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_51),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_76),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_33),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_66),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_106),
.Y(n_214)
);

BUFx2_ASAP7_75t_SL g215 ( 
.A(n_45),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_90),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_163),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_31),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_74),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_75),
.Y(n_220)
);

BUFx2_ASAP7_75t_SL g221 ( 
.A(n_182),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_103),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_17),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_19),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_69),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_148),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_97),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_143),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_78),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_86),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_111),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_82),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_135),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_164),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_99),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_116),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_58),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_151),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_114),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_132),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_85),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_139),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_60),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_190),
.Y(n_244)
);

INVxp67_ASAP7_75t_SL g245 ( 
.A(n_153),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_23),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_168),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_146),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_149),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_61),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_79),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g252 ( 
.A(n_63),
.B(n_147),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_22),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_173),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_165),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_40),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_83),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_107),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_115),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_184),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_194),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_175),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_126),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_27),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_160),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_140),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_28),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_192),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_18),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g270 ( 
.A(n_121),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_46),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_89),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_54),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_88),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_124),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_120),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_150),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_112),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_197),
.Y(n_279)
);

BUFx5_ASAP7_75t_L g280 ( 
.A(n_133),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_3),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_129),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_169),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_33),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_67),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_68),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_131),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_170),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_142),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_84),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_119),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_122),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_92),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_174),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_20),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_19),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_29),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_43),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_179),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_96),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_53),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_128),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_62),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_109),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_4),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_2),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_65),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_172),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_55),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_152),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_195),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_108),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_141),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_145),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_134),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_104),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_59),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_127),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_72),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_166),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_177),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_5),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_117),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_100),
.Y(n_324)
);

BUFx5_ASAP7_75t_L g325 ( 
.A(n_185),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_4),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_38),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_191),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_7),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_80),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_2),
.Y(n_331)
);

INVx5_ASAP7_75t_L g332 ( 
.A(n_206),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_205),
.B(n_327),
.Y(n_333)
);

CKINVDCx6p67_ASAP7_75t_R g334 ( 
.A(n_212),
.Y(n_334)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_329),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_206),
.Y(n_336)
);

AND2x4_ASAP7_75t_L g337 ( 
.A(n_204),
.B(n_0),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_222),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_198),
.Y(n_339)
);

INVxp33_ASAP7_75t_SL g340 ( 
.A(n_331),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_209),
.Y(n_341)
);

AND2x6_ASAP7_75t_L g342 ( 
.A(n_222),
.B(n_41),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_224),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_280),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_218),
.Y(n_345)
);

OA21x2_ASAP7_75t_L g346 ( 
.A1(n_200),
.A2(n_1),
.B(n_6),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_222),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_280),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_233),
.Y(n_349)
);

AND2x4_ASAP7_75t_L g350 ( 
.A(n_213),
.B(n_8),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_223),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_233),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_326),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_270),
.B(n_9),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_233),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_264),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_280),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_280),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_236),
.B(n_13),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_267),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_325),
.Y(n_361)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_269),
.Y(n_362)
);

INVx4_ASAP7_75t_L g363 ( 
.A(n_254),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_281),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_254),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_246),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_366)
);

AND2x6_ASAP7_75t_L g367 ( 
.A(n_254),
.B(n_42),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_325),
.Y(n_368)
);

OAI21x1_ASAP7_75t_L g369 ( 
.A1(n_207),
.A2(n_47),
.B(n_44),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_325),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_216),
.B(n_16),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_295),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_325),
.Y(n_373)
);

INVx5_ASAP7_75t_L g374 ( 
.A(n_255),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_201),
.Y(n_375)
);

INVx4_ASAP7_75t_L g376 ( 
.A(n_255),
.Y(n_376)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_226),
.B(n_20),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_203),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_272),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_202),
.B(n_21),
.Y(n_380)
);

INVx4_ASAP7_75t_L g381 ( 
.A(n_272),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_211),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_214),
.Y(n_383)
);

OAI21x1_ASAP7_75t_L g384 ( 
.A1(n_208),
.A2(n_49),
.B(n_48),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_253),
.B(n_24),
.Y(n_385)
);

AND2x4_ASAP7_75t_L g386 ( 
.A(n_227),
.B(n_25),
.Y(n_386)
);

INVx5_ASAP7_75t_L g387 ( 
.A(n_272),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_231),
.B(n_26),
.Y(n_388)
);

OA21x2_ASAP7_75t_L g389 ( 
.A1(n_219),
.A2(n_26),
.B(n_27),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_256),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_199),
.Y(n_391)
);

INVx5_ASAP7_75t_L g392 ( 
.A(n_289),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_289),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_289),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_284),
.A2(n_30),
.B1(n_32),
.B2(n_34),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_296),
.A2(n_297),
.B1(n_306),
.B2(n_305),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_248),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_285),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_286),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_241),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_325),
.Y(n_401)
);

BUFx8_ASAP7_75t_L g402 ( 
.A(n_325),
.Y(n_402)
);

INVx6_ASAP7_75t_L g403 ( 
.A(n_252),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_303),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_321),
.B(n_35),
.Y(n_405)
);

OA21x2_ASAP7_75t_L g406 ( 
.A1(n_230),
.A2(n_36),
.B(n_38),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_304),
.B(n_319),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_234),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_322),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_237),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_304),
.B(n_36),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_238),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_210),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_242),
.B(n_39),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_243),
.B(n_39),
.Y(n_415)
);

INVx5_ASAP7_75t_L g416 ( 
.A(n_215),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_244),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_247),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_249),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_257),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_258),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_259),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_265),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_266),
.B(n_50),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_282),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_268),
.Y(n_426)
);

OA21x2_ASAP7_75t_L g427 ( 
.A1(n_274),
.A2(n_52),
.B(n_56),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_275),
.B(n_57),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_279),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_283),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_287),
.B(n_64),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_336),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_333),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_336),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g435 ( 
.A(n_391),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_390),
.B(n_263),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_407),
.B(n_245),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_400),
.Y(n_438)
);

OAI21x1_ASAP7_75t_L g439 ( 
.A1(n_369),
.A2(n_291),
.B(n_290),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_338),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_338),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_413),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_347),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_425),
.Y(n_444)
);

AO21x2_ASAP7_75t_L g445 ( 
.A1(n_380),
.A2(n_245),
.B(n_293),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_334),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_345),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_347),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_349),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_351),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_349),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_349),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_352),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_355),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_409),
.B(n_292),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_355),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_355),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_365),
.Y(n_458)
);

OR2x6_ASAP7_75t_L g459 ( 
.A(n_354),
.B(n_221),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_396),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_379),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_379),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_340),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_379),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_393),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_402),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_402),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_393),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_375),
.B(n_330),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_394),
.Y(n_470)
);

INVx4_ASAP7_75t_L g471 ( 
.A(n_342),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_394),
.Y(n_472)
);

NOR2xp67_ASAP7_75t_L g473 ( 
.A(n_416),
.B(n_332),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_416),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_335),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_403),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_412),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_417),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_418),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_335),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g481 ( 
.A(n_419),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_421),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_422),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_363),
.Y(n_484)
);

INVx4_ASAP7_75t_L g485 ( 
.A(n_342),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_378),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_481),
.Y(n_487)
);

INVx2_ASAP7_75t_SL g488 ( 
.A(n_476),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_437),
.B(n_359),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_486),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_451),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_484),
.B(n_424),
.Y(n_492)
);

NOR2x1p5_ASAP7_75t_L g493 ( 
.A(n_466),
.B(n_411),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_454),
.Y(n_494)
);

BUFx5_ASAP7_75t_L g495 ( 
.A(n_477),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_470),
.Y(n_496)
);

INVxp67_ASAP7_75t_SL g497 ( 
.A(n_475),
.Y(n_497)
);

BUFx5_ASAP7_75t_L g498 ( 
.A(n_478),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_445),
.B(n_428),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_445),
.B(n_428),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_432),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_434),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_443),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_458),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_436),
.B(n_431),
.Y(n_505)
);

NOR3xp33_ASAP7_75t_L g506 ( 
.A(n_460),
.B(n_395),
.C(n_366),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_458),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_455),
.B(n_385),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_L g509 ( 
.A1(n_459),
.A2(n_386),
.B1(n_388),
.B2(n_377),
.Y(n_509)
);

INVx8_ASAP7_75t_L g510 ( 
.A(n_438),
.Y(n_510)
);

BUFx5_ASAP7_75t_L g511 ( 
.A(n_479),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_433),
.B(n_371),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_464),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_469),
.B(n_374),
.Y(n_514)
);

AND2x6_ASAP7_75t_L g515 ( 
.A(n_435),
.B(n_337),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_440),
.Y(n_516)
);

BUFx5_ASAP7_75t_L g517 ( 
.A(n_482),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_441),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_469),
.B(n_374),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_480),
.Y(n_520)
);

NAND3xp33_ASAP7_75t_L g521 ( 
.A(n_447),
.B(n_405),
.C(n_350),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_448),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_439),
.A2(n_384),
.B(n_427),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_449),
.B(n_387),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_452),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_453),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_450),
.B(n_350),
.Y(n_527)
);

AO221x1_ASAP7_75t_L g528 ( 
.A1(n_459),
.A2(n_299),
.B1(n_307),
.B2(n_301),
.C(n_298),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_456),
.B(n_392),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_457),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_442),
.B(n_414),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_461),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_483),
.B(n_415),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_462),
.Y(n_534)
);

NAND2x1_ASAP7_75t_L g535 ( 
.A(n_471),
.B(n_342),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_465),
.B(n_363),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_468),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_489),
.A2(n_463),
.B1(n_485),
.B2(n_471),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_490),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_505),
.B(n_485),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_520),
.B(n_339),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_494),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_492),
.A2(n_500),
.B(n_499),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_496),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_488),
.B(n_467),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_510),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_491),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_487),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_502),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_506),
.A2(n_346),
.B1(n_406),
.B2(n_389),
.Y(n_550)
);

O2A1O1Ixp33_ASAP7_75t_L g551 ( 
.A1(n_508),
.A2(n_426),
.B(n_423),
.C(n_383),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_504),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_SL g553 ( 
.A1(n_521),
.A2(n_353),
.B1(n_444),
.B2(n_446),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_527),
.B(n_509),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_512),
.B(n_397),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_523),
.A2(n_535),
.B(n_519),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_531),
.B(n_474),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_526),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_L g559 ( 
.A1(n_528),
.A2(n_346),
.B1(n_406),
.B2(n_389),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_533),
.B(n_343),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_522),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_530),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_515),
.B(n_497),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_515),
.B(n_398),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_516),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_515),
.B(n_398),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_518),
.Y(n_567)
);

INVx5_ASAP7_75t_L g568 ( 
.A(n_526),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_507),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_514),
.B(n_398),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_525),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_534),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_495),
.B(n_399),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_495),
.B(n_498),
.Y(n_574)
);

INVx5_ASAP7_75t_L g575 ( 
.A(n_526),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_495),
.B(n_399),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_498),
.B(n_404),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_513),
.Y(n_578)
);

BUFx12f_ASAP7_75t_L g579 ( 
.A(n_493),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_498),
.B(n_404),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_532),
.B(n_360),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_537),
.Y(n_582)
);

INVxp67_ASAP7_75t_SL g583 ( 
.A(n_536),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_501),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_498),
.B(n_404),
.Y(n_585)
);

BUFx10_ASAP7_75t_L g586 ( 
.A(n_503),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_511),
.B(n_472),
.Y(n_587)
);

INVx5_ASAP7_75t_L g588 ( 
.A(n_511),
.Y(n_588)
);

INVx5_ASAP7_75t_L g589 ( 
.A(n_511),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_517),
.B(n_217),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_517),
.B(n_309),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_524),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_529),
.B(n_220),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_546),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_588),
.A2(n_589),
.B(n_543),
.Y(n_595)
);

O2A1O1Ixp33_ASAP7_75t_L g596 ( 
.A1(n_554),
.A2(n_408),
.B(n_410),
.C(n_382),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_588),
.A2(n_427),
.B(n_473),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_581),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_560),
.B(n_364),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_539),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_588),
.A2(n_315),
.B(n_314),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_581),
.Y(n_602)
);

AOI21xp5_ASAP7_75t_L g603 ( 
.A1(n_589),
.A2(n_323),
.B(n_316),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_538),
.A2(n_228),
.B1(n_229),
.B2(n_225),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_548),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_555),
.B(n_232),
.Y(n_606)
);

INVx8_ASAP7_75t_L g607 ( 
.A(n_579),
.Y(n_607)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_574),
.A2(n_348),
.B(n_344),
.Y(n_608)
);

A2O1A1Ixp33_ASAP7_75t_L g609 ( 
.A1(n_540),
.A2(n_430),
.B(n_358),
.C(n_361),
.Y(n_609)
);

AOI22x1_ASAP7_75t_L g610 ( 
.A1(n_556),
.A2(n_239),
.B1(n_240),
.B2(n_235),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_545),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_560),
.B(n_372),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_563),
.B(n_250),
.Y(n_613)
);

OAI21x1_ASAP7_75t_L g614 ( 
.A1(n_587),
.A2(n_368),
.B(n_357),
.Y(n_614)
);

A2O1A1Ixp33_ASAP7_75t_SL g615 ( 
.A1(n_550),
.A2(n_430),
.B(n_370),
.C(n_401),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_542),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_583),
.B(n_251),
.Y(n_617)
);

O2A1O1Ixp33_ASAP7_75t_L g618 ( 
.A1(n_551),
.A2(n_373),
.B(n_341),
.C(n_356),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_561),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_562),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_578),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_558),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_564),
.A2(n_261),
.B(n_260),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_572),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_565),
.Y(n_625)
);

A2O1A1Ixp33_ASAP7_75t_SL g626 ( 
.A1(n_559),
.A2(n_362),
.B(n_367),
.C(n_262),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_565),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_567),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_567),
.Y(n_629)
);

NOR2xp67_ASAP7_75t_SL g630 ( 
.A(n_568),
.B(n_271),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_566),
.A2(n_276),
.B(n_273),
.Y(n_631)
);

A2O1A1Ixp33_ASAP7_75t_SL g632 ( 
.A1(n_571),
.A2(n_308),
.B(n_277),
.C(n_278),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_592),
.B(n_544),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_541),
.B(n_420),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_578),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_547),
.Y(n_636)
);

BUFx2_ASAP7_75t_L g637 ( 
.A(n_541),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_582),
.Y(n_638)
);

A2O1A1Ixp33_ASAP7_75t_SL g639 ( 
.A1(n_571),
.A2(n_311),
.B(n_288),
.C(n_328),
.Y(n_639)
);

A2O1A1Ixp33_ASAP7_75t_L g640 ( 
.A1(n_584),
.A2(n_313),
.B(n_294),
.C(n_324),
.Y(n_640)
);

OAI21x1_ASAP7_75t_L g641 ( 
.A1(n_614),
.A2(n_576),
.B(n_573),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_625),
.Y(n_642)
);

OAI21x1_ASAP7_75t_L g643 ( 
.A1(n_595),
.A2(n_580),
.B(n_577),
.Y(n_643)
);

OA21x2_ASAP7_75t_L g644 ( 
.A1(n_609),
.A2(n_591),
.B(n_585),
.Y(n_644)
);

AOI21x1_ASAP7_75t_L g645 ( 
.A1(n_613),
.A2(n_597),
.B(n_590),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_594),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_622),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_629),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_615),
.A2(n_575),
.B(n_570),
.Y(n_649)
);

INVx1_ASAP7_75t_SL g650 ( 
.A(n_605),
.Y(n_650)
);

AOI22x1_ASAP7_75t_L g651 ( 
.A1(n_608),
.A2(n_549),
.B1(n_552),
.B2(n_569),
.Y(n_651)
);

INVx6_ASAP7_75t_L g652 ( 
.A(n_607),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_622),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_620),
.Y(n_654)
);

AO21x2_ASAP7_75t_L g655 ( 
.A1(n_626),
.A2(n_593),
.B(n_557),
.Y(n_655)
);

AO21x2_ASAP7_75t_L g656 ( 
.A1(n_606),
.A2(n_586),
.B(n_429),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_611),
.B(n_553),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_627),
.Y(n_658)
);

AOI22x1_ASAP7_75t_L g659 ( 
.A1(n_628),
.A2(n_317),
.B1(n_300),
.B2(n_302),
.Y(n_659)
);

INVx8_ASAP7_75t_L g660 ( 
.A(n_599),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_635),
.Y(n_661)
);

BUFx4f_ASAP7_75t_L g662 ( 
.A(n_635),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_621),
.Y(n_663)
);

AOI22x1_ASAP7_75t_L g664 ( 
.A1(n_600),
.A2(n_320),
.B1(n_310),
.B2(n_312),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_619),
.Y(n_665)
);

INVx6_ASAP7_75t_L g666 ( 
.A(n_599),
.Y(n_666)
);

OAI21x1_ASAP7_75t_L g667 ( 
.A1(n_610),
.A2(n_70),
.B(n_71),
.Y(n_667)
);

INVx6_ASAP7_75t_L g668 ( 
.A(n_612),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g669 ( 
.A(n_637),
.B(n_420),
.Y(n_669)
);

AOI22x1_ASAP7_75t_L g670 ( 
.A1(n_624),
.A2(n_636),
.B1(n_638),
.B2(n_616),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_598),
.Y(n_671)
);

AO21x2_ASAP7_75t_L g672 ( 
.A1(n_617),
.A2(n_73),
.B(n_77),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_602),
.Y(n_673)
);

AOI22x1_ASAP7_75t_L g674 ( 
.A1(n_634),
.A2(n_601),
.B1(n_603),
.B2(n_623),
.Y(n_674)
);

OR2x6_ASAP7_75t_L g675 ( 
.A(n_633),
.B(n_429),
.Y(n_675)
);

OAI21x1_ASAP7_75t_L g676 ( 
.A1(n_596),
.A2(n_81),
.B(n_87),
.Y(n_676)
);

INVx5_ASAP7_75t_L g677 ( 
.A(n_630),
.Y(n_677)
);

OAI21x1_ASAP7_75t_L g678 ( 
.A1(n_631),
.A2(n_93),
.B(n_94),
.Y(n_678)
);

OAI21x1_ASAP7_75t_L g679 ( 
.A1(n_618),
.A2(n_95),
.B(n_98),
.Y(n_679)
);

OA21x2_ASAP7_75t_L g680 ( 
.A1(n_641),
.A2(n_640),
.B(n_604),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_665),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_642),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_658),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_658),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_673),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_657),
.A2(n_318),
.B1(n_381),
.B2(n_376),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_670),
.Y(n_687)
);

OR2x6_ASAP7_75t_L g688 ( 
.A(n_660),
.B(n_381),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_670),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_647),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_648),
.Y(n_691)
);

AOI21x1_ASAP7_75t_L g692 ( 
.A1(n_645),
.A2(n_639),
.B(n_632),
.Y(n_692)
);

INVx5_ASAP7_75t_L g693 ( 
.A(n_661),
.Y(n_693)
);

OAI21x1_ASAP7_75t_L g694 ( 
.A1(n_643),
.A2(n_101),
.B(n_102),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_654),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_663),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_651),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_671),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_646),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_651),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_669),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_644),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_650),
.B(n_105),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_653),
.Y(n_704)
);

OAI22xp33_ASAP7_75t_L g705 ( 
.A1(n_675),
.A2(n_668),
.B1(n_666),
.B2(n_677),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_666),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_644),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_652),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_662),
.Y(n_709)
);

AOI21x1_ASAP7_75t_L g710 ( 
.A1(n_649),
.A2(n_123),
.B(n_125),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_709),
.B(n_677),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_701),
.B(n_656),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_681),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_682),
.B(n_655),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_SL g715 ( 
.A(n_699),
.B(n_655),
.Y(n_715)
);

O2A1O1Ixp33_ASAP7_75t_SL g716 ( 
.A1(n_705),
.A2(n_659),
.B(n_664),
.C(n_676),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_703),
.B(n_672),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_708),
.B(n_678),
.Y(n_718)
);

XNOR2xp5_ASAP7_75t_L g719 ( 
.A(n_706),
.B(n_674),
.Y(n_719)
);

NAND3xp33_ASAP7_75t_L g720 ( 
.A(n_686),
.B(n_667),
.C(n_679),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_682),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_695),
.B(n_130),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_683),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_693),
.Y(n_724)
);

AO31x2_ASAP7_75t_L g725 ( 
.A1(n_697),
.A2(n_136),
.A3(n_137),
.B(n_138),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_684),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_691),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_685),
.Y(n_728)
);

AO31x2_ASAP7_75t_L g729 ( 
.A1(n_697),
.A2(n_155),
.A3(n_156),
.B(n_157),
.Y(n_729)
);

OR2x2_ASAP7_75t_L g730 ( 
.A(n_704),
.B(n_158),
.Y(n_730)
);

AO31x2_ASAP7_75t_L g731 ( 
.A1(n_700),
.A2(n_159),
.A3(n_161),
.B(n_162),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_688),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_721),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_713),
.B(n_707),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_723),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_726),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_714),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_728),
.B(n_702),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_727),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_712),
.B(n_698),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_717),
.B(n_689),
.Y(n_741)
);

BUFx2_ASAP7_75t_SL g742 ( 
.A(n_732),
.Y(n_742)
);

OA21x2_ASAP7_75t_L g743 ( 
.A1(n_720),
.A2(n_700),
.B(n_689),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_725),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_719),
.B(n_687),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_729),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_731),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_731),
.Y(n_748)
);

BUFx2_ASAP7_75t_L g749 ( 
.A(n_715),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_718),
.Y(n_750)
);

AO21x2_ASAP7_75t_L g751 ( 
.A1(n_716),
.A2(n_710),
.B(n_692),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_724),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_722),
.B(n_696),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_730),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_711),
.B(n_680),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_741),
.B(n_680),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_735),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_737),
.B(n_694),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_736),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_745),
.B(n_690),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_754),
.B(n_740),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_734),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_734),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_738),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_742),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_750),
.Y(n_766)
);

OR2x2_ASAP7_75t_L g767 ( 
.A(n_761),
.B(n_755),
.Y(n_767)
);

INVx1_ASAP7_75t_SL g768 ( 
.A(n_765),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_756),
.B(n_749),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_759),
.Y(n_770)
);

OR2x2_ASAP7_75t_L g771 ( 
.A(n_762),
.B(n_763),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_762),
.B(n_744),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_757),
.Y(n_773)
);

OR2x2_ASAP7_75t_L g774 ( 
.A(n_767),
.B(n_766),
.Y(n_774)
);

OR2x2_ASAP7_75t_L g775 ( 
.A(n_769),
.B(n_764),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_768),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_773),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_777),
.Y(n_778)
);

XOR2x2_ASAP7_75t_L g779 ( 
.A(n_776),
.B(n_760),
.Y(n_779)
);

OR2x2_ASAP7_75t_L g780 ( 
.A(n_774),
.B(n_771),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_778),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_780),
.B(n_775),
.Y(n_782)
);

INVx1_ASAP7_75t_SL g783 ( 
.A(n_779),
.Y(n_783)
);

INVx1_ASAP7_75t_SL g784 ( 
.A(n_783),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_782),
.B(n_770),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_784),
.B(n_781),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_785),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_787),
.B(n_772),
.Y(n_788)
);

AOI211xp5_ASAP7_75t_L g789 ( 
.A1(n_786),
.A2(n_753),
.B(n_752),
.C(n_758),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_788),
.Y(n_790)
);

NOR2x1_ASAP7_75t_SL g791 ( 
.A(n_789),
.B(n_751),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_790),
.Y(n_792)
);

NAND2x1p5_ASAP7_75t_SL g793 ( 
.A(n_791),
.B(n_739),
.Y(n_793)
);

OAI211xp5_ASAP7_75t_SL g794 ( 
.A1(n_792),
.A2(n_739),
.B(n_733),
.C(n_747),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_794),
.A2(n_793),
.B1(n_746),
.B2(n_748),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_795),
.B(n_743),
.Y(n_796)
);

CKINVDCx20_ASAP7_75t_R g797 ( 
.A(n_796),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_SL g798 ( 
.A1(n_797),
.A2(n_743),
.B1(n_176),
.B2(n_178),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_798),
.B(n_180),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_R g800 ( 
.A1(n_799),
.A2(n_181),
.B1(n_183),
.B2(n_186),
.Y(n_800)
);

OR2x6_ASAP7_75t_L g801 ( 
.A(n_800),
.B(n_188),
.Y(n_801)
);

AOI31xp33_ASAP7_75t_L g802 ( 
.A1(n_801),
.A2(n_196),
.A3(n_189),
.B(n_193),
.Y(n_802)
);


endmodule