module real_jpeg_33899_n_13 (n_329, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_329;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx2_ASAP7_75t_L g86 ( 
.A(n_0),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_0),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_0),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_0),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_1),
.A2(n_170),
.B1(n_172),
.B2(n_173),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_1),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_1),
.A2(n_172),
.B1(n_216),
.B2(n_221),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_1),
.A2(n_172),
.B1(n_262),
.B2(n_264),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_2),
.Y(n_122)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_2),
.Y(n_161)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_3),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_3),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_4),
.A2(n_75),
.B1(n_78),
.B2(n_81),
.Y(n_74)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_4),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_5),
.A2(n_144),
.B1(n_147),
.B2(n_148),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_5),
.Y(n_147)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_6),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_7),
.B(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_7),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_7),
.B(n_127),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_7),
.A2(n_110),
.B1(n_206),
.B2(n_209),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_7),
.B(n_154),
.Y(n_236)
);

OAI21xp33_ASAP7_75t_L g270 ( 
.A1(n_7),
.A2(n_142),
.B(n_250),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_8),
.Y(n_131)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_10),
.A2(n_48),
.B1(n_52),
.B2(n_57),
.Y(n_47)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_10),
.A2(n_57),
.B1(n_239),
.B2(n_245),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_11),
.Y(n_108)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_11),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_11),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_11),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_12),
.A2(n_60),
.B1(n_65),
.B2(n_66),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_12),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_12),
.A2(n_65),
.B1(n_94),
.B2(n_97),
.Y(n_93)
);

OAI22x1_ASAP7_75t_SL g178 ( 
.A1(n_12),
.A2(n_65),
.B1(n_179),
.B2(n_184),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_228),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_227),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_202),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_17),
.B(n_202),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_123),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_71),
.B2(n_72),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI21xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_47),
.B(n_58),
.Y(n_20)
);

OAI22xp33_ASAP7_75t_L g214 ( 
.A1(n_21),
.A2(n_47),
.B1(n_215),
.B2(n_224),
.Y(n_214)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_21),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_38),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

OAI22x1_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_26),
.B1(n_30),
.B2(n_34),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_24),
.Y(n_146)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_25),
.Y(n_292)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_L g297 ( 
.A(n_32),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_41),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_46),
.Y(n_318)
);

INVx3_ASAP7_75t_SL g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_55),
.Y(n_302)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_58),
.B(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_70),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_59),
.B(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_64),
.Y(n_167)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_70),
.Y(n_224)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_99),
.Y(n_72)
);

XNOR2x1_ASAP7_75t_L g226 ( 
.A(n_73),
.B(n_99),
.Y(n_226)
);

OA21x2_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_82),
.B(n_87),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_74),
.A2(n_142),
.B1(n_143),
.B2(n_150),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_77),
.Y(n_278)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_80),
.Y(n_307)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_86),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_87),
.A2(n_261),
.B(n_265),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_93),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_88),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_88),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_91),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx8_ASAP7_75t_L g252 ( 
.A(n_92),
.Y(n_252)
);

NAND2xp33_ASAP7_75t_SL g250 ( 
.A(n_93),
.B(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_96),
.Y(n_249)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_104),
.B1(n_109),
.B2(n_114),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_107),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_108),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_108),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_110),
.B(n_224),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_110),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_110),
.B(n_300),
.Y(n_299)
);

OAI21xp33_ASAP7_75t_SL g315 ( 
.A1(n_110),
.A2(n_299),
.B(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_116),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_117),
.Y(n_187)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_122),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_122),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_152),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_140),
.B2(n_141),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_132),
.B1(n_135),
.B2(n_138),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_134),
.Y(n_176)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_137),
.Y(n_208)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_142),
.A2(n_238),
.B(n_250),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_151),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_168),
.B(n_177),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_154),
.B(n_178),
.Y(n_212)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

AND2x4_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_189),
.Y(n_188)
);

AOI22x1_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_159),
.B1(n_162),
.B2(n_165),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_158),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_188),
.Y(n_177)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_188),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_194),
.B1(n_197),
.B2(n_200),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_213),
.C(n_225),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_203),
.B(n_214),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B(n_212),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_SL g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_215),
.A2(n_224),
.B(n_233),
.Y(n_232)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_220),
.Y(n_312)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_225),
.A2(n_226),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OAI321xp33_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_256),
.A3(n_320),
.B1(n_326),
.B2(n_327),
.C(n_329),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_253),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_230),
.B(n_253),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_235),
.C(n_237),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_232),
.A2(n_235),
.B1(n_236),
.B2(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_232),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_234),
.B(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_237),
.Y(n_323)
);

INVxp33_ASAP7_75t_SL g282 ( 
.A(n_238),
.Y(n_282)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_241),
.Y(n_264)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_244),
.Y(n_263)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_280),
.B(n_319),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_269),
.B(n_279),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_259),
.B(n_260),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_261),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_277),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_285),
.Y(n_280)
);

NOR2xp67_ASAP7_75t_L g319 ( 
.A(n_281),
.B(n_285),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_313),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_286),
.B(n_313),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_298),
.B1(n_303),
.B2(n_308),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_293),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_309),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

BUFx4f_ASAP7_75t_SL g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NOR2xp67_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_322),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);


endmodule