module fake_jpeg_13125_n_353 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_353);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_353;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g105 ( 
.A(n_45),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_51),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_29),
.B(n_8),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_53),
.B(n_39),
.Y(n_81)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_18),
.B(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_0),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_21),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_64),
.Y(n_70)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

NAND2x1_ASAP7_75t_SL g64 ( 
.A(n_26),
.B(n_9),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_21),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_40),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_50),
.B1(n_51),
.B2(n_66),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_71),
.A2(n_80),
.B1(n_69),
.B2(n_31),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_18),
.B1(n_41),
.B2(n_36),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_73),
.A2(n_85),
.B1(n_103),
.B2(n_111),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_45),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_74),
.B(n_78),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_39),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_79),
.B(n_81),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_18),
.B1(n_41),
.B2(n_31),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_29),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_82),
.B(n_87),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_107),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_60),
.A2(n_41),
.B1(n_22),
.B2(n_35),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_19),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_44),
.B(n_19),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_59),
.A2(n_27),
.B1(n_21),
.B2(n_35),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_93),
.A2(n_61),
.B1(n_49),
.B2(n_34),
.Y(n_124)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_45),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_98),
.Y(n_143)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

INVx3_ASAP7_75t_SL g135 ( 
.A(n_100),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_48),
.B(n_24),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_101),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_24),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_102),
.B(n_109),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_47),
.A2(n_22),
.B1(n_35),
.B2(n_32),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_37),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_67),
.B(n_37),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_52),
.A2(n_22),
.B1(n_32),
.B2(n_28),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_84),
.A2(n_62),
.B1(n_32),
.B2(n_21),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_115),
.A2(n_118),
.B1(n_121),
.B2(n_128),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_70),
.A2(n_21),
.B1(n_27),
.B2(n_28),
.Y(n_118)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_122),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_34),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_123),
.B(n_138),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_SL g167 ( 
.A1(n_124),
.A2(n_105),
.B(n_95),
.C(n_108),
.Y(n_167)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_126),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

INVx3_ASAP7_75t_SL g158 ( 
.A(n_127),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_83),
.B1(n_106),
.B2(n_94),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_129),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_L g130 ( 
.A1(n_89),
.A2(n_49),
.B1(n_38),
.B2(n_40),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_130),
.A2(n_137),
.B1(n_99),
.B2(n_90),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_112),
.A2(n_30),
.B1(n_38),
.B2(n_40),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_131),
.A2(n_147),
.B1(n_149),
.B2(n_96),
.Y(n_166)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_72),
.Y(n_132)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_132),
.Y(n_173)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_134),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_30),
.B1(n_42),
.B2(n_38),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_76),
.B(n_0),
.Y(n_138)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_142),
.Y(n_185)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_76),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_144),
.B(n_145),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_94),
.B(n_104),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_100),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_152),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_77),
.A2(n_40),
.B1(n_42),
.B2(n_2),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_77),
.A2(n_42),
.B1(n_1),
.B2(n_2),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_113),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_150),
.A2(n_154),
.B1(n_110),
.B2(n_96),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_104),
.B(n_3),
.Y(n_151)
);

A2O1A1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_151),
.A2(n_105),
.B(n_4),
.C(n_7),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_86),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_92),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_141),
.A2(n_108),
.B1(n_95),
.B2(n_114),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_155),
.A2(n_159),
.B1(n_169),
.B2(n_182),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_123),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_161),
.B(n_164),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_86),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_162),
.B(n_165),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_136),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_75),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_166),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_167),
.B(n_175),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_154),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_141),
.A2(n_114),
.B1(n_75),
.B2(n_110),
.Y(n_169)
);

AO22x1_ASAP7_75t_L g177 ( 
.A1(n_130),
.A2(n_99),
.B1(n_90),
.B2(n_4),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_177),
.B(n_135),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_145),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_179),
.B(n_188),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_117),
.A2(n_6),
.B(n_7),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_180),
.A2(n_187),
.B(n_189),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_143),
.A2(n_99),
.B(n_90),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_181),
.A2(n_146),
.B(n_133),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_116),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_182)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_126),
.Y(n_184)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_184),
.Y(n_206)
);

AOI32xp33_ASAP7_75t_L g186 ( 
.A1(n_117),
.A2(n_9),
.A3(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_186)
);

OR2x2_ASAP7_75t_SL g204 ( 
.A(n_186),
.B(n_187),
.Y(n_204)
);

AOI32xp33_ASAP7_75t_L g187 ( 
.A1(n_116),
.A2(n_13),
.A3(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_148),
.Y(n_188)
);

AOI32xp33_ASAP7_75t_L g189 ( 
.A1(n_148),
.A2(n_14),
.A3(n_15),
.B1(n_17),
.B2(n_138),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_153),
.A2(n_17),
.B1(n_115),
.B2(n_151),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_190),
.A2(n_135),
.B1(n_158),
.B2(n_168),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_191),
.A2(n_202),
.B(n_212),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_193),
.Y(n_250)
);

AND2x2_ASAP7_75t_SL g194 ( 
.A(n_179),
.B(n_119),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_194),
.Y(n_237)
);

INVxp33_ASAP7_75t_L g195 ( 
.A(n_160),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_195),
.B(n_196),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_176),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_161),
.B(n_148),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_197),
.B(n_211),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_143),
.C(n_119),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_200),
.C(n_173),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_129),
.C(n_181),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_201),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_163),
.A2(n_144),
.B1(n_127),
.B2(n_125),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_204),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_185),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_207),
.B(n_213),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_163),
.A2(n_122),
.B1(n_127),
.B2(n_152),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_209),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_189),
.A2(n_122),
.B1(n_120),
.B2(n_132),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_182),
.B(n_140),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_180),
.B(n_134),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_185),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_218),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_156),
.Y(n_215)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_215),
.Y(n_246)
);

NAND2x1_ASAP7_75t_SL g216 ( 
.A(n_171),
.B(n_142),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_216),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_156),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_175),
.A2(n_190),
.B1(n_159),
.B2(n_177),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_223),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_178),
.B(n_135),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_178),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_177),
.A2(n_167),
.B1(n_157),
.B2(n_183),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_212),
.Y(n_244)
);

MAJx2_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_220),
.C(n_205),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_226),
.B(n_228),
.C(n_239),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_157),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_216),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_232),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_216),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_249),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_194),
.B(n_173),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_251),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_196),
.B(n_183),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_207),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_218),
.Y(n_258)
);

NAND2xp67_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_191),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_245),
.B(n_247),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_192),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_170),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_215),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_200),
.B(n_167),
.C(n_171),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_197),
.B(n_167),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_199),
.B(n_167),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_217),
.Y(n_265)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_201),
.Y(n_253)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_253),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_255),
.B(n_261),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_238),
.A2(n_221),
.B1(n_208),
.B2(n_203),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_257),
.A2(n_275),
.B1(n_234),
.B2(n_237),
.Y(n_279)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_258),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_192),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_259),
.B(n_228),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_225),
.A2(n_202),
.B(n_213),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_260),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_238),
.A2(n_219),
.B1(n_224),
.B2(n_223),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_235),
.A2(n_219),
.B1(n_210),
.B2(n_211),
.Y(n_262)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_262),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_225),
.A2(n_199),
.B(n_217),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_263),
.A2(n_274),
.B(n_230),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_233),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_267),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_271),
.Y(n_282)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_243),
.Y(n_270)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_270),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_248),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_240),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_244),
.A2(n_210),
.B1(n_217),
.B2(n_209),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_234),
.A2(n_204),
.B1(n_215),
.B2(n_158),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_241),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_239),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_278),
.B(n_268),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_279),
.A2(n_281),
.B1(n_261),
.B2(n_275),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_274),
.A2(n_257),
.B1(n_263),
.B2(n_227),
.Y(n_281)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_283),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_284),
.B(n_291),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_254),
.B(n_236),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_294),
.C(n_268),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_260),
.A2(n_232),
.B(n_231),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_289),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_206),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_290),
.B(n_292),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_256),
.A2(n_237),
.B(n_227),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_293),
.A2(n_271),
.B(n_267),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_254),
.B(n_226),
.C(n_252),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_295),
.Y(n_296)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_296),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_297),
.B(n_300),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_298),
.A2(n_306),
.B1(n_307),
.B2(n_287),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_303),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_283),
.Y(n_302)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_302),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_266),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_277),
.A2(n_266),
.B1(n_255),
.B2(n_273),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_277),
.A2(n_265),
.B1(n_264),
.B2(n_251),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_278),
.B(n_280),
.C(n_288),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_297),
.C(n_300),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_283),
.Y(n_310)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_310),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_316),
.Y(n_323)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_304),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_315),
.A2(n_286),
.B1(n_264),
.B2(n_305),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_280),
.Y(n_316)
);

OAI21xp33_ASAP7_75t_L g318 ( 
.A1(n_308),
.A2(n_295),
.B(n_272),
.Y(n_318)
);

MAJx2_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_299),
.C(n_301),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_320),
.C(n_317),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_303),
.B(n_293),
.Y(n_320)
);

NAND2xp33_ASAP7_75t_SL g321 ( 
.A(n_305),
.B(n_291),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_321),
.A2(n_289),
.B(n_282),
.Y(n_332)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_324),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_325),
.B(n_332),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_316),
.B(n_286),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_326),
.B(n_330),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_322),
.A2(n_313),
.B1(n_298),
.B2(n_315),
.Y(n_327)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_327),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_328),
.B(n_329),
.C(n_331),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_307),
.C(n_285),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_312),
.A2(n_287),
.B1(n_306),
.B2(n_285),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_281),
.C(n_279),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_323),
.B(n_314),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_333),
.B(n_335),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_323),
.B(n_292),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_329),
.B(n_311),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_337),
.B(n_320),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_336),
.B(n_325),
.C(n_331),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_341),
.B(n_342),
.Y(n_348)
);

AOI322xp5_ASAP7_75t_L g342 ( 
.A1(n_340),
.A2(n_328),
.A3(n_311),
.B1(n_253),
.B2(n_229),
.C1(n_269),
.C2(n_250),
.Y(n_342)
);

AOI322xp5_ASAP7_75t_L g344 ( 
.A1(n_334),
.A2(n_339),
.A3(n_336),
.B1(n_338),
.B2(n_333),
.C1(n_229),
.C2(n_246),
.Y(n_344)
);

NAND3xp33_ASAP7_75t_SL g346 ( 
.A(n_344),
.B(n_345),
.C(n_338),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_346),
.A2(n_347),
.B(n_341),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_343),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_349),
.A2(n_348),
.B(n_246),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_350),
.A2(n_193),
.B(n_206),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_351),
.A2(n_193),
.B(n_184),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_352),
.B(n_158),
.Y(n_353)
);


endmodule