module fake_jpeg_674_n_229 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_229);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_36),
.B(n_38),
.Y(n_95)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_3),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g82 ( 
.A(n_39),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_25),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_60),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_15),
.B(n_3),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_51),
.B(n_59),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_35),
.B(n_3),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_52),
.B(n_62),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_61),
.Y(n_71)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_17),
.B(n_4),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_67),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_64),
.B(n_65),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_66),
.B(n_6),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_69),
.Y(n_90)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_19),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_40),
.A2(n_22),
.B1(n_32),
.B2(n_26),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_78),
.A2(n_86),
.B1(n_10),
.B2(n_11),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_52),
.A2(n_22),
.B1(n_32),
.B2(n_26),
.Y(n_86)
);

NAND2x1_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_53),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_105),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_38),
.A2(n_31),
.B1(n_34),
.B2(n_25),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_89),
.A2(n_94),
.B1(n_106),
.B2(n_11),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_100),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_51),
.A2(n_34),
.B1(n_27),
.B2(n_7),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_36),
.B(n_27),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_59),
.B(n_5),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_101),
.B(n_102),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_60),
.B(n_5),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_62),
.B(n_66),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_104),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_64),
.B(n_6),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_65),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_98),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_41),
.C(n_43),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_130),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_97),
.A2(n_45),
.B(n_46),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_110),
.A2(n_123),
.B(n_87),
.Y(n_140)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_108),
.Y(n_111)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_108),
.Y(n_112)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_90),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_126),
.Y(n_142)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_9),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_117),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_77),
.B(n_10),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_118),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_119),
.A2(n_82),
.B1(n_88),
.B2(n_99),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_SL g144 ( 
.A1(n_120),
.A2(n_124),
.B(n_99),
.Y(n_144)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_77),
.A2(n_11),
.B(n_103),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_96),
.A2(n_85),
.B1(n_92),
.B2(n_73),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

NOR2xp67_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_103),
.Y(n_126)
);

AND2x2_ASAP7_75t_SL g127 ( 
.A(n_81),
.B(n_91),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_129),
.Y(n_145)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_81),
.Y(n_128)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_75),
.Y(n_129)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_133),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_71),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g135 ( 
.A(n_98),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_135),
.A2(n_88),
.B1(n_92),
.B2(n_87),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_136),
.Y(n_169)
);

AO22x1_ASAP7_75t_L g138 ( 
.A1(n_111),
.A2(n_96),
.B1(n_74),
.B2(n_75),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_139),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_134),
.A2(n_79),
.B1(n_83),
.B2(n_84),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_141),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_112),
.A2(n_79),
.B1(n_72),
.B2(n_80),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_150),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_121),
.A2(n_84),
.B1(n_74),
.B2(n_82),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_148),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_99),
.B(n_72),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_127),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_110),
.A2(n_80),
.B1(n_99),
.B2(n_129),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_158),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_119),
.A2(n_116),
.B1(n_117),
.B2(n_109),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_151),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_162),
.Y(n_183)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_152),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_165),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_142),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_114),
.C(n_123),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_153),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_167),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_131),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_173),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_113),
.Y(n_171)
);

A2O1A1O1Ixp25_ASAP7_75t_L g182 ( 
.A1(n_171),
.A2(n_149),
.B(n_130),
.C(n_138),
.D(n_157),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_172),
.A2(n_140),
.B(n_145),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_133),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_153),
.B(n_130),
.Y(n_174)
);

AOI322xp5_ASAP7_75t_SL g184 ( 
.A1(n_174),
.A2(n_138),
.A3(n_148),
.B1(n_127),
.B2(n_141),
.C1(n_135),
.C2(n_137),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_177),
.C(n_187),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_160),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_184),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_161),
.A2(n_156),
.B(n_147),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_161),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_171),
.B(n_166),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_159),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_168),
.A2(n_146),
.B1(n_149),
.B2(n_158),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_181),
.A2(n_188),
.B1(n_155),
.B2(n_163),
.Y(n_193)
);

AOI322xp5_ASAP7_75t_L g192 ( 
.A1(n_182),
.A2(n_164),
.A3(n_165),
.B1(n_172),
.B2(n_163),
.C1(n_159),
.C2(n_162),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_157),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_168),
.A2(n_155),
.B1(n_125),
.B2(n_154),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_189),
.A2(n_185),
.B(n_177),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_183),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_194),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_192),
.B(n_185),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_193),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_180),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_199),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_186),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_197),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_188),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_169),
.C(n_115),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_181),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_204),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_187),
.Y(n_204)
);

MAJx2_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_175),
.C(n_195),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_207),
.B(n_198),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_200),
.B(n_202),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_209),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_205),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_211),
.A2(n_207),
.B(n_182),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_190),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_213),
.C(n_190),
.Y(n_214)
);

MAJx2_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_154),
.C(n_128),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_215),
.A2(n_137),
.B1(n_118),
.B2(n_122),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_210),
.A2(n_199),
.B(n_189),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_217),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_205),
.C(n_178),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_213),
.C(n_193),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_221),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_220),
.B(n_135),
.Y(n_225)
);

OAI21x1_ASAP7_75t_L g223 ( 
.A1(n_222),
.A2(n_132),
.B(n_125),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_225),
.Y(n_227)
);

BUFx24_ASAP7_75t_SL g226 ( 
.A(n_224),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_226),
.A2(n_219),
.B(n_221),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_227),
.Y(n_229)
);


endmodule