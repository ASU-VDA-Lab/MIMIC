module real_aes_4519_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_503;
wire n_287;
wire n_357;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_582;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_85;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_150;
wire n_147;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_589;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_L g247 ( .A(n_0), .B(n_248), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_1), .Y(n_268) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_2), .Y(n_80) );
O2A1O1Ixp33_ASAP7_75t_SL g332 ( .A1(n_2), .A2(n_263), .B(n_333), .C(n_334), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_3), .B(n_148), .Y(n_147) );
OAI22xp33_ASAP7_75t_L g254 ( .A1(n_4), .A2(n_61), .B1(n_252), .B2(n_255), .Y(n_254) );
INVx1_ASAP7_75t_SL g186 ( .A(n_5), .Y(n_186) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_6), .Y(n_291) );
INVx1_ASAP7_75t_L g159 ( .A(n_7), .Y(n_159) );
OAI22xp5_ASAP7_75t_L g323 ( .A1(n_8), .A2(n_51), .B1(n_237), .B2(n_255), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_9), .Y(n_363) );
INVx1_ASAP7_75t_L g108 ( .A(n_10), .Y(n_108) );
INVxp67_ASAP7_75t_L g155 ( .A(n_10), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_10), .B(n_54), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g322 ( .A1(n_11), .A2(n_45), .B1(n_252), .B2(n_269), .Y(n_322) );
OA21x2_ASAP7_75t_L g224 ( .A1(n_12), .A2(n_50), .B(n_225), .Y(n_224) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_12), .A2(n_50), .B(n_225), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g103 ( .A(n_13), .B(n_92), .Y(n_103) );
AOI22xp33_ASAP7_75t_L g130 ( .A1(n_14), .A2(n_52), .B1(n_131), .B2(n_133), .Y(n_130) );
AOI22xp33_ASAP7_75t_L g85 ( .A1(n_15), .A2(n_72), .B1(n_86), .B2(n_111), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_16), .Y(n_284) );
BUFx3_ASAP7_75t_L g198 ( .A(n_17), .Y(n_198) );
AOI22xp33_ASAP7_75t_L g134 ( .A1(n_18), .A2(n_55), .B1(n_135), .B2(n_138), .Y(n_134) );
O2A1O1Ixp33_ASAP7_75t_L g338 ( .A1(n_19), .A2(n_256), .B(n_339), .C(n_340), .Y(n_338) );
OAI22xp33_ASAP7_75t_SL g251 ( .A1(n_20), .A2(n_33), .B1(n_231), .B2(n_252), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g230 ( .A1(n_21), .A2(n_26), .B1(n_231), .B2(n_233), .Y(n_230) );
BUFx6f_ASAP7_75t_L g92 ( .A(n_22), .Y(n_92) );
O2A1O1Ixp5_ASAP7_75t_L g302 ( .A1(n_23), .A2(n_263), .B(n_303), .C(n_304), .Y(n_302) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_23), .Y(n_604) );
XOR2xp5_ASAP7_75t_L g609 ( .A(n_24), .B(n_82), .Y(n_609) );
INVx1_ASAP7_75t_L g93 ( .A(n_25), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_25), .B(n_53), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_27), .B(n_241), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g305 ( .A(n_28), .Y(n_305) );
AOI221xp5_ASAP7_75t_L g163 ( .A1(n_29), .A2(n_65), .B1(n_164), .B2(n_166), .C(n_168), .Y(n_163) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_30), .Y(n_187) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_31), .Y(n_336) );
INVx1_ASAP7_75t_L g169 ( .A(n_32), .Y(n_169) );
INVx1_ASAP7_75t_L g225 ( .A(n_34), .Y(n_225) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_35), .Y(n_209) );
AND2x4_ASAP7_75t_L g226 ( .A(n_35), .B(n_207), .Y(n_226) );
AND2x4_ASAP7_75t_L g258 ( .A(n_35), .B(n_207), .Y(n_258) );
INVx1_ASAP7_75t_L g143 ( .A(n_36), .Y(n_143) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_37), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_38), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_L g287 ( .A1(n_39), .A2(n_263), .B(n_288), .C(n_290), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_40), .Y(n_311) );
INVx2_ASAP7_75t_L g368 ( .A(n_41), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_42), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_43), .B(n_272), .Y(n_271) );
AOI22xp5_ASAP7_75t_L g235 ( .A1(n_44), .A2(n_59), .B1(n_236), .B2(n_238), .Y(n_235) );
OA22x2_ASAP7_75t_L g98 ( .A1(n_46), .A2(n_54), .B1(n_92), .B2(n_96), .Y(n_98) );
INVx1_ASAP7_75t_L g118 ( .A(n_46), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_47), .Y(n_270) );
HB1xp67_ASAP7_75t_L g183 ( .A(n_48), .Y(n_183) );
NAND2xp33_ASAP7_75t_R g326 ( .A(n_49), .B(n_224), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_49), .A2(n_75), .B1(n_241), .B2(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g110 ( .A(n_53), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_53), .B(n_116), .Y(n_178) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_53), .Y(n_201) );
OAI21xp33_ASAP7_75t_L g119 ( .A1(n_54), .A2(n_60), .B(n_120), .Y(n_119) );
AOI22xp33_ASAP7_75t_L g121 ( .A1(n_56), .A2(n_64), .B1(n_122), .B2(n_126), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_57), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g364 ( .A(n_58), .Y(n_364) );
INVx1_ASAP7_75t_L g95 ( .A(n_60), .Y(n_95) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_60), .B(n_71), .Y(n_176) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_62), .Y(n_232) );
INVx1_ASAP7_75t_L g234 ( .A(n_62), .Y(n_234) );
BUFx5_ASAP7_75t_L g252 ( .A(n_62), .Y(n_252) );
INVx2_ASAP7_75t_L g344 ( .A(n_63), .Y(n_344) );
INVx2_ASAP7_75t_L g293 ( .A(n_66), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g341 ( .A(n_67), .Y(n_341) );
INVx2_ASAP7_75t_SL g207 ( .A(n_68), .Y(n_207) );
HB1xp67_ASAP7_75t_L g181 ( .A(n_69), .Y(n_181) );
INVx1_ASAP7_75t_L g309 ( .A(n_70), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g101 ( .A(n_71), .B(n_102), .Y(n_101) );
INVx2_ASAP7_75t_L g315 ( .A(n_73), .Y(n_315) );
OAI21xp33_ASAP7_75t_SL g282 ( .A1(n_74), .A2(n_252), .B(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_75), .B(n_241), .Y(n_358) );
INVxp67_ASAP7_75t_SL g392 ( .A(n_75), .Y(n_392) );
INVx1_ASAP7_75t_L g162 ( .A(n_76), .Y(n_162) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_193), .B1(n_210), .B2(n_594), .C(n_602), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_180), .Y(n_78) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_80), .A2(n_81), .B1(n_82), .B2(n_179), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_80), .Y(n_179) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_81), .A2(n_82), .B1(n_604), .B2(n_605), .Y(n_603) );
INVx1_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
NAND4xp75_ASAP7_75t_L g83 ( .A(n_84), .B(n_129), .C(n_141), .D(n_163), .Y(n_83) );
AND2x2_ASAP7_75t_L g84 ( .A(n_85), .B(n_121), .Y(n_84) );
BUFx12f_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AND2x4_ASAP7_75t_L g87 ( .A(n_88), .B(n_99), .Y(n_87) );
AND2x4_ASAP7_75t_L g123 ( .A(n_88), .B(n_124), .Y(n_123) );
AND2x4_ASAP7_75t_L g135 ( .A(n_88), .B(n_136), .Y(n_135) );
AND2x4_ASAP7_75t_L g138 ( .A(n_88), .B(n_139), .Y(n_138) );
AND2x4_ASAP7_75t_L g88 ( .A(n_89), .B(n_97), .Y(n_88) );
AND2x2_ASAP7_75t_L g146 ( .A(n_89), .B(n_98), .Y(n_146) );
INVx1_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
AND2x2_ASAP7_75t_L g132 ( .A(n_90), .B(n_98), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g90 ( .A(n_91), .B(n_94), .Y(n_90) );
NAND2xp33_ASAP7_75t_L g91 ( .A(n_92), .B(n_93), .Y(n_91) );
INVx2_ASAP7_75t_L g96 ( .A(n_92), .Y(n_96) );
INVx3_ASAP7_75t_L g102 ( .A(n_92), .Y(n_102) );
NAND2xp33_ASAP7_75t_L g109 ( .A(n_92), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g120 ( .A(n_92), .Y(n_120) );
HB1xp67_ASAP7_75t_L g151 ( .A(n_92), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_93), .B(n_118), .Y(n_117) );
INVxp67_ASAP7_75t_L g202 ( .A(n_93), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g94 ( .A(n_95), .B(n_96), .Y(n_94) );
OAI21xp5_ASAP7_75t_L g154 ( .A1(n_95), .A2(n_120), .B(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
AND2x2_ASAP7_75t_L g153 ( .A(n_98), .B(n_154), .Y(n_153) );
AND2x4_ASAP7_75t_L g113 ( .A(n_99), .B(n_114), .Y(n_113) );
AND2x4_ASAP7_75t_L g131 ( .A(n_99), .B(n_132), .Y(n_131) );
AND2x4_ASAP7_75t_L g99 ( .A(n_100), .B(n_104), .Y(n_99) );
OR2x2_ASAP7_75t_L g125 ( .A(n_100), .B(n_105), .Y(n_125) );
AND2x4_ASAP7_75t_L g136 ( .A(n_100), .B(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g140 ( .A(n_100), .Y(n_140) );
AND2x2_ASAP7_75t_L g149 ( .A(n_100), .B(n_150), .Y(n_149) );
AND2x4_ASAP7_75t_L g100 ( .A(n_101), .B(n_103), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_102), .B(n_108), .Y(n_107) );
INVxp67_ASAP7_75t_L g116 ( .A(n_102), .Y(n_116) );
NAND3xp33_ASAP7_75t_L g177 ( .A(n_103), .B(n_115), .C(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g137 ( .A(n_106), .Y(n_137) );
AND2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_109), .Y(n_106) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx8_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x4_ASAP7_75t_L g128 ( .A(n_114), .B(n_124), .Y(n_128) );
AND2x4_ASAP7_75t_L g161 ( .A(n_114), .B(n_139), .Y(n_161) );
AND2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_119), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
HB1xp67_ASAP7_75t_L g203 ( .A(n_118), .Y(n_203) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x4_ASAP7_75t_L g133 ( .A(n_124), .B(n_132), .Y(n_133) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx3_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx6_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_134), .Y(n_129) );
AND2x4_ASAP7_75t_L g158 ( .A(n_132), .B(n_136), .Y(n_158) );
AND2x2_ASAP7_75t_L g165 ( .A(n_132), .B(n_139), .Y(n_165) );
AND2x4_ASAP7_75t_L g145 ( .A(n_136), .B(n_146), .Y(n_145) );
AND2x4_ASAP7_75t_L g139 ( .A(n_137), .B(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g167 ( .A(n_139), .B(n_146), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_142), .B(n_156), .Y(n_141) );
OAI21xp33_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_144), .B(n_147), .Y(n_142) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x4_ASAP7_75t_L g148 ( .A(n_149), .B(n_153), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
INVx1_ASAP7_75t_L g173 ( .A(n_151), .Y(n_173) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_152), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_159), .B1(n_160), .B2(n_162), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
HB1xp67_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
HB1xp67_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AO21x2_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_177), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_175), .B(n_176), .Y(n_174) );
AOI22xp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B1(n_191), .B2(n_192), .Y(n_180) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_181), .Y(n_191) );
CKINVDCx16_ASAP7_75t_R g192 ( .A(n_182), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B1(n_185), .B2(n_190), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_183), .Y(n_190) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
OAI22xp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B1(n_188), .B2(n_189), .Y(n_185) );
INVx1_ASAP7_75t_L g188 ( .A(n_186), .Y(n_188) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_187), .Y(n_189) );
BUFx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_196), .B(n_204), .Y(n_195) );
INVxp67_ASAP7_75t_SL g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g607 ( .A(n_197), .B(n_204), .Y(n_607) );
AOI211xp5_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_200), .C(n_203), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_201), .B(n_202), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_205), .B(n_208), .Y(n_204) );
OR2x2_ASAP7_75t_L g611 ( .A(n_205), .B(n_209), .Y(n_611) );
INVx1_ASAP7_75t_L g614 ( .A(n_205), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_205), .B(n_208), .Y(n_615) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
HB1xp67_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx2_ASAP7_75t_SL g211 ( .A(n_212), .Y(n_211) );
AND2x4_ASAP7_75t_L g212 ( .A(n_213), .B(n_464), .Y(n_212) );
AND4x1_ASAP7_75t_L g213 ( .A(n_214), .B(n_412), .C(n_432), .D(n_444), .Y(n_213) );
AOI311xp33_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_294), .A3(n_327), .B(n_345), .C(n_382), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_217), .B(n_274), .Y(n_216) );
AND2x4_ASAP7_75t_L g217 ( .A(n_218), .B(n_244), .Y(n_217) );
INVx3_ASAP7_75t_L g381 ( .A(n_218), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_218), .B(n_405), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_218), .B(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g534 ( .A(n_218), .B(n_518), .Y(n_534) );
INVx3_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g423 ( .A(n_219), .B(n_349), .Y(n_423) );
INVx1_ASAP7_75t_L g486 ( .A(n_219), .Y(n_486) );
AND2x2_ASAP7_75t_L g528 ( .A(n_219), .B(n_259), .Y(n_528) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g504 ( .A(n_220), .Y(n_504) );
OAI21x1_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_227), .B(n_240), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_222), .B(n_226), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_222), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
BUFx3_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g280 ( .A(n_224), .Y(n_280) );
INVx1_ASAP7_75t_L g316 ( .A(n_224), .Y(n_316) );
INVx2_ASAP7_75t_L g377 ( .A(n_224), .Y(n_377) );
AND2x2_ASAP7_75t_L g279 ( .A(n_226), .B(n_280), .Y(n_279) );
INVx4_ASAP7_75t_L g312 ( .A(n_226), .Y(n_312) );
INVx1_ASAP7_75t_L g399 ( .A(n_227), .Y(n_399) );
OA22x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_230), .B1(n_235), .B2(n_239), .Y(n_227) );
INVx4_ASAP7_75t_L g601 ( .A(n_228), .Y(n_601) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g239 ( .A(n_229), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_229), .B(n_251), .Y(n_250) );
INVx3_ASAP7_75t_L g256 ( .A(n_229), .Y(n_256) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_229), .Y(n_263) );
INVx4_ASAP7_75t_L g286 ( .A(n_229), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_229), .B(n_309), .Y(n_308) );
INVx2_ASAP7_75t_SL g238 ( .A(n_231), .Y(n_238) );
AOI22xp33_ASAP7_75t_SL g264 ( .A1(n_231), .A2(n_252), .B1(n_265), .B2(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g335 ( .A(n_231), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g362 ( .A1(n_231), .A2(n_252), .B1(n_363), .B2(n_364), .Y(n_362) );
INVx6_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx2_ASAP7_75t_L g255 ( .A(n_232), .Y(n_255) );
INVx2_ASAP7_75t_L g269 ( .A(n_232), .Y(n_269) );
INVx3_ASAP7_75t_L g289 ( .A(n_232), .Y(n_289) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_233), .B(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_233), .B(n_341), .Y(n_340) );
AOI22xp5_ASAP7_75t_L g366 ( .A1(n_233), .A2(n_269), .B1(n_367), .B2(n_368), .Y(n_366) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx2_ASAP7_75t_L g237 ( .A(n_234), .Y(n_237) );
INVx1_ASAP7_75t_L g333 ( .A(n_236), .Y(n_333) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g402 ( .A(n_240), .Y(n_402) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g248 ( .A(n_242), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_242), .B(n_258), .Y(n_257) );
NOR2xp33_ASAP7_75t_SL g343 ( .A(n_242), .B(n_344), .Y(n_343) );
INVx4_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g273 ( .A(n_243), .Y(n_273) );
BUFx3_ASAP7_75t_L g401 ( .A(n_243), .Y(n_401) );
AND2x2_ASAP7_75t_L g515 ( .A(n_244), .B(n_381), .Y(n_515) );
INVx1_ASAP7_75t_SL g539 ( .A(n_244), .Y(n_539) );
AND2x2_ASAP7_75t_L g552 ( .A(n_244), .B(n_503), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_244), .B(n_347), .Y(n_553) );
AND2x4_ASAP7_75t_L g244 ( .A(n_245), .B(n_259), .Y(n_244) );
AND2x2_ASAP7_75t_L g436 ( .A(n_245), .B(n_277), .Y(n_436) );
INVx3_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g349 ( .A(n_246), .Y(n_349) );
NAND2xp33_ASAP7_75t_R g395 ( .A(n_246), .B(n_277), .Y(n_395) );
AND2x2_ASAP7_75t_L g405 ( .A(n_246), .B(n_259), .Y(n_405) );
INVx1_ASAP7_75t_L g476 ( .A(n_246), .Y(n_476) );
AND2x2_ASAP7_75t_L g518 ( .A(n_246), .B(n_277), .Y(n_518) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_246), .Y(n_545) );
AND2x4_ASAP7_75t_L g246 ( .A(n_247), .B(n_249), .Y(n_246) );
INVx2_ASAP7_75t_L g261 ( .A(n_248), .Y(n_261) );
NOR2xp33_ASAP7_75t_SL g342 ( .A(n_248), .B(n_312), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_253), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g267 ( .A1(n_252), .A2(n_268), .B1(n_269), .B2(n_270), .Y(n_267) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_252), .B(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_252), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_252), .B(n_311), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_256), .B(n_257), .Y(n_253) );
OAI221xp5_ASAP7_75t_L g262 ( .A1(n_256), .A2(n_258), .B1(n_263), .B2(n_264), .C(n_267), .Y(n_262) );
INVx1_ASAP7_75t_L g325 ( .A(n_258), .Y(n_325) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_258), .Y(n_389) );
OR2x2_ASAP7_75t_L g397 ( .A(n_259), .B(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g485 ( .A(n_259), .B(n_486), .Y(n_485) );
OA21x2_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_262), .B(n_271), .Y(n_259) );
OA21x2_ASAP7_75t_L g351 ( .A1(n_260), .A2(n_262), .B(n_271), .Y(n_351) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g391 ( .A(n_261), .B(n_392), .Y(n_391) );
AOI22xp5_ASAP7_75t_L g321 ( .A1(n_263), .A2(n_286), .B1(n_322), .B2(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g369 ( .A(n_263), .Y(n_369) );
OAI22xp33_ASAP7_75t_L g390 ( .A1(n_263), .A2(n_286), .B1(n_362), .B2(n_366), .Y(n_390) );
INVx1_ASAP7_75t_L g339 ( .A(n_269), .Y(n_339) );
NOR2xp67_ASAP7_75t_L g324 ( .A(n_272), .B(n_325), .Y(n_324) );
INVx3_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_273), .B(n_293), .Y(n_292) );
BUFx3_ASAP7_75t_L g313 ( .A(n_273), .Y(n_313) );
AND2x2_ASAP7_75t_L g548 ( .A(n_274), .B(n_529), .Y(n_548) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g557 ( .A(n_275), .B(n_495), .Y(n_557) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g404 ( .A(n_276), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g498 ( .A(n_276), .Y(n_498) );
AND2x2_ASAP7_75t_L g503 ( .A(n_276), .B(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
BUFx2_ASAP7_75t_L g347 ( .A(n_277), .Y(n_347) );
INVx2_ASAP7_75t_L g418 ( .A(n_277), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_277), .B(n_351), .Y(n_421) );
INVx1_ASAP7_75t_L g448 ( .A(n_277), .Y(n_448) );
OR2x2_ASAP7_75t_L g455 ( .A(n_277), .B(n_349), .Y(n_455) );
AND2x2_ASAP7_75t_L g489 ( .A(n_277), .B(n_490), .Y(n_489) );
INVx3_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AOI21x1_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_281), .B(n_292), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_285), .B(n_287), .Y(n_281) );
AOI221xp5_ASAP7_75t_L g360 ( .A1(n_285), .A2(n_312), .B1(n_361), .B2(n_365), .C(n_369), .Y(n_360) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g306 ( .A1(n_286), .A2(n_307), .B1(n_308), .B2(n_310), .Y(n_306) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g303 ( .A(n_289), .Y(n_303) );
INVx1_ASAP7_75t_L g307 ( .A(n_289), .Y(n_307) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
BUFx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_296), .B(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g472 ( .A(n_297), .B(n_409), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_317), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_298), .B(n_357), .Y(n_580) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g459 ( .A(n_299), .B(n_319), .Y(n_459) );
AND2x2_ASAP7_75t_L g480 ( .A(n_299), .B(n_373), .Y(n_480) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
BUFx2_ASAP7_75t_R g354 ( .A(n_300), .Y(n_354) );
INVx2_ASAP7_75t_L g411 ( .A(n_300), .Y(n_411) );
AND2x2_ASAP7_75t_L g461 ( .A(n_300), .B(n_462), .Y(n_461) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_300), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_300), .B(n_330), .Y(n_509) );
AND2x2_ASAP7_75t_L g514 ( .A(n_300), .B(n_430), .Y(n_514) );
AO21x2_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_313), .B(n_314), .Y(n_300) );
NOR3xp33_ASAP7_75t_L g301 ( .A(n_302), .B(n_306), .C(n_312), .Y(n_301) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_305), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g359 ( .A(n_313), .B(n_360), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x4_ASAP7_75t_L g410 ( .A(n_318), .B(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g583 ( .A(n_318), .B(n_430), .Y(n_583) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g386 ( .A(n_319), .B(n_387), .Y(n_386) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_319), .Y(n_427) );
INVx1_ASAP7_75t_L g462 ( .A(n_319), .Y(n_462) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_326), .Y(n_319) );
AND2x2_ASAP7_75t_L g374 ( .A(n_320), .B(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_324), .Y(n_320) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx2_ASAP7_75t_SL g479 ( .A(n_329), .Y(n_479) );
INVx1_ASAP7_75t_L g501 ( .A(n_329), .Y(n_501) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g356 ( .A(n_330), .B(n_357), .Y(n_356) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_330), .Y(n_378) );
INVx1_ASAP7_75t_L g385 ( .A(n_330), .Y(n_385) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_330), .Y(n_409) );
AND2x4_ASAP7_75t_L g414 ( .A(n_330), .B(n_387), .Y(n_414) );
INVx2_ASAP7_75t_L g430 ( .A(n_330), .Y(n_430) );
AND2x2_ASAP7_75t_L g440 ( .A(n_330), .B(n_357), .Y(n_440) );
AO31x2_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_337), .A3(n_342), .B(n_343), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_339), .Y(n_598) );
OAI22xp33_ASAP7_75t_SL g345 ( .A1(n_346), .A2(n_352), .B1(n_370), .B2(n_379), .Y(n_345) );
NAND2x1p5_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
AND2x2_ASAP7_75t_L g380 ( .A(n_348), .B(n_381), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_348), .A2(n_433), .B1(n_437), .B2(n_443), .Y(n_432) );
AND2x4_ASAP7_75t_L g529 ( .A(n_348), .B(n_530), .Y(n_529) );
NAND2x1p5_ASAP7_75t_L g574 ( .A(n_348), .B(n_497), .Y(n_574) );
AND2x4_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
AND2x4_ASAP7_75t_L g495 ( .A(n_350), .B(n_398), .Y(n_495) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g490 ( .A(n_351), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_355), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x4_ASAP7_75t_L g564 ( .A(n_355), .B(n_461), .Y(n_564) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g468 ( .A(n_356), .B(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_357), .B(n_411), .Y(n_431) );
AND2x2_ASAP7_75t_L g463 ( .A(n_357), .B(n_385), .Y(n_463) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
AND2x2_ASAP7_75t_L g373 ( .A(n_359), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AOI21xp33_ASAP7_75t_L g587 ( .A1(n_370), .A2(n_588), .B(n_591), .Y(n_587) );
HB1xp67_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_378), .Y(n_371) );
OR2x2_ASAP7_75t_L g550 ( .A(n_372), .B(n_385), .Y(n_550) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g571 ( .A(n_373), .Y(n_571) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g445 ( .A(n_381), .B(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g522 ( .A(n_381), .B(n_405), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_393), .B1(n_403), .B2(n_406), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
AND2x4_ASAP7_75t_L g507 ( .A(n_386), .B(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g513 ( .A(n_386), .B(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g451 ( .A(n_387), .Y(n_451) );
OAI21x1_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_390), .B(n_391), .Y(n_387) );
AND2x2_ASAP7_75t_L g595 ( .A(n_389), .B(n_596), .Y(n_595) );
INVxp67_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_396), .B(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g592 ( .A(n_396), .B(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g456 ( .A(n_397), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_400), .B(n_402), .Y(n_398) );
INVx3_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NAND2xp33_ASAP7_75t_L g532 ( .A(n_403), .B(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx3_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_408), .B(n_410), .Y(n_407) );
INVxp67_ASAP7_75t_L g524 ( .A(n_408), .Y(n_524) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g413 ( .A(n_410), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g439 ( .A(n_410), .B(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g446 ( .A(n_410), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g520 ( .A(n_410), .B(n_479), .Y(n_520) );
OAI31xp33_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_415), .A3(n_417), .B(n_419), .Y(n_412) );
INVx2_ASAP7_75t_L g424 ( .A(n_413), .Y(n_424) );
INVx2_ASAP7_75t_SL g442 ( .A(n_414), .Y(n_442) );
AND2x2_ASAP7_75t_L g458 ( .A(n_414), .B(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g555 ( .A(n_414), .B(n_469), .Y(n_555) );
AND2x4_ASAP7_75t_L g575 ( .A(n_414), .B(n_461), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_414), .B(n_426), .Y(n_590) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
A2O1A1Ixp33_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_422), .B(n_424), .C(n_425), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
NOR2xp67_ASAP7_75t_L g475 ( .A(n_421), .B(n_476), .Y(n_475) );
OAI22xp33_ASAP7_75t_L g452 ( .A1(n_422), .A2(n_453), .B1(n_457), .B2(n_460), .Y(n_452) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g443 ( .A(n_425), .Y(n_443) );
OR2x2_ASAP7_75t_L g425 ( .A(n_426), .B(n_428), .Y(n_425) );
OR2x2_ASAP7_75t_L g441 ( .A(n_426), .B(n_442), .Y(n_441) );
AOI322xp5_ASAP7_75t_L g525 ( .A1(n_426), .A2(n_449), .A3(n_526), .B1(n_529), .B2(n_531), .C1(n_532), .C2(n_535), .Y(n_525) );
INVx2_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g586 ( .A(n_428), .Y(n_586) );
OR2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_431), .Y(n_428) );
INVx1_ASAP7_75t_L g562 ( .A(n_429), .Y(n_562) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g584 ( .A(n_431), .Y(n_584) );
INVxp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g493 ( .A(n_436), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_441), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g535 ( .A(n_440), .B(n_461), .Y(n_535) );
INVx2_ASAP7_75t_L g541 ( .A(n_441), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_449), .B(n_452), .Y(n_444) );
INVx1_ASAP7_75t_L g511 ( .A(n_446), .Y(n_511) );
INVx1_ASAP7_75t_L g483 ( .A(n_447), .Y(n_483) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_448), .B(n_490), .Y(n_568) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_450), .B(n_492), .Y(n_531) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_456), .Y(n_453) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g593 ( .A(n_455), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_456), .A2(n_582), .B1(n_585), .B2(n_586), .Y(n_581) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g561 ( .A(n_459), .B(n_562), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_460), .A2(n_478), .B1(n_481), .B2(n_487), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_463), .Y(n_460) );
INVx2_ASAP7_75t_SL g492 ( .A(n_461), .Y(n_492) );
NOR2xp67_ASAP7_75t_L g464 ( .A(n_465), .B(n_546), .Y(n_464) );
NAND4xp25_ASAP7_75t_L g465 ( .A(n_466), .B(n_505), .C(n_525), .D(n_536), .Y(n_465) );
NOR3xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_477), .C(n_491), .Y(n_466) );
AOI21xp33_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_471), .B(n_473), .Y(n_467) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx2_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
NAND2x1p5_ASAP7_75t_SL g478 ( .A(n_479), .B(n_480), .Y(n_478) );
INVx1_ASAP7_75t_L g499 ( .A(n_480), .Y(n_499) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_480), .Y(n_558) );
INVxp33_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
NOR2x1_ASAP7_75t_L g482 ( .A(n_483), .B(n_484), .Y(n_482) );
INVx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
OAI322xp33_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_493), .A3(n_494), .B1(n_496), .B2(n_499), .C1(n_500), .C2(n_502), .Y(n_491) );
OR2x2_ASAP7_75t_L g523 ( .A(n_492), .B(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g506 ( .A(n_494), .Y(n_506) );
INVx2_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_495), .B(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g540 ( .A(n_497), .Y(n_540) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
OAI21xp33_ASAP7_75t_L g510 ( .A1(n_501), .A2(n_511), .B(n_512), .Y(n_510) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g530 ( .A(n_504), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_504), .B(n_545), .Y(n_544) );
AOI221x1_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_507), .B1(n_510), .B2(n_515), .C(n_516), .Y(n_505) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
OR2x2_ASAP7_75t_L g570 ( .A(n_509), .B(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_513), .A2(n_548), .B(n_549), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_519), .B1(n_521), .B2(n_523), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_518), .B(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_520), .A2(n_537), .B1(n_541), .B2(n_542), .Y(n_536) );
OAI221xp5_ASAP7_75t_SL g576 ( .A1(n_521), .A2(n_570), .B1(n_577), .B2(n_578), .C(n_581), .Y(n_576) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_539), .B(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g543 ( .A(n_540), .B(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_544), .Y(n_577) );
INVxp67_ASAP7_75t_L g567 ( .A(n_545), .Y(n_567) );
NAND3xp33_ASAP7_75t_L g546 ( .A(n_547), .B(n_556), .C(n_572), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_551), .B1(n_553), .B2(n_554), .Y(n_549) );
INVxp67_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AOI221xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_558), .B1(n_559), .B2(n_565), .C(n_569), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_563), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
INVx1_ASAP7_75t_L g585 ( .A(n_568), .Y(n_585) );
AOI211xp5_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_575), .B(n_576), .C(n_587), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
BUFx4f_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
OA21x2_ASAP7_75t_L g613 ( .A1(n_596), .A2(n_614), .B(n_615), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_599), .Y(n_596) );
CKINVDCx16_ASAP7_75t_R g597 ( .A(n_598), .Y(n_597) );
CKINVDCx20_ASAP7_75t_R g599 ( .A(n_600), .Y(n_599) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
OAI222xp33_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_606), .B1(n_608), .B2(n_610), .C1(n_612), .C2(n_616), .Y(n_602) );
CKINVDCx20_ASAP7_75t_R g605 ( .A(n_604), .Y(n_605) );
INVx1_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
BUFx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
endmodule