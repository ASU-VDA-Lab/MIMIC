module fake_netlist_5_405_n_1148 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_1148);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_1148;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_1126;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_1141;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_928;
wire n_1139;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_721;
wire n_998;
wire n_841;
wire n_1050;
wire n_1099;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_245;
wire n_501;
wire n_823;
wire n_725;
wire n_983;
wire n_1128;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_1112;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_1120;
wire n_915;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_864;
wire n_859;
wire n_1110;
wire n_951;
wire n_1121;
wire n_821;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_949;
wire n_854;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_946;
wire n_417;
wire n_1048;
wire n_932;
wire n_612;
wire n_1001;
wire n_385;
wire n_498;
wire n_516;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_1118;
wire n_509;
wire n_568;
wire n_947;
wire n_373;
wire n_820;
wire n_757;
wire n_1090;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_1024;
wire n_556;
wire n_1063;
wire n_1107;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_1143;
wire n_804;
wire n_867;
wire n_1124;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_1104;
wire n_563;
wire n_756;
wire n_1145;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_394;
wire n_250;
wire n_579;
wire n_992;
wire n_1049;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_1135;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_406;
wire n_519;
wire n_470;
wire n_919;
wire n_782;
wire n_908;
wire n_1108;
wire n_325;
wire n_449;
wire n_1073;
wire n_1100;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_291;
wire n_1147;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_976;
wire n_1096;
wire n_1095;
wire n_234;
wire n_343;
wire n_428;
wire n_308;
wire n_379;
wire n_267;
wire n_570;
wire n_457;
wire n_514;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_1142;
wire n_660;
wire n_223;
wire n_1114;
wire n_1129;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_995;
wire n_961;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_1062;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_922;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_816;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_680;
wire n_974;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_1119;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_1064;
wire n_923;
wire n_772;
wire n_691;
wire n_1134;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_342;
wire n_482;
wire n_517;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_236;
wire n_1069;
wire n_1075;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_477;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_990;
wire n_836;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_1113;
wire n_652;
wire n_778;
wire n_1111;
wire n_1122;
wire n_306;
wire n_1093;
wire n_722;
wire n_907;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_1102;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_1015;
wire n_1000;
wire n_891;
wire n_1140;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_1058;
wire n_362;
wire n_876;
wire n_332;
wire n_1053;
wire n_1101;
wire n_273;
wire n_585;
wire n_349;
wire n_1106;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_1014;
wire n_917;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_1052;
wire n_963;
wire n_954;
wire n_627;
wire n_1116;
wire n_767;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_1091;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_1059;
wire n_1084;
wire n_1131;
wire n_1133;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_607;
wire n_575;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_707;
wire n_710;
wire n_795;
wire n_695;
wire n_832;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_1072;
wire n_1130;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_1027;
wire n_971;
wire n_490;
wire n_805;
wire n_910;
wire n_326;
wire n_794;
wire n_996;
wire n_921;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_572;
wire n_366;
wire n_712;
wire n_754;
wire n_847;
wire n_936;
wire n_815;
wire n_1136;
wire n_246;
wire n_596;
wire n_1125;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_1109;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_1080;
wire n_266;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_1038;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_811;
wire n_766;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_1092;
wire n_238;
wire n_1117;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_1138;
wire n_536;
wire n_531;
wire n_1004;
wire n_935;
wire n_242;
wire n_817;
wire n_1032;
wire n_360;
wire n_594;
wire n_764;
wire n_872;
wire n_1056;
wire n_960;
wire n_890;
wire n_759;
wire n_1018;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_1123;
wire n_985;
wire n_904;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_1144;
wire n_1137;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_183),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_58),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_156),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_41),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_122),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_81),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_70),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_150),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_97),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_62),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_190),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_145),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_107),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_7),
.Y(n_235)
);

BUFx5_ASAP7_75t_L g236 ( 
.A(n_67),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_159),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_44),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_217),
.Y(n_239)
);

INVxp67_ASAP7_75t_SL g240 ( 
.A(n_144),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_174),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_215),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_57),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_113),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_102),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_128),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_202),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_77),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_124),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_180),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_23),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_152),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_170),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_198),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_188),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_115),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_17),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_23),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_28),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_37),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_54),
.Y(n_261)
);

BUFx8_ASAP7_75t_SL g262 ( 
.A(n_173),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_136),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_151),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_78),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_155),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_92),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_16),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_139),
.Y(n_269)
);

INVxp33_ASAP7_75t_SL g270 ( 
.A(n_52),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_18),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_117),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_42),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_197),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_141),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_206),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_104),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_68),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_207),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_108),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_74),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_132),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_209),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_20),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_171),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_2),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_86),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_204),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_13),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_172),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_120),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_59),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_46),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_50),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_257),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_251),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_286),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_228),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_228),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_222),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_231),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_235),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_258),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_268),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_284),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_238),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_262),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_223),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_236),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_289),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_233),
.Y(n_311)
);

INVxp33_ASAP7_75t_L g312 ( 
.A(n_262),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_234),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_239),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_236),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_278),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_241),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_242),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_236),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_271),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_255),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_259),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_237),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_266),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g325 ( 
.A(n_271),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_272),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_236),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_275),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_283),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_285),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_287),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_294),
.Y(n_332)
);

INVxp33_ASAP7_75t_SL g333 ( 
.A(n_221),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_231),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_294),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_246),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_246),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_247),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_260),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_260),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_263),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_224),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_236),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_298),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_300),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_299),
.Y(n_346)
);

OAI22x1_ASAP7_75t_R g347 ( 
.A1(n_295),
.A2(n_310),
.B1(n_338),
.B2(n_323),
.Y(n_347)
);

BUFx8_ASAP7_75t_L g348 ( 
.A(n_325),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_301),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_323),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_342),
.B(n_282),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_301),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_309),
.Y(n_353)
);

OAI21x1_ASAP7_75t_L g354 ( 
.A1(n_343),
.A2(n_291),
.B(n_263),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_341),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_341),
.Y(n_356)
);

INVx5_ASAP7_75t_L g357 ( 
.A(n_309),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_316),
.A2(n_270),
.B1(n_279),
.B2(n_252),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_342),
.B(n_292),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_332),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_308),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_311),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_315),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_331),
.B(n_291),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_296),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_335),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_336),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_333),
.B(n_225),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_339),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_302),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_340),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_315),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_307),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_333),
.B(n_293),
.Y(n_374)
);

BUFx2_ASAP7_75t_L g375 ( 
.A(n_302),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_319),
.Y(n_376)
);

CKINVDCx8_ASAP7_75t_R g377 ( 
.A(n_307),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_316),
.B(n_320),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_343),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_319),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_303),
.B(n_226),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_297),
.Y(n_382)
);

OAI21x1_ASAP7_75t_L g383 ( 
.A1(n_327),
.A2(n_240),
.B(n_236),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_313),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_334),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_306),
.B(n_290),
.Y(n_386)
);

OA21x2_ASAP7_75t_L g387 ( 
.A1(n_327),
.A2(n_229),
.B(n_227),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_303),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_304),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_304),
.B(n_230),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_305),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_337),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_338),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_328),
.B(n_288),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_314),
.Y(n_395)
);

OAI21x1_ASAP7_75t_L g396 ( 
.A1(n_330),
.A2(n_243),
.B(n_232),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_317),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_318),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_348),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_372),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_348),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_348),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_389),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_345),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_389),
.Y(n_405)
);

NAND2xp33_ASAP7_75t_R g406 ( 
.A(n_375),
.B(n_0),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_393),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_393),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_375),
.Y(n_409)
);

INVx2_ASAP7_75t_SL g410 ( 
.A(n_392),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_R g411 ( 
.A(n_373),
.B(n_377),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_350),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_373),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_377),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_347),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_390),
.Y(n_416)
);

INVx2_ASAP7_75t_SL g417 ( 
.A(n_391),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_376),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_388),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_388),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_370),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_372),
.Y(n_422)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_385),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_362),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_372),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_372),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_368),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_353),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_374),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_384),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_395),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_358),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_381),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_378),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_395),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_386),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_365),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_351),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_359),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_394),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_344),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_376),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_365),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_344),
.Y(n_444)
);

BUFx2_ASAP7_75t_L g445 ( 
.A(n_385),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_346),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_379),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_379),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_346),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_361),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_372),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_382),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_361),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_364),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_397),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_397),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_398),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_398),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_382),
.B(n_312),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_360),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_371),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_371),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_387),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_360),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_371),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_366),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_371),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_366),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_387),
.B(n_353),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_349),
.B(n_321),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_367),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_367),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_371),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_R g474 ( 
.A(n_349),
.B(n_295),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_436),
.B(n_387),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_423),
.B(n_326),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_470),
.B(n_369),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_446),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_431),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_428),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_445),
.B(n_369),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_435),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_428),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_410),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_463),
.B(n_353),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_437),
.Y(n_486)
);

AND2x2_ASAP7_75t_SL g487 ( 
.A(n_432),
.B(n_310),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_438),
.B(n_253),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_443),
.B(n_383),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g490 ( 
.A(n_474),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_427),
.B(n_261),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_452),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_455),
.B(n_322),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_418),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_L g495 ( 
.A1(n_469),
.A2(n_396),
.B1(n_383),
.B2(n_354),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_404),
.B(n_352),
.Y(n_496)
);

INVxp67_ASAP7_75t_SL g497 ( 
.A(n_425),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_424),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_412),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g500 ( 
.A(n_411),
.Y(n_500)
);

AND2x2_ASAP7_75t_SL g501 ( 
.A(n_409),
.B(n_281),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_418),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_440),
.B(n_442),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_442),
.B(n_363),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_429),
.B(n_244),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_447),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_430),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_447),
.B(n_363),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_460),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_464),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_416),
.B(n_245),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_411),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_441),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_456),
.B(n_248),
.Y(n_514)
);

INVx1_ASAP7_75t_SL g515 ( 
.A(n_474),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_448),
.A2(n_396),
.B1(n_462),
.B2(n_461),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_454),
.B(n_249),
.Y(n_517)
);

BUFx8_ASAP7_75t_SL g518 ( 
.A(n_415),
.Y(n_518)
);

OAI21xp33_ASAP7_75t_L g519 ( 
.A1(n_457),
.A2(n_329),
.B(n_324),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_466),
.Y(n_520)
);

INVx6_ASAP7_75t_L g521 ( 
.A(n_425),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_458),
.B(n_417),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_468),
.B(n_352),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_471),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_472),
.Y(n_525)
);

INVx6_ASAP7_75t_L g526 ( 
.A(n_425),
.Y(n_526)
);

AND2x6_ASAP7_75t_L g527 ( 
.A(n_422),
.B(n_426),
.Y(n_527)
);

INVx4_ASAP7_75t_L g528 ( 
.A(n_425),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_448),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_450),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_453),
.Y(n_531)
);

INVx5_ASAP7_75t_L g532 ( 
.A(n_451),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_444),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_400),
.B(n_363),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_451),
.B(n_380),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_449),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_465),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_451),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_467),
.Y(n_539)
);

AND2x6_ASAP7_75t_L g540 ( 
.A(n_473),
.B(n_451),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_407),
.Y(n_541)
);

AO22x2_ASAP7_75t_L g542 ( 
.A1(n_406),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_419),
.B(n_420),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_SL g544 ( 
.A(n_433),
.B(n_250),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_421),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_403),
.B(n_356),
.Y(n_546)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_414),
.Y(n_547)
);

INVxp67_ASAP7_75t_SL g548 ( 
.A(n_406),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_405),
.B(n_439),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_459),
.B(n_356),
.Y(n_550)
);

INVxp67_ASAP7_75t_SL g551 ( 
.A(n_434),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_413),
.A2(n_274),
.B1(n_256),
.B2(n_264),
.Y(n_552)
);

AND3x4_ASAP7_75t_L g553 ( 
.A(n_408),
.B(n_1),
.C(n_3),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_399),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_401),
.A2(n_354),
.B1(n_355),
.B2(n_380),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_SL g556 ( 
.A(n_402),
.B(n_254),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_431),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_463),
.A2(n_355),
.B1(n_380),
.B2(n_276),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_436),
.B(n_355),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_460),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_479),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_482),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_529),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_488),
.B(n_265),
.Y(n_564)
);

AND2x6_ASAP7_75t_L g565 ( 
.A(n_489),
.B(n_355),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_486),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_506),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_506),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_494),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_503),
.B(n_355),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_507),
.B(n_25),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_502),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_475),
.A2(n_280),
.B1(n_277),
.B2(n_273),
.Y(n_573)
);

AND2x6_ASAP7_75t_L g574 ( 
.A(n_489),
.B(n_26),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_557),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_496),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_503),
.B(n_267),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_481),
.B(n_27),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_475),
.A2(n_269),
.B1(n_357),
.B2(n_109),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_500),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_548),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_559),
.B(n_357),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_559),
.B(n_357),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_499),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_496),
.Y(n_585)
);

BUFx4f_ASAP7_75t_L g586 ( 
.A(n_530),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_537),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_476),
.B(n_3),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_539),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_548),
.B(n_4),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_522),
.B(n_4),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_511),
.B(n_5),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_480),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_477),
.B(n_357),
.Y(n_594)
);

BUFx8_ASAP7_75t_L g595 ( 
.A(n_554),
.Y(n_595)
);

OR2x2_ASAP7_75t_SL g596 ( 
.A(n_531),
.B(n_5),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_483),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_523),
.B(n_357),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_504),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_SL g600 ( 
.A1(n_487),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_504),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_523),
.B(n_6),
.Y(n_602)
);

BUFx4f_ASAP7_75t_L g603 ( 
.A(n_533),
.Y(n_603)
);

INVx4_ASAP7_75t_L g604 ( 
.A(n_492),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_492),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_508),
.Y(n_606)
);

NOR3xp33_ASAP7_75t_L g607 ( 
.A(n_491),
.B(n_8),
.C(n_9),
.Y(n_607)
);

AND2x6_ASAP7_75t_L g608 ( 
.A(n_485),
.B(n_29),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_478),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_508),
.Y(n_610)
);

AND2x2_ASAP7_75t_SL g611 ( 
.A(n_501),
.B(n_9),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_505),
.B(n_10),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_520),
.B(n_10),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_550),
.Y(n_614)
);

NAND2x1p5_ASAP7_75t_L g615 ( 
.A(n_520),
.B(n_30),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_493),
.B(n_11),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_492),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_498),
.B(n_31),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_498),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_538),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_498),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_535),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_546),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_497),
.B(n_11),
.Y(n_624)
);

NAND2x1p5_ASAP7_75t_L g625 ( 
.A(n_560),
.B(n_32),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_513),
.B(n_536),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_534),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_535),
.Y(n_628)
);

AO22x2_ASAP7_75t_L g629 ( 
.A1(n_553),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_570),
.A2(n_497),
.B(n_532),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_627),
.B(n_509),
.Y(n_631)
);

NOR3xp33_ASAP7_75t_L g632 ( 
.A(n_564),
.B(n_517),
.C(n_545),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_614),
.B(n_510),
.Y(n_633)
);

OAI21xp5_ASAP7_75t_L g634 ( 
.A1(n_628),
.A2(n_601),
.B(n_599),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_601),
.B(n_485),
.Y(n_635)
);

O2A1O1Ixp5_ASAP7_75t_L g636 ( 
.A1(n_592),
.A2(n_612),
.B(n_624),
.C(n_577),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_582),
.A2(n_532),
.B(n_528),
.Y(n_637)
);

INVx11_ASAP7_75t_L g638 ( 
.A(n_595),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_563),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_583),
.A2(n_532),
.B(n_528),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_594),
.A2(n_534),
.B(n_558),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_623),
.B(n_560),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_581),
.B(n_524),
.Y(n_643)
);

AND2x2_ASAP7_75t_SL g644 ( 
.A(n_611),
.B(n_607),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_L g645 ( 
.A1(n_628),
.A2(n_495),
.B(n_516),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_606),
.B(n_525),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_598),
.A2(n_610),
.B(n_622),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_616),
.B(n_490),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_578),
.A2(n_555),
.B(n_514),
.Y(n_649)
);

AOI21x1_ASAP7_75t_L g650 ( 
.A1(n_620),
.A2(n_527),
.B(n_540),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_578),
.A2(n_544),
.B(n_484),
.Y(n_651)
);

OAI22xp5_ASAP7_75t_L g652 ( 
.A1(n_590),
.A2(n_542),
.B1(n_490),
.B2(n_515),
.Y(n_652)
);

INVxp67_ASAP7_75t_L g653 ( 
.A(n_591),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_605),
.A2(n_544),
.B(n_526),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_617),
.A2(n_526),
.B(n_521),
.Y(n_655)
);

AOI21x1_ASAP7_75t_L g656 ( 
.A1(n_619),
.A2(n_527),
.B(n_540),
.Y(n_656)
);

AOI21xp33_ASAP7_75t_L g657 ( 
.A1(n_602),
.A2(n_542),
.B(n_519),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_561),
.B(n_515),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_586),
.B(n_545),
.Y(n_659)
);

OAI21xp5_ASAP7_75t_L g660 ( 
.A1(n_579),
.A2(n_552),
.B(n_527),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_604),
.A2(n_521),
.B(n_519),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_604),
.A2(n_540),
.B(n_551),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_618),
.A2(n_540),
.B(n_552),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_L g664 ( 
.A1(n_618),
.A2(n_543),
.B(n_556),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_588),
.B(n_549),
.Y(n_665)
);

OAI21xp5_ASAP7_75t_L g666 ( 
.A1(n_573),
.A2(n_566),
.B(n_562),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_567),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_575),
.A2(n_512),
.B1(n_547),
.B2(n_541),
.Y(n_668)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_585),
.A2(n_547),
.B1(n_556),
.B2(n_527),
.Y(n_669)
);

OAI21x1_ASAP7_75t_L g670 ( 
.A1(n_568),
.A2(n_34),
.B(n_33),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_626),
.B(n_12),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_621),
.B(n_14),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_587),
.B(n_15),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_571),
.A2(n_36),
.B(n_35),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_571),
.A2(n_39),
.B(n_38),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_569),
.Y(n_676)
);

OAI321xp33_ASAP7_75t_L g677 ( 
.A1(n_600),
.A2(n_15),
.A3(n_16),
.B1(n_17),
.B2(n_18),
.C(n_19),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g678 ( 
.A1(n_576),
.A2(n_129),
.B(n_220),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_586),
.B(n_518),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_574),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_629),
.A2(n_589),
.B1(n_603),
.B2(n_596),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_603),
.B(n_626),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_593),
.A2(n_127),
.B(n_218),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_597),
.B(n_19),
.Y(n_684)
);

BUFx12f_ASAP7_75t_L g685 ( 
.A(n_595),
.Y(n_685)
);

OAI22xp5_ASAP7_75t_L g686 ( 
.A1(n_629),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_613),
.B(n_40),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_572),
.Y(n_688)
);

OAI21xp5_ASAP7_75t_L g689 ( 
.A1(n_565),
.A2(n_130),
.B(n_216),
.Y(n_689)
);

AO21x1_ASAP7_75t_L g690 ( 
.A1(n_615),
.A2(n_21),
.B(n_22),
.Y(n_690)
);

INVxp67_ASAP7_75t_L g691 ( 
.A(n_609),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_665),
.B(n_580),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_648),
.B(n_608),
.Y(n_693)
);

OAI21xp33_ASAP7_75t_L g694 ( 
.A1(n_631),
.A2(n_584),
.B(n_625),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_658),
.B(n_608),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_644),
.B(n_574),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_646),
.B(n_608),
.Y(n_697)
);

BUFx12f_ASAP7_75t_L g698 ( 
.A(n_685),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_682),
.B(n_574),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_645),
.A2(n_565),
.B(n_574),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_680),
.Y(n_701)
);

O2A1O1Ixp33_ASAP7_75t_L g702 ( 
.A1(n_686),
.A2(n_608),
.B(n_24),
.C(n_565),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_632),
.B(n_565),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_R g704 ( 
.A(n_680),
.B(n_691),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_639),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_676),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_671),
.B(n_24),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_651),
.A2(n_43),
.B1(n_45),
.B2(n_47),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_664),
.B(n_48),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_635),
.B(n_49),
.Y(n_710)
);

OAI21xp5_ASAP7_75t_L g711 ( 
.A1(n_636),
.A2(n_51),
.B(n_53),
.Y(n_711)
);

O2A1O1Ixp33_ASAP7_75t_L g712 ( 
.A1(n_686),
.A2(n_55),
.B(n_56),
.C(n_60),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_659),
.Y(n_713)
);

A2O1A1Ixp33_ASAP7_75t_L g714 ( 
.A1(n_649),
.A2(n_61),
.B(n_63),
.C(n_64),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_688),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_667),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_643),
.Y(n_717)
);

INVxp67_ASAP7_75t_L g718 ( 
.A(n_633),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_653),
.B(n_65),
.Y(n_719)
);

OAI22xp5_ASAP7_75t_L g720 ( 
.A1(n_635),
.A2(n_66),
.B1(n_69),
.B2(n_71),
.Y(n_720)
);

BUFx4_ASAP7_75t_SL g721 ( 
.A(n_638),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_668),
.Y(n_722)
);

NAND3xp33_ASAP7_75t_SL g723 ( 
.A(n_690),
.B(n_219),
.C(n_73),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_652),
.B(n_72),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_L g725 ( 
.A1(n_641),
.A2(n_75),
.B(n_76),
.Y(n_725)
);

O2A1O1Ixp33_ASAP7_75t_L g726 ( 
.A1(n_681),
.A2(n_79),
.B(n_80),
.C(n_82),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_634),
.Y(n_727)
);

OAI22x1_ASAP7_75t_L g728 ( 
.A1(n_687),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_728)
);

AOI21x1_ASAP7_75t_L g729 ( 
.A1(n_630),
.A2(n_87),
.B(n_88),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_652),
.B(n_89),
.Y(n_730)
);

NAND3xp33_ASAP7_75t_L g731 ( 
.A(n_666),
.B(n_90),
.C(n_91),
.Y(n_731)
);

AOI21xp5_ASAP7_75t_L g732 ( 
.A1(n_663),
.A2(n_93),
.B(n_94),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_657),
.B(n_95),
.Y(n_733)
);

AO31x2_ASAP7_75t_L g734 ( 
.A1(n_647),
.A2(n_96),
.A3(n_98),
.B(n_99),
.Y(n_734)
);

OR2x6_ASAP7_75t_L g735 ( 
.A(n_662),
.B(n_100),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_681),
.B(n_668),
.Y(n_736)
);

BUFx2_ASAP7_75t_L g737 ( 
.A(n_672),
.Y(n_737)
);

O2A1O1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_677),
.A2(n_101),
.B(n_103),
.C(n_105),
.Y(n_738)
);

BUFx2_ASAP7_75t_L g739 ( 
.A(n_673),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_684),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_657),
.B(n_106),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_660),
.A2(n_110),
.B(n_111),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_669),
.B(n_112),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_661),
.B(n_114),
.Y(n_744)
);

A2O1A1Ixp33_ASAP7_75t_L g745 ( 
.A1(n_689),
.A2(n_116),
.B(n_118),
.C(n_119),
.Y(n_745)
);

BUFx3_ASAP7_75t_L g746 ( 
.A(n_670),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_637),
.A2(n_121),
.B(n_123),
.Y(n_747)
);

OAI22xp5_ASAP7_75t_L g748 ( 
.A1(n_654),
.A2(n_125),
.B1(n_126),
.B2(n_131),
.Y(n_748)
);

A2O1A1Ixp33_ASAP7_75t_L g749 ( 
.A1(n_674),
.A2(n_133),
.B(n_134),
.C(n_135),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_705),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_706),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_692),
.B(n_679),
.Y(n_752)
);

BUFx12f_ASAP7_75t_L g753 ( 
.A(n_698),
.Y(n_753)
);

BUFx4f_ASAP7_75t_SL g754 ( 
.A(n_717),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_717),
.Y(n_755)
);

CKINVDCx20_ASAP7_75t_R g756 ( 
.A(n_704),
.Y(n_756)
);

BUFx12f_ASAP7_75t_L g757 ( 
.A(n_717),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_716),
.Y(n_758)
);

BUFx12f_ASAP7_75t_L g759 ( 
.A(n_713),
.Y(n_759)
);

CKINVDCx20_ASAP7_75t_R g760 ( 
.A(n_722),
.Y(n_760)
);

CKINVDCx11_ASAP7_75t_R g761 ( 
.A(n_721),
.Y(n_761)
);

OR2x2_ASAP7_75t_L g762 ( 
.A(n_718),
.B(n_642),
.Y(n_762)
);

NAND2x1p5_ASAP7_75t_L g763 ( 
.A(n_699),
.B(n_650),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_736),
.A2(n_675),
.B1(n_678),
.B2(n_683),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_715),
.Y(n_765)
);

OR2x2_ASAP7_75t_L g766 ( 
.A(n_739),
.B(n_655),
.Y(n_766)
);

BUFx10_ASAP7_75t_L g767 ( 
.A(n_713),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_713),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_699),
.Y(n_769)
);

INVx5_ASAP7_75t_L g770 ( 
.A(n_735),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_719),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_701),
.Y(n_772)
);

BUFx2_ASAP7_75t_L g773 ( 
.A(n_696),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_707),
.B(n_737),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_740),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_695),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_701),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_703),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_724),
.B(n_137),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_727),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_727),
.Y(n_781)
);

BUFx3_ASAP7_75t_L g782 ( 
.A(n_735),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_728),
.Y(n_783)
);

CKINVDCx20_ASAP7_75t_R g784 ( 
.A(n_693),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_697),
.Y(n_785)
);

BUFx2_ASAP7_75t_L g786 ( 
.A(n_743),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_730),
.Y(n_787)
);

INVx8_ASAP7_75t_L g788 ( 
.A(n_694),
.Y(n_788)
);

INVx1_ASAP7_75t_SL g789 ( 
.A(n_710),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_733),
.B(n_640),
.Y(n_790)
);

INVx1_ASAP7_75t_SL g791 ( 
.A(n_741),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_734),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_729),
.Y(n_793)
);

INVx1_ASAP7_75t_SL g794 ( 
.A(n_744),
.Y(n_794)
);

INVx5_ASAP7_75t_SL g795 ( 
.A(n_726),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_746),
.Y(n_796)
);

BUFx3_ASAP7_75t_L g797 ( 
.A(n_734),
.Y(n_797)
);

INVx1_ASAP7_75t_SL g798 ( 
.A(n_709),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_734),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_723),
.Y(n_800)
);

INVx6_ASAP7_75t_L g801 ( 
.A(n_702),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_708),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_738),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_731),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_711),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_714),
.Y(n_806)
);

NAND2x1p5_ASAP7_75t_L g807 ( 
.A(n_732),
.B(n_656),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_748),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_720),
.Y(n_809)
);

OR2x2_ASAP7_75t_L g810 ( 
.A(n_700),
.B(n_138),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_747),
.Y(n_811)
);

BUFx4_ASAP7_75t_SL g812 ( 
.A(n_712),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_749),
.Y(n_813)
);

BUFx12f_ASAP7_75t_L g814 ( 
.A(n_745),
.Y(n_814)
);

INVx6_ASAP7_75t_L g815 ( 
.A(n_742),
.Y(n_815)
);

A2O1A1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_805),
.A2(n_725),
.B(n_142),
.C(n_143),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_750),
.Y(n_817)
);

AND2x4_ASAP7_75t_L g818 ( 
.A(n_782),
.B(n_140),
.Y(n_818)
);

O2A1O1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_805),
.A2(n_146),
.B(n_147),
.C(n_148),
.Y(n_819)
);

AO31x2_ASAP7_75t_L g820 ( 
.A1(n_799),
.A2(n_149),
.A3(n_153),
.B(n_154),
.Y(n_820)
);

CKINVDCx9p33_ASAP7_75t_R g821 ( 
.A(n_773),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_781),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_757),
.Y(n_823)
);

AO21x2_ASAP7_75t_L g824 ( 
.A1(n_792),
.A2(n_157),
.B(n_158),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_780),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_801),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_791),
.B(n_163),
.Y(n_827)
);

OAI21x1_ASAP7_75t_L g828 ( 
.A1(n_807),
.A2(n_164),
.B(n_165),
.Y(n_828)
);

OAI21x1_ASAP7_75t_L g829 ( 
.A1(n_807),
.A2(n_166),
.B(n_167),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_751),
.Y(n_830)
);

INVx1_ASAP7_75t_SL g831 ( 
.A(n_774),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_758),
.Y(n_832)
);

OAI21x1_ASAP7_75t_L g833 ( 
.A1(n_811),
.A2(n_168),
.B(n_169),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_778),
.B(n_175),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_765),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_SL g836 ( 
.A1(n_787),
.A2(n_176),
.B(n_177),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_772),
.Y(n_837)
);

OAI21xp5_ASAP7_75t_L g838 ( 
.A1(n_803),
.A2(n_178),
.B(n_179),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_775),
.Y(n_839)
);

OA21x2_ASAP7_75t_L g840 ( 
.A1(n_793),
.A2(n_181),
.B(n_182),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_772),
.Y(n_841)
);

A2O1A1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_779),
.A2(n_184),
.B(n_185),
.C(n_186),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_772),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_801),
.A2(n_187),
.B1(n_189),
.B2(n_191),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_777),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_766),
.Y(n_846)
);

OR2x2_ASAP7_75t_L g847 ( 
.A(n_791),
.B(n_192),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_777),
.Y(n_848)
);

OA21x2_ASAP7_75t_L g849 ( 
.A1(n_790),
.A2(n_194),
.B(n_195),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_794),
.A2(n_196),
.B(n_199),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_796),
.Y(n_851)
);

OAI21x1_ASAP7_75t_L g852 ( 
.A1(n_764),
.A2(n_200),
.B(n_201),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_771),
.Y(n_853)
);

AND2x4_ASAP7_75t_L g854 ( 
.A(n_755),
.B(n_203),
.Y(n_854)
);

AND2x4_ASAP7_75t_L g855 ( 
.A(n_769),
.B(n_205),
.Y(n_855)
);

A2O1A1Ixp33_ASAP7_75t_L g856 ( 
.A1(n_770),
.A2(n_208),
.B(n_210),
.C(n_211),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_789),
.B(n_794),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_796),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_754),
.Y(n_859)
);

NOR2x1_ASAP7_75t_R g860 ( 
.A(n_761),
.B(n_212),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_797),
.Y(n_861)
);

AOI222xp33_ASAP7_75t_L g862 ( 
.A1(n_809),
.A2(n_213),
.B1(n_214),
.B2(n_814),
.C1(n_801),
.C2(n_786),
.Y(n_862)
);

OAI21x1_ASAP7_75t_L g863 ( 
.A1(n_764),
.A2(n_790),
.B(n_763),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_776),
.B(n_785),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_783),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_770),
.A2(n_789),
.B(n_798),
.Y(n_866)
);

OAI21xp5_ASAP7_75t_L g867 ( 
.A1(n_808),
.A2(n_798),
.B(n_810),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_762),
.Y(n_868)
);

OAI21x1_ASAP7_75t_L g869 ( 
.A1(n_763),
.A2(n_815),
.B(n_770),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_800),
.B(n_770),
.Y(n_870)
);

OA21x2_ASAP7_75t_L g871 ( 
.A1(n_815),
.A2(n_795),
.B(n_800),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_754),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_752),
.B(n_784),
.Y(n_873)
);

CKINVDCx6p67_ASAP7_75t_R g874 ( 
.A(n_761),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_822),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_817),
.B(n_769),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_846),
.B(n_769),
.Y(n_877)
);

BUFx2_ASAP7_75t_L g878 ( 
.A(n_861),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_830),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_832),
.Y(n_880)
);

OA21x2_ASAP7_75t_L g881 ( 
.A1(n_863),
.A2(n_815),
.B(n_812),
.Y(n_881)
);

INVx2_ASAP7_75t_SL g882 ( 
.A(n_839),
.Y(n_882)
);

OAI21x1_ASAP7_75t_L g883 ( 
.A1(n_869),
.A2(n_852),
.B(n_828),
.Y(n_883)
);

CKINVDCx11_ASAP7_75t_R g884 ( 
.A(n_874),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_825),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_835),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_857),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_862),
.A2(n_802),
.B1(n_806),
.B2(n_800),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_857),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_849),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_851),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_849),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_849),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_871),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_858),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_820),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_871),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_868),
.Y(n_898)
);

AOI21x1_ASAP7_75t_L g899 ( 
.A1(n_870),
.A2(n_812),
.B(n_795),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_820),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_845),
.Y(n_901)
);

HB1xp67_ASAP7_75t_SL g902 ( 
.A(n_823),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_848),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_820),
.Y(n_904)
);

NAND2x1p5_ASAP7_75t_L g905 ( 
.A(n_870),
.B(n_804),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_865),
.B(n_804),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_853),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_824),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_831),
.B(n_867),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_840),
.Y(n_910)
);

AO21x2_ASAP7_75t_L g911 ( 
.A1(n_866),
.A2(n_795),
.B(n_804),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_853),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_824),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_833),
.Y(n_914)
);

OAI21x1_ASAP7_75t_L g915 ( 
.A1(n_829),
.A2(n_788),
.B(n_806),
.Y(n_915)
);

INVx4_ASAP7_75t_L g916 ( 
.A(n_853),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_853),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_875),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_875),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_875),
.B(n_873),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_SL g921 ( 
.A1(n_888),
.A2(n_862),
.B(n_838),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_884),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_887),
.B(n_867),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_898),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_878),
.Y(n_925)
);

AOI222xp33_ASAP7_75t_L g926 ( 
.A1(n_909),
.A2(n_838),
.B1(n_860),
.B2(n_826),
.C1(n_844),
.C2(n_842),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_885),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_909),
.B(n_866),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_879),
.B(n_841),
.Y(n_929)
);

HB1xp67_ASAP7_75t_L g930 ( 
.A(n_878),
.Y(n_930)
);

INVx3_ASAP7_75t_L g931 ( 
.A(n_894),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_R g932 ( 
.A(n_902),
.B(n_756),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_879),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_880),
.B(n_864),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_R g935 ( 
.A(n_899),
.B(n_760),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_880),
.B(n_843),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_906),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_894),
.Y(n_938)
);

OAI22xp33_ASAP7_75t_SL g939 ( 
.A1(n_905),
.A2(n_827),
.B1(n_847),
.B2(n_850),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_886),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_899),
.A2(n_850),
.B(n_856),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_889),
.B(n_843),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_894),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_886),
.Y(n_944)
);

BUFx2_ASAP7_75t_L g945 ( 
.A(n_897),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_891),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_905),
.B(n_827),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_889),
.B(n_837),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_891),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_918),
.Y(n_950)
);

OR2x6_ASAP7_75t_L g951 ( 
.A(n_941),
.B(n_905),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_945),
.B(n_897),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_933),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_933),
.Y(n_954)
);

NOR2x1p5_ASAP7_75t_L g955 ( 
.A(n_922),
.B(n_753),
.Y(n_955)
);

INVxp67_ASAP7_75t_SL g956 ( 
.A(n_925),
.Y(n_956)
);

OA21x2_ASAP7_75t_L g957 ( 
.A1(n_945),
.A2(n_892),
.B(n_893),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_940),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_931),
.B(n_897),
.Y(n_959)
);

OR2x2_ASAP7_75t_L g960 ( 
.A(n_928),
.B(n_900),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_940),
.Y(n_961)
);

HB1xp67_ASAP7_75t_L g962 ( 
.A(n_918),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_944),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_919),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_919),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_944),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_931),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_946),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_946),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_927),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_949),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_920),
.B(n_882),
.Y(n_972)
);

AND2x4_ASAP7_75t_SL g973 ( 
.A(n_924),
.B(n_894),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_953),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_954),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_957),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_957),
.Y(n_977)
);

INVxp67_ASAP7_75t_L g978 ( 
.A(n_951),
.Y(n_978)
);

AOI21x1_ASAP7_75t_L g979 ( 
.A1(n_959),
.A2(n_947),
.B(n_930),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_960),
.B(n_923),
.Y(n_980)
);

BUFx2_ASAP7_75t_L g981 ( 
.A(n_956),
.Y(n_981)
);

AOI22xp33_ASAP7_75t_L g982 ( 
.A1(n_951),
.A2(n_926),
.B1(n_939),
.B2(n_921),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_968),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_969),
.Y(n_984)
);

A2O1A1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_973),
.A2(n_921),
.B(n_819),
.C(n_856),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_957),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_951),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_959),
.B(n_920),
.Y(n_988)
);

BUFx2_ASAP7_75t_L g989 ( 
.A(n_952),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_952),
.B(n_934),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_976),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_989),
.B(n_934),
.Y(n_992)
);

BUFx2_ASAP7_75t_L g993 ( 
.A(n_981),
.Y(n_993)
);

OR2x2_ASAP7_75t_L g994 ( 
.A(n_980),
.B(n_972),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_974),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_975),
.Y(n_996)
);

OAI321xp33_ASAP7_75t_L g997 ( 
.A1(n_982),
.A2(n_826),
.A3(n_844),
.B1(n_894),
.B2(n_819),
.C(n_906),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_976),
.Y(n_998)
);

OR2x2_ASAP7_75t_L g999 ( 
.A(n_978),
.B(n_971),
.Y(n_999)
);

HB1xp67_ASAP7_75t_L g1000 ( 
.A(n_983),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_984),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_978),
.B(n_967),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_993),
.B(n_987),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_1000),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_1002),
.B(n_987),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_1002),
.B(n_987),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_992),
.B(n_987),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_994),
.B(n_990),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_995),
.B(n_982),
.Y(n_1009)
);

INVxp67_ASAP7_75t_SL g1010 ( 
.A(n_991),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_1003),
.B(n_955),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_1004),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_1007),
.B(n_996),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_1005),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_1009),
.B(n_1001),
.Y(n_1015)
);

HB1xp67_ASAP7_75t_L g1016 ( 
.A(n_1005),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_1010),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_SL g1018 ( 
.A(n_1011),
.B(n_922),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_1017),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_1016),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_1012),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_1014),
.Y(n_1022)
);

INVx1_ASAP7_75t_SL g1023 ( 
.A(n_1013),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1015),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_1015),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_1011),
.B(n_1005),
.Y(n_1026)
);

HB1xp67_ASAP7_75t_L g1027 ( 
.A(n_1016),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_1011),
.B(n_1006),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_1026),
.B(n_1006),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_1027),
.B(n_1000),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_1028),
.B(n_1006),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_1018),
.B(n_1008),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1027),
.Y(n_1033)
);

BUFx2_ASAP7_75t_L g1034 ( 
.A(n_1020),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1022),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1019),
.Y(n_1036)
);

OR2x2_ASAP7_75t_L g1037 ( 
.A(n_1023),
.B(n_999),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1034),
.B(n_1025),
.Y(n_1038)
);

OAI21xp33_ASAP7_75t_SL g1039 ( 
.A1(n_1032),
.A2(n_1025),
.B(n_1010),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1033),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_1029),
.B(n_1024),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_1031),
.B(n_1021),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_1030),
.A2(n_997),
.B(n_985),
.C(n_998),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1030),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_1037),
.B(n_991),
.Y(n_1045)
);

XNOR2xp5_ASAP7_75t_L g1046 ( 
.A(n_1035),
.B(n_939),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_1042),
.B(n_1036),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_1041),
.B(n_988),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_1045),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1038),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_1040),
.B(n_998),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_1044),
.B(n_979),
.Y(n_1052)
);

OR2x2_ASAP7_75t_L g1053 ( 
.A(n_1043),
.B(n_986),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1039),
.B(n_958),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1049),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_1048),
.B(n_1046),
.Y(n_1056)
);

NAND2xp33_ASAP7_75t_L g1057 ( 
.A(n_1053),
.B(n_932),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_1050),
.B(n_937),
.Y(n_1058)
);

INVxp67_ASAP7_75t_L g1059 ( 
.A(n_1051),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1047),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_1054),
.B(n_977),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_1052),
.B(n_977),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1048),
.B(n_986),
.Y(n_1063)
);

NOR3xp33_ASAP7_75t_L g1064 ( 
.A(n_1055),
.B(n_985),
.C(n_818),
.Y(n_1064)
);

NAND4xp75_ASAP7_75t_L g1065 ( 
.A(n_1060),
.B(n_859),
.C(n_872),
.D(n_834),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_1059),
.B(n_1057),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_1058),
.B(n_823),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1056),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1061),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_1063),
.B(n_823),
.Y(n_1070)
);

NAND4xp25_ASAP7_75t_L g1071 ( 
.A(n_1062),
.B(n_818),
.C(n_842),
.D(n_836),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_1059),
.B(n_823),
.Y(n_1072)
);

AOI221xp5_ASAP7_75t_L g1073 ( 
.A1(n_1072),
.A2(n_816),
.B1(n_935),
.B2(n_768),
.C(n_967),
.Y(n_1073)
);

AOI21xp33_ASAP7_75t_L g1074 ( 
.A1(n_1068),
.A2(n_759),
.B(n_854),
.Y(n_1074)
);

NAND3xp33_ASAP7_75t_SL g1075 ( 
.A(n_1066),
.B(n_816),
.C(n_937),
.Y(n_1075)
);

NAND4xp75_ASAP7_75t_L g1076 ( 
.A(n_1069),
.B(n_881),
.C(n_948),
.D(n_942),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1070),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_1064),
.A2(n_894),
.B1(n_938),
.B2(n_931),
.Y(n_1078)
);

AOI21xp33_ASAP7_75t_SL g1079 ( 
.A1(n_1067),
.A2(n_855),
.B(n_854),
.Y(n_1079)
);

CKINVDCx20_ASAP7_75t_R g1080 ( 
.A(n_1077),
.Y(n_1080)
);

INVx1_ASAP7_75t_SL g1081 ( 
.A(n_1074),
.Y(n_1081)
);

O2A1O1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_1075),
.A2(n_1071),
.B(n_1065),
.C(n_855),
.Y(n_1082)
);

OAI21xp33_ASAP7_75t_L g1083 ( 
.A1(n_1078),
.A2(n_973),
.B(n_967),
.Y(n_1083)
);

AOI221xp5_ASAP7_75t_L g1084 ( 
.A1(n_1079),
.A2(n_1073),
.B1(n_1076),
.B2(n_938),
.C(n_943),
.Y(n_1084)
);

INVx2_ASAP7_75t_SL g1085 ( 
.A(n_1077),
.Y(n_1085)
);

AND5x1_ASAP7_75t_L g1086 ( 
.A(n_1073),
.B(n_821),
.C(n_767),
.D(n_938),
.E(n_943),
.Y(n_1086)
);

OAI221xp5_ASAP7_75t_SL g1087 ( 
.A1(n_1077),
.A2(n_943),
.B1(n_913),
.B2(n_908),
.C(n_966),
.Y(n_1087)
);

NAND4xp25_ASAP7_75t_SL g1088 ( 
.A(n_1077),
.B(n_963),
.C(n_961),
.D(n_942),
.Y(n_1088)
);

OAI22xp33_ASAP7_75t_SL g1089 ( 
.A1(n_1085),
.A2(n_913),
.B1(n_908),
.B2(n_837),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1080),
.B(n_1081),
.Y(n_1090)
);

OAI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_1084),
.A2(n_771),
.B1(n_788),
.B2(n_962),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_1083),
.A2(n_771),
.B1(n_911),
.B2(n_917),
.Y(n_1092)
);

NOR2x1_ASAP7_75t_L g1093 ( 
.A(n_1082),
.B(n_1088),
.Y(n_1093)
);

NOR2x1_ASAP7_75t_L g1094 ( 
.A(n_1086),
.B(n_911),
.Y(n_1094)
);

NAND2xp33_ASAP7_75t_L g1095 ( 
.A(n_1087),
.B(n_962),
.Y(n_1095)
);

XNOR2xp5_ASAP7_75t_L g1096 ( 
.A(n_1080),
.B(n_911),
.Y(n_1096)
);

NOR2x1_ASAP7_75t_L g1097 ( 
.A(n_1080),
.B(n_916),
.Y(n_1097)
);

AOI311xp33_ASAP7_75t_L g1098 ( 
.A1(n_1084),
.A2(n_895),
.A3(n_904),
.B(n_896),
.C(n_900),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1090),
.Y(n_1099)
);

NAND3xp33_ASAP7_75t_L g1100 ( 
.A(n_1093),
.B(n_1097),
.C(n_1096),
.Y(n_1100)
);

NOR2xp67_ASAP7_75t_L g1101 ( 
.A(n_1092),
.B(n_965),
.Y(n_1101)
);

OAI211xp5_ASAP7_75t_L g1102 ( 
.A1(n_1094),
.A2(n_788),
.B(n_965),
.C(n_916),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1091),
.A2(n_895),
.B(n_901),
.Y(n_1103)
);

NOR3xp33_ASAP7_75t_L g1104 ( 
.A(n_1095),
.B(n_916),
.C(n_913),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1089),
.Y(n_1105)
);

INVxp33_ASAP7_75t_L g1106 ( 
.A(n_1098),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_1097),
.B(n_948),
.Y(n_1107)
);

NOR2xp67_ASAP7_75t_L g1108 ( 
.A(n_1090),
.B(n_916),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_1097),
.Y(n_1109)
);

HB1xp67_ASAP7_75t_L g1110 ( 
.A(n_1097),
.Y(n_1110)
);

NOR2x1p5_ASAP7_75t_L g1111 ( 
.A(n_1090),
.B(n_912),
.Y(n_1111)
);

INVx1_ASAP7_75t_SL g1112 ( 
.A(n_1109),
.Y(n_1112)
);

INVx1_ASAP7_75t_SL g1113 ( 
.A(n_1110),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1099),
.A2(n_903),
.B(n_901),
.Y(n_1114)
);

BUFx2_ASAP7_75t_L g1115 ( 
.A(n_1111),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1100),
.Y(n_1116)
);

INVx3_ASAP7_75t_SL g1117 ( 
.A(n_1105),
.Y(n_1117)
);

BUFx2_ASAP7_75t_L g1118 ( 
.A(n_1107),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_1108),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1101),
.B(n_767),
.Y(n_1120)
);

OAI22x1_ASAP7_75t_L g1121 ( 
.A1(n_1117),
.A2(n_1112),
.B1(n_1113),
.B2(n_1118),
.Y(n_1121)
);

AO22x2_ASAP7_75t_L g1122 ( 
.A1(n_1116),
.A2(n_1104),
.B1(n_1102),
.B2(n_1106),
.Y(n_1122)
);

OA22x2_ASAP7_75t_L g1123 ( 
.A1(n_1119),
.A2(n_1103),
.B1(n_907),
.B2(n_964),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_1120),
.A2(n_907),
.B1(n_917),
.B2(n_950),
.Y(n_1124)
);

XOR2x2_ASAP7_75t_L g1125 ( 
.A(n_1115),
.B(n_881),
.Y(n_1125)
);

AO22x2_ASAP7_75t_L g1126 ( 
.A1(n_1114),
.A2(n_917),
.B1(n_964),
.B2(n_950),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1118),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1112),
.A2(n_912),
.B1(n_936),
.B2(n_970),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1121),
.Y(n_1129)
);

NOR2x1_ASAP7_75t_L g1130 ( 
.A(n_1127),
.B(n_908),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1122),
.A2(n_913),
.B(n_908),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1129),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1132),
.A2(n_1125),
.B1(n_1123),
.B2(n_1131),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1133),
.Y(n_1134)
);

AOI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_1134),
.A2(n_1130),
.B1(n_1126),
.B2(n_1124),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1134),
.A2(n_1128),
.B1(n_970),
.B2(n_912),
.Y(n_1136)
);

AOI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1134),
.A2(n_936),
.B1(n_912),
.B2(n_929),
.Y(n_1137)
);

XNOR2xp5_ASAP7_75t_SL g1138 ( 
.A(n_1135),
.B(n_821),
.Y(n_1138)
);

AOI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1136),
.A2(n_912),
.B1(n_929),
.B2(n_881),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_R g1140 ( 
.A1(n_1137),
.A2(n_949),
.B1(n_882),
.B2(n_910),
.Y(n_1140)
);

XNOR2xp5_ASAP7_75t_L g1141 ( 
.A(n_1138),
.B(n_915),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1139),
.A2(n_912),
.B1(n_903),
.B2(n_892),
.Y(n_1142)
);

AOI22xp5_ASAP7_75t_SL g1143 ( 
.A1(n_1140),
.A2(n_910),
.B1(n_876),
.B2(n_881),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1141),
.A2(n_915),
.B(n_876),
.Y(n_1144)
);

AO21x2_ASAP7_75t_L g1145 ( 
.A1(n_1143),
.A2(n_890),
.B(n_893),
.Y(n_1145)
);

OAI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1142),
.A2(n_883),
.B(n_914),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1144),
.A2(n_914),
.B(n_877),
.Y(n_1147)
);

AOI211xp5_ASAP7_75t_L g1148 ( 
.A1(n_1147),
.A2(n_1146),
.B(n_1145),
.C(n_813),
.Y(n_1148)
);


endmodule