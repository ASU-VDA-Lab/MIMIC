module real_jpeg_16641_n_32 (n_17, n_199, n_8, n_0, n_21, n_2, n_188, n_29, n_196, n_191, n_10, n_31, n_9, n_201, n_12, n_24, n_189, n_6, n_190, n_28, n_194, n_192, n_198, n_23, n_11, n_14, n_25, n_195, n_7, n_22, n_18, n_3, n_193, n_197, n_5, n_4, n_1, n_26, n_27, n_20, n_19, n_200, n_30, n_16, n_15, n_13, n_32);

input n_17;
input n_199;
input n_8;
input n_0;
input n_21;
input n_2;
input n_188;
input n_29;
input n_196;
input n_191;
input n_10;
input n_31;
input n_9;
input n_201;
input n_12;
input n_24;
input n_189;
input n_6;
input n_190;
input n_28;
input n_194;
input n_192;
input n_198;
input n_23;
input n_11;
input n_14;
input n_25;
input n_195;
input n_7;
input n_22;
input n_18;
input n_3;
input n_193;
input n_197;
input n_5;
input n_4;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_200;
input n_30;
input n_16;
input n_15;
input n_13;

output n_32;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_150;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

AOI21x1_ASAP7_75t_L g110 ( 
.A1(n_0),
.A2(n_111),
.B(n_122),
.Y(n_110)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_0),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_1),
.B(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_1),
.Y(n_146)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_2),
.Y(n_104)
);

AOI322xp5_ASAP7_75t_SL g141 ( 
.A1(n_2),
.A2(n_93),
.A3(n_103),
.B1(n_106),
.B2(n_142),
.C1(n_144),
.C2(n_199),
.Y(n_141)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_3),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_SL g123 ( 
.A(n_3),
.B(n_113),
.C(n_119),
.Y(n_123)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_4),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_5),
.Y(n_149)
);

MAJx2_ASAP7_75t_L g108 ( 
.A(n_6),
.B(n_109),
.C(n_136),
.Y(n_108)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_7),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_7),
.B(n_96),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_8),
.Y(n_68)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_9),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_10),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_11),
.B(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_11),
.Y(n_160)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_12),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_12),
.B(n_82),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_13),
.B(n_47),
.C(n_172),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_15),
.Y(n_177)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_16),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_17),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_18),
.B(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_18),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_19),
.Y(n_184)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_21),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_22),
.A2(n_34),
.B1(n_35),
.B2(n_42),
.Y(n_33)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_22),
.A2(n_45),
.B1(n_178),
.B2(n_180),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_22),
.B(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_23),
.B(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_23),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_24),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_24),
.B(n_60),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_25),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_26),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_26),
.B(n_89),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_27),
.B(n_49),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_28),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_29),
.Y(n_61)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_31),
.B(n_114),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_43),
.Y(n_32)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_37),
.B(n_168),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_37),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_37),
.B(n_177),
.Y(n_176)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_38),
.Y(n_185)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_39),
.B(n_181),
.Y(n_180)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_40),
.B(n_107),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

BUFx4f_ASAP7_75t_SL g76 ( 
.A(n_41),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_42),
.A2(n_44),
.B1(n_182),
.B2(n_186),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_46),
.C(n_175),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_42),
.B(n_179),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_51),
.B(n_52),
.C(n_171),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_165),
.B(n_170),
.Y(n_52)
);

OAI31xp33_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_78),
.A3(n_147),
.B(n_151),
.Y(n_53)
);

NAND3xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_65),
.C(n_71),
.Y(n_54)
);

AOI321xp33_ASAP7_75t_L g151 ( 
.A1(n_55),
.A2(n_65),
.A3(n_152),
.B1(n_153),
.B2(n_156),
.C(n_200),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

OAI322xp33_ASAP7_75t_L g156 ( 
.A1(n_56),
.A2(n_66),
.A3(n_157),
.B1(n_162),
.B2(n_163),
.C1(n_164),
.C2(n_201),
.Y(n_156)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_57),
.Y(n_163)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_59),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_67),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_97),
.Y(n_96)
);

NAND3xp33_ASAP7_75t_L g157 ( 
.A(n_71),
.B(n_158),
.C(n_159),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_77),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_72),
.B(n_77),
.Y(n_152)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AOI31xp67_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_87),
.A3(n_108),
.B(n_138),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NOR3xp33_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_92),
.C(n_98),
.Y(n_87)
);

NOR3xp33_ASAP7_75t_L g142 ( 
.A(n_88),
.B(n_100),
.C(n_143),
.Y(n_142)
);

NOR2x1_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_91),
.B(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_91),
.B(n_137),
.Y(n_136)
);

OAI321xp33_ASAP7_75t_L g138 ( 
.A1(n_92),
.A2(n_98),
.A3(n_139),
.B1(n_140),
.B2(n_141),
.C(n_198),
.Y(n_138)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_130),
.C(n_131),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_117),
.C(n_118),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NOR2x1_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B(n_125),
.Y(n_122)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_129),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_169),
.Y(n_170)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_183),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_188),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_189),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_190),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_191),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_192),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_193),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_194),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_195),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_196),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_197),
.Y(n_137)
);


endmodule