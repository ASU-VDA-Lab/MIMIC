module fake_jpeg_8193_n_296 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_296);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_296;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_152;
wire n_73;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_33),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_0),
.Y(n_48)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_43),
.Y(n_51)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_27),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_23),
.B1(n_28),
.B2(n_29),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_47),
.A2(n_49),
.B1(n_61),
.B2(n_62),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_54),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_42),
.A2(n_23),
.B1(n_26),
.B2(n_24),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_23),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_52),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_28),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_53),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_21),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_58),
.Y(n_82)
);

INVxp33_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_44),
.B1(n_42),
.B2(n_26),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_44),
.A2(n_18),
.B1(n_28),
.B2(n_22),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_68),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_35),
.B1(n_26),
.B2(n_24),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_66),
.A2(n_69),
.B1(n_70),
.B2(n_21),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_0),
.Y(n_83)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_38),
.A2(n_35),
.B1(n_18),
.B2(n_17),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_38),
.A2(n_35),
.B1(n_18),
.B2(n_17),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_72),
.Y(n_110)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_80),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_62),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_75),
.B(n_81),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_57),
.A2(n_21),
.B1(n_31),
.B2(n_30),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_77),
.A2(n_90),
.B1(n_102),
.B2(n_107),
.Y(n_129)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_51),
.Y(n_81)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_85),
.A2(n_9),
.B1(n_16),
.B2(n_15),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_31),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_86),
.A2(n_88),
.B(n_34),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

BUFx24_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_31),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_46),
.B(n_34),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_94),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_46),
.A2(n_30),
.B1(n_33),
.B2(n_25),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

FAx1_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_33),
.CI(n_1),
.CON(n_93),
.SN(n_93)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_52),
.Y(n_128)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_53),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_97),
.Y(n_114)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_98),
.Y(n_122)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_100),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_54),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_104),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_58),
.A2(n_30),
.B1(n_33),
.B2(n_29),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_106),
.Y(n_125)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_56),
.A2(n_32),
.B1(n_20),
.B2(n_22),
.Y(n_107)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_94),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_76),
.A2(n_48),
.B(n_64),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_102),
.C(n_88),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_48),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_120),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_52),
.Y(n_120)
);

NOR3xp33_ASAP7_75t_SL g156 ( 
.A(n_123),
.B(n_107),
.C(n_15),
.Y(n_156)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_127),
.B(n_133),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_93),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_86),
.B(n_88),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_137),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_131),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_19),
.Y(n_132)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_85),
.A2(n_19),
.B1(n_32),
.B2(n_20),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_134),
.A2(n_137),
.B1(n_129),
.B2(n_133),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_136),
.A2(n_11),
.B1(n_12),
.B2(n_15),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_86),
.B(n_0),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_67),
.Y(n_138)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_SL g176 ( 
.A1(n_140),
.A2(n_156),
.B(n_165),
.Y(n_176)
);

AO22x1_ASAP7_75t_L g141 ( 
.A1(n_129),
.A2(n_93),
.B1(n_84),
.B2(n_90),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_141),
.B(n_142),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_142),
.A2(n_118),
.B(n_117),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_144),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_79),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_151),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_119),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_149),
.B(n_157),
.Y(n_188)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_150),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_109),
.C(n_92),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_154),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_87),
.Y(n_154)
);

INVx11_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_155),
.A2(n_126),
.B1(n_73),
.B2(n_122),
.Y(n_195)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_131),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_160),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_99),
.B1(n_108),
.B2(n_107),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_159),
.A2(n_161),
.B1(n_116),
.B2(n_118),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_127),
.B(n_103),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_135),
.A2(n_107),
.B1(n_78),
.B2(n_97),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_73),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_166),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_114),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_163),
.A2(n_113),
.B1(n_138),
.B2(n_117),
.Y(n_170)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_111),
.Y(n_166)
);

FAx1_ASAP7_75t_SL g167 ( 
.A(n_115),
.B(n_105),
.CI(n_54),
.CON(n_167),
.SN(n_167)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_168),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_132),
.B(n_92),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_114),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_125),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_170),
.A2(n_172),
.B1(n_174),
.B2(n_182),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_159),
.A2(n_135),
.B1(n_136),
.B2(n_120),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_147),
.A2(n_145),
.B1(n_141),
.B2(n_161),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_144),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_184),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_112),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_181),
.A2(n_196),
.B(n_198),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_140),
.A2(n_113),
.B1(n_123),
.B2(n_111),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_155),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_185),
.A2(n_190),
.B1(n_112),
.B2(n_124),
.Y(n_213)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_153),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_189),
.Y(n_214)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_139),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_141),
.A2(n_139),
.B1(n_142),
.B2(n_151),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_150),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_191),
.B(n_194),
.Y(n_211)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_192),
.Y(n_204)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_197),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_143),
.Y(n_194)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_195),
.Y(n_205)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_154),
.Y(n_197)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_208),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_148),
.C(n_164),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_206),
.C(n_209),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_188),
.B(n_146),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_216),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_178),
.Y(n_206)
);

MAJx2_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_167),
.C(n_164),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_207),
.B(n_213),
.Y(n_234)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_183),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_167),
.Y(n_209)
);

OA21x2_ASAP7_75t_L g210 ( 
.A1(n_193),
.A2(n_156),
.B(n_112),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_210),
.A2(n_217),
.B(n_212),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_171),
.B(n_124),
.C(n_125),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_197),
.C(n_186),
.Y(n_223)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_177),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_198),
.A2(n_112),
.B(n_1),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_217),
.A2(n_173),
.B(n_179),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_175),
.B(n_126),
.Y(n_218)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_218),
.Y(n_225)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_183),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_184),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_54),
.Y(n_221)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_221),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_230),
.C(n_232),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_224),
.A2(n_204),
.B(n_8),
.Y(n_255)
);

A2O1A1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_226),
.A2(n_210),
.B(n_214),
.C(n_202),
.Y(n_246)
);

AO22x1_ASAP7_75t_L g227 ( 
.A1(n_207),
.A2(n_176),
.B1(n_172),
.B2(n_182),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_238),
.Y(n_241)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_185),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_181),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_216),
.B(n_189),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_233),
.B(n_240),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_213),
.A2(n_181),
.B1(n_191),
.B2(n_194),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_236),
.A2(n_237),
.B1(n_205),
.B2(n_208),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_205),
.A2(n_180),
.B1(n_112),
.B2(n_121),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_214),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_98),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_219),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_200),
.B(n_91),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_220),
.Y(n_242)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_242),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_243),
.A2(n_246),
.B1(n_253),
.B2(n_238),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_199),
.Y(n_244)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_244),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_237),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_254),
.Y(n_259)
);

NOR3xp33_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_210),
.C(n_219),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_226),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_235),
.Y(n_251)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_251),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_234),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_236),
.A2(n_204),
.B1(n_211),
.B2(n_180),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_215),
.C(n_201),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_255),
.A2(n_9),
.B(n_13),
.Y(n_266)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_256),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_245),
.A2(n_239),
.B1(n_225),
.B2(n_234),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_258),
.A2(n_261),
.B1(n_249),
.B2(n_254),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_227),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_260),
.B(n_265),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_267),
.Y(n_277)
);

OAI21xp33_ASAP7_75t_L g265 ( 
.A1(n_241),
.A2(n_232),
.B(n_230),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_266),
.A2(n_246),
.B(n_241),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_222),
.Y(n_267)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_268),
.Y(n_278)
);

OAI221xp5_ASAP7_75t_L g269 ( 
.A1(n_259),
.A2(n_255),
.B1(n_253),
.B2(n_243),
.C(n_252),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_276),
.Y(n_279)
);

NAND3xp33_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_223),
.C(n_248),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_272),
.B(n_264),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_273),
.A2(n_266),
.B(n_7),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_8),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_275),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_262),
.B(n_8),
.Y(n_275)
);

OAI221xp5_ASAP7_75t_L g276 ( 
.A1(n_265),
.A2(n_13),
.B1(n_7),
.B2(n_9),
.C(n_4),
.Y(n_276)
);

INVxp67_ASAP7_75t_SL g280 ( 
.A(n_272),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_10),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_282),
.A2(n_270),
.B1(n_271),
.B2(n_277),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_267),
.C(n_263),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_283),
.A2(n_5),
.B(n_10),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_284),
.A2(n_5),
.B1(n_10),
.B2(n_13),
.Y(n_287)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_285),
.Y(n_290)
);

A2O1A1O1Ixp25_ASAP7_75t_L g286 ( 
.A1(n_279),
.A2(n_7),
.B(n_12),
.C(n_11),
.D(n_4),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_289),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_288),
.C(n_281),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_291),
.A2(n_278),
.B1(n_279),
.B2(n_289),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_293),
.B(n_294),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_290),
.A2(n_292),
.B(n_2),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_0),
.Y(n_296)
);


endmodule