module fake_aes_11803_n_38 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_10, n_8, n_0, n_38);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_10;
input n_8;
input n_0;
output n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_17;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
BUFx6f_ASAP7_75t_L g15 ( .A(n_13), .Y(n_15) );
NAND2xp5_ASAP7_75t_SL g16 ( .A(n_5), .B(n_14), .Y(n_16) );
INVxp67_ASAP7_75t_L g17 ( .A(n_6), .Y(n_17) );
AND2x2_ASAP7_75t_L g18 ( .A(n_4), .B(n_8), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_1), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_7), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_0), .Y(n_21) );
AND3x2_ASAP7_75t_SL g22 ( .A(n_20), .B(n_0), .C(n_1), .Y(n_22) );
AOI22xp5_ASAP7_75t_L g23 ( .A1(n_21), .A2(n_19), .B1(n_18), .B2(n_17), .Y(n_23) );
BUFx3_ASAP7_75t_L g24 ( .A(n_15), .Y(n_24) );
OAI21x1_ASAP7_75t_L g25 ( .A1(n_23), .A2(n_20), .B(n_16), .Y(n_25) );
OAI21x1_ASAP7_75t_L g26 ( .A1(n_23), .A2(n_16), .B(n_15), .Y(n_26) );
INVx2_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
AND2x4_ASAP7_75t_L g28 ( .A(n_27), .B(n_25), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_28), .B(n_25), .Y(n_29) );
AOI32xp33_ASAP7_75t_L g30 ( .A1(n_28), .A2(n_22), .A3(n_24), .B1(n_4), .B2(n_2), .Y(n_30) );
NAND2xp5_ASAP7_75t_L g31 ( .A(n_30), .B(n_28), .Y(n_31) );
AOI211xp5_ASAP7_75t_L g32 ( .A1(n_29), .A2(n_15), .B(n_3), .C(n_2), .Y(n_32) );
INVx2_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
AOI221xp5_ASAP7_75t_L g34 ( .A1(n_32), .A2(n_15), .B1(n_3), .B2(n_10), .C(n_11), .Y(n_34) );
AOI21xp33_ASAP7_75t_SL g35 ( .A1(n_33), .A2(n_9), .B(n_12), .Y(n_35) );
INVx1_ASAP7_75t_L g36 ( .A(n_34), .Y(n_36) );
INVx2_ASAP7_75t_L g37 ( .A(n_36), .Y(n_37) );
NOR2xp67_ASAP7_75t_L g38 ( .A(n_37), .B(n_35), .Y(n_38) );
endmodule