module real_jpeg_26031_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_49;
wire n_10;
wire n_68;
wire n_83;
wire n_78;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_61;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_16;

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_0),
.B(n_15),
.C(n_34),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_0),
.A2(n_31),
.B1(n_40),
.B2(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_0),
.A2(n_14),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_0),
.B(n_74),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_3),
.A2(n_15),
.B1(n_21),
.B2(n_22),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_3),
.A2(n_22),
.B1(n_31),
.B2(n_40),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_4),
.A2(n_15),
.B1(n_21),
.B2(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_5),
.A2(n_31),
.B1(n_40),
.B2(n_48),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_5),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_5),
.A2(n_15),
.B1(n_21),
.B2(n_48),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_67),
.Y(n_9)
);

AOI21xp5_ASAP7_75t_L g10 ( 
.A1(n_11),
.A2(n_49),
.B(n_66),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_28),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_12),
.B(n_28),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_19),
.B1(n_23),
.B2(n_25),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_14),
.B(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_14),
.A2(n_26),
.B(n_62),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_16),
.Y(n_14)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_15),
.A2(n_21),
.B1(n_34),
.B2(n_41),
.Y(n_42)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_20),
.A2(n_53),
.B(n_54),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_21),
.B(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_35),
.B2(n_36),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_30),
.B(n_35),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_34),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_31),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_31),
.A2(n_40),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

BUFx4f_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_43),
.B(n_45),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_38),
.B(n_47),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_42),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_42),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_44),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_42),
.A2(n_80),
.B(n_81),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_57),
.B(n_65),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_52),
.Y(n_65)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_83),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_69),
.B(n_70),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_82),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_78),
.B2(n_79),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);


endmodule