module fake_netlist_5_949_n_569 (n_82, n_10, n_24, n_83, n_61, n_75, n_65, n_78, n_74, n_57, n_37, n_31, n_13, n_66, n_60, n_16, n_43, n_0, n_58, n_9, n_69, n_18, n_42, n_22, n_1, n_45, n_46, n_21, n_38, n_80, n_4, n_35, n_73, n_17, n_19, n_30, n_5, n_33, n_14, n_84, n_23, n_29, n_79, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_62, n_71, n_59, n_26, n_55, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_36, n_76, n_27, n_64, n_77, n_81, n_28, n_70, n_68, n_72, n_32, n_41, n_56, n_51, n_63, n_11, n_7, n_15, n_48, n_50, n_52, n_569);

input n_82;
input n_10;
input n_24;
input n_83;
input n_61;
input n_75;
input n_65;
input n_78;
input n_74;
input n_57;
input n_37;
input n_31;
input n_13;
input n_66;
input n_60;
input n_16;
input n_43;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_42;
input n_22;
input n_1;
input n_45;
input n_46;
input n_21;
input n_38;
input n_80;
input n_4;
input n_35;
input n_73;
input n_17;
input n_19;
input n_30;
input n_5;
input n_33;
input n_14;
input n_84;
input n_23;
input n_29;
input n_79;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_62;
input n_71;
input n_59;
input n_26;
input n_55;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_36;
input n_76;
input n_27;
input n_64;
input n_77;
input n_81;
input n_28;
input n_70;
input n_68;
input n_72;
input n_32;
input n_41;
input n_56;
input n_51;
input n_63;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;

output n_569;

wire n_137;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_444;
wire n_469;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_418;
wire n_248;
wire n_136;
wire n_124;
wire n_146;
wire n_86;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_408;
wire n_376;
wire n_503;
wire n_127;
wire n_235;
wire n_226;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_452;
wire n_397;
wire n_525;
wire n_111;
wire n_493;
wire n_483;
wire n_544;
wire n_155;
wire n_552;
wire n_547;
wire n_116;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_139;
wire n_105;
wire n_280;
wire n_378;
wire n_551;
wire n_382;
wire n_554;
wire n_254;
wire n_302;
wire n_265;
wire n_526;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_173;
wire n_198;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_321;
wire n_292;
wire n_100;
wire n_455;
wire n_417;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_507;
wire n_119;
wire n_497;
wire n_559;
wire n_275;
wire n_252;
wire n_295;
wire n_133;
wire n_330;
wire n_508;
wire n_506;
wire n_509;
wire n_568;
wire n_147;
wire n_373;
wire n_307;
wire n_439;
wire n_87;
wire n_150;
wire n_530;
wire n_556;
wire n_106;
wire n_209;
wire n_259;
wire n_448;
wire n_375;
wire n_301;
wire n_93;
wire n_186;
wire n_537;
wire n_134;
wire n_191;
wire n_492;
wire n_563;
wire n_171;
wire n_153;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_320;
wire n_518;
wire n_505;
wire n_286;
wire n_122;
wire n_282;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_132;
wire n_90;
wire n_546;
wire n_101;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_152;
wire n_540;
wire n_317;
wire n_323;
wire n_195;
wire n_356;
wire n_227;
wire n_271;
wire n_94;
wire n_335;
wire n_123;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_297;
wire n_156;
wire n_225;
wire n_377;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_131;
wire n_192;
wire n_223;
wire n_392;
wire n_158;
wire n_138;
wire n_264;
wire n_109;
wire n_472;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_95;
wire n_183;
wire n_185;
wire n_243;
wire n_398;
wire n_396;
wire n_347;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_459;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_221;
wire n_178;
wire n_386;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_104;
wire n_415;
wire n_141;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_336;
wire n_145;
wire n_521;
wire n_337;
wire n_430;
wire n_313;
wire n_88;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_311;
wire n_208;
wire n_142;
wire n_214;
wire n_328;
wire n_140;
wire n_299;
wire n_303;
wire n_369;
wire n_296;
wire n_241;
wire n_357;
wire n_184;
wire n_446;
wire n_445;
wire n_144;
wire n_114;
wire n_96;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_129;
wire n_342;
wire n_482;
wire n_517;
wire n_98;
wire n_361;
wire n_464;
wire n_363;
wire n_413;
wire n_402;
wire n_197;
wire n_107;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_384;
wire n_460;
wire n_277;
wire n_92;
wire n_338;
wire n_149;
wire n_477;
wire n_461;
wire n_333;
wire n_309;
wire n_512;
wire n_462;
wire n_130;
wire n_322;
wire n_567;
wire n_258;
wire n_151;
wire n_306;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_474;
wire n_112;
wire n_542;
wire n_85;
wire n_488;
wire n_463;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_489;
wire n_310;
wire n_504;
wire n_511;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_102;
wire n_273;
wire n_349;
wire n_270;
wire n_230;
wire n_118;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_206;
wire n_172;
wire n_217;
wire n_440;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_365;
wire n_91;
wire n_176;
wire n_557;
wire n_182;
wire n_143;
wire n_354;
wire n_480;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_180;
wire n_560;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_108;
wire n_487;
wire n_495;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_405;
wire n_359;
wire n_490;
wire n_117;
wire n_326;
wire n_233;
wire n_404;
wire n_205;
wire n_366;
wire n_113;
wire n_246;
wire n_179;
wire n_125;
wire n_410;
wire n_558;
wire n_269;
wire n_529;
wire n_128;
wire n_285;
wire n_412;
wire n_120;
wire n_232;
wire n_327;
wire n_135;
wire n_126;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_565;
wire n_426;
wire n_520;
wire n_566;
wire n_409;
wire n_500;
wire n_562;
wire n_154;
wire n_148;
wire n_300;
wire n_435;
wire n_159;
wire n_334;
wire n_541;
wire n_391;
wire n_434;
wire n_539;
wire n_175;
wire n_538;
wire n_262;
wire n_238;
wire n_99;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_121;
wire n_242;
wire n_360;
wire n_200;
wire n_162;
wire n_222;
wire n_89;
wire n_438;
wire n_115;
wire n_324;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_103;
wire n_348;
wire n_97;
wire n_166;
wire n_424;
wire n_256;
wire n_305;
wire n_533;
wire n_278;
wire n_110;

INVx1_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

CKINVDCx5p33_ASAP7_75t_R g86 ( 
.A(n_62),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVxp67_ASAP7_75t_SL g89 ( 
.A(n_20),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

INVxp33_ASAP7_75t_SL g91 ( 
.A(n_65),
.Y(n_91)
);

INVxp67_ASAP7_75t_SL g92 ( 
.A(n_64),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_83),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_28),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_2),
.Y(n_97)
);

INVxp67_ASAP7_75t_SL g98 ( 
.A(n_53),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_17),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_9),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_39),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_19),
.Y(n_103)
);

CKINVDCx5p33_ASAP7_75t_R g104 ( 
.A(n_72),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_44),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_6),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_1),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

CKINVDCx5p33_ASAP7_75t_R g109 ( 
.A(n_50),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_37),
.B(n_71),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_1),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_0),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

INVxp67_ASAP7_75t_SL g114 ( 
.A(n_4),
.Y(n_114)
);

INVxp67_ASAP7_75t_SL g115 ( 
.A(n_30),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_12),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_15),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_33),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_16),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_35),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_25),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_9),
.Y(n_122)
);

INVxp33_ASAP7_75t_L g123 ( 
.A(n_13),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_82),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_52),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_67),
.Y(n_126)
);

INVx4_ASAP7_75t_R g127 ( 
.A(n_48),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_4),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_18),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_36),
.Y(n_132)
);

INVxp33_ASAP7_75t_SL g133 ( 
.A(n_26),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_49),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_75),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_55),
.Y(n_136)
);

INVx2_ASAP7_75t_SL g137 ( 
.A(n_76),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_56),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_0),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_32),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_2),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_41),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_59),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_60),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_80),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_47),
.Y(n_147)
);

INVxp67_ASAP7_75t_SL g148 ( 
.A(n_21),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_77),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_45),
.Y(n_150)
);

INVxp67_ASAP7_75t_SL g151 ( 
.A(n_51),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_31),
.Y(n_152)
);

INVxp67_ASAP7_75t_SL g153 ( 
.A(n_79),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_11),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_23),
.Y(n_155)
);

INVxp33_ASAP7_75t_SL g156 ( 
.A(n_42),
.Y(n_156)
);

INVxp33_ASAP7_75t_L g157 ( 
.A(n_73),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_5),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_43),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_22),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_7),
.Y(n_161)
);

INVxp33_ASAP7_75t_L g162 ( 
.A(n_69),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_68),
.Y(n_163)
);

INVxp67_ASAP7_75t_SL g164 ( 
.A(n_10),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_6),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_145),
.B(n_123),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_107),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_101),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_165),
.Y(n_169)
);

AND2x4_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_3),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_123),
.B(n_8),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_113),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_165),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_101),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_165),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_106),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_111),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_112),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_107),
.B(n_8),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_122),
.Y(n_181)
);

NOR2x1_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_14),
.Y(n_182)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_113),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_142),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_135),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_97),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_87),
.B(n_66),
.Y(n_190)
);

AND2x6_ASAP7_75t_L g191 ( 
.A(n_113),
.B(n_24),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_85),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_97),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_88),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_157),
.B(n_27),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_113),
.Y(n_196)
);

AND2x4_ASAP7_75t_L g197 ( 
.A(n_87),
.B(n_34),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_93),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_94),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_125),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_157),
.B(n_40),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_99),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_125),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_141),
.B(n_137),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_102),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_129),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_141),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_105),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_108),
.Y(n_209)
);

NAND2xp33_ASAP7_75t_SL g210 ( 
.A(n_162),
.B(n_129),
.Y(n_210)
);

OA21x2_ASAP7_75t_L g211 ( 
.A1(n_116),
.A2(n_54),
.B(n_134),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_136),
.Y(n_212)
);

AND2x4_ASAP7_75t_L g213 ( 
.A(n_100),
.B(n_130),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_114),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_126),
.B(n_150),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_118),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_119),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_121),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_124),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_91),
.B(n_156),
.Y(n_220)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_110),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_128),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_90),
.B(n_164),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_89),
.B(n_148),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_92),
.B(n_151),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_136),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_131),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_98),
.B(n_153),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_132),
.Y(n_229)
);

BUFx6f_ASAP7_75t_SL g230 ( 
.A(n_138),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_96),
.B(n_120),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_139),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_143),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_146),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_147),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_149),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_152),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_154),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_163),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_169),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_166),
.B(n_91),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_210),
.A2(n_135),
.B1(n_133),
.B2(n_156),
.Y(n_242)
);

AND2x4_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_115),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_173),
.Y(n_244)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_191),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_213),
.A2(n_133),
.B1(n_117),
.B2(n_103),
.Y(n_246)
);

OR2x6_ASAP7_75t_L g247 ( 
.A(n_220),
.B(n_160),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_212),
.B(n_155),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_175),
.Y(n_249)
);

BUFx8_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_220),
.B(n_86),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_95),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_176),
.Y(n_253)
);

NOR2xp67_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_104),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_200),
.B(n_109),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_226),
.Y(n_256)
);

NOR2xp67_ASAP7_75t_L g257 ( 
.A(n_214),
.B(n_144),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_172),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_213),
.B(n_127),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_221),
.A2(n_214),
.B1(n_170),
.B2(n_215),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_200),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_224),
.B(n_228),
.Y(n_262)
);

NOR3xp33_ASAP7_75t_L g263 ( 
.A(n_171),
.B(n_167),
.C(n_228),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_170),
.B(n_197),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_200),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_206),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_223),
.B(n_225),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_203),
.B(n_207),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_223),
.B(n_225),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_203),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_197),
.B(n_203),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_167),
.A2(n_180),
.B1(n_206),
.B2(n_195),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_207),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_172),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_168),
.B(n_174),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_172),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_189),
.B(n_204),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_207),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_188),
.B(n_204),
.Y(n_279)
);

INVxp67_ASAP7_75t_SL g280 ( 
.A(n_190),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_192),
.B(n_202),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_196),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_201),
.B(n_190),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_183),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_189),
.B(n_234),
.Y(n_285)
);

OAI221xp5_ASAP7_75t_L g286 ( 
.A1(n_177),
.A2(n_178),
.B1(n_186),
.B2(n_181),
.C(n_185),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_230),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_183),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_194),
.A2(n_216),
.B(n_237),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_218),
.Y(n_290)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_199),
.B(n_233),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_218),
.B(n_227),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_229),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_218),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_227),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_184),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_232),
.Y(n_297)
);

INVxp33_ASAP7_75t_L g298 ( 
.A(n_179),
.Y(n_298)
);

BUFx12f_ASAP7_75t_L g299 ( 
.A(n_250),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_279),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_285),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_268),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_290),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_268),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_263),
.A2(n_238),
.B1(n_219),
.B2(n_236),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_258),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_267),
.B(n_182),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_274),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_291),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_276),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_261),
.Y(n_311)
);

AND2x4_ASAP7_75t_L g312 ( 
.A(n_275),
.B(n_187),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_265),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_270),
.Y(n_314)
);

OR2x6_ASAP7_75t_L g315 ( 
.A(n_247),
.B(n_266),
.Y(n_315)
);

AOI211xp5_ASAP7_75t_L g316 ( 
.A1(n_269),
.A2(n_209),
.B(n_222),
.C(n_198),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_280),
.B(n_235),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_273),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_257),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_242),
.A2(n_205),
.B1(n_208),
.B2(n_217),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_260),
.B(n_227),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_246),
.B(n_193),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_278),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_290),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_283),
.B(n_191),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_288),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_277),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_262),
.B(n_191),
.Y(n_328)
);

O2A1O1Ixp33_ASAP7_75t_L g329 ( 
.A1(n_239),
.A2(n_211),
.B(n_264),
.C(n_289),
.Y(n_329)
);

OR2x6_ASAP7_75t_L g330 ( 
.A(n_247),
.B(n_211),
.Y(n_330)
);

INVx2_ASAP7_75t_SL g331 ( 
.A(n_247),
.Y(n_331)
);

INVx2_ASAP7_75t_SL g332 ( 
.A(n_256),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_290),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_242),
.A2(n_272),
.B1(n_241),
.B2(n_251),
.Y(n_334)
);

A2O1A1Ixp33_ASAP7_75t_L g335 ( 
.A1(n_271),
.A2(n_248),
.B(n_289),
.C(n_243),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_243),
.B(n_254),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_255),
.B(n_292),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_298),
.B(n_252),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_272),
.A2(n_259),
.B1(n_286),
.B2(n_296),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_255),
.B(n_284),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_282),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_281),
.B(n_253),
.Y(n_342)
);

AND2x4_ASAP7_75t_L g343 ( 
.A(n_244),
.B(n_240),
.Y(n_343)
);

AOI221xp5_ASAP7_75t_L g344 ( 
.A1(n_293),
.A2(n_297),
.B1(n_249),
.B2(n_287),
.C(n_294),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_245),
.B(n_294),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_294),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_250),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_295),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_245),
.B(n_295),
.Y(n_349)
);

BUFx2_ASAP7_75t_SL g350 ( 
.A(n_295),
.Y(n_350)
);

OR2x2_ASAP7_75t_L g351 ( 
.A(n_277),
.B(n_212),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_280),
.B(n_267),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_268),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_280),
.B(n_267),
.Y(n_354)
);

INVx2_ASAP7_75t_SL g355 ( 
.A(n_301),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g356 ( 
.A1(n_354),
.A2(n_352),
.B1(n_330),
.B2(n_328),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_338),
.B(n_332),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_324),
.Y(n_358)
);

INVx3_ASAP7_75t_SL g359 ( 
.A(n_315),
.Y(n_359)
);

O2A1O1Ixp33_ASAP7_75t_L g360 ( 
.A1(n_335),
.A2(n_329),
.B(n_307),
.C(n_322),
.Y(n_360)
);

NAND3xp33_ASAP7_75t_L g361 ( 
.A(n_316),
.B(n_305),
.C(n_353),
.Y(n_361)
);

BUFx10_ASAP7_75t_L g362 ( 
.A(n_312),
.Y(n_362)
);

A2O1A1Ixp33_ASAP7_75t_L g363 ( 
.A1(n_334),
.A2(n_304),
.B(n_302),
.C(n_325),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_337),
.A2(n_336),
.B(n_349),
.Y(n_364)
);

A2O1A1Ixp33_ASAP7_75t_L g365 ( 
.A1(n_334),
.A2(n_342),
.B(n_317),
.C(n_316),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_305),
.A2(n_339),
.B1(n_331),
.B2(n_351),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_327),
.B(n_309),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_345),
.A2(n_340),
.B(n_321),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_300),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_341),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_330),
.A2(n_339),
.B(n_320),
.Y(n_371)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_306),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_333),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_312),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_315),
.Y(n_375)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_308),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_326),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_320),
.A2(n_330),
.B1(n_319),
.B2(n_318),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_346),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_310),
.Y(n_380)
);

OR2x6_ASAP7_75t_L g381 ( 
.A(n_299),
.B(n_347),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_303),
.Y(n_382)
);

INVx2_ASAP7_75t_SL g383 ( 
.A(n_348),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_311),
.B(n_313),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_344),
.B(n_314),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_323),
.Y(n_386)
);

INVx3_ASAP7_75t_SL g387 ( 
.A(n_303),
.Y(n_387)
);

OR2x2_ASAP7_75t_SL g388 ( 
.A(n_350),
.B(n_188),
.Y(n_388)
);

AND2x4_ASAP7_75t_L g389 ( 
.A(n_302),
.B(n_304),
.Y(n_389)
);

BUFx12f_ASAP7_75t_L g390 ( 
.A(n_299),
.Y(n_390)
);

NAND2x1p5_ASAP7_75t_L g391 ( 
.A(n_301),
.B(n_332),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_343),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_352),
.B(n_354),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_299),
.Y(n_394)
);

NAND2x1p5_ASAP7_75t_L g395 ( 
.A(n_301),
.B(n_332),
.Y(n_395)
);

NAND2x1p5_ASAP7_75t_L g396 ( 
.A(n_301),
.B(n_332),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_338),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_338),
.B(n_267),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_352),
.B(n_354),
.Y(n_399)
);

BUFx12f_ASAP7_75t_L g400 ( 
.A(n_299),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_327),
.Y(n_401)
);

OR2x2_ASAP7_75t_L g402 ( 
.A(n_327),
.B(n_188),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_352),
.B(n_354),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_343),
.Y(n_404)
);

AND2x2_ASAP7_75t_SL g405 ( 
.A(n_334),
.B(n_263),
.Y(n_405)
);

BUFx4f_ASAP7_75t_SL g406 ( 
.A(n_299),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_306),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_338),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_352),
.B(n_354),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_329),
.A2(n_335),
.B(n_328),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_338),
.B(n_267),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_338),
.B(n_267),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_343),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_343),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_302),
.B(n_304),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_302),
.B(n_304),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_343),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_386),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_398),
.B(n_411),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_387),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_412),
.B(n_399),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_390),
.Y(n_422)
);

AO31x2_ASAP7_75t_L g423 ( 
.A1(n_363),
.A2(n_366),
.A3(n_365),
.B(n_399),
.Y(n_423)
);

OR2x6_ASAP7_75t_L g424 ( 
.A(n_371),
.B(n_368),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_370),
.Y(n_425)
);

OAI22xp33_ASAP7_75t_L g426 ( 
.A1(n_393),
.A2(n_409),
.B1(n_403),
.B2(n_371),
.Y(n_426)
);

INVx2_ASAP7_75t_SL g427 ( 
.A(n_389),
.Y(n_427)
);

AO21x2_ASAP7_75t_L g428 ( 
.A1(n_410),
.A2(n_360),
.B(n_364),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_372),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_405),
.B(n_416),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_404),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_413),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_414),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_389),
.B(n_415),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_392),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_417),
.Y(n_436)
);

OAI21x1_ASAP7_75t_L g437 ( 
.A1(n_356),
.A2(n_382),
.B(n_384),
.Y(n_437)
);

AOI21x1_ASAP7_75t_L g438 ( 
.A1(n_380),
.A2(n_416),
.B(n_415),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_377),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_397),
.B(n_408),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_376),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_376),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_407),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_400),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_374),
.B(n_385),
.Y(n_445)
);

INVxp33_ASAP7_75t_L g446 ( 
.A(n_367),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_407),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_383),
.Y(n_448)
);

OR2x6_ASAP7_75t_L g449 ( 
.A(n_391),
.B(n_396),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_374),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_379),
.Y(n_451)
);

OA21x2_ASAP7_75t_L g452 ( 
.A1(n_361),
.A2(n_378),
.B(n_366),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g453 ( 
.A(n_401),
.Y(n_453)
);

AOI222xp33_ASAP7_75t_L g454 ( 
.A1(n_369),
.A2(n_361),
.B1(n_401),
.B2(n_357),
.C1(n_375),
.C2(n_359),
.Y(n_454)
);

OR2x6_ASAP7_75t_L g455 ( 
.A(n_395),
.B(n_355),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_378),
.B(n_362),
.Y(n_456)
);

OA21x2_ASAP7_75t_L g457 ( 
.A1(n_402),
.A2(n_369),
.B(n_388),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_358),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_358),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_373),
.Y(n_460)
);

OR2x6_ASAP7_75t_L g461 ( 
.A(n_381),
.B(n_373),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_381),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_381),
.B(n_394),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_406),
.B(n_398),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_386),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_387),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_386),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_398),
.B(n_411),
.Y(n_468)
);

INVx4_ASAP7_75t_L g469 ( 
.A(n_420),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_421),
.B(n_419),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_425),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_453),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_421),
.B(n_419),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_418),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_434),
.B(n_430),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_426),
.B(n_468),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_465),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_467),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g479 ( 
.A(n_453),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_439),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_468),
.B(n_445),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_430),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_445),
.B(n_452),
.Y(n_483)
);

INVx5_ASAP7_75t_SL g484 ( 
.A(n_420),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_434),
.B(n_427),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_452),
.B(n_423),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_423),
.B(n_424),
.Y(n_487)
);

OAI31xp33_ASAP7_75t_L g488 ( 
.A1(n_446),
.A2(n_456),
.A3(n_464),
.B(n_435),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_466),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_456),
.A2(n_427),
.B1(n_424),
.B2(n_454),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_423),
.B(n_424),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_450),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_L g493 ( 
.A1(n_470),
.A2(n_424),
.B1(n_446),
.B2(n_457),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_472),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_472),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_474),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_470),
.B(n_473),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_473),
.B(n_441),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_471),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_481),
.B(n_440),
.Y(n_500)
);

AOI222xp33_ASAP7_75t_L g501 ( 
.A1(n_481),
.A2(n_433),
.B1(n_432),
.B2(n_431),
.C1(n_464),
.C2(n_436),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_482),
.B(n_448),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_477),
.Y(n_503)
);

OAI221xp5_ASAP7_75t_L g504 ( 
.A1(n_490),
.A2(n_457),
.B1(n_451),
.B2(n_449),
.C(n_448),
.Y(n_504)
);

OAI211xp5_ASAP7_75t_SL g505 ( 
.A1(n_488),
.A2(n_462),
.B(n_443),
.C(n_447),
.Y(n_505)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_476),
.B(n_428),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_478),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_482),
.B(n_483),
.Y(n_508)
);

OAI31xp33_ASAP7_75t_SL g509 ( 
.A1(n_483),
.A2(n_437),
.A3(n_460),
.B(n_459),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_487),
.B(n_442),
.Y(n_510)
);

OAI222xp33_ASAP7_75t_L g511 ( 
.A1(n_479),
.A2(n_449),
.B1(n_455),
.B2(n_461),
.C1(n_438),
.C2(n_442),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_487),
.B(n_429),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_494),
.Y(n_513)
);

AOI31xp33_ASAP7_75t_L g514 ( 
.A1(n_501),
.A2(n_422),
.A3(n_444),
.B(n_463),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_500),
.B(n_475),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_497),
.B(n_491),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_497),
.B(n_491),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_495),
.B(n_475),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_494),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_496),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_503),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_507),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_502),
.B(n_475),
.Y(n_523)
);

OR2x2_ASAP7_75t_L g524 ( 
.A(n_508),
.B(n_486),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_498),
.B(n_479),
.Y(n_525)
);

INVx1_ASAP7_75t_SL g526 ( 
.A(n_510),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_498),
.B(n_492),
.Y(n_527)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_510),
.Y(n_528)
);

INVxp67_ASAP7_75t_SL g529 ( 
.A(n_512),
.Y(n_529)
);

OAI22xp33_ASAP7_75t_L g530 ( 
.A1(n_504),
.A2(n_449),
.B1(n_455),
.B2(n_457),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_519),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_514),
.B(n_458),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_520),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_527),
.B(n_512),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_516),
.B(n_517),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_523),
.B(n_469),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_525),
.B(n_493),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_515),
.B(n_499),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_521),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_535),
.B(n_516),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_534),
.B(n_513),
.Y(n_541)
);

OR2x2_ASAP7_75t_L g542 ( 
.A(n_531),
.B(n_524),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_531),
.B(n_513),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_533),
.B(n_506),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_539),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_538),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_537),
.Y(n_547)
);

OR2x2_ASAP7_75t_L g548 ( 
.A(n_532),
.B(n_524),
.Y(n_548)
);

NAND3xp33_ASAP7_75t_L g549 ( 
.A(n_547),
.B(n_536),
.C(n_509),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_548),
.B(n_530),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_542),
.Y(n_551)
);

AOI221xp5_ASAP7_75t_SL g552 ( 
.A1(n_543),
.A2(n_541),
.B1(n_546),
.B2(n_545),
.C(n_544),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_540),
.B(n_518),
.Y(n_553)
);

AOI211xp5_ASAP7_75t_SL g554 ( 
.A1(n_544),
.A2(n_511),
.B(n_529),
.C(n_505),
.Y(n_554)
);

NOR3xp33_ASAP7_75t_L g555 ( 
.A(n_547),
.B(n_469),
.C(n_485),
.Y(n_555)
);

NOR2x1_ASAP7_75t_L g556 ( 
.A(n_549),
.B(n_522),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_551),
.Y(n_557)
);

AOI221xp5_ASAP7_75t_L g558 ( 
.A1(n_552),
.A2(n_526),
.B1(n_517),
.B2(n_528),
.C(n_489),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_550),
.Y(n_559)
);

NAND3xp33_ASAP7_75t_L g560 ( 
.A(n_556),
.B(n_554),
.C(n_555),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_559),
.B(n_553),
.Y(n_561)
);

NAND2x1_ASAP7_75t_SL g562 ( 
.A(n_557),
.B(n_463),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_560),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_562),
.Y(n_564)
);

NOR3x2_ASAP7_75t_L g565 ( 
.A(n_563),
.B(n_422),
.C(n_444),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_565),
.B(n_561),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_566),
.A2(n_564),
.B(n_558),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_567),
.Y(n_568)
);

AOI211xp5_ASAP7_75t_L g569 ( 
.A1(n_568),
.A2(n_489),
.B(n_484),
.C(n_480),
.Y(n_569)
);


endmodule