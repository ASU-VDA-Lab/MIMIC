module fake_netlist_5_1953_n_1933 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1933);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1933;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_174;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_990;
wire n_836;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_177;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_1089;
wire n_927;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g158 ( 
.A(n_85),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_114),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_9),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_98),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_19),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_102),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_30),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_100),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_21),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_4),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_82),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_106),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_150),
.Y(n_170)
);

BUFx10_ASAP7_75t_L g171 ( 
.A(n_23),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_10),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_50),
.Y(n_173)
);

BUFx10_ASAP7_75t_L g174 ( 
.A(n_62),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_113),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_140),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_47),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_4),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_79),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_105),
.Y(n_180)
);

BUFx10_ASAP7_75t_L g181 ( 
.A(n_136),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_86),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_130),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_75),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_115),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_83),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_58),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_48),
.Y(n_188)
);

BUFx8_ASAP7_75t_SL g189 ( 
.A(n_22),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_52),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_27),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_81),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_68),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_42),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_21),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_127),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_17),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_91),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_90),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_41),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_78),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_40),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_26),
.Y(n_203)
);

BUFx8_ASAP7_75t_SL g204 ( 
.A(n_22),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_64),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_14),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_93),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_155),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_7),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_34),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_128),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_31),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_147),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_2),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_123),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_51),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_53),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_129),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_71),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_139),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_5),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_46),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_17),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_59),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_87),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_73),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_125),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_80),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_151),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_135),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_28),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_1),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_133),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_33),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_35),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_10),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_138),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_32),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_19),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_143),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_43),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_57),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_36),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_49),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_5),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_33),
.Y(n_246)
);

INVxp67_ASAP7_75t_SL g247 ( 
.A(n_25),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_61),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_76),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_6),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_110),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_41),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_117),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_119),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_156),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_6),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_54),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_42),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_84),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_103),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_20),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_12),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_152),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_39),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_101),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_112),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_63),
.Y(n_267)
);

CKINVDCx12_ASAP7_75t_R g268 ( 
.A(n_31),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_153),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_96),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_146),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_7),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_20),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_120),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_8),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_97),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_2),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_28),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_116),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_56),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_94),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_149),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_11),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_92),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_111),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_24),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_157),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_132),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_8),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_37),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_77),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_27),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_142),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_36),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_37),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_40),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_107),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_23),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_30),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_137),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_126),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_13),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_3),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_109),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_1),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_121),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_99),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_69),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_134),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_88),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_32),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_154),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_29),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_191),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_189),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_159),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_204),
.Y(n_317)
);

INVxp33_ASAP7_75t_SL g318 ( 
.A(n_162),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_191),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_191),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_183),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_185),
.Y(n_322)
);

INVxp33_ASAP7_75t_SL g323 ( 
.A(n_162),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_191),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_196),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_199),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_205),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_207),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_193),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_198),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_268),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_191),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_273),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_217),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_273),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_283),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_283),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_286),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_286),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_167),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_167),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_215),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_278),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_230),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_278),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_222),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_160),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_172),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_211),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_313),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_214),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_282),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_211),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_225),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_194),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_197),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_177),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_293),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_212),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_221),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_226),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_233),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_232),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_238),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_239),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_237),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_227),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_245),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_293),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_250),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_241),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_242),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_253),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_258),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_249),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_254),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_255),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_277),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_257),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_290),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_259),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_305),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_311),
.Y(n_383)
);

INVxp33_ASAP7_75t_L g384 ( 
.A(n_158),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_260),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_202),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_202),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g388 ( 
.A(n_161),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_174),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_325),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_321),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_314),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_314),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_353),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_319),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_388),
.B(n_163),
.Y(n_396)
);

CKINVDCx11_ASAP7_75t_R g397 ( 
.A(n_322),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_349),
.B(n_369),
.Y(n_398)
);

OA21x2_ASAP7_75t_L g399 ( 
.A1(n_319),
.A2(n_180),
.B(n_179),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_329),
.B(n_176),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_353),
.B(n_256),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_357),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_320),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_320),
.B(n_163),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_324),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_324),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_332),
.Y(n_407)
);

AND2x6_ASAP7_75t_L g408 ( 
.A(n_332),
.B(n_179),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_335),
.Y(n_409)
);

OAI21x1_ASAP7_75t_L g410 ( 
.A1(n_335),
.A2(n_188),
.B(n_180),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_348),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_333),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_348),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_351),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_365),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_330),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_350),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_350),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_355),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_316),
.A2(n_296),
.B1(n_234),
.B2(n_236),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_358),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_333),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_355),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_336),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_356),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_356),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_359),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_358),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_359),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_360),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_360),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_340),
.B(n_188),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_336),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_337),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_340),
.B(n_256),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_363),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_337),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_338),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_338),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_363),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_341),
.B(n_343),
.Y(n_441)
);

AND2x6_ASAP7_75t_L g442 ( 
.A(n_389),
.B(n_208),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_364),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_339),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_331),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_339),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_326),
.B(n_168),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_364),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_368),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_368),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_341),
.B(n_208),
.Y(n_451)
);

BUFx12f_ASAP7_75t_L g452 ( 
.A(n_315),
.Y(n_452)
);

OA21x2_ASAP7_75t_L g453 ( 
.A1(n_370),
.A2(n_218),
.B(n_216),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_389),
.B(n_174),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_327),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_370),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_318),
.B(n_174),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_374),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_393),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_392),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_428),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_410),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_392),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_400),
.B(n_328),
.Y(n_464)
);

INVx2_ASAP7_75t_SL g465 ( 
.A(n_428),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_391),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_398),
.B(n_342),
.Y(n_467)
);

NOR2x1p5_ASAP7_75t_L g468 ( 
.A(n_390),
.B(n_317),
.Y(n_468)
);

AOI22xp33_ASAP7_75t_L g469 ( 
.A1(n_398),
.A2(n_375),
.B1(n_384),
.B2(n_323),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_447),
.B(n_334),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_411),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_411),
.Y(n_472)
);

AOI22xp33_ASAP7_75t_L g473 ( 
.A1(n_432),
.A2(n_451),
.B1(n_401),
.B2(n_453),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_393),
.Y(n_474)
);

BUFx6f_ASAP7_75t_SL g475 ( 
.A(n_394),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_421),
.B(n_346),
.Y(n_476)
);

AND2x6_ASAP7_75t_L g477 ( 
.A(n_401),
.B(n_216),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_410),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_455),
.B(n_354),
.Y(n_479)
);

OR2x6_ASAP7_75t_L g480 ( 
.A(n_452),
.B(n_345),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_410),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_392),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_403),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_403),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_405),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_413),
.Y(n_486)
);

BUFx10_ASAP7_75t_L g487 ( 
.A(n_414),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_421),
.B(n_361),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_396),
.B(n_371),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_405),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_435),
.B(n_386),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_396),
.B(n_373),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_404),
.B(n_381),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_404),
.B(n_385),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_397),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_406),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_406),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_394),
.Y(n_498)
);

AO21x2_ASAP7_75t_L g499 ( 
.A1(n_457),
.A2(n_184),
.B(n_165),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_407),
.Y(n_500)
);

NAND3xp33_ASAP7_75t_L g501 ( 
.A(n_420),
.B(n_347),
.C(n_200),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_394),
.B(n_263),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_407),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_432),
.A2(n_218),
.B1(n_309),
.B2(n_240),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_393),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_393),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_453),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_422),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_422),
.Y(n_509)
);

NAND2xp33_ASAP7_75t_SL g510 ( 
.A(n_435),
.B(n_164),
.Y(n_510)
);

INVx4_ASAP7_75t_L g511 ( 
.A(n_453),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_413),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_442),
.B(n_265),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_417),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_395),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_395),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_445),
.A2(n_372),
.B1(n_379),
.B2(n_377),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_417),
.Y(n_518)
);

BUFx10_ASAP7_75t_L g519 ( 
.A(n_414),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_395),
.Y(n_520)
);

AO21x2_ASAP7_75t_L g521 ( 
.A1(n_454),
.A2(n_187),
.B(n_186),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_418),
.Y(n_522)
);

BUFx10_ASAP7_75t_L g523 ( 
.A(n_415),
.Y(n_523)
);

INVx4_ASAP7_75t_L g524 ( 
.A(n_453),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_422),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_422),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_442),
.B(n_266),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_432),
.B(n_386),
.Y(n_528)
);

INVxp33_ASAP7_75t_L g529 ( 
.A(n_415),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_442),
.Y(n_530)
);

INVx5_ASAP7_75t_L g531 ( 
.A(n_408),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_395),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_416),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_445),
.B(n_367),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_422),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_422),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_422),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_432),
.A2(n_240),
.B1(n_309),
.B2(n_270),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_418),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_437),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_437),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_419),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_420),
.B(n_376),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_402),
.Y(n_544)
);

AND2x6_ASAP7_75t_L g545 ( 
.A(n_451),
.B(n_270),
.Y(n_545)
);

OR2x2_ASAP7_75t_L g546 ( 
.A(n_441),
.B(n_387),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_402),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_452),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_453),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_451),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_437),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_437),
.Y(n_552)
);

NAND2xp33_ASAP7_75t_SL g553 ( 
.A(n_441),
.B(n_164),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_419),
.B(n_362),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_423),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_423),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_451),
.B(n_366),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_425),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_437),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_425),
.B(n_344),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_437),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_426),
.B(n_374),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_426),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_427),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_452),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_427),
.B(n_352),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_442),
.B(n_271),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_429),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_429),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_442),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_430),
.Y(n_571)
);

INVxp33_ASAP7_75t_L g572 ( 
.A(n_430),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_442),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_442),
.B(n_274),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_437),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_446),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_442),
.A2(n_383),
.B1(n_382),
.B2(n_380),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_431),
.B(n_378),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_446),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_442),
.B(n_201),
.Y(n_580)
);

OR2x6_ASAP7_75t_L g581 ( 
.A(n_431),
.B(n_387),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_436),
.Y(n_582)
);

NAND3xp33_ASAP7_75t_L g583 ( 
.A(n_436),
.B(n_262),
.C(n_235),
.Y(n_583)
);

AND2x6_ASAP7_75t_L g584 ( 
.A(n_440),
.B(n_213),
.Y(n_584)
);

INVx1_ASAP7_75t_SL g585 ( 
.A(n_440),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_443),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_446),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_443),
.B(n_181),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_449),
.B(n_168),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_446),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_438),
.B(n_219),
.Y(n_591)
);

OAI22xp33_ASAP7_75t_SL g592 ( 
.A1(n_449),
.A2(n_247),
.B1(n_234),
.B2(n_166),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_450),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_450),
.B(n_181),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_456),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_438),
.B(n_220),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_446),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_446),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_456),
.B(n_169),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_446),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_438),
.B(n_224),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_448),
.B(n_169),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_448),
.B(n_170),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_438),
.B(n_228),
.Y(n_604)
);

INVx8_ASAP7_75t_L g605 ( 
.A(n_408),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_399),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_448),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_444),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_550),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_473),
.B(n_229),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_550),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_533),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_498),
.B(n_378),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_533),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_507),
.B(n_399),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_471),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_544),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_507),
.B(n_399),
.Y(n_618)
);

AND2x4_ASAP7_75t_L g619 ( 
.A(n_498),
.B(n_528),
.Y(n_619)
);

BUFx4f_ASAP7_75t_L g620 ( 
.A(n_480),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_528),
.B(n_380),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_460),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_472),
.Y(n_623)
);

NAND3x1_ASAP7_75t_L g624 ( 
.A(n_517),
.B(n_382),
.C(n_383),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_489),
.A2(n_288),
.B1(n_173),
.B2(n_175),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_460),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_486),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_585),
.B(n_171),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_492),
.B(n_210),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_463),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_512),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_514),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_463),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_507),
.B(n_399),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_482),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_465),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_507),
.B(n_399),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_518),
.Y(n_638)
);

NOR3xp33_ASAP7_75t_L g639 ( 
.A(n_592),
.B(n_279),
.C(n_267),
.Y(n_639)
);

NAND3xp33_ASAP7_75t_L g640 ( 
.A(n_522),
.B(n_269),
.C(n_312),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_544),
.Y(n_641)
);

NOR2x1p5_ASAP7_75t_L g642 ( 
.A(n_565),
.B(n_166),
.Y(n_642)
);

NAND2x1p5_ASAP7_75t_L g643 ( 
.A(n_530),
.B(n_244),
.Y(n_643)
);

AND2x4_ASAP7_75t_L g644 ( 
.A(n_562),
.B(n_458),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_562),
.B(n_458),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_507),
.B(n_248),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_562),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_539),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_578),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_482),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_542),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_555),
.Y(n_652)
);

INVxp67_ASAP7_75t_L g653 ( 
.A(n_554),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_556),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_608),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_578),
.B(n_458),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_558),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_563),
.Y(n_658)
);

NAND2x1p5_ASAP7_75t_L g659 ( 
.A(n_530),
.B(n_251),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_572),
.B(n_465),
.Y(n_660)
);

HB1xp67_ASAP7_75t_L g661 ( 
.A(n_461),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_578),
.Y(n_662)
);

BUFx10_ASAP7_75t_L g663 ( 
.A(n_534),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_549),
.B(n_280),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_549),
.B(n_287),
.Y(n_665)
);

INVx4_ASAP7_75t_L g666 ( 
.A(n_549),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_564),
.B(n_409),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_568),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_569),
.B(n_409),
.Y(n_669)
);

AOI22x1_ASAP7_75t_L g670 ( 
.A1(n_511),
.A2(n_304),
.B1(n_310),
.B2(n_308),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_467),
.B(n_171),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_572),
.B(n_170),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_571),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_487),
.Y(n_674)
);

AND2x4_ASAP7_75t_L g675 ( 
.A(n_582),
.B(n_444),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_586),
.B(n_444),
.Y(n_676)
);

INVx5_ASAP7_75t_L g677 ( 
.A(n_462),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_593),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_595),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_496),
.Y(n_680)
);

AND2x4_ASAP7_75t_L g681 ( 
.A(n_581),
.B(n_444),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_496),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_459),
.Y(n_683)
);

OAI22xp5_ASAP7_75t_L g684 ( 
.A1(n_469),
.A2(n_178),
.B1(n_289),
.B2(n_292),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_459),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_459),
.Y(n_686)
);

INVx4_ASAP7_75t_L g687 ( 
.A(n_549),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_608),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_467),
.A2(n_297),
.B1(n_175),
.B2(n_182),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_549),
.B(n_173),
.Y(n_690)
);

AND2x4_ASAP7_75t_L g691 ( 
.A(n_581),
.B(n_412),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_474),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_529),
.B(n_171),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_474),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_474),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_487),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_606),
.B(n_408),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_570),
.Y(n_698)
);

INVx4_ASAP7_75t_SL g699 ( 
.A(n_545),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_483),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_505),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_505),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_495),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_581),
.B(n_412),
.Y(n_704)
);

AND2x6_ASAP7_75t_L g705 ( 
.A(n_606),
.B(n_412),
.Y(n_705)
);

NAND3x1_ASAP7_75t_L g706 ( 
.A(n_560),
.B(n_243),
.C(n_178),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_505),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_570),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_515),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_483),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_515),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_515),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_493),
.B(n_182),
.Y(n_713)
);

INVx8_ASAP7_75t_L g714 ( 
.A(n_480),
.Y(n_714)
);

BUFx2_ASAP7_75t_L g715 ( 
.A(n_547),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_516),
.Y(n_716)
);

INVx1_ASAP7_75t_SL g717 ( 
.A(n_487),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_484),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_494),
.B(n_190),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_516),
.Y(n_720)
);

INVx4_ASAP7_75t_L g721 ( 
.A(n_462),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_484),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_485),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_516),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_529),
.B(n_243),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_520),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_511),
.B(n_408),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_520),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_SL g729 ( 
.A1(n_547),
.A2(n_298),
.B1(n_289),
.B2(n_292),
.Y(n_729)
);

NAND2x1p5_ASAP7_75t_L g730 ( 
.A(n_511),
.B(n_424),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_520),
.Y(n_731)
);

AND2x4_ASAP7_75t_L g732 ( 
.A(n_581),
.B(n_424),
.Y(n_732)
);

AND2x2_ASAP7_75t_SL g733 ( 
.A(n_566),
.B(n_181),
.Y(n_733)
);

NAND3xp33_ASAP7_75t_L g734 ( 
.A(n_504),
.B(n_538),
.C(n_591),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_485),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_524),
.B(n_408),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_462),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_532),
.Y(n_738)
);

A2O1A1Ixp33_ASAP7_75t_L g739 ( 
.A1(n_589),
.A2(n_439),
.B(n_434),
.C(n_433),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_532),
.Y(n_740)
);

BUFx10_ASAP7_75t_L g741 ( 
.A(n_495),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_532),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_506),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_524),
.B(n_408),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_524),
.A2(n_236),
.B1(n_295),
.B2(n_275),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_491),
.B(n_424),
.Y(n_746)
);

AND2x4_ASAP7_75t_L g747 ( 
.A(n_491),
.B(n_583),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_462),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_490),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_490),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_466),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_506),
.Y(n_752)
);

AND2x4_ASAP7_75t_L g753 ( 
.A(n_521),
.B(n_433),
.Y(n_753)
);

AOI22xp5_ASAP7_75t_L g754 ( 
.A1(n_499),
.A2(n_285),
.B1(n_192),
.B2(n_276),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_519),
.B(n_243),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_497),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_519),
.B(n_523),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_SL g758 ( 
.A(n_475),
.B(n_190),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_497),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_476),
.B(n_192),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_500),
.B(n_408),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_462),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_477),
.A2(n_302),
.B1(n_294),
.B2(n_295),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_500),
.B(n_408),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_557),
.B(n_275),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_478),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_503),
.Y(n_767)
);

NAND2x1p5_ASAP7_75t_L g768 ( 
.A(n_531),
.B(n_433),
.Y(n_768)
);

INVx1_ASAP7_75t_SL g769 ( 
.A(n_519),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_503),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_607),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_546),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_523),
.Y(n_773)
);

HB1xp67_ASAP7_75t_L g774 ( 
.A(n_546),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_478),
.B(n_276),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_535),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_478),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_535),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_478),
.B(n_408),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_535),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_478),
.B(n_434),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_655),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_766),
.B(n_499),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_629),
.B(n_499),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_644),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_629),
.A2(n_713),
.B1(n_719),
.B2(n_747),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_647),
.B(n_649),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_636),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_766),
.B(n_477),
.Y(n_789)
);

CKINVDCx20_ASAP7_75t_R g790 ( 
.A(n_612),
.Y(n_790)
);

CKINVDCx20_ASAP7_75t_R g791 ( 
.A(n_751),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_666),
.B(n_687),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_653),
.B(n_543),
.Y(n_793)
);

NAND3xp33_ASAP7_75t_SL g794 ( 
.A(n_653),
.B(n_565),
.C(n_548),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_636),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_644),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_688),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_666),
.B(n_477),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_687),
.B(n_477),
.Y(n_799)
);

BUFx3_ASAP7_75t_L g800 ( 
.A(n_614),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_645),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_737),
.B(n_477),
.Y(n_802)
);

INVx2_ASAP7_75t_SL g803 ( 
.A(n_628),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_647),
.B(n_488),
.Y(n_804)
);

AND2x6_ASAP7_75t_SL g805 ( 
.A(n_713),
.B(n_480),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_698),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_703),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_698),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_737),
.B(n_477),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_737),
.B(n_602),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_661),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_748),
.B(n_603),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_663),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_773),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_645),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_719),
.B(n_660),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_660),
.B(n_599),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_656),
.Y(n_818)
);

NOR3xp33_ASAP7_75t_SL g819 ( 
.A(n_729),
.B(n_303),
.C(n_302),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_760),
.B(n_521),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_733),
.B(n_479),
.Y(n_821)
);

AND2x6_ASAP7_75t_L g822 ( 
.A(n_777),
.B(n_481),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_656),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_661),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_647),
.B(n_523),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_707),
.Y(n_826)
);

BUFx3_ASAP7_75t_L g827 ( 
.A(n_617),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_707),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_649),
.B(n_502),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_743),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_662),
.B(n_480),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_621),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_619),
.B(n_468),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_752),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_746),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_649),
.B(n_677),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_663),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_746),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_700),
.Y(n_839)
);

INVx5_ASAP7_75t_L g840 ( 
.A(n_705),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_760),
.B(n_521),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_R g842 ( 
.A(n_758),
.B(n_548),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_677),
.B(n_619),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_621),
.B(n_470),
.Y(n_844)
);

HB1xp67_ASAP7_75t_L g845 ( 
.A(n_774),
.Y(n_845)
);

INVx2_ASAP7_75t_SL g846 ( 
.A(n_693),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_741),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_R g848 ( 
.A(n_758),
.B(n_553),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_698),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_681),
.B(n_501),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_748),
.B(n_481),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_681),
.B(n_588),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_610),
.A2(n_545),
.B1(n_584),
.B2(n_553),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_677),
.B(n_464),
.Y(n_854)
);

INVx5_ASAP7_75t_L g855 ( 
.A(n_705),
.Y(n_855)
);

AOI22xp5_ASAP7_75t_L g856 ( 
.A1(n_747),
.A2(n_545),
.B1(n_475),
.B2(n_573),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_671),
.B(n_594),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_680),
.B(n_481),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_677),
.B(n_510),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_682),
.B(n_481),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_710),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_756),
.Y(n_862)
);

AND2x2_ASAP7_75t_SL g863 ( 
.A(n_620),
.B(n_577),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_774),
.B(n_475),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_718),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_613),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_708),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_748),
.B(n_481),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_767),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_762),
.B(n_596),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_770),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_772),
.B(n_613),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_691),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_725),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_609),
.A2(n_545),
.B1(n_573),
.B2(n_584),
.Y(n_875)
);

NAND2x1p5_ASAP7_75t_L g876 ( 
.A(n_721),
.B(n_531),
.Y(n_876)
);

INVx3_ASAP7_75t_SL g877 ( 
.A(n_741),
.Y(n_877)
);

INVx3_ASAP7_75t_L g878 ( 
.A(n_708),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_762),
.B(n_601),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_708),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_722),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_611),
.A2(n_545),
.B1(n_584),
.B2(n_513),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_672),
.B(n_545),
.Y(n_883)
);

BUFx3_ASAP7_75t_L g884 ( 
.A(n_641),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_723),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_610),
.A2(n_584),
.B1(n_527),
.B2(n_574),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_672),
.B(n_510),
.Y(n_887)
);

INVxp67_ASAP7_75t_L g888 ( 
.A(n_755),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_691),
.B(n_508),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_762),
.B(n_604),
.Y(n_890)
);

INVx5_ASAP7_75t_L g891 ( 
.A(n_705),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_735),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_749),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_721),
.B(n_584),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_615),
.B(n_584),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_615),
.B(n_552),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_750),
.Y(n_897)
);

INVxp67_ASAP7_75t_L g898 ( 
.A(n_765),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_775),
.A2(n_567),
.B1(n_580),
.B2(n_552),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_759),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_704),
.Y(n_901)
);

CKINVDCx8_ASAP7_75t_R g902 ( 
.A(n_715),
.Y(n_902)
);

INVx4_ASAP7_75t_L g903 ( 
.A(n_705),
.Y(n_903)
);

OAI22xp5_ASAP7_75t_L g904 ( 
.A1(n_745),
.A2(n_294),
.B1(n_298),
.B2(n_299),
.Y(n_904)
);

AOI22xp5_ASAP7_75t_L g905 ( 
.A1(n_775),
.A2(n_559),
.B1(n_552),
.B2(n_598),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_616),
.B(n_623),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_704),
.B(n_281),
.Y(n_907)
);

NOR3xp33_ASAP7_75t_SL g908 ( 
.A(n_684),
.B(n_299),
.C(n_303),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_683),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_732),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_675),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_625),
.B(n_281),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_627),
.B(n_559),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_690),
.A2(n_559),
.B1(n_600),
.B2(n_598),
.Y(n_914)
);

AO22x1_ASAP7_75t_L g915 ( 
.A1(n_639),
.A2(n_203),
.B1(n_195),
.B2(n_209),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_674),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_618),
.B(n_508),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_675),
.Y(n_918)
);

CKINVDCx8_ASAP7_75t_R g919 ( 
.A(n_714),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_717),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_685),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_732),
.B(n_284),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_618),
.B(n_509),
.Y(n_923)
);

AND2x6_ASAP7_75t_SL g924 ( 
.A(n_757),
.B(n_206),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_634),
.B(n_509),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_634),
.B(n_525),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_686),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_637),
.B(n_525),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_631),
.B(n_526),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_676),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_632),
.B(n_526),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_717),
.B(n_284),
.Y(n_932)
);

INVx5_ASAP7_75t_L g933 ( 
.A(n_753),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_676),
.Y(n_934)
);

AND2x4_ASAP7_75t_L g935 ( 
.A(n_638),
.B(n_536),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_648),
.B(n_536),
.Y(n_936)
);

INVx2_ASAP7_75t_SL g937 ( 
.A(n_696),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_651),
.B(n_537),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_692),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_769),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_652),
.B(n_654),
.Y(n_941)
);

AND2x4_ASAP7_75t_L g942 ( 
.A(n_657),
.B(n_537),
.Y(n_942)
);

O2A1O1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_690),
.A2(n_575),
.B(n_600),
.C(n_597),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_637),
.B(n_540),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_714),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_763),
.B(n_285),
.Y(n_946)
);

INVx1_ASAP7_75t_SL g947 ( 
.A(n_769),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_781),
.B(n_540),
.Y(n_948)
);

INVx6_ASAP7_75t_L g949 ( 
.A(n_642),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_694),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_695),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_701),
.Y(n_952)
);

INVxp67_ASAP7_75t_SL g953 ( 
.A(n_730),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_702),
.Y(n_954)
);

INVxp67_ASAP7_75t_SL g955 ( 
.A(n_730),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_709),
.Y(n_956)
);

INVx2_ASAP7_75t_SL g957 ( 
.A(n_667),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_781),
.B(n_541),
.Y(n_958)
);

NOR2xp67_ASAP7_75t_L g959 ( 
.A(n_754),
.B(n_541),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_711),
.Y(n_960)
);

NOR2x2_ASAP7_75t_L g961 ( 
.A(n_745),
.B(n_684),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_667),
.Y(n_962)
);

INVx1_ASAP7_75t_SL g963 ( 
.A(n_624),
.Y(n_963)
);

CKINVDCx16_ASAP7_75t_R g964 ( 
.A(n_689),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_712),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_716),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_720),
.B(n_551),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_724),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_726),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_728),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_763),
.B(n_288),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_658),
.B(n_551),
.Y(n_972)
);

NAND2x1p5_ASAP7_75t_L g973 ( 
.A(n_620),
.B(n_531),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_668),
.B(n_291),
.Y(n_974)
);

OR2x2_ASAP7_75t_L g975 ( 
.A(n_816),
.B(n_673),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_786),
.B(n_678),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_833),
.B(n_679),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_849),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_933),
.B(n_731),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_849),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_849),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_835),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_880),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_830),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_933),
.B(n_669),
.Y(n_985)
);

HB1xp67_ASAP7_75t_L g986 ( 
.A(n_788),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_793),
.B(n_639),
.Y(n_987)
);

AND3x2_ASAP7_75t_SL g988 ( 
.A(n_961),
.B(n_706),
.C(n_771),
.Y(n_988)
);

INVx2_ASAP7_75t_SL g989 ( 
.A(n_827),
.Y(n_989)
);

AOI221xp5_ASAP7_75t_L g990 ( 
.A1(n_904),
.A2(n_640),
.B1(n_231),
.B2(n_246),
.C(n_252),
.Y(n_990)
);

NAND2x1_ASAP7_75t_L g991 ( 
.A(n_903),
.B(n_738),
.Y(n_991)
);

BUFx3_ASAP7_75t_L g992 ( 
.A(n_791),
.Y(n_992)
);

OAI21xp33_ASAP7_75t_L g993 ( 
.A1(n_912),
.A2(n_669),
.B(n_261),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_810),
.A2(n_665),
.B(n_646),
.Y(n_994)
);

OR2x6_ASAP7_75t_L g995 ( 
.A(n_800),
.B(n_714),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_884),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_866),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_833),
.B(n_699),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_838),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_940),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_814),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_880),
.Y(n_1002)
);

AOI22xp33_ASAP7_75t_L g1003 ( 
.A1(n_946),
.A2(n_670),
.B1(n_753),
.B2(n_734),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_933),
.B(n_740),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_834),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_831),
.B(n_699),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_880),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_782),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_933),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_817),
.B(n_784),
.Y(n_1010)
);

AOI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_821),
.A2(n_665),
.B1(n_664),
.B2(n_646),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_845),
.Y(n_1012)
);

HB1xp67_ASAP7_75t_L g1013 ( 
.A(n_811),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_901),
.B(n_910),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_898),
.B(n_664),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_797),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_862),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_795),
.B(n_742),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_839),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_831),
.B(n_699),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_920),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_945),
.Y(n_1022)
);

NAND2xp33_ASAP7_75t_L g1023 ( 
.A(n_901),
.B(n_643),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_917),
.B(n_697),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_901),
.B(n_643),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_869),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_945),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_910),
.B(n_659),
.Y(n_1028)
);

INVx1_ASAP7_75t_SL g1029 ( 
.A(n_947),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_945),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_790),
.Y(n_1031)
);

CKINVDCx20_ASAP7_75t_R g1032 ( 
.A(n_807),
.Y(n_1032)
);

AOI22x1_ASAP7_75t_L g1033 ( 
.A1(n_826),
.A2(n_659),
.B1(n_778),
.B2(n_776),
.Y(n_1033)
);

HB1xp67_ASAP7_75t_L g1034 ( 
.A(n_824),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_861),
.Y(n_1035)
);

BUFx12f_ASAP7_75t_L g1036 ( 
.A(n_847),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_871),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_889),
.Y(n_1038)
);

BUFx12f_ASAP7_75t_L g1039 ( 
.A(n_949),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_910),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_917),
.B(n_697),
.Y(n_1041)
);

NOR2x1p5_ASAP7_75t_L g1042 ( 
.A(n_794),
.B(n_727),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_923),
.B(n_622),
.Y(n_1043)
);

AND2x6_ASAP7_75t_L g1044 ( 
.A(n_856),
.B(n_727),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_906),
.Y(n_1045)
);

INVx4_ASAP7_75t_L g1046 ( 
.A(n_930),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_930),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_923),
.B(n_626),
.Y(n_1048)
);

BUFx3_ASAP7_75t_L g1049 ( 
.A(n_902),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_925),
.B(n_630),
.Y(n_1050)
);

INVx1_ASAP7_75t_SL g1051 ( 
.A(n_947),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_865),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_925),
.B(n_633),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_863),
.A2(n_734),
.B1(n_779),
.B2(n_736),
.Y(n_1054)
);

AND2x4_ASAP7_75t_L g1055 ( 
.A(n_832),
.B(n_779),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_885),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_926),
.B(n_635),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_941),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_893),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_931),
.Y(n_1060)
);

INVx4_ASAP7_75t_L g1061 ( 
.A(n_930),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_936),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_926),
.B(n_650),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_929),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_928),
.B(n_736),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_887),
.A2(n_744),
.B1(n_640),
.B2(n_739),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_928),
.B(n_744),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_938),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_889),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_972),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_850),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_944),
.B(n_780),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_873),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_919),
.Y(n_1074)
);

INVx4_ASAP7_75t_L g1075 ( 
.A(n_806),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_944),
.B(n_761),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_810),
.B(n_761),
.Y(n_1077)
);

BUFx4f_ASAP7_75t_L g1078 ( 
.A(n_877),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_881),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_844),
.B(n_764),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_844),
.B(n_764),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_806),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_812),
.B(n_587),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_820),
.A2(n_561),
.B(n_575),
.C(n_597),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_812),
.B(n_579),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_929),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_803),
.B(n_223),
.Y(n_1087)
);

BUFx12f_ASAP7_75t_L g1088 ( 
.A(n_949),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_892),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_R g1090 ( 
.A(n_813),
.B(n_837),
.Y(n_1090)
);

INVx3_ASAP7_75t_SL g1091 ( 
.A(n_937),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_897),
.Y(n_1092)
);

AOI211xp5_ASAP7_75t_L g1093 ( 
.A1(n_904),
.A2(n_264),
.B(n_272),
.C(n_291),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_852),
.B(n_590),
.Y(n_1094)
);

INVx4_ASAP7_75t_L g1095 ( 
.A(n_808),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_888),
.B(n_310),
.Y(n_1096)
);

INVxp67_ASAP7_75t_SL g1097 ( 
.A(n_792),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_896),
.B(n_561),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_896),
.B(n_576),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_841),
.B(n_576),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_935),
.Y(n_1101)
);

INVx3_ASAP7_75t_L g1102 ( 
.A(n_808),
.Y(n_1102)
);

INVxp67_ASAP7_75t_SL g1103 ( 
.A(n_851),
.Y(n_1103)
);

BUFx8_ASAP7_75t_L g1104 ( 
.A(n_916),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_852),
.B(n_590),
.Y(n_1105)
);

AO22x1_ASAP7_75t_L g1106 ( 
.A1(n_963),
.A2(n_297),
.B1(n_300),
.B2(n_301),
.Y(n_1106)
);

HB1xp67_ASAP7_75t_L g1107 ( 
.A(n_850),
.Y(n_1107)
);

AND2x4_ASAP7_75t_L g1108 ( 
.A(n_957),
.B(n_587),
.Y(n_1108)
);

NAND2xp33_ASAP7_75t_L g1109 ( 
.A(n_840),
.B(n_768),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_857),
.A2(n_579),
.B(n_300),
.C(n_301),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_948),
.B(n_768),
.Y(n_1111)
);

OR2x2_ASAP7_75t_L g1112 ( 
.A(n_846),
.B(n_434),
.Y(n_1112)
);

HB1xp67_ASAP7_75t_L g1113 ( 
.A(n_874),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_900),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_867),
.Y(n_1115)
);

BUFx8_ASAP7_75t_SL g1116 ( 
.A(n_962),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_948),
.B(n_439),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_932),
.B(n_439),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_962),
.B(n_308),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_958),
.B(n_605),
.Y(n_1120)
);

BUFx4f_ASAP7_75t_L g1121 ( 
.A(n_867),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_911),
.B(n_65),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_935),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_958),
.B(n_858),
.Y(n_1124)
);

NOR2xp67_ASAP7_75t_L g1125 ( 
.A(n_974),
.B(n_306),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_860),
.B(n_605),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_878),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_984),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1017),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_1029),
.Y(n_1130)
);

INVx2_ASAP7_75t_SL g1131 ( 
.A(n_1001),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_1009),
.Y(n_1132)
);

OR2x2_ASAP7_75t_L g1133 ( 
.A(n_1029),
.B(n_964),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_1026),
.Y(n_1134)
);

AND2x2_ASAP7_75t_SL g1135 ( 
.A(n_1078),
.B(n_864),
.Y(n_1135)
);

OAI221xp5_ASAP7_75t_L g1136 ( 
.A1(n_1093),
.A2(n_990),
.B1(n_993),
.B2(n_908),
.C(n_987),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1045),
.B(n_963),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1037),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1124),
.A2(n_792),
.B(n_953),
.Y(n_1139)
);

CKINVDCx11_ASAP7_75t_R g1140 ( 
.A(n_1032),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_1011),
.A2(n_959),
.B(n_883),
.C(n_971),
.Y(n_1141)
);

BUFx4f_ASAP7_75t_SL g1142 ( 
.A(n_1039),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1079),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_1022),
.Y(n_1144)
);

O2A1O1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_976),
.A2(n_872),
.B(n_907),
.C(n_922),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_998),
.B(n_918),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1005),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_1009),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1089),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_1022),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1124),
.A2(n_955),
.B(n_994),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_1022),
.Y(n_1152)
);

BUFx12f_ASAP7_75t_L g1153 ( 
.A(n_1088),
.Y(n_1153)
);

CKINVDCx20_ASAP7_75t_R g1154 ( 
.A(n_992),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_1027),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1058),
.B(n_819),
.Y(n_1156)
);

INVx3_ASAP7_75t_L g1157 ( 
.A(n_1006),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1092),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1114),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1071),
.B(n_934),
.Y(n_1160)
);

INVxp67_ASAP7_75t_L g1161 ( 
.A(n_1012),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1010),
.B(n_878),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1010),
.B(n_785),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1060),
.B(n_796),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1008),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_990),
.A2(n_848),
.B1(n_823),
.B2(n_815),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1016),
.Y(n_1167)
);

AOI33xp33_ASAP7_75t_L g1168 ( 
.A1(n_1087),
.A2(n_968),
.A3(n_966),
.B1(n_927),
.B2(n_921),
.B3(n_960),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1019),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_996),
.Y(n_1170)
);

INVxp67_ASAP7_75t_SL g1171 ( 
.A(n_986),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1051),
.B(n_842),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_1000),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1035),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1052),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1056),
.Y(n_1176)
);

BUFx2_ASAP7_75t_SL g1177 ( 
.A(n_989),
.Y(n_1177)
);

NAND2x1p5_ASAP7_75t_L g1178 ( 
.A(n_1046),
.B(n_840),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_1107),
.A2(n_801),
.B1(n_818),
.B2(n_942),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_975),
.B(n_942),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1059),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_999),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_1051),
.Y(n_1183)
);

AOI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1015),
.A2(n_825),
.B1(n_804),
.B2(n_854),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1112),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_976),
.A2(n_855),
.B1(n_840),
.B2(n_891),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_982),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_994),
.A2(n_851),
.B(n_868),
.Y(n_1188)
);

NOR2x1_ASAP7_75t_R g1189 ( 
.A(n_1036),
.B(n_859),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_1021),
.B(n_840),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_998),
.B(n_787),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_1027),
.Y(n_1192)
);

AND2x6_ASAP7_75t_L g1193 ( 
.A(n_1006),
.B(n_783),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_997),
.B(n_915),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1064),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1018),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_1013),
.B(n_805),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1062),
.B(n_909),
.Y(n_1198)
);

AOI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1100),
.A2(n_829),
.B(n_783),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1125),
.A2(n_977),
.B1(n_1042),
.B2(n_1055),
.Y(n_1200)
);

INVx8_ASAP7_75t_L g1201 ( 
.A(n_1020),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1086),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_1034),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_1020),
.Y(n_1204)
);

BUFx2_ASAP7_75t_L g1205 ( 
.A(n_1104),
.Y(n_1205)
);

BUFx3_ASAP7_75t_L g1206 ( 
.A(n_1104),
.Y(n_1206)
);

AND2x4_ASAP7_75t_L g1207 ( 
.A(n_977),
.B(n_939),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1101),
.Y(n_1208)
);

OAI211xp5_ASAP7_75t_L g1209 ( 
.A1(n_1096),
.A2(n_853),
.B(n_950),
.C(n_951),
.Y(n_1209)
);

INVx3_ASAP7_75t_L g1210 ( 
.A(n_1038),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1123),
.Y(n_1211)
);

AOI221xp5_ASAP7_75t_L g1212 ( 
.A1(n_1106),
.A2(n_306),
.B1(n_307),
.B2(n_969),
.C(n_970),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1103),
.A2(n_855),
.B1(n_891),
.B2(n_903),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1055),
.A2(n_952),
.B1(n_965),
.B2(n_956),
.Y(n_1214)
);

AOI221xp5_ASAP7_75t_L g1215 ( 
.A1(n_1054),
.A2(n_307),
.B1(n_954),
.B2(n_913),
.C(n_943),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1118),
.B(n_828),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1038),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1069),
.Y(n_1218)
);

BUFx8_ASAP7_75t_L g1219 ( 
.A(n_1074),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_1090),
.Y(n_1220)
);

BUFx12f_ASAP7_75t_L g1221 ( 
.A(n_1074),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1113),
.B(n_924),
.Y(n_1222)
);

INVx1_ASAP7_75t_SL g1223 ( 
.A(n_1091),
.Y(n_1223)
);

OAI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1103),
.A2(n_891),
.B1(n_855),
.B2(n_868),
.Y(n_1224)
);

OR2x2_ASAP7_75t_L g1225 ( 
.A(n_1073),
.B(n_967),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_1027),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1030),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1069),
.A2(n_843),
.B1(n_895),
.B2(n_891),
.Y(n_1228)
);

A2O1A1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_1110),
.A2(n_875),
.B(n_886),
.C(n_882),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1094),
.B(n_967),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1080),
.A2(n_895),
.B1(n_855),
.B2(n_879),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1083),
.Y(n_1232)
);

AOI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1054),
.A2(n_870),
.B1(n_879),
.B2(n_890),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1082),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_1074),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1023),
.A2(n_799),
.B(n_798),
.Y(n_1236)
);

OAI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1078),
.A2(n_894),
.B1(n_799),
.B2(n_798),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1120),
.A2(n_870),
.B(n_890),
.Y(n_1238)
);

BUFx4_ASAP7_75t_SL g1239 ( 
.A(n_1031),
.Y(n_1239)
);

INVx5_ASAP7_75t_L g1240 ( 
.A(n_980),
.Y(n_1240)
);

AOI21xp33_ASAP7_75t_L g1241 ( 
.A1(n_1066),
.A2(n_899),
.B(n_914),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1049),
.B(n_836),
.Y(n_1242)
);

AOI221xp5_ASAP7_75t_L g1243 ( 
.A1(n_1066),
.A2(n_789),
.B1(n_894),
.B2(n_809),
.C(n_802),
.Y(n_1243)
);

AOI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1068),
.A2(n_905),
.B1(n_789),
.B2(n_809),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1083),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1085),
.Y(n_1246)
);

AND2x6_ASAP7_75t_L g1247 ( 
.A(n_1122),
.B(n_802),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_1082),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_995),
.B(n_822),
.Y(n_1249)
);

INVx2_ASAP7_75t_SL g1250 ( 
.A(n_1030),
.Y(n_1250)
);

AOI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1070),
.A2(n_1081),
.B1(n_1122),
.B2(n_1044),
.Y(n_1251)
);

BUFx2_ASAP7_75t_L g1252 ( 
.A(n_1116),
.Y(n_1252)
);

NAND3xp33_ASAP7_75t_L g1253 ( 
.A(n_1003),
.B(n_531),
.C(n_3),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1120),
.A2(n_876),
.B(n_973),
.Y(n_1254)
);

NOR2xp67_ASAP7_75t_L g1255 ( 
.A(n_1046),
.B(n_66),
.Y(n_1255)
);

OR2x2_ASAP7_75t_L g1256 ( 
.A(n_1094),
.B(n_973),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1024),
.B(n_822),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_SL g1258 ( 
.A(n_1061),
.B(n_822),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_1030),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1085),
.Y(n_1260)
);

BUFx2_ASAP7_75t_L g1261 ( 
.A(n_980),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1109),
.A2(n_876),
.B(n_605),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_980),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_981),
.Y(n_1264)
);

OR2x6_ASAP7_75t_L g1265 ( 
.A(n_995),
.B(n_605),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_SL g1266 ( 
.A1(n_1097),
.A2(n_822),
.B1(n_9),
.B2(n_11),
.Y(n_1266)
);

AND2x4_ASAP7_75t_L g1267 ( 
.A(n_995),
.B(n_60),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1044),
.A2(n_531),
.B1(n_12),
.B2(n_13),
.Y(n_1268)
);

A2O1A1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1077),
.A2(n_0),
.B(n_14),
.C(n_15),
.Y(n_1269)
);

INVx4_ASAP7_75t_L g1270 ( 
.A(n_1040),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_1061),
.B(n_148),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1108),
.Y(n_1272)
);

O2A1O1Ixp5_ASAP7_75t_SL g1273 ( 
.A1(n_1119),
.A2(n_1100),
.B(n_1014),
.C(n_1025),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1108),
.Y(n_1274)
);

BUFx3_ASAP7_75t_L g1275 ( 
.A(n_981),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1024),
.B(n_0),
.Y(n_1276)
);

BUFx8_ASAP7_75t_SL g1277 ( 
.A(n_1040),
.Y(n_1277)
);

OR2x2_ASAP7_75t_L g1278 ( 
.A(n_1105),
.B(n_15),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1041),
.B(n_16),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1065),
.A2(n_70),
.B(n_144),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_SL g1281 ( 
.A1(n_988),
.A2(n_16),
.B1(n_18),
.B2(n_24),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1102),
.Y(n_1282)
);

A2O1A1Ixp33_ASAP7_75t_L g1283 ( 
.A1(n_1253),
.A2(n_1136),
.B(n_1241),
.C(n_1229),
.Y(n_1283)
);

NOR2x1_ASAP7_75t_SL g1284 ( 
.A(n_1253),
.B(n_1028),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1129),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1137),
.B(n_1077),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_1249),
.B(n_1105),
.Y(n_1287)
);

OA21x2_ASAP7_75t_L g1288 ( 
.A1(n_1241),
.A2(n_1084),
.B(n_1117),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1160),
.B(n_1040),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_1201),
.Y(n_1290)
);

AO21x2_ASAP7_75t_L g1291 ( 
.A1(n_1151),
.A2(n_1117),
.B(n_1098),
.Y(n_1291)
);

OR2x2_ASAP7_75t_L g1292 ( 
.A(n_1133),
.B(n_978),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1188),
.A2(n_1033),
.B(n_1098),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1134),
.Y(n_1294)
);

INVx3_ASAP7_75t_L g1295 ( 
.A(n_1201),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1254),
.A2(n_1099),
.B(n_1072),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1238),
.A2(n_1099),
.B(n_1072),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1236),
.A2(n_1053),
.B(n_1050),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1128),
.Y(n_1299)
);

BUFx6f_ASAP7_75t_L g1300 ( 
.A(n_1201),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1251),
.A2(n_1121),
.B1(n_985),
.B2(n_1065),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1138),
.Y(n_1302)
);

A2O1A1Ixp33_ASAP7_75t_L g1303 ( 
.A1(n_1145),
.A2(n_1067),
.B(n_1041),
.C(n_1076),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1199),
.A2(n_1053),
.B(n_1063),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1158),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_1140),
.Y(n_1306)
);

NAND3xp33_ASAP7_75t_L g1307 ( 
.A(n_1269),
.B(n_1047),
.C(n_979),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1156),
.B(n_978),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1143),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1251),
.A2(n_1121),
.B1(n_1067),
.B2(n_979),
.Y(n_1310)
);

OA21x2_ASAP7_75t_L g1311 ( 
.A1(n_1141),
.A2(n_1057),
.B(n_1050),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1139),
.A2(n_1048),
.B(n_1057),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1149),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1159),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1182),
.Y(n_1315)
);

AND2x4_ASAP7_75t_L g1316 ( 
.A(n_1249),
.B(n_1102),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1273),
.A2(n_1063),
.B(n_1043),
.Y(n_1317)
);

BUFx6f_ASAP7_75t_L g1318 ( 
.A(n_1240),
.Y(n_1318)
);

INVx4_ASAP7_75t_L g1319 ( 
.A(n_1240),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1167),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1232),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1180),
.B(n_1047),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1213),
.A2(n_1224),
.B(n_1186),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1213),
.A2(n_1048),
.B(n_1043),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1174),
.Y(n_1325)
);

AO21x2_ASAP7_75t_L g1326 ( 
.A1(n_1237),
.A2(n_1111),
.B(n_1076),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1175),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1200),
.A2(n_1004),
.B1(n_1047),
.B2(n_1126),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1224),
.A2(n_991),
.B(n_1111),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1172),
.B(n_1216),
.Y(n_1330)
);

NOR2xp67_ASAP7_75t_SL g1331 ( 
.A(n_1153),
.B(n_981),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1245),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_SL g1333 ( 
.A1(n_1276),
.A2(n_1279),
.B(n_1184),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1187),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1186),
.A2(n_1126),
.B(n_1004),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1262),
.A2(n_1075),
.B(n_1095),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1246),
.Y(n_1337)
);

AOI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1276),
.A2(n_1044),
.B(n_988),
.Y(n_1338)
);

BUFx2_ASAP7_75t_L g1339 ( 
.A(n_1173),
.Y(n_1339)
);

NOR2xp67_ASAP7_75t_L g1340 ( 
.A(n_1220),
.B(n_1161),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_1277),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1260),
.Y(n_1342)
);

AND2x4_ASAP7_75t_L g1343 ( 
.A(n_1265),
.B(n_1002),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1183),
.B(n_1127),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1257),
.A2(n_1002),
.B(n_1007),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1163),
.A2(n_1075),
.B(n_1095),
.Y(n_1346)
);

OR2x2_ASAP7_75t_L g1347 ( 
.A(n_1130),
.B(n_1007),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1202),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1257),
.A2(n_1044),
.B(n_1115),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1165),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1208),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1169),
.Y(n_1352)
);

AOI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1222),
.A2(n_1127),
.B1(n_1115),
.B2(n_1082),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1176),
.Y(n_1354)
);

INVx3_ASAP7_75t_L g1355 ( 
.A(n_1157),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1170),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1185),
.B(n_1127),
.Y(n_1357)
);

OAI222xp33_ASAP7_75t_L g1358 ( 
.A1(n_1268),
.A2(n_18),
.B1(n_25),
.B2(n_26),
.C1(n_29),
.C2(n_34),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1281),
.A2(n_1115),
.B1(n_983),
.B2(n_39),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1225),
.Y(n_1360)
);

INVxp67_ASAP7_75t_SL g1361 ( 
.A(n_1162),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1243),
.A2(n_1280),
.B(n_1233),
.Y(n_1362)
);

AND2x4_ASAP7_75t_L g1363 ( 
.A(n_1265),
.B(n_983),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1198),
.Y(n_1364)
);

CKINVDCx12_ASAP7_75t_R g1365 ( 
.A(n_1189),
.Y(n_1365)
);

AND2x4_ASAP7_75t_L g1366 ( 
.A(n_1265),
.B(n_983),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1171),
.B(n_35),
.Y(n_1367)
);

O2A1O1Ixp5_ASAP7_75t_L g1368 ( 
.A1(n_1209),
.A2(n_38),
.B(n_44),
.C(n_45),
.Y(n_1368)
);

CKINVDCx14_ASAP7_75t_R g1369 ( 
.A(n_1252),
.Y(n_1369)
);

INVx1_ASAP7_75t_SL g1370 ( 
.A(n_1223),
.Y(n_1370)
);

CKINVDCx20_ASAP7_75t_R g1371 ( 
.A(n_1219),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1281),
.A2(n_1266),
.B1(n_1279),
.B2(n_1196),
.Y(n_1372)
);

AO21x2_ASAP7_75t_L g1373 ( 
.A1(n_1233),
.A2(n_1184),
.B(n_1162),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1181),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1198),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1244),
.A2(n_1231),
.B(n_1228),
.Y(n_1376)
);

OA21x2_ASAP7_75t_L g1377 ( 
.A1(n_1215),
.A2(n_38),
.B(n_55),
.Y(n_1377)
);

AO21x2_ASAP7_75t_L g1378 ( 
.A1(n_1244),
.A2(n_67),
.B(n_72),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1163),
.A2(n_145),
.B(n_89),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1147),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1166),
.A2(n_74),
.B(n_95),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1132),
.A2(n_104),
.B(n_108),
.Y(n_1382)
);

AO21x2_ASAP7_75t_L g1383 ( 
.A1(n_1190),
.A2(n_118),
.B(n_122),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1164),
.Y(n_1384)
);

AOI211xp5_ASAP7_75t_L g1385 ( 
.A1(n_1197),
.A2(n_124),
.B(n_131),
.C(n_141),
.Y(n_1385)
);

BUFx8_ASAP7_75t_L g1386 ( 
.A(n_1205),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1164),
.Y(n_1387)
);

AO31x2_ASAP7_75t_L g1388 ( 
.A1(n_1282),
.A2(n_1217),
.A3(n_1218),
.B(n_1274),
.Y(n_1388)
);

INVx2_ASAP7_75t_SL g1389 ( 
.A(n_1219),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1230),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1207),
.B(n_1168),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1132),
.A2(n_1148),
.B(n_1210),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1148),
.A2(n_1210),
.B(n_1178),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1195),
.Y(n_1394)
);

O2A1O1Ixp33_ASAP7_75t_SL g1395 ( 
.A1(n_1256),
.A2(n_1212),
.B(n_1272),
.C(n_1278),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1211),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1207),
.B(n_1203),
.Y(n_1397)
);

OR2x6_ASAP7_75t_L g1398 ( 
.A(n_1267),
.B(n_1221),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1214),
.A2(n_1255),
.B(n_1179),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1194),
.B(n_1146),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1146),
.B(n_1242),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1255),
.A2(n_1248),
.B(n_1234),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_1154),
.B(n_1191),
.Y(n_1403)
);

OR2x6_ASAP7_75t_L g1404 ( 
.A(n_1267),
.B(n_1177),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1193),
.Y(n_1405)
);

BUFx6f_ASAP7_75t_L g1406 ( 
.A(n_1240),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1234),
.A2(n_1248),
.B(n_1204),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1135),
.B(n_1157),
.Y(n_1408)
);

OAI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1247),
.A2(n_1193),
.B(n_1191),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1204),
.A2(n_1193),
.B(n_1247),
.Y(n_1410)
);

INVx1_ASAP7_75t_SL g1411 ( 
.A(n_1223),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1263),
.Y(n_1412)
);

INVx3_ASAP7_75t_L g1413 ( 
.A(n_1270),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1247),
.A2(n_1193),
.B1(n_1271),
.B2(n_1206),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1235),
.A2(n_1250),
.B1(n_1261),
.B2(n_1131),
.Y(n_1415)
);

AOI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1271),
.A2(n_1247),
.B(n_1258),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1258),
.A2(n_1189),
.B(n_1270),
.Y(n_1417)
);

NAND2x1_ASAP7_75t_L g1418 ( 
.A(n_1263),
.B(n_1264),
.Y(n_1418)
);

O2A1O1Ixp33_ASAP7_75t_SL g1419 ( 
.A1(n_1263),
.A2(n_1264),
.B(n_1144),
.C(n_1150),
.Y(n_1419)
);

OA21x2_ASAP7_75t_L g1420 ( 
.A1(n_1264),
.A2(n_1192),
.B(n_1144),
.Y(n_1420)
);

AO21x2_ASAP7_75t_L g1421 ( 
.A1(n_1144),
.A2(n_1226),
.B(n_1150),
.Y(n_1421)
);

BUFx3_ASAP7_75t_L g1422 ( 
.A(n_1142),
.Y(n_1422)
);

OAI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1275),
.A2(n_1239),
.B(n_1152),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1150),
.A2(n_1152),
.B(n_1155),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1152),
.A2(n_1155),
.B(n_1192),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1259),
.B(n_1155),
.Y(n_1426)
);

NAND2x1p5_ASAP7_75t_L g1427 ( 
.A(n_1192),
.B(n_1259),
.Y(n_1427)
);

INVx3_ASAP7_75t_L g1428 ( 
.A(n_1226),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1259),
.A2(n_1226),
.B(n_1227),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1227),
.B(n_1137),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1390),
.B(n_1227),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1359),
.A2(n_1372),
.B1(n_1283),
.B2(n_1398),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1361),
.B(n_1364),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1390),
.B(n_1401),
.Y(n_1434)
);

INVxp33_ASAP7_75t_L g1435 ( 
.A(n_1403),
.Y(n_1435)
);

OA21x2_ASAP7_75t_L g1436 ( 
.A1(n_1293),
.A2(n_1323),
.B(n_1317),
.Y(n_1436)
);

INVx4_ASAP7_75t_L g1437 ( 
.A(n_1318),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_SL g1438 ( 
.A1(n_1381),
.A2(n_1284),
.B1(n_1377),
.B2(n_1362),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_1318),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1330),
.B(n_1430),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1360),
.B(n_1292),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1359),
.A2(n_1372),
.B1(n_1333),
.B2(n_1391),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1361),
.B(n_1375),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1294),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1299),
.Y(n_1445)
);

OR2x6_ASAP7_75t_L g1446 ( 
.A(n_1409),
.B(n_1416),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1400),
.B(n_1289),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1302),
.Y(n_1448)
);

INVx1_ASAP7_75t_SL g1449 ( 
.A(n_1347),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1309),
.Y(n_1450)
);

INVx4_ASAP7_75t_L g1451 ( 
.A(n_1318),
.Y(n_1451)
);

INVx6_ASAP7_75t_L g1452 ( 
.A(n_1386),
.Y(n_1452)
);

INVx4_ASAP7_75t_L g1453 ( 
.A(n_1318),
.Y(n_1453)
);

INVx4_ASAP7_75t_L g1454 ( 
.A(n_1406),
.Y(n_1454)
);

OR2x6_ASAP7_75t_L g1455 ( 
.A(n_1410),
.B(n_1405),
.Y(n_1455)
);

OAI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1283),
.A2(n_1303),
.B(n_1368),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1294),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1313),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_SL g1459 ( 
.A1(n_1377),
.A2(n_1378),
.B1(n_1301),
.B2(n_1408),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1384),
.B(n_1387),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1310),
.A2(n_1398),
.B1(n_1308),
.B2(n_1403),
.Y(n_1461)
);

NAND2xp33_ASAP7_75t_R g1462 ( 
.A(n_1306),
.B(n_1398),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1305),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1305),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1350),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1315),
.Y(n_1466)
);

BUFx12f_ASAP7_75t_L g1467 ( 
.A(n_1306),
.Y(n_1467)
);

BUFx10_ASAP7_75t_L g1468 ( 
.A(n_1344),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1320),
.Y(n_1469)
);

AND2x4_ASAP7_75t_L g1470 ( 
.A(n_1343),
.B(n_1363),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1378),
.A2(n_1339),
.B1(n_1377),
.B2(n_1373),
.Y(n_1471)
);

OR2x6_ASAP7_75t_L g1472 ( 
.A(n_1410),
.B(n_1405),
.Y(n_1472)
);

INVx2_ASAP7_75t_SL g1473 ( 
.A(n_1356),
.Y(n_1473)
);

AO21x2_ASAP7_75t_L g1474 ( 
.A1(n_1293),
.A2(n_1303),
.B(n_1317),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1350),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_1371),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_SL g1477 ( 
.A1(n_1404),
.A2(n_1373),
.B1(n_1399),
.B2(n_1379),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_L g1478 ( 
.A(n_1406),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1321),
.B(n_1332),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1357),
.B(n_1286),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1352),
.Y(n_1481)
);

BUFx12f_ASAP7_75t_L g1482 ( 
.A(n_1386),
.Y(n_1482)
);

AOI221xp5_ASAP7_75t_L g1483 ( 
.A1(n_1358),
.A2(n_1395),
.B1(n_1368),
.B2(n_1385),
.C(n_1411),
.Y(n_1483)
);

INVx4_ASAP7_75t_SL g1484 ( 
.A(n_1422),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1325),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1322),
.B(n_1287),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1307),
.A2(n_1404),
.B1(n_1287),
.B2(n_1370),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1404),
.A2(n_1287),
.B1(n_1328),
.B2(n_1414),
.Y(n_1488)
);

AOI21xp33_ASAP7_75t_L g1489 ( 
.A1(n_1326),
.A2(n_1311),
.B(n_1376),
.Y(n_1489)
);

AOI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1395),
.A2(n_1365),
.B1(n_1371),
.B2(n_1397),
.Y(n_1490)
);

NOR2x1_ASAP7_75t_R g1491 ( 
.A(n_1422),
.B(n_1341),
.Y(n_1491)
);

AOI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1336),
.A2(n_1346),
.B(n_1311),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1327),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1344),
.B(n_1352),
.Y(n_1494)
);

OAI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1353),
.A2(n_1356),
.B1(n_1340),
.B2(n_1338),
.Y(n_1495)
);

OR2x6_ASAP7_75t_L g1496 ( 
.A(n_1349),
.B(n_1323),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1285),
.B(n_1314),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1348),
.B(n_1351),
.Y(n_1498)
);

CKINVDCx11_ASAP7_75t_R g1499 ( 
.A(n_1341),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1334),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_SL g1501 ( 
.A1(n_1399),
.A2(n_1376),
.B1(n_1383),
.B2(n_1386),
.Y(n_1501)
);

OAI211xp5_ASAP7_75t_L g1502 ( 
.A1(n_1367),
.A2(n_1414),
.B(n_1396),
.C(n_1394),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_L g1503 ( 
.A(n_1369),
.B(n_1316),
.Y(n_1503)
);

CKINVDCx9p33_ASAP7_75t_R g1504 ( 
.A(n_1426),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1354),
.Y(n_1505)
);

AOI221xp5_ASAP7_75t_L g1506 ( 
.A1(n_1415),
.A2(n_1380),
.B1(n_1331),
.B2(n_1321),
.C(n_1342),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1354),
.B(n_1374),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1332),
.B(n_1337),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1374),
.B(n_1316),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1337),
.B(n_1342),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1388),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1369),
.A2(n_1389),
.B1(n_1406),
.B2(n_1311),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1316),
.B(n_1355),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1345),
.Y(n_1514)
);

INVx4_ASAP7_75t_L g1515 ( 
.A(n_1406),
.Y(n_1515)
);

BUFx2_ASAP7_75t_L g1516 ( 
.A(n_1420),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1355),
.A2(n_1363),
.B1(n_1366),
.B2(n_1319),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1412),
.B(n_1295),
.Y(n_1518)
);

BUFx8_ASAP7_75t_L g1519 ( 
.A(n_1290),
.Y(n_1519)
);

INVx3_ASAP7_75t_L g1520 ( 
.A(n_1290),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1363),
.A2(n_1366),
.B1(n_1319),
.B2(n_1423),
.Y(n_1521)
);

AND2x4_ASAP7_75t_L g1522 ( 
.A(n_1343),
.B(n_1366),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1388),
.B(n_1428),
.Y(n_1523)
);

OAI21x1_ASAP7_75t_L g1524 ( 
.A1(n_1329),
.A2(n_1296),
.B(n_1335),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1388),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1407),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1428),
.Y(n_1527)
);

OR2x6_ASAP7_75t_L g1528 ( 
.A(n_1329),
.B(n_1335),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1383),
.A2(n_1343),
.B1(n_1326),
.B2(n_1300),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_SL g1530 ( 
.A1(n_1417),
.A2(n_1382),
.B1(n_1290),
.B2(n_1300),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1421),
.B(n_1420),
.Y(n_1531)
);

NAND3xp33_ASAP7_75t_SL g1532 ( 
.A(n_1418),
.B(n_1427),
.C(n_1382),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1304),
.B(n_1324),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1421),
.B(n_1420),
.Y(n_1534)
);

A2O1A1Ixp33_ASAP7_75t_L g1535 ( 
.A1(n_1312),
.A2(n_1324),
.B(n_1298),
.C(n_1297),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1297),
.B(n_1296),
.Y(n_1536)
);

OAI21x1_ASAP7_75t_L g1537 ( 
.A1(n_1298),
.A2(n_1304),
.B(n_1392),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1295),
.B(n_1427),
.Y(n_1538)
);

OAI21xp33_ASAP7_75t_L g1539 ( 
.A1(n_1413),
.A2(n_1402),
.B(n_1290),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1300),
.A2(n_1413),
.B1(n_1291),
.B2(n_1288),
.Y(n_1540)
);

INVxp67_ASAP7_75t_L g1541 ( 
.A(n_1424),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1392),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1300),
.A2(n_1291),
.B1(n_1288),
.B2(n_1393),
.Y(n_1543)
);

OAI221xp5_ASAP7_75t_L g1544 ( 
.A1(n_1288),
.A2(n_1419),
.B1(n_1393),
.B2(n_1425),
.C(n_1429),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1419),
.B(n_1429),
.Y(n_1545)
);

OAI21x1_ASAP7_75t_L g1546 ( 
.A1(n_1293),
.A2(n_1329),
.B(n_1296),
.Y(n_1546)
);

CKINVDCx8_ASAP7_75t_R g1547 ( 
.A(n_1306),
.Y(n_1547)
);

INVx3_ASAP7_75t_L g1548 ( 
.A(n_1290),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1390),
.B(n_1401),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1294),
.Y(n_1550)
);

O2A1O1Ixp33_ASAP7_75t_L g1551 ( 
.A1(n_1283),
.A2(n_629),
.B(n_653),
.C(n_1136),
.Y(n_1551)
);

OR2x6_ASAP7_75t_L g1552 ( 
.A(n_1409),
.B(n_1416),
.Y(n_1552)
);

CKINVDCx16_ASAP7_75t_R g1553 ( 
.A(n_1467),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1432),
.A2(n_1442),
.B1(n_1456),
.B2(n_1483),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_1499),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1433),
.B(n_1443),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1498),
.Y(n_1557)
);

NOR2x1_ASAP7_75t_L g1558 ( 
.A(n_1532),
.B(n_1495),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_1523),
.B(n_1449),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1480),
.B(n_1440),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1551),
.A2(n_1456),
.B(n_1483),
.Y(n_1561)
);

O2A1O1Ixp33_ASAP7_75t_L g1562 ( 
.A1(n_1432),
.A2(n_1502),
.B(n_1512),
.C(n_1471),
.Y(n_1562)
);

OR2x6_ASAP7_75t_L g1563 ( 
.A(n_1446),
.B(n_1552),
.Y(n_1563)
);

CKINVDCx16_ASAP7_75t_R g1564 ( 
.A(n_1482),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1461),
.A2(n_1490),
.B1(n_1438),
.B2(n_1435),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1497),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_R g1567 ( 
.A(n_1476),
.B(n_1547),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_R g1568 ( 
.A(n_1462),
.B(n_1452),
.Y(n_1568)
);

NOR2x1p5_ASAP7_75t_L g1569 ( 
.A(n_1520),
.B(n_1548),
.Y(n_1569)
);

NAND2xp33_ASAP7_75t_R g1570 ( 
.A(n_1520),
.B(n_1548),
.Y(n_1570)
);

OAI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1490),
.A2(n_1487),
.B1(n_1488),
.B2(n_1452),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_R g1572 ( 
.A(n_1519),
.B(n_1473),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1434),
.B(n_1549),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1447),
.B(n_1486),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_SL g1575 ( 
.A1(n_1512),
.A2(n_1521),
.B1(n_1552),
.B2(n_1446),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1445),
.Y(n_1576)
);

AND2x4_ASAP7_75t_SL g1577 ( 
.A(n_1468),
.B(n_1494),
.Y(n_1577)
);

AND2x4_ASAP7_75t_SL g1578 ( 
.A(n_1468),
.B(n_1513),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_1484),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1448),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1433),
.B(n_1443),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1460),
.B(n_1479),
.Y(n_1582)
);

NAND2xp33_ASAP7_75t_R g1583 ( 
.A(n_1470),
.B(n_1522),
.Y(n_1583)
);

AOI21xp33_ASAP7_75t_L g1584 ( 
.A1(n_1459),
.A2(n_1477),
.B(n_1501),
.Y(n_1584)
);

BUFx4f_ASAP7_75t_SL g1585 ( 
.A(n_1519),
.Y(n_1585)
);

NOR3xp33_ASAP7_75t_SL g1586 ( 
.A(n_1521),
.B(n_1539),
.C(n_1517),
.Y(n_1586)
);

NAND2xp33_ASAP7_75t_R g1587 ( 
.A(n_1470),
.B(n_1522),
.Y(n_1587)
);

BUFx3_ASAP7_75t_L g1588 ( 
.A(n_1503),
.Y(n_1588)
);

A2O1A1Ixp33_ASAP7_75t_L g1589 ( 
.A1(n_1492),
.A2(n_1539),
.B(n_1489),
.C(n_1506),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1450),
.Y(n_1590)
);

OAI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1449),
.A2(n_1529),
.B1(n_1552),
.B2(n_1446),
.Y(n_1591)
);

INVx2_ASAP7_75t_SL g1592 ( 
.A(n_1484),
.Y(n_1592)
);

NAND2xp33_ASAP7_75t_SL g1593 ( 
.A(n_1439),
.B(n_1478),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1458),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1509),
.B(n_1441),
.Y(n_1595)
);

OAI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1460),
.A2(n_1517),
.B1(n_1530),
.B2(n_1518),
.Y(n_1596)
);

OAI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1466),
.A2(n_1469),
.B1(n_1500),
.B2(n_1485),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1479),
.B(n_1510),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1444),
.Y(n_1599)
);

NAND2x1p5_ASAP7_75t_L g1600 ( 
.A(n_1526),
.B(n_1516),
.Y(n_1600)
);

AO31x2_ASAP7_75t_L g1601 ( 
.A1(n_1535),
.A2(n_1533),
.A3(n_1514),
.B(n_1511),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1493),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_R g1603 ( 
.A(n_1439),
.B(n_1478),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1525),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_R g1605 ( 
.A(n_1439),
.B(n_1478),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1457),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1508),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1431),
.B(n_1507),
.Y(n_1608)
);

OA21x2_ASAP7_75t_L g1609 ( 
.A1(n_1489),
.A2(n_1546),
.B(n_1524),
.Y(n_1609)
);

CKINVDCx20_ASAP7_75t_R g1610 ( 
.A(n_1504),
.Y(n_1610)
);

BUFx12f_ASAP7_75t_L g1611 ( 
.A(n_1437),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1538),
.B(n_1550),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1508),
.Y(n_1613)
);

NAND2xp33_ASAP7_75t_R g1614 ( 
.A(n_1531),
.B(n_1534),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1510),
.B(n_1464),
.Y(n_1615)
);

CKINVDCx16_ASAP7_75t_R g1616 ( 
.A(n_1437),
.Y(n_1616)
);

NOR3xp33_ASAP7_75t_SL g1617 ( 
.A(n_1544),
.B(n_1545),
.C(n_1533),
.Y(n_1617)
);

AND2x4_ASAP7_75t_L g1618 ( 
.A(n_1455),
.B(n_1472),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1463),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1465),
.A2(n_1505),
.B1(n_1481),
.B2(n_1475),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1527),
.Y(n_1621)
);

INVx3_ASAP7_75t_L g1622 ( 
.A(n_1451),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_1451),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1455),
.B(n_1472),
.Y(n_1624)
);

CKINVDCx16_ASAP7_75t_R g1625 ( 
.A(n_1453),
.Y(n_1625)
);

OAI21xp33_ASAP7_75t_L g1626 ( 
.A1(n_1540),
.A2(n_1543),
.B(n_1536),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1541),
.Y(n_1627)
);

OR2x6_ASAP7_75t_L g1628 ( 
.A(n_1496),
.B(n_1472),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1580),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1602),
.Y(n_1630)
);

BUFx3_ASAP7_75t_L g1631 ( 
.A(n_1600),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1604),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1563),
.B(n_1436),
.Y(n_1633)
);

HB1xp67_ASAP7_75t_L g1634 ( 
.A(n_1559),
.Y(n_1634)
);

AND2x4_ASAP7_75t_L g1635 ( 
.A(n_1618),
.B(n_1455),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1556),
.B(n_1542),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1601),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1601),
.Y(n_1638)
);

AND2x4_ASAP7_75t_L g1639 ( 
.A(n_1618),
.B(n_1496),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1563),
.B(n_1436),
.Y(n_1640)
);

OAI221xp5_ASAP7_75t_L g1641 ( 
.A1(n_1561),
.A2(n_1496),
.B1(n_1544),
.B2(n_1528),
.C(n_1545),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1604),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1563),
.B(n_1528),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1573),
.B(n_1528),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1624),
.B(n_1474),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1628),
.B(n_1474),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1559),
.B(n_1537),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1576),
.Y(n_1648)
);

BUFx3_ASAP7_75t_L g1649 ( 
.A(n_1600),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1601),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1628),
.B(n_1453),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1590),
.Y(n_1652)
);

INVx5_ASAP7_75t_L g1653 ( 
.A(n_1628),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1594),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1601),
.Y(n_1655)
);

OR2x6_ASAP7_75t_SL g1656 ( 
.A(n_1591),
.B(n_1491),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1617),
.B(n_1454),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1597),
.Y(n_1658)
);

OAI221xp5_ASAP7_75t_L g1659 ( 
.A1(n_1554),
.A2(n_1454),
.B1(n_1515),
.B2(n_1562),
.C(n_1584),
.Y(n_1659)
);

INVx2_ASAP7_75t_SL g1660 ( 
.A(n_1627),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1597),
.Y(n_1661)
);

BUFx2_ASAP7_75t_L g1662 ( 
.A(n_1617),
.Y(n_1662)
);

BUFx2_ASAP7_75t_L g1663 ( 
.A(n_1557),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1599),
.Y(n_1664)
);

INVx5_ASAP7_75t_L g1665 ( 
.A(n_1622),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1615),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1556),
.B(n_1515),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1615),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1581),
.B(n_1613),
.Y(n_1669)
);

BUFx2_ASAP7_75t_L g1670 ( 
.A(n_1566),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1581),
.B(n_1626),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1607),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1575),
.B(n_1609),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1575),
.B(n_1609),
.Y(n_1674)
);

AOI31xp33_ASAP7_75t_L g1675 ( 
.A1(n_1554),
.A2(n_1584),
.A3(n_1558),
.B(n_1565),
.Y(n_1675)
);

INVx3_ASAP7_75t_L g1676 ( 
.A(n_1606),
.Y(n_1676)
);

OAI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1675),
.A2(n_1662),
.B1(n_1659),
.B2(n_1610),
.Y(n_1677)
);

NAND3xp33_ASAP7_75t_L g1678 ( 
.A(n_1675),
.B(n_1562),
.C(n_1589),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1662),
.A2(n_1571),
.B1(n_1596),
.B2(n_1588),
.Y(n_1679)
);

NAND4xp25_ASAP7_75t_L g1680 ( 
.A(n_1671),
.B(n_1620),
.C(n_1614),
.D(n_1582),
.Y(n_1680)
);

OA21x2_ASAP7_75t_L g1681 ( 
.A1(n_1637),
.A2(n_1586),
.B(n_1582),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1634),
.B(n_1608),
.Y(n_1682)
);

NAND3xp33_ASAP7_75t_L g1683 ( 
.A(n_1659),
.B(n_1586),
.C(n_1620),
.Y(n_1683)
);

OAI221xp5_ASAP7_75t_SL g1684 ( 
.A1(n_1671),
.A2(n_1592),
.B1(n_1560),
.B2(n_1598),
.C(n_1574),
.Y(n_1684)
);

NAND3xp33_ASAP7_75t_L g1685 ( 
.A(n_1658),
.B(n_1621),
.C(n_1623),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1667),
.B(n_1564),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1667),
.B(n_1595),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1669),
.B(n_1612),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1658),
.A2(n_1577),
.B1(n_1568),
.B2(n_1611),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1645),
.B(n_1578),
.Y(n_1690)
);

OAI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1656),
.A2(n_1641),
.B1(n_1585),
.B2(n_1579),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1669),
.B(n_1598),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1666),
.B(n_1619),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1645),
.B(n_1625),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1666),
.B(n_1616),
.Y(n_1695)
);

NAND3xp33_ASAP7_75t_L g1696 ( 
.A(n_1661),
.B(n_1641),
.C(n_1673),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1668),
.B(n_1569),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1668),
.B(n_1622),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1663),
.B(n_1553),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1645),
.B(n_1605),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1663),
.B(n_1603),
.Y(n_1701)
);

OA211x2_ASAP7_75t_L g1702 ( 
.A1(n_1656),
.A2(n_1585),
.B(n_1593),
.C(n_1572),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1673),
.B(n_1567),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1673),
.B(n_1555),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1674),
.B(n_1583),
.Y(n_1705)
);

OA211x2_ASAP7_75t_L g1706 ( 
.A1(n_1656),
.A2(n_1570),
.B(n_1587),
.C(n_1636),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1670),
.B(n_1661),
.Y(n_1707)
);

OA21x2_ASAP7_75t_L g1708 ( 
.A1(n_1637),
.A2(n_1638),
.B(n_1650),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1674),
.B(n_1670),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1672),
.B(n_1636),
.Y(n_1710)
);

NAND4xp25_ASAP7_75t_L g1711 ( 
.A(n_1674),
.B(n_1657),
.C(n_1672),
.D(n_1640),
.Y(n_1711)
);

OA21x2_ASAP7_75t_L g1712 ( 
.A1(n_1637),
.A2(n_1650),
.B(n_1655),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1648),
.B(n_1654),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1635),
.B(n_1644),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1635),
.B(n_1644),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1648),
.B(n_1654),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1635),
.B(n_1639),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1632),
.Y(n_1718)
);

OAI21xp5_ASAP7_75t_SL g1719 ( 
.A1(n_1657),
.A2(n_1643),
.B(n_1639),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1652),
.B(n_1676),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1711),
.B(n_1647),
.Y(n_1721)
);

HB1xp67_ASAP7_75t_L g1722 ( 
.A(n_1709),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1717),
.B(n_1643),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1718),
.B(n_1632),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1717),
.B(n_1643),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1707),
.B(n_1709),
.Y(n_1726)
);

BUFx2_ASAP7_75t_L g1727 ( 
.A(n_1681),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1705),
.B(n_1715),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1718),
.B(n_1642),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1708),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1708),
.Y(n_1731)
);

HB1xp67_ASAP7_75t_L g1732 ( 
.A(n_1720),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1710),
.Y(n_1733)
);

INVx3_ASAP7_75t_L g1734 ( 
.A(n_1708),
.Y(n_1734)
);

AND2x4_ASAP7_75t_L g1735 ( 
.A(n_1714),
.B(n_1653),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1692),
.B(n_1642),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1693),
.B(n_1716),
.Y(n_1737)
);

AND2x4_ASAP7_75t_L g1738 ( 
.A(n_1714),
.B(n_1653),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1713),
.B(n_1652),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1688),
.B(n_1629),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1696),
.B(n_1647),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1708),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1696),
.B(n_1676),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1680),
.B(n_1687),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1719),
.B(n_1676),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1698),
.B(n_1629),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1705),
.B(n_1630),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1715),
.B(n_1639),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1694),
.B(n_1700),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1712),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1712),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1694),
.B(n_1639),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1681),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1700),
.B(n_1639),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1712),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1681),
.B(n_1676),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1703),
.B(n_1653),
.Y(n_1757)
);

BUFx2_ASAP7_75t_L g1758 ( 
.A(n_1722),
.Y(n_1758)
);

HB1xp67_ASAP7_75t_L g1759 ( 
.A(n_1733),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1744),
.B(n_1703),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1734),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1724),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1734),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1724),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1735),
.B(n_1653),
.Y(n_1765)
);

AND2x4_ASAP7_75t_L g1766 ( 
.A(n_1735),
.B(n_1653),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1729),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1757),
.B(n_1704),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1757),
.B(n_1704),
.Y(n_1769)
);

INVx1_ASAP7_75t_SL g1770 ( 
.A(n_1727),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1744),
.B(n_1697),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1729),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1728),
.B(n_1681),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1747),
.B(n_1682),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1728),
.B(n_1690),
.Y(n_1775)
);

INVx2_ASAP7_75t_SL g1776 ( 
.A(n_1735),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1726),
.B(n_1684),
.Y(n_1777)
);

OR2x2_ASAP7_75t_L g1778 ( 
.A(n_1726),
.B(n_1695),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1739),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1723),
.B(n_1690),
.Y(n_1780)
);

OR2x2_ASAP7_75t_L g1781 ( 
.A(n_1743),
.B(n_1664),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1747),
.B(n_1737),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1743),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1741),
.B(n_1721),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1739),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1737),
.B(n_1630),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1723),
.B(n_1682),
.Y(n_1787)
);

INVx3_ASAP7_75t_L g1788 ( 
.A(n_1734),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1749),
.B(n_1699),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1746),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1735),
.B(n_1653),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1734),
.Y(n_1792)
);

BUFx3_ASAP7_75t_L g1793 ( 
.A(n_1727),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1730),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1725),
.B(n_1748),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1725),
.B(n_1686),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1746),
.Y(n_1797)
);

NOR2xp67_ASAP7_75t_R g1798 ( 
.A(n_1753),
.B(n_1702),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1736),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1793),
.Y(n_1800)
);

OAI322xp33_ASAP7_75t_L g1801 ( 
.A1(n_1784),
.A2(n_1741),
.A3(n_1678),
.B1(n_1677),
.B2(n_1721),
.C1(n_1691),
.C2(n_1756),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1760),
.B(n_1749),
.Y(n_1802)
);

NOR2x1p5_ASAP7_75t_L g1803 ( 
.A(n_1771),
.B(n_1678),
.Y(n_1803)
);

AOI22xp5_ASAP7_75t_L g1804 ( 
.A1(n_1768),
.A2(n_1683),
.B1(n_1769),
.B2(n_1789),
.Y(n_1804)
);

OAI32xp33_ASAP7_75t_L g1805 ( 
.A1(n_1777),
.A2(n_1745),
.A3(n_1756),
.B1(n_1683),
.B2(n_1679),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1758),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1758),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1768),
.B(n_1754),
.Y(n_1808)
);

XNOR2xp5_ASAP7_75t_L g1809 ( 
.A(n_1769),
.B(n_1702),
.Y(n_1809)
);

OA222x2_ASAP7_75t_L g1810 ( 
.A1(n_1793),
.A2(n_1745),
.B1(n_1631),
.B2(n_1649),
.C1(n_1706),
.C2(n_1701),
.Y(n_1810)
);

INVxp67_ASAP7_75t_L g1811 ( 
.A(n_1793),
.Y(n_1811)
);

OR2x2_ASAP7_75t_L g1812 ( 
.A(n_1784),
.B(n_1740),
.Y(n_1812)
);

OAI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1777),
.A2(n_1685),
.B1(n_1706),
.B2(n_1653),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1788),
.Y(n_1814)
);

AOI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1796),
.A2(n_1738),
.B1(n_1685),
.B2(n_1657),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1795),
.B(n_1738),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1759),
.B(n_1732),
.Y(n_1817)
);

OR2x2_ASAP7_75t_L g1818 ( 
.A(n_1778),
.B(n_1740),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1781),
.Y(n_1819)
);

NAND3xp33_ASAP7_75t_L g1820 ( 
.A(n_1783),
.B(n_1689),
.C(n_1736),
.Y(n_1820)
);

OA222x2_ASAP7_75t_L g1821 ( 
.A1(n_1798),
.A2(n_1631),
.B1(n_1649),
.B2(n_1755),
.C1(n_1751),
.C2(n_1750),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1796),
.B(n_1754),
.Y(n_1822)
);

AOI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1776),
.A2(n_1738),
.B1(n_1752),
.B2(n_1651),
.Y(n_1823)
);

OAI22xp5_ASAP7_75t_L g1824 ( 
.A1(n_1778),
.A2(n_1752),
.B1(n_1738),
.B2(n_1748),
.Y(n_1824)
);

AOI22xp5_ASAP7_75t_L g1825 ( 
.A1(n_1776),
.A2(n_1651),
.B1(n_1646),
.B2(n_1633),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1788),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1795),
.B(n_1633),
.Y(n_1827)
);

NOR2xp67_ASAP7_75t_SL g1828 ( 
.A(n_1798),
.B(n_1665),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1775),
.B(n_1635),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1782),
.B(n_1660),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1781),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1774),
.B(n_1782),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1775),
.B(n_1635),
.Y(n_1833)
);

AOI22xp33_ASAP7_75t_L g1834 ( 
.A1(n_1770),
.A2(n_1633),
.B1(n_1640),
.B2(n_1638),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1803),
.B(n_1787),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1806),
.Y(n_1836)
);

OAI211xp5_ASAP7_75t_SL g1837 ( 
.A1(n_1804),
.A2(n_1770),
.B(n_1797),
.C(n_1790),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1807),
.Y(n_1838)
);

OR2x2_ASAP7_75t_L g1839 ( 
.A(n_1802),
.B(n_1799),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1811),
.Y(n_1840)
);

NOR2xp67_ASAP7_75t_SL g1841 ( 
.A(n_1820),
.B(n_1800),
.Y(n_1841)
);

HB1xp67_ASAP7_75t_L g1842 ( 
.A(n_1811),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1800),
.Y(n_1843)
);

NOR2xp33_ASAP7_75t_SL g1844 ( 
.A(n_1813),
.B(n_1765),
.Y(n_1844)
);

OAI21xp5_ASAP7_75t_L g1845 ( 
.A1(n_1813),
.A2(n_1765),
.B(n_1791),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1817),
.B(n_1799),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1819),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1831),
.Y(n_1848)
);

INVxp67_ASAP7_75t_SL g1849 ( 
.A(n_1814),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1830),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1812),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1818),
.B(n_1797),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1822),
.B(n_1790),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1808),
.Y(n_1854)
);

OAI21xp5_ASAP7_75t_L g1855 ( 
.A1(n_1805),
.A2(n_1765),
.B(n_1791),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1832),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1810),
.B(n_1787),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1816),
.B(n_1833),
.Y(n_1858)
);

INVxp67_ASAP7_75t_SL g1859 ( 
.A(n_1814),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1858),
.Y(n_1860)
);

AOI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1841),
.A2(n_1809),
.B1(n_1815),
.B2(n_1823),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1842),
.Y(n_1862)
);

AOI332xp33_ASAP7_75t_L g1863 ( 
.A1(n_1840),
.A2(n_1856),
.A3(n_1838),
.B1(n_1836),
.B2(n_1851),
.B3(n_1848),
.C1(n_1847),
.C2(n_1843),
.Y(n_1863)
);

INVxp33_ASAP7_75t_L g1864 ( 
.A(n_1835),
.Y(n_1864)
);

AOI22xp33_ASAP7_75t_L g1865 ( 
.A1(n_1857),
.A2(n_1801),
.B1(n_1765),
.B2(n_1791),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1842),
.Y(n_1866)
);

NAND3xp33_ASAP7_75t_L g1867 ( 
.A(n_1844),
.B(n_1828),
.C(n_1834),
.Y(n_1867)
);

NOR2xp33_ASAP7_75t_L g1868 ( 
.A(n_1837),
.B(n_1824),
.Y(n_1868)
);

AOI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1857),
.A2(n_1791),
.B1(n_1766),
.B2(n_1816),
.Y(n_1869)
);

HB1xp67_ASAP7_75t_L g1870 ( 
.A(n_1849),
.Y(n_1870)
);

AOI21xp33_ASAP7_75t_L g1871 ( 
.A1(n_1855),
.A2(n_1834),
.B(n_1826),
.Y(n_1871)
);

INVx2_ASAP7_75t_SL g1872 ( 
.A(n_1858),
.Y(n_1872)
);

OAI21xp33_ASAP7_75t_L g1873 ( 
.A1(n_1854),
.A2(n_1825),
.B(n_1773),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1849),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1850),
.B(n_1829),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1853),
.B(n_1785),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1859),
.B(n_1779),
.Y(n_1877)
);

AND2x4_ASAP7_75t_L g1878 ( 
.A(n_1859),
.B(n_1766),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1870),
.Y(n_1879)
);

OAI22xp5_ASAP7_75t_L g1880 ( 
.A1(n_1865),
.A2(n_1845),
.B1(n_1846),
.B2(n_1839),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1870),
.Y(n_1881)
);

AOI221xp5_ASAP7_75t_L g1882 ( 
.A1(n_1868),
.A2(n_1852),
.B1(n_1821),
.B2(n_1772),
.C(n_1767),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_SL g1883 ( 
.A(n_1867),
.B(n_1852),
.Y(n_1883)
);

O2A1O1Ixp33_ASAP7_75t_L g1884 ( 
.A1(n_1862),
.A2(n_1826),
.B(n_1773),
.C(n_1764),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1874),
.Y(n_1885)
);

OAI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1861),
.A2(n_1766),
.B1(n_1827),
.B2(n_1780),
.Y(n_1886)
);

NAND3x1_ASAP7_75t_SL g1887 ( 
.A(n_1875),
.B(n_1827),
.C(n_1780),
.Y(n_1887)
);

NAND2x1p5_ASAP7_75t_L g1888 ( 
.A(n_1878),
.B(n_1766),
.Y(n_1888)
);

AOI22xp5_ASAP7_75t_L g1889 ( 
.A1(n_1872),
.A2(n_1779),
.B1(n_1785),
.B2(n_1767),
.Y(n_1889)
);

OAI222xp33_ASAP7_75t_L g1890 ( 
.A1(n_1883),
.A2(n_1869),
.B1(n_1866),
.B2(n_1860),
.C1(n_1878),
.C2(n_1876),
.Y(n_1890)
);

OAI21xp5_ASAP7_75t_SL g1891 ( 
.A1(n_1882),
.A2(n_1864),
.B(n_1871),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1881),
.B(n_1873),
.Y(n_1892)
);

NAND3xp33_ASAP7_75t_L g1893 ( 
.A(n_1879),
.B(n_1871),
.C(n_1877),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1885),
.Y(n_1894)
);

OAI21xp33_ASAP7_75t_SL g1895 ( 
.A1(n_1880),
.A2(n_1877),
.B(n_1889),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1886),
.B(n_1764),
.Y(n_1896)
);

INVx1_ASAP7_75t_SL g1897 ( 
.A(n_1888),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1884),
.B(n_1772),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1887),
.B(n_1762),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1894),
.Y(n_1900)
);

INVx2_ASAP7_75t_SL g1901 ( 
.A(n_1897),
.Y(n_1901)
);

OAI21xp33_ASAP7_75t_L g1902 ( 
.A1(n_1891),
.A2(n_1863),
.B(n_1762),
.Y(n_1902)
);

NOR2x1_ASAP7_75t_L g1903 ( 
.A(n_1893),
.B(n_1788),
.Y(n_1903)
);

AOI211x1_ASAP7_75t_L g1904 ( 
.A1(n_1890),
.A2(n_1786),
.B(n_1751),
.C(n_1755),
.Y(n_1904)
);

OAI211xp5_ASAP7_75t_SL g1905 ( 
.A1(n_1902),
.A2(n_1895),
.B(n_1892),
.C(n_1901),
.Y(n_1905)
);

OAI31xp33_ASAP7_75t_L g1906 ( 
.A1(n_1900),
.A2(n_1899),
.A3(n_1898),
.B(n_1896),
.Y(n_1906)
);

NAND3xp33_ASAP7_75t_L g1907 ( 
.A(n_1904),
.B(n_1794),
.C(n_1792),
.Y(n_1907)
);

OAI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1903),
.A2(n_1788),
.B1(n_1786),
.B2(n_1761),
.Y(n_1908)
);

NOR3x1_ASAP7_75t_L g1909 ( 
.A(n_1901),
.B(n_1750),
.C(n_1660),
.Y(n_1909)
);

AOI21xp33_ASAP7_75t_L g1910 ( 
.A1(n_1901),
.A2(n_1794),
.B(n_1792),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1909),
.Y(n_1911)
);

NOR2x1_ASAP7_75t_L g1912 ( 
.A(n_1905),
.B(n_1792),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1907),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1906),
.B(n_1794),
.Y(n_1914)
);

OR2x2_ASAP7_75t_L g1915 ( 
.A(n_1910),
.B(n_1763),
.Y(n_1915)
);

AOI22xp5_ASAP7_75t_L g1916 ( 
.A1(n_1911),
.A2(n_1908),
.B1(n_1763),
.B2(n_1761),
.Y(n_1916)
);

AOI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1913),
.A2(n_1763),
.B1(n_1761),
.B2(n_1742),
.Y(n_1917)
);

CKINVDCx20_ASAP7_75t_R g1918 ( 
.A(n_1914),
.Y(n_1918)
);

NOR2x1_ASAP7_75t_L g1919 ( 
.A(n_1918),
.B(n_1912),
.Y(n_1919)
);

HB1xp67_ASAP7_75t_L g1920 ( 
.A(n_1919),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1920),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1920),
.B(n_1916),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1922),
.Y(n_1923)
);

AOI22xp33_ASAP7_75t_L g1924 ( 
.A1(n_1921),
.A2(n_1915),
.B1(n_1917),
.B2(n_1742),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1923),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1924),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1925),
.Y(n_1927)
);

OAI22xp5_ASAP7_75t_SL g1928 ( 
.A1(n_1927),
.A2(n_1926),
.B1(n_1742),
.B2(n_1731),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1928),
.Y(n_1929)
);

OAI21xp5_ASAP7_75t_L g1930 ( 
.A1(n_1929),
.A2(n_1731),
.B(n_1730),
.Y(n_1930)
);

AOI22xp33_ASAP7_75t_L g1931 ( 
.A1(n_1930),
.A2(n_1731),
.B1(n_1730),
.B2(n_1631),
.Y(n_1931)
);

OAI22xp5_ASAP7_75t_L g1932 ( 
.A1(n_1931),
.A2(n_1665),
.B1(n_1649),
.B2(n_1660),
.Y(n_1932)
);

AOI211xp5_ASAP7_75t_L g1933 ( 
.A1(n_1932),
.A2(n_1651),
.B(n_1640),
.C(n_1646),
.Y(n_1933)
);


endmodule