module fake_jpeg_25157_n_186 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_186);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx5_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_4),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_30),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_18),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_24),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_33),
.A2(n_30),
.B1(n_24),
.B2(n_25),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_27),
.A2(n_19),
.B1(n_15),
.B2(n_13),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_27),
.B1(n_30),
.B2(n_17),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_26),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_18),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_37),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_41),
.B(n_25),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_50),
.Y(n_58)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_44),
.B(n_45),
.Y(n_61)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVxp67_ASAP7_75t_SL g47 ( 
.A(n_38),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_24),
.B1(n_19),
.B2(n_27),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_48),
.A2(n_53),
.B1(n_23),
.B2(n_28),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_49),
.A2(n_37),
.B1(n_42),
.B2(n_34),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_35),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_51),
.A2(n_23),
.B1(n_28),
.B2(n_34),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_25),
.Y(n_52)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_42),
.A2(n_27),
.B1(n_30),
.B2(n_15),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_54),
.A2(n_30),
.B1(n_39),
.B2(n_40),
.Y(n_63)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_20),
.Y(n_56)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_59),
.A2(n_65),
.B1(n_51),
.B2(n_37),
.Y(n_82)
);

NOR2x1_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_33),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_62),
.B(n_51),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_39),
.B1(n_40),
.B2(n_46),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_66),
.A2(n_45),
.B1(n_53),
.B2(n_44),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_37),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_SL g79 ( 
.A(n_67),
.B(n_50),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_56),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_68),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_85),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_52),
.Y(n_74)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_75),
.B(n_76),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_64),
.B(n_43),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_77),
.A2(n_81),
.B1(n_82),
.B2(n_66),
.Y(n_94)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_84),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_67),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_62),
.Y(n_98)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_89),
.B(n_90),
.Y(n_105)
);

A2O1A1O1Ixp25_ASAP7_75t_L g90 ( 
.A1(n_79),
.A2(n_58),
.B(n_61),
.C(n_47),
.D(n_45),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_64),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_95),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_61),
.C(n_58),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_97),
.C(n_31),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_26),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_57),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_59),
.B(n_45),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_36),
.B(n_34),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_57),
.C(n_65),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_90),
.Y(n_113)
);

BUFx12_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_72),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_102),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_60),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_110),
.Y(n_117)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_97),
.A2(n_62),
.B1(n_84),
.B2(n_78),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_36),
.B1(n_28),
.B2(n_23),
.Y(n_128)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_107),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_88),
.B(n_73),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_108),
.A2(n_39),
.B1(n_70),
.B2(n_42),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_75),
.B1(n_73),
.B2(n_85),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_109),
.A2(n_98),
.B1(n_54),
.B2(n_42),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_113),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_114),
.A2(n_128),
.B1(n_55),
.B2(n_26),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_116),
.A2(n_122),
.B1(n_108),
.B2(n_23),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_106),
.A2(n_70),
.B1(n_28),
.B2(n_23),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_123),
.B(n_124),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_26),
.C(n_36),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_110),
.C(n_99),
.Y(n_132)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_18),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_101),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_132),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_105),
.C(n_113),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_133),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_131),
.A2(n_140),
.B1(n_114),
.B2(n_120),
.Y(n_147)
);

OAI322xp33_ASAP7_75t_L g133 ( 
.A1(n_127),
.A2(n_99),
.A3(n_108),
.B1(n_16),
.B2(n_22),
.C1(n_12),
.C2(n_18),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_26),
.C(n_29),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_134),
.Y(n_146)
);

NAND3xp33_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_10),
.C(n_11),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_135),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_22),
.Y(n_136)
);

BUFx24_ASAP7_75t_SL g144 ( 
.A(n_136),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_22),
.Y(n_137)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_26),
.C(n_29),
.Y(n_138)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_141),
.A2(n_124),
.B(n_119),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_143),
.B(n_7),
.Y(n_161)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_132),
.A2(n_125),
.B(n_128),
.C(n_16),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_17),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_139),
.A2(n_138),
.B1(n_137),
.B2(n_134),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_152),
.A2(n_55),
.B1(n_17),
.B2(n_8),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_150),
.B(n_136),
.Y(n_153)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_154),
.B(n_157),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_142),
.B(n_129),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_158),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_29),
.C(n_31),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_146),
.A2(n_143),
.B1(n_151),
.B2(n_144),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_159),
.A2(n_7),
.B(n_9),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_29),
.C(n_31),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_160),
.A2(n_161),
.B(n_0),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_156),
.A2(n_145),
.B1(n_149),
.B2(n_29),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_164),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_12),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_31),
.C(n_12),
.Y(n_172)
);

NOR2xp67_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_158),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_169),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_162),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_174),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_175),
.C(n_0),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_6),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_31),
.C(n_6),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_167),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_179),
.Y(n_181)
);

AOI322xp5_ASAP7_75t_L g178 ( 
.A1(n_173),
.A2(n_163),
.A3(n_6),
.B1(n_8),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_178)
);

AOI322xp5_ASAP7_75t_L g182 ( 
.A1(n_178),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_0),
.C1(n_1),
.C2(n_2),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_177),
.A2(n_4),
.B(n_9),
.Y(n_180)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_180),
.Y(n_183)
);

AOI321xp33_ASAP7_75t_L g184 ( 
.A1(n_182),
.A2(n_1),
.A3(n_2),
.B1(n_11),
.B2(n_150),
.C(n_80),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_181),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_183),
.Y(n_186)
);


endmodule