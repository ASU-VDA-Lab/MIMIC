module real_aes_8787_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g105 ( .A(n_0), .B(n_83), .C(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g122 ( .A(n_0), .Y(n_122) );
A2O1A1Ixp33_ASAP7_75t_L g237 ( .A1(n_1), .A2(n_139), .B(n_143), .C(n_238), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_2), .A2(n_175), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g463 ( .A(n_3), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_4), .B(n_215), .Y(n_272) );
AOI21xp33_ASAP7_75t_L g490 ( .A1(n_5), .A2(n_175), .B(n_491), .Y(n_490) );
AND2x6_ASAP7_75t_L g139 ( .A(n_6), .B(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g198 ( .A(n_7), .Y(n_198) );
INVx1_ASAP7_75t_L g104 ( .A(n_8), .Y(n_104) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_8), .B(n_40), .Y(n_123) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_9), .A2(n_174), .B(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_10), .B(n_151), .Y(n_242) );
INVx1_ASAP7_75t_L g495 ( .A(n_11), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_12), .B(n_209), .Y(n_518) );
INVx1_ASAP7_75t_L g159 ( .A(n_13), .Y(n_159) );
INVx1_ASAP7_75t_L g540 ( .A(n_14), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_15), .A2(n_149), .B(n_223), .C(n_225), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_16), .B(n_215), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_17), .B(n_474), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_18), .B(n_175), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_19), .B(n_188), .Y(n_187) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_20), .A2(n_209), .B(n_210), .C(n_212), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_21), .B(n_215), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_22), .B(n_151), .Y(n_259) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_23), .A2(n_183), .B(n_225), .C(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_24), .B(n_151), .Y(n_150) );
CKINVDCx16_ASAP7_75t_R g255 ( .A(n_25), .Y(n_255) );
INVx1_ASAP7_75t_L g147 ( .A(n_26), .Y(n_147) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_27), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_28), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_29), .B(n_151), .Y(n_464) );
INVx1_ASAP7_75t_L g181 ( .A(n_30), .Y(n_181) );
INVx1_ASAP7_75t_L g485 ( .A(n_31), .Y(n_485) );
INVx2_ASAP7_75t_L g137 ( .A(n_32), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g245 ( .A(n_33), .Y(n_245) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_34), .A2(n_209), .B(n_268), .C(n_270), .Y(n_267) );
AOI222xp33_ASAP7_75t_L g450 ( .A1(n_35), .A2(n_87), .B1(n_451), .B2(n_732), .C1(n_735), .C2(n_736), .Y(n_450) );
INVxp67_ASAP7_75t_L g182 ( .A(n_36), .Y(n_182) );
A2O1A1Ixp33_ASAP7_75t_L g142 ( .A1(n_37), .A2(n_143), .B(n_146), .C(n_154), .Y(n_142) );
CKINVDCx14_ASAP7_75t_R g266 ( .A(n_38), .Y(n_266) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_39), .A2(n_139), .B(n_143), .C(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_40), .B(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g484 ( .A(n_41), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g195 ( .A1(n_42), .A2(n_196), .B(n_197), .C(n_199), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_43), .B(n_151), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_44), .B(n_447), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g124 ( .A1(n_45), .A2(n_125), .B1(n_126), .B2(n_445), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_45), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g161 ( .A(n_46), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_47), .Y(n_177) );
INVx1_ASAP7_75t_L g207 ( .A(n_48), .Y(n_207) );
CKINVDCx16_ASAP7_75t_R g486 ( .A(n_49), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_50), .B(n_175), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_51), .A2(n_143), .B1(n_212), .B2(n_483), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_52), .Y(n_512) );
CKINVDCx16_ASAP7_75t_R g460 ( .A(n_53), .Y(n_460) );
CKINVDCx14_ASAP7_75t_R g194 ( .A(n_54), .Y(n_194) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_55), .A2(n_196), .B(n_270), .C(n_494), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_56), .Y(n_533) );
INVx1_ASAP7_75t_L g492 ( .A(n_57), .Y(n_492) );
INVx1_ASAP7_75t_L g140 ( .A(n_58), .Y(n_140) );
INVx1_ASAP7_75t_L g158 ( .A(n_59), .Y(n_158) );
INVx1_ASAP7_75t_SL g269 ( .A(n_60), .Y(n_269) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_61), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_62), .B(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g258 ( .A(n_63), .Y(n_258) );
A2O1A1Ixp33_ASAP7_75t_SL g473 ( .A1(n_64), .A2(n_270), .B(n_474), .C(n_475), .Y(n_473) );
INVxp67_ASAP7_75t_L g476 ( .A(n_65), .Y(n_476) );
INVx1_ASAP7_75t_L g108 ( .A(n_66), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_67), .A2(n_175), .B(n_193), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g262 ( .A(n_68), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_69), .A2(n_175), .B(n_220), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_70), .Y(n_488) );
INVx1_ASAP7_75t_L g527 ( .A(n_71), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_72), .A2(n_174), .B(n_176), .Y(n_173) );
CKINVDCx16_ASAP7_75t_R g141 ( .A(n_73), .Y(n_141) );
INVx1_ASAP7_75t_L g221 ( .A(n_74), .Y(n_221) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_75), .A2(n_139), .B(n_143), .C(n_529), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_76), .A2(n_175), .B(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g224 ( .A(n_77), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_78), .B(n_148), .Y(n_509) );
INVx2_ASAP7_75t_L g156 ( .A(n_79), .Y(n_156) );
INVx1_ASAP7_75t_L g239 ( .A(n_80), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_81), .B(n_474), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_L g461 ( .A1(n_82), .A2(n_139), .B(n_143), .C(n_462), .Y(n_461) );
OR2x2_ASAP7_75t_L g119 ( .A(n_83), .B(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g728 ( .A(n_83), .Y(n_728) );
OR2x2_ASAP7_75t_L g731 ( .A(n_83), .B(n_121), .Y(n_731) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_84), .A2(n_143), .B(n_257), .C(n_260), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_85), .B(n_155), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_86), .Y(n_467) );
CKINVDCx14_ASAP7_75t_R g735 ( .A(n_87), .Y(n_735) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_88), .A2(n_139), .B(n_143), .C(n_516), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_89), .Y(n_522) );
INVx1_ASAP7_75t_L g472 ( .A(n_90), .Y(n_472) );
CKINVDCx16_ASAP7_75t_R g537 ( .A(n_91), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_92), .B(n_148), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_93), .B(n_163), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_94), .B(n_163), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_95), .A2(n_100), .B1(n_109), .B2(n_741), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_96), .B(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g211 ( .A(n_97), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_98), .A2(n_175), .B(n_471), .Y(n_470) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
CKINVDCx6p67_ASAP7_75t_R g742 ( .A(n_101), .Y(n_742) );
CKINVDCx9p33_ASAP7_75t_R g101 ( .A(n_102), .Y(n_101) );
NOR2xp33_ASAP7_75t_L g102 ( .A(n_103), .B(n_105), .Y(n_102) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
OA21x2_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_115), .B(n_449), .Y(n_109) );
BUFx2_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_SL g740 ( .A(n_113), .Y(n_740) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
OAI21xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_124), .B(n_446), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_119), .Y(n_448) );
NOR2x2_ASAP7_75t_L g738 ( .A(n_120), .B(n_728), .Y(n_738) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g727 ( .A(n_121), .B(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
HB1xp67_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OAI22xp5_ASAP7_75t_SL g451 ( .A1(n_127), .A2(n_452), .B1(n_725), .B2(n_729), .Y(n_451) );
INVx1_ASAP7_75t_SL g734 ( .A(n_127), .Y(n_734) );
OR5x1_ASAP7_75t_L g127 ( .A(n_128), .B(n_339), .C(n_403), .D(n_419), .E(n_434), .Y(n_127) );
NAND4xp25_ASAP7_75t_L g128 ( .A(n_129), .B(n_273), .C(n_300), .D(n_323), .Y(n_128) );
AOI21xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_216), .B(n_227), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g130 ( .A(n_131), .B(n_165), .Y(n_130) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx3_ASAP7_75t_SL g250 ( .A(n_132), .Y(n_250) );
AND2x4_ASAP7_75t_L g286 ( .A(n_132), .B(n_275), .Y(n_286) );
OR2x2_ASAP7_75t_L g296 ( .A(n_132), .B(n_252), .Y(n_296) );
OR2x2_ASAP7_75t_L g342 ( .A(n_132), .B(n_168), .Y(n_342) );
AND2x2_ASAP7_75t_L g356 ( .A(n_132), .B(n_251), .Y(n_356) );
AND2x2_ASAP7_75t_L g399 ( .A(n_132), .B(n_289), .Y(n_399) );
AND2x2_ASAP7_75t_L g406 ( .A(n_132), .B(n_263), .Y(n_406) );
AND2x2_ASAP7_75t_L g425 ( .A(n_132), .B(n_315), .Y(n_425) );
AND2x2_ASAP7_75t_L g443 ( .A(n_132), .B(n_285), .Y(n_443) );
OR2x6_ASAP7_75t_L g132 ( .A(n_133), .B(n_160), .Y(n_132) );
O2A1O1Ixp33_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_141), .B(n_142), .C(n_155), .Y(n_133) );
OAI21xp5_ASAP7_75t_L g235 ( .A1(n_134), .A2(n_236), .B(n_237), .Y(n_235) );
OAI21xp5_ASAP7_75t_L g254 ( .A1(n_134), .A2(n_255), .B(n_256), .Y(n_254) );
OAI21xp5_ASAP7_75t_L g459 ( .A1(n_134), .A2(n_460), .B(n_461), .Y(n_459) );
OAI22xp33_ASAP7_75t_L g481 ( .A1(n_134), .A2(n_185), .B1(n_482), .B2(n_486), .Y(n_481) );
OAI21xp5_ASAP7_75t_L g526 ( .A1(n_134), .A2(n_527), .B(n_528), .Y(n_526) );
NAND2x1p5_ASAP7_75t_L g134 ( .A(n_135), .B(n_139), .Y(n_134) );
AND2x4_ASAP7_75t_L g175 ( .A(n_135), .B(n_139), .Y(n_175) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_138), .Y(n_135) );
INVx1_ASAP7_75t_L g153 ( .A(n_136), .Y(n_153) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g144 ( .A(n_137), .Y(n_144) );
INVx1_ASAP7_75t_L g213 ( .A(n_137), .Y(n_213) );
INVx1_ASAP7_75t_L g145 ( .A(n_138), .Y(n_145) );
INVx3_ASAP7_75t_L g149 ( .A(n_138), .Y(n_149) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_138), .Y(n_151) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_138), .Y(n_184) );
INVx1_ASAP7_75t_L g474 ( .A(n_138), .Y(n_474) );
BUFx3_ASAP7_75t_L g154 ( .A(n_139), .Y(n_154) );
INVx4_ASAP7_75t_SL g185 ( .A(n_139), .Y(n_185) );
INVx5_ASAP7_75t_L g178 ( .A(n_143), .Y(n_178) );
AND2x6_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
BUFx3_ASAP7_75t_L g200 ( .A(n_144), .Y(n_200) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_144), .Y(n_271) );
O2A1O1Ixp33_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_150), .C(n_152), .Y(n_146) );
OAI22xp33_ASAP7_75t_L g180 ( .A1(n_148), .A2(n_181), .B1(n_182), .B2(n_183), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_L g462 ( .A1(n_148), .A2(n_463), .B(n_464), .C(n_465), .Y(n_462) );
INVx5_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_149), .B(n_198), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_149), .B(n_476), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_149), .B(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g196 ( .A(n_151), .Y(n_196) );
INVx4_ASAP7_75t_L g209 ( .A(n_151), .Y(n_209) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_153), .B(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g189 ( .A(n_155), .Y(n_189) );
OA21x2_ASAP7_75t_L g191 ( .A1(n_155), .A2(n_192), .B(n_201), .Y(n_191) );
INVx1_ASAP7_75t_L g234 ( .A(n_155), .Y(n_234) );
OA21x2_ASAP7_75t_L g534 ( .A1(n_155), .A2(n_535), .B(n_541), .Y(n_534) );
AND2x2_ASAP7_75t_SL g155 ( .A(n_156), .B(n_157), .Y(n_155) );
AND2x2_ASAP7_75t_L g164 ( .A(n_156), .B(n_157), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
INVx3_ASAP7_75t_L g215 ( .A(n_162), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_162), .B(n_245), .Y(n_244) );
AO21x2_ASAP7_75t_L g253 ( .A1(n_162), .A2(n_254), .B(n_261), .Y(n_253) );
NOR2xp33_ASAP7_75t_SL g511 ( .A(n_162), .B(n_512), .Y(n_511) );
INVx4_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
HB1xp67_ASAP7_75t_L g204 ( .A(n_163), .Y(n_204) );
OA21x2_ASAP7_75t_L g469 ( .A1(n_163), .A2(n_470), .B(n_477), .Y(n_469) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g171 ( .A(n_164), .Y(n_171) );
INVx1_ASAP7_75t_L g408 ( .A(n_165), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_166), .B(n_190), .Y(n_165) );
AND2x2_ASAP7_75t_L g318 ( .A(n_166), .B(n_251), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_166), .B(n_338), .Y(n_337) );
AOI32xp33_ASAP7_75t_L g351 ( .A1(n_166), .A2(n_352), .A3(n_355), .B1(n_357), .B2(n_361), .Y(n_351) );
AND2x2_ASAP7_75t_L g421 ( .A(n_166), .B(n_315), .Y(n_421) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_SL g167 ( .A(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g285 ( .A(n_168), .B(n_252), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_168), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g327 ( .A(n_168), .B(n_274), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_168), .B(n_406), .Y(n_405) );
AO21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_172), .B(n_186), .Y(n_168) );
INVx1_ASAP7_75t_L g290 ( .A(n_169), .Y(n_290) );
AO21x2_ASAP7_75t_L g525 ( .A1(n_169), .A2(n_526), .B(n_532), .Y(n_525) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AOI21xp5_ASAP7_75t_SL g505 ( .A1(n_170), .A2(n_506), .B(n_507), .Y(n_505) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AO21x2_ASAP7_75t_L g458 ( .A1(n_171), .A2(n_459), .B(n_466), .Y(n_458) );
AO21x2_ASAP7_75t_L g480 ( .A1(n_171), .A2(n_481), .B(n_487), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_171), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
OA21x2_ASAP7_75t_L g289 ( .A1(n_173), .A2(n_187), .B(n_290), .Y(n_289) );
BUFx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_SL g176 ( .A1(n_177), .A2(n_178), .B(n_179), .C(n_185), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_SL g193 ( .A1(n_178), .A2(n_185), .B(n_194), .C(n_195), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_SL g206 ( .A1(n_178), .A2(n_185), .B(n_207), .C(n_208), .Y(n_206) );
O2A1O1Ixp33_ASAP7_75t_SL g220 ( .A1(n_178), .A2(n_185), .B(n_221), .C(n_222), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_L g265 ( .A1(n_178), .A2(n_185), .B(n_266), .C(n_267), .Y(n_265) );
O2A1O1Ixp33_ASAP7_75t_L g471 ( .A1(n_178), .A2(n_185), .B(n_472), .C(n_473), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_178), .A2(n_185), .B(n_492), .C(n_493), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_L g536 ( .A1(n_178), .A2(n_185), .B(n_537), .C(n_538), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_183), .B(n_211), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_183), .B(n_224), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_183), .B(n_540), .Y(n_539) );
INVx4_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g241 ( .A(n_184), .Y(n_241) );
OAI22xp5_ASAP7_75t_SL g483 ( .A1(n_184), .A2(n_241), .B1(n_484), .B2(n_485), .Y(n_483) );
INVx1_ASAP7_75t_L g260 ( .A(n_185), .Y(n_260) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_189), .B(n_262), .Y(n_261) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_189), .A2(n_514), .B(n_521), .Y(n_513) );
AND2x2_ASAP7_75t_L g292 ( .A(n_190), .B(n_231), .Y(n_292) );
AND2x2_ASAP7_75t_L g368 ( .A(n_190), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_SL g440 ( .A(n_190), .Y(n_440) );
AND2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_202), .Y(n_190) );
OR2x2_ASAP7_75t_L g230 ( .A(n_191), .B(n_203), .Y(n_230) );
AND2x2_ASAP7_75t_L g247 ( .A(n_191), .B(n_248), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_191), .B(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g299 ( .A(n_191), .Y(n_299) );
AND2x2_ASAP7_75t_L g326 ( .A(n_191), .B(n_203), .Y(n_326) );
BUFx3_ASAP7_75t_L g329 ( .A(n_191), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_191), .B(n_304), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_191), .B(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g243 ( .A(n_199), .Y(n_243) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g225 ( .A(n_200), .Y(n_225) );
INVx2_ASAP7_75t_L g280 ( .A(n_202), .Y(n_280) );
AND2x2_ASAP7_75t_L g298 ( .A(n_202), .B(n_278), .Y(n_298) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g309 ( .A(n_203), .B(n_218), .Y(n_309) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_203), .Y(n_322) );
OA21x2_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B(n_214), .Y(n_203) );
OA21x2_ASAP7_75t_L g218 ( .A1(n_204), .A2(n_219), .B(n_226), .Y(n_218) );
OA21x2_ASAP7_75t_L g263 ( .A1(n_204), .A2(n_264), .B(n_272), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_209), .B(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g465 ( .A(n_212), .Y(n_465) );
INVx3_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
OA21x2_ASAP7_75t_L g489 ( .A1(n_215), .A2(n_490), .B(n_496), .Y(n_489) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_217), .B(n_329), .Y(n_379) );
HB1xp67_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx1_ASAP7_75t_SL g248 ( .A(n_218), .Y(n_248) );
NAND3xp33_ASAP7_75t_L g297 ( .A(n_218), .B(n_298), .C(n_299), .Y(n_297) );
OR2x2_ASAP7_75t_L g305 ( .A(n_218), .B(n_278), .Y(n_305) );
AND2x2_ASAP7_75t_L g325 ( .A(n_218), .B(n_278), .Y(n_325) );
AND2x2_ASAP7_75t_L g369 ( .A(n_218), .B(n_233), .Y(n_369) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_246), .B(n_249), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_229), .B(n_231), .Y(n_228) );
AND2x2_ASAP7_75t_L g444 ( .A(n_229), .B(n_369), .Y(n_444) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_230), .A2(n_342), .B1(n_384), .B2(n_386), .Y(n_383) );
OR2x2_ASAP7_75t_L g390 ( .A(n_230), .B(n_305), .Y(n_390) );
OR2x2_ASAP7_75t_L g414 ( .A(n_230), .B(n_415), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_230), .B(n_334), .Y(n_427) );
AND2x2_ASAP7_75t_L g320 ( .A(n_231), .B(n_321), .Y(n_320) );
AOI21xp5_ASAP7_75t_L g407 ( .A1(n_231), .A2(n_393), .B(n_408), .Y(n_407) );
AOI32xp33_ASAP7_75t_L g428 ( .A1(n_231), .A2(n_318), .A3(n_429), .B1(n_431), .B2(n_432), .Y(n_428) );
OR2x2_ASAP7_75t_L g439 ( .A(n_231), .B(n_440), .Y(n_439) );
CKINVDCx16_ASAP7_75t_R g231 ( .A(n_232), .Y(n_231) );
OR2x2_ASAP7_75t_L g307 ( .A(n_232), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_232), .B(n_321), .Y(n_386) );
BUFx3_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx4_ASAP7_75t_L g278 ( .A(n_233), .Y(n_278) );
AND2x2_ASAP7_75t_L g344 ( .A(n_233), .B(n_309), .Y(n_344) );
AND3x2_ASAP7_75t_L g353 ( .A(n_233), .B(n_247), .C(n_354), .Y(n_353) );
AO21x2_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_244), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_234), .B(n_467), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_234), .B(n_522), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_234), .B(n_533), .Y(n_532) );
O2A1O1Ixp5_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_240), .B(n_242), .C(n_243), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_L g257 ( .A1(n_240), .A2(n_243), .B(n_258), .C(n_259), .Y(n_257) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_243), .A2(n_509), .B(n_510), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_243), .A2(n_530), .B(n_531), .Y(n_529) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g279 ( .A(n_248), .B(n_280), .Y(n_279) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_248), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_248), .B(n_278), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
AND2x2_ASAP7_75t_L g274 ( .A(n_250), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g314 ( .A(n_250), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g332 ( .A(n_250), .B(n_263), .Y(n_332) );
AND2x2_ASAP7_75t_L g350 ( .A(n_250), .B(n_252), .Y(n_350) );
OR2x2_ASAP7_75t_L g364 ( .A(n_250), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g410 ( .A(n_250), .B(n_338), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_251), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_263), .Y(n_251) );
AND2x2_ASAP7_75t_L g311 ( .A(n_252), .B(n_289), .Y(n_311) );
OR2x2_ASAP7_75t_L g365 ( .A(n_252), .B(n_289), .Y(n_365) );
AND2x2_ASAP7_75t_L g418 ( .A(n_252), .B(n_275), .Y(n_418) );
INVx2_ASAP7_75t_SL g252 ( .A(n_253), .Y(n_252) );
BUFx2_ASAP7_75t_L g316 ( .A(n_253), .Y(n_316) );
AND2x2_ASAP7_75t_L g338 ( .A(n_253), .B(n_263), .Y(n_338) );
INVx2_ASAP7_75t_L g275 ( .A(n_263), .Y(n_275) );
INVx1_ASAP7_75t_L g295 ( .A(n_263), .Y(n_295) );
INVx3_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_271), .Y(n_519) );
AOI211xp5_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_276), .B(n_281), .C(n_293), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_274), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g437 ( .A(n_274), .Y(n_437) );
AND2x2_ASAP7_75t_L g315 ( .A(n_275), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_279), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_278), .B(n_279), .Y(n_287) );
INVx1_ASAP7_75t_L g372 ( .A(n_278), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_278), .B(n_299), .Y(n_396) );
AND2x2_ASAP7_75t_L g412 ( .A(n_278), .B(n_326), .Y(n_412) );
NAND2xp5_ASAP7_75t_SL g394 ( .A(n_279), .B(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g303 ( .A(n_280), .Y(n_303) );
OAI22xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_287), .B1(n_288), .B2(n_291), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_284), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_285), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g310 ( .A(n_286), .B(n_311), .Y(n_310) );
AOI221xp5_ASAP7_75t_SL g375 ( .A1(n_286), .A2(n_328), .B1(n_376), .B2(n_381), .C(n_383), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_286), .B(n_349), .Y(n_382) );
INVx1_ASAP7_75t_L g442 ( .A(n_288), .Y(n_442) );
BUFx3_ASAP7_75t_L g349 ( .A(n_289), .Y(n_349) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AOI21xp33_ASAP7_75t_SL g293 ( .A1(n_294), .A2(n_296), .B(n_297), .Y(n_293) );
INVx1_ASAP7_75t_L g358 ( .A(n_295), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_295), .B(n_349), .Y(n_402) );
INVx1_ASAP7_75t_L g359 ( .A(n_296), .Y(n_359) );
NAND2xp5_ASAP7_75t_SL g360 ( .A(n_296), .B(n_349), .Y(n_360) );
INVxp67_ASAP7_75t_L g380 ( .A(n_298), .Y(n_380) );
AND2x2_ASAP7_75t_L g321 ( .A(n_299), .B(n_322), .Y(n_321) );
O2A1O1Ixp33_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_306), .B(n_310), .C(n_312), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx1_ASAP7_75t_SL g335 ( .A(n_303), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_304), .B(n_335), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_304), .B(n_326), .Y(n_377) );
INVx2_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g312 ( .A1(n_307), .A2(n_313), .B1(n_317), .B2(n_319), .Y(n_312) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g328 ( .A(n_309), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g373 ( .A(n_309), .B(n_374), .Y(n_373) );
OAI21xp33_ASAP7_75t_L g376 ( .A1(n_311), .A2(n_377), .B(n_378), .Y(n_376) );
INVx1_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
AOI221xp5_ASAP7_75t_L g323 ( .A1(n_315), .A2(n_324), .B1(n_327), .B2(n_328), .C(n_330), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_315), .B(n_349), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_315), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g431 ( .A(n_321), .Y(n_431) );
INVxp67_ASAP7_75t_L g354 ( .A(n_322), .Y(n_354) );
INVx1_ASAP7_75t_L g361 ( .A(n_324), .Y(n_361) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
AND2x2_ASAP7_75t_L g400 ( .A(n_325), .B(n_329), .Y(n_400) );
INVx1_ASAP7_75t_L g374 ( .A(n_329), .Y(n_374) );
NAND2xp5_ASAP7_75t_SL g404 ( .A(n_329), .B(n_344), .Y(n_404) );
OAI32xp33_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_333), .A3(n_335), .B1(n_336), .B2(n_337), .Y(n_330) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx2_ASAP7_75t_SL g343 ( .A(n_338), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_338), .B(n_370), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_338), .B(n_399), .Y(n_430) );
NAND2x1p5_ASAP7_75t_L g438 ( .A(n_338), .B(n_349), .Y(n_438) );
NAND5xp2_ASAP7_75t_L g339 ( .A(n_340), .B(n_362), .C(n_375), .D(n_387), .E(n_388), .Y(n_339) );
AOI221xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_344), .B1(n_345), .B2(n_347), .C(n_351), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp33_ASAP7_75t_SL g366 ( .A(n_346), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_349), .B(n_418), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_350), .A2(n_363), .B1(n_366), .B2(n_370), .Y(n_362) );
INVx2_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
OAI211xp5_ASAP7_75t_SL g357 ( .A1(n_353), .A2(n_358), .B(n_359), .C(n_360), .Y(n_357) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_SL g385 ( .A(n_365), .Y(n_385) );
INVx1_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_374), .B(n_423), .Y(n_433) );
OR2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AOI222xp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_391), .B1(n_393), .B2(n_397), .C1(n_400), .C2(n_401), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
OAI221xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_405), .B1(n_407), .B2(n_409), .C(n_411), .Y(n_403) );
INVx1_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
OAI21xp33_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_413), .B(n_416), .Y(n_411) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g423 ( .A(n_415), .Y(n_423) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OAI221xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_422), .B1(n_424), .B2(n_426), .C(n_428), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
INVxp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
A2O1A1Ixp33_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_438), .B(n_439), .C(n_441), .Y(n_434) );
INVxp67_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OAI21xp33_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_443), .B(n_444), .Y(n_441) );
NAND3xp33_ASAP7_75t_L g449 ( .A(n_446), .B(n_450), .C(n_739), .Y(n_449) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g733 ( .A(n_452), .Y(n_733) );
OR4x1_ASAP7_75t_L g452 ( .A(n_453), .B(n_614), .C(n_674), .D(n_701), .Y(n_452) );
NAND4xp25_ASAP7_75t_SL g453 ( .A(n_454), .B(n_562), .C(n_593), .D(n_610), .Y(n_453) );
O2A1O1Ixp33_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_497), .B(n_499), .C(n_542), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_456), .B(n_478), .Y(n_455) );
INVx1_ASAP7_75t_L g604 ( .A(n_456), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_456), .A2(n_645), .B1(n_693), .B2(n_723), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_468), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_457), .B(n_549), .Y(n_548) );
OR2x2_ASAP7_75t_L g555 ( .A(n_457), .B(n_480), .Y(n_555) );
AND2x2_ASAP7_75t_L g597 ( .A(n_457), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_457), .B(n_498), .Y(n_609) );
INVx1_ASAP7_75t_L g649 ( .A(n_457), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_457), .B(n_703), .Y(n_702) );
INVx3_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g577 ( .A(n_458), .B(n_480), .Y(n_577) );
INVx3_ASAP7_75t_L g581 ( .A(n_458), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_458), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g668 ( .A(n_468), .B(n_489), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_468), .B(n_581), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_468), .B(n_696), .Y(n_695) );
INVx3_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g498 ( .A(n_469), .B(n_480), .Y(n_498) );
INVx1_ASAP7_75t_L g550 ( .A(n_469), .Y(n_550) );
BUFx2_ASAP7_75t_L g554 ( .A(n_469), .Y(n_554) );
AND2x2_ASAP7_75t_L g598 ( .A(n_469), .B(n_479), .Y(n_598) );
OR2x2_ASAP7_75t_L g637 ( .A(n_469), .B(n_479), .Y(n_637) );
AND2x2_ASAP7_75t_L g662 ( .A(n_469), .B(n_489), .Y(n_662) );
AND2x2_ASAP7_75t_L g721 ( .A(n_469), .B(n_551), .Y(n_721) );
INVx1_ASAP7_75t_L g696 ( .A(n_478), .Y(n_696) );
OR2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_489), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_479), .B(n_489), .Y(n_582) );
AND2x2_ASAP7_75t_L g592 ( .A(n_479), .B(n_581), .Y(n_592) );
BUFx2_ASAP7_75t_L g603 ( .A(n_479), .Y(n_603) );
INVx3_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_L g625 ( .A(n_480), .B(n_489), .Y(n_625) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_480), .Y(n_680) );
AND2x2_ASAP7_75t_SL g497 ( .A(n_489), .B(n_498), .Y(n_497) );
INVx1_ASAP7_75t_SL g551 ( .A(n_489), .Y(n_551) );
BUFx2_ASAP7_75t_L g576 ( .A(n_489), .Y(n_576) );
INVx2_ASAP7_75t_L g595 ( .A(n_489), .Y(n_595) );
AND2x2_ASAP7_75t_L g657 ( .A(n_489), .B(n_581), .Y(n_657) );
AOI321xp33_ASAP7_75t_L g676 ( .A1(n_497), .A2(n_677), .A3(n_678), .B1(n_679), .B2(n_681), .C(n_682), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_498), .B(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_498), .B(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g670 ( .A(n_498), .B(n_649), .Y(n_670) );
AND2x2_ASAP7_75t_L g703 ( .A(n_498), .B(n_595), .Y(n_703) );
INVx1_ASAP7_75t_SL g499 ( .A(n_500), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_523), .Y(n_500) );
OR2x2_ASAP7_75t_L g605 ( .A(n_501), .B(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_513), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx3_ASAP7_75t_L g557 ( .A(n_504), .Y(n_557) );
AND2x2_ASAP7_75t_L g567 ( .A(n_504), .B(n_525), .Y(n_567) );
AND2x2_ASAP7_75t_L g572 ( .A(n_504), .B(n_547), .Y(n_572) );
INVx1_ASAP7_75t_L g589 ( .A(n_504), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_504), .B(n_570), .Y(n_608) );
AND2x2_ASAP7_75t_L g613 ( .A(n_504), .B(n_546), .Y(n_613) );
OR2x2_ASAP7_75t_L g645 ( .A(n_504), .B(n_634), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_504), .B(n_558), .Y(n_684) );
AND2x2_ASAP7_75t_L g718 ( .A(n_504), .B(n_544), .Y(n_718) );
OR2x6_ASAP7_75t_L g504 ( .A(n_505), .B(n_511), .Y(n_504) );
INVx1_ASAP7_75t_L g545 ( .A(n_513), .Y(n_545) );
INVx2_ASAP7_75t_L g560 ( .A(n_513), .Y(n_560) );
AND2x2_ASAP7_75t_L g600 ( .A(n_513), .B(n_571), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_513), .B(n_547), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_520), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B(n_519), .Y(n_516) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g706 ( .A(n_524), .B(n_557), .Y(n_706) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_534), .Y(n_524) );
INVx2_ASAP7_75t_L g547 ( .A(n_525), .Y(n_547) );
AND2x2_ASAP7_75t_L g700 ( .A(n_525), .B(n_560), .Y(n_700) );
AND2x2_ASAP7_75t_L g546 ( .A(n_534), .B(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g561 ( .A(n_534), .Y(n_561) );
INVx1_ASAP7_75t_L g571 ( .A(n_534), .Y(n_571) );
OAI22xp33_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_548), .B1(n_552), .B2(n_556), .Y(n_542) );
OAI22xp33_ASAP7_75t_L g697 ( .A1(n_543), .A2(n_661), .B1(n_698), .B2(n_699), .Y(n_697) );
INVx1_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
INVx1_ASAP7_75t_L g612 ( .A(n_545), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_546), .B(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g607 ( .A(n_547), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_547), .B(n_560), .Y(n_634) );
INVx1_ASAP7_75t_L g650 ( .A(n_547), .Y(n_650) );
AND2x2_ASAP7_75t_L g591 ( .A(n_549), .B(n_592), .Y(n_591) );
INVx3_ASAP7_75t_SL g630 ( .A(n_549), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_549), .B(n_555), .Y(n_707) );
AND2x4_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
INVx1_ASAP7_75t_L g716 ( .A(n_552), .Y(n_716) );
OR2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_555), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_553), .B(n_649), .Y(n_691) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx3_ASAP7_75t_SL g596 ( .A(n_555), .Y(n_596) );
NAND2x1_ASAP7_75t_SL g556 ( .A(n_557), .B(n_558), .Y(n_556) );
AND2x2_ASAP7_75t_L g617 ( .A(n_557), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g624 ( .A(n_557), .B(n_561), .Y(n_624) );
AND2x2_ASAP7_75t_L g629 ( .A(n_557), .B(n_570), .Y(n_629) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_557), .Y(n_678) );
OAI311xp33_ASAP7_75t_L g701 ( .A1(n_558), .A2(n_702), .A3(n_704), .B1(n_705), .C1(n_715), .Y(n_701) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
OR2x2_ASAP7_75t_L g714 ( .A(n_559), .B(n_587), .Y(n_714) );
OR2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
AND2x2_ASAP7_75t_L g570 ( .A(n_560), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g618 ( .A(n_560), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g673 ( .A(n_560), .Y(n_673) );
INVx1_ASAP7_75t_L g566 ( .A(n_561), .Y(n_566) );
INVx1_ASAP7_75t_L g586 ( .A(n_561), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_561), .B(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g619 ( .A(n_561), .Y(n_619) );
AOI221xp5_ASAP7_75t_SL g562 ( .A1(n_563), .A2(n_565), .B1(n_573), .B2(n_578), .C(n_583), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_568), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
INVx4_ASAP7_75t_L g587 ( .A(n_567), .Y(n_587) );
AND2x2_ASAP7_75t_L g681 ( .A(n_567), .B(n_600), .Y(n_681) );
AND2x2_ASAP7_75t_L g688 ( .A(n_567), .B(n_570), .Y(n_688) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_570), .B(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g599 ( .A(n_572), .B(n_600), .Y(n_599) );
INVx1_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_575), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g724 ( .A(n_577), .B(n_668), .Y(n_724) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g709 ( .A(n_581), .B(n_637), .Y(n_709) );
OAI211xp5_ASAP7_75t_L g674 ( .A1(n_582), .A2(n_675), .B(n_676), .C(n_689), .Y(n_674) );
AOI21xp33_ASAP7_75t_SL g583 ( .A1(n_584), .A2(n_588), .B(n_590), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NOR2xp67_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
INVx1_ASAP7_75t_L g653 ( .A(n_587), .Y(n_653) );
OAI221xp5_ASAP7_75t_L g682 ( .A1(n_588), .A2(n_683), .B1(n_684), .B2(n_685), .C(n_686), .Y(n_682) );
AND2x2_ASAP7_75t_L g659 ( .A(n_589), .B(n_600), .Y(n_659) );
AND2x2_ASAP7_75t_L g712 ( .A(n_589), .B(n_607), .Y(n_712) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_592), .B(n_630), .Y(n_654) );
O2A1O1Ixp33_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_597), .B(n_599), .C(n_601), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
AND2x2_ASAP7_75t_L g640 ( .A(n_595), .B(n_598), .Y(n_640) );
OR2x2_ASAP7_75t_L g683 ( .A(n_595), .B(n_637), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_596), .B(n_662), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_596), .B(n_668), .Y(n_667) );
INVx1_ASAP7_75t_SL g627 ( .A(n_597), .Y(n_627) );
INVx1_ASAP7_75t_L g693 ( .A(n_600), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_605), .B1(n_608), .B2(n_609), .Y(n_601) );
INVx1_ASAP7_75t_L g616 ( .A(n_602), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_603), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g679 ( .A(n_604), .B(n_680), .Y(n_679) );
INVxp67_ASAP7_75t_L g665 ( .A(n_606), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_607), .B(n_693), .Y(n_692) );
OAI22xp33_ASAP7_75t_L g666 ( .A1(n_608), .A2(n_667), .B1(n_669), .B2(n_671), .Y(n_666) );
INVx1_ASAP7_75t_L g675 ( .A(n_611), .Y(n_675) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
AND2x2_ASAP7_75t_L g717 ( .A(n_612), .B(n_712), .Y(n_717) );
AOI222xp33_ASAP7_75t_L g646 ( .A1(n_613), .A2(n_647), .B1(n_650), .B2(n_651), .C1(n_654), .C2(n_655), .Y(n_646) );
NAND4xp25_ASAP7_75t_SL g614 ( .A(n_615), .B(n_635), .C(n_646), .D(n_658), .Y(n_614) );
AOI221xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_617), .B1(n_620), .B2(n_625), .C(n_626), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_618), .B(n_653), .Y(n_652) );
INVxp67_ASAP7_75t_L g644 ( .A(n_619), .Y(n_644) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_620), .A2(n_690), .B1(n_692), .B2(n_694), .C(n_697), .Y(n_689) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g632 ( .A(n_624), .B(n_633), .Y(n_632) );
OAI21xp33_ASAP7_75t_L g686 ( .A1(n_625), .A2(n_687), .B(n_688), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_628), .B1(n_630), .B2(n_631), .Y(n_626) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OAI21xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_638), .B(n_641), .Y(n_635) );
INVxp67_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .Y(n_642) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g677 ( .A(n_648), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_649), .B(n_668), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_649), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_653), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_SL g685 ( .A(n_657), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_660), .B1(n_663), .B2(n_665), .C(n_666), .Y(n_658) );
INVxp67_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AOI222xp33_ASAP7_75t_L g705 ( .A1(n_668), .A2(n_706), .B1(n_707), .B2(n_708), .C1(n_710), .C2(n_713), .Y(n_705) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_672), .B(n_712), .Y(n_711) );
INVxp67_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g704 ( .A(n_678), .Y(n_704) );
INVxp67_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVxp33_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AOI221xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_717), .B1(n_718), .B2(n_719), .C(n_722), .Y(n_715) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVxp67_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
OAI22xp5_ASAP7_75t_SL g732 ( .A1(n_725), .A2(n_731), .B1(n_733), .B2(n_734), .Y(n_732) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
INVx3_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_742), .Y(n_741) );
endmodule