module fake_jpeg_27953_n_250 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_250);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_250;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_36),
.B(n_19),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_37),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx4_ASAP7_75t_SL g75 ( 
.A(n_39),
.Y(n_75)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_46),
.Y(n_62)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_30),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_24),
.B1(n_22),
.B2(n_33),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_48),
.A2(n_58),
.B1(n_63),
.B2(n_21),
.Y(n_98)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_47),
.A2(n_32),
.B1(n_31),
.B2(n_25),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_52),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_45),
.Y(n_54)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_37),
.B(n_30),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_56),
.B(n_71),
.Y(n_103)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_47),
.A2(n_32),
.B1(n_31),
.B2(n_25),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_72),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_34),
.B1(n_33),
.B2(n_32),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_70),
.Y(n_84)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_38),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_37),
.B(n_34),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_74),
.A2(n_42),
.B1(n_40),
.B2(n_38),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_78),
.A2(n_107),
.B1(n_59),
.B2(n_27),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_SL g81 ( 
.A(n_72),
.B(n_20),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_23),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_46),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_82),
.B(n_89),
.Y(n_111)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_88),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_41),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_85),
.B(n_86),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_41),
.Y(n_86)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_18),
.Y(n_89)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_93),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_18),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_99),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_53),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_95),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_98),
.A2(n_105),
.B1(n_65),
.B2(n_54),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_28),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_28),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_49),
.B(n_39),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_102),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_50),
.B(n_28),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_65),
.A2(n_40),
.B1(n_42),
.B2(n_21),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_50),
.B(n_14),
.Y(n_107)
);

NOR2x1_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_39),
.Y(n_108)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_109),
.A2(n_115),
.B1(n_116),
.B2(n_119),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_97),
.A2(n_54),
.B1(n_64),
.B2(n_68),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_98),
.A2(n_81),
.B1(n_77),
.B2(n_106),
.Y(n_116)
);

NAND2x1_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_101),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_117),
.A2(n_124),
.B(n_90),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_2),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_105),
.A2(n_69),
.B1(n_57),
.B2(n_55),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_45),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_128),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_87),
.A2(n_23),
.B(n_26),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_59),
.B1(n_75),
.B2(n_27),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_126),
.A2(n_130),
.B1(n_80),
.B2(n_94),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_127),
.B(n_133),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_79),
.B(n_19),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_76),
.B(n_27),
.C(n_19),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_92),
.C(n_91),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_83),
.A2(n_35),
.B1(n_26),
.B2(n_4),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_90),
.A2(n_35),
.B1(n_3),
.B2(n_4),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_130),
.Y(n_143)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_103),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_134),
.B(n_9),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_135),
.A2(n_143),
.B1(n_155),
.B2(n_158),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_113),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_136),
.B(n_145),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_141),
.C(n_124),
.Y(n_168)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_148),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_123),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_139),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_96),
.C(n_76),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_80),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_128),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_146),
.B(n_147),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_78),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_104),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_149),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_151),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_96),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_153),
.A2(n_121),
.B(n_114),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_154),
.Y(n_177)
);

AO21x2_ASAP7_75t_L g155 ( 
.A1(n_117),
.A2(n_109),
.B(n_126),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_88),
.Y(n_156)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_156),
.Y(n_162)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_114),
.Y(n_157)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_157),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_111),
.B(n_8),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_2),
.Y(n_159)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_159),
.Y(n_166)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_160),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_173),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_117),
.C(n_129),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_3),
.C(n_5),
.Y(n_194)
);

NOR3xp33_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_121),
.C(n_132),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_182),
.Y(n_183)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_175),
.Y(n_190)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_137),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_179),
.B(n_181),
.Y(n_195)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_141),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_138),
.Y(n_185)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_185),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_171),
.A2(n_144),
.B1(n_155),
.B2(n_148),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_186),
.A2(n_189),
.B1(n_192),
.B2(n_162),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_163),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_187),
.Y(n_208)
);

AOI322xp5_ASAP7_75t_L g188 ( 
.A1(n_173),
.A2(n_155),
.A3(n_153),
.B1(n_140),
.B2(n_159),
.C1(n_158),
.C2(n_150),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_178),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_161),
.A2(n_155),
.B1(n_152),
.B2(n_143),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_176),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_191),
.A2(n_196),
.B(n_197),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_161),
.A2(n_155),
.B1(n_157),
.B2(n_12),
.Y(n_192)
);

A2O1A1O1Ixp25_ASAP7_75t_L g193 ( 
.A1(n_168),
.A2(n_16),
.B(n_11),
.C(n_12),
.D(n_13),
.Y(n_193)
);

A2O1A1O1Ixp25_ASAP7_75t_L g214 ( 
.A1(n_193),
.A2(n_14),
.B(n_177),
.C(n_6),
.D(n_7),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_178),
.C(n_166),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_164),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_198),
.Y(n_202)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_199),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_180),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_200),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_203),
.A2(n_214),
.B1(n_166),
.B2(n_192),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_195),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_209),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_212),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_170),
.Y(n_207)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_207),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_182),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_190),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_204),
.A2(n_191),
.B1(n_179),
.B2(n_162),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_218),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_184),
.C(n_197),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_220),
.C(n_224),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_208),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_219),
.B(n_201),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_212),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_209),
.A2(n_186),
.B1(n_175),
.B2(n_174),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_225),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_190),
.C(n_199),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_227),
.B(n_230),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_222),
.A2(n_206),
.B(n_211),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_228),
.A2(n_227),
.B(n_230),
.Y(n_238)
);

MAJx2_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_224),
.C(n_217),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_229),
.B(n_218),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_219),
.B(n_202),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_223),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_232),
.B(n_181),
.Y(n_236)
);

MAJx2_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_238),
.C(n_165),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_226),
.A2(n_193),
.B1(n_214),
.B2(n_167),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_239),
.Y(n_243)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_236),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_165),
.Y(n_239)
);

AOI21x1_ASAP7_75t_L g240 ( 
.A1(n_237),
.A2(n_233),
.B(n_194),
.Y(n_240)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_240),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_242),
.A2(n_234),
.B(n_5),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_245),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_243),
.Y(n_246)
);

OAI21x1_ASAP7_75t_SL g247 ( 
.A1(n_246),
.A2(n_241),
.B(n_6),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_247),
.A2(n_244),
.B1(n_3),
.B2(n_7),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_248),
.Y(n_250)
);


endmodule