module fake_jpeg_9681_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_21),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_37),
.B(n_42),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_0),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_0),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_18),
.C(n_32),
.Y(n_68)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_19),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_68),
.Y(n_80)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_60),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_46),
.A2(n_27),
.B1(n_28),
.B2(n_25),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_28),
.B1(n_46),
.B2(n_48),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx6_ASAP7_75t_SL g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

NAND3xp33_ASAP7_75t_SL g62 ( 
.A(n_41),
.B(n_19),
.C(n_35),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_47),
.Y(n_96)
);

CKINVDCx9p33_ASAP7_75t_R g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_64),
.B(n_67),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_42),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_44),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_74),
.B(n_78),
.C(n_83),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_75),
.A2(n_82),
.B1(n_70),
.B2(n_53),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_44),
.Y(n_78)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_84),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_48),
.B1(n_28),
.B2(n_25),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_42),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_55),
.A2(n_19),
.B1(n_30),
.B2(n_32),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_91),
.B1(n_95),
.B2(n_31),
.Y(n_102)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

BUFx2_ASAP7_75t_SL g107 ( 
.A(n_87),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_53),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_93),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_55),
.A2(n_30),
.B1(n_18),
.B2(n_23),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_67),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_96),
.A2(n_93),
.B(n_84),
.Y(n_129)
);

AO22x2_ASAP7_75t_L g97 ( 
.A1(n_50),
.A2(n_38),
.B1(n_43),
.B2(n_45),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_97),
.A2(n_45),
.B1(n_56),
.B2(n_69),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_17),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_99),
.Y(n_127)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_100),
.B(n_117),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx11_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_102),
.A2(n_105),
.B1(n_129),
.B2(n_97),
.Y(n_130)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_106),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_76),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_109),
.Y(n_148)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_110),
.Y(n_131)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_70),
.B1(n_99),
.B2(n_75),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_76),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_90),
.A2(n_53),
.B1(n_70),
.B2(n_39),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_119),
.A2(n_79),
.B1(n_51),
.B2(n_81),
.Y(n_151)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_86),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_125),
.Y(n_140)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_126),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_130),
.A2(n_137),
.B1(n_66),
.B2(n_111),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_74),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_139),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_80),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_134),
.A2(n_149),
.B(n_37),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_78),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_80),
.C(n_51),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_142),
.B(n_147),
.C(n_153),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_83),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_104),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_105),
.B(n_80),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_100),
.B(n_72),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_151),
.A2(n_121),
.B1(n_112),
.B2(n_126),
.Y(n_171)
);

AND2x6_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_15),
.Y(n_152)
);

AOI32xp33_ASAP7_75t_L g159 ( 
.A1(n_152),
.A2(n_144),
.A3(n_140),
.B1(n_33),
.B2(n_34),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_39),
.Y(n_153)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_165),
.Y(n_190)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_160),
.Y(n_193)
);

OAI32xp33_ASAP7_75t_L g158 ( 
.A1(n_147),
.A2(n_128),
.A3(n_113),
.B1(n_119),
.B2(n_115),
.Y(n_158)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

NAND3xp33_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_10),
.C(n_15),
.Y(n_184)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_151),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_162),
.B(n_173),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_101),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_168),
.C(n_172),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_135),
.A2(n_29),
.B(n_49),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_164),
.A2(n_167),
.B(n_179),
.Y(n_195)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_135),
.A2(n_49),
.B(n_20),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_40),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_169),
.B(n_24),
.Y(n_200)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_176),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_171),
.A2(n_174),
.B1(n_177),
.B2(n_150),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_104),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_137),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_26),
.Y(n_212)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_155),
.A2(n_145),
.B1(n_136),
.B2(n_146),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_116),
.Y(n_178)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_154),
.A2(n_107),
.B(n_120),
.Y(n_179)
);

OA21x2_ASAP7_75t_L g180 ( 
.A1(n_154),
.A2(n_155),
.B(n_134),
.Y(n_180)
);

AO21x1_ASAP7_75t_L g204 ( 
.A1(n_180),
.A2(n_181),
.B(n_58),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_152),
.A2(n_57),
.B(n_59),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_138),
.B(n_103),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_183),
.B(n_131),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_184),
.B(n_201),
.Y(n_220)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_170),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_185),
.B(n_87),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_187),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_175),
.A2(n_138),
.B1(n_146),
.B2(n_132),
.Y(n_188)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_188),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_162),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_189),
.B(n_205),
.Y(n_235)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_191),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_157),
.A2(n_111),
.B1(n_148),
.B2(n_109),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_194),
.A2(n_166),
.B1(n_158),
.B2(n_31),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_173),
.A2(n_150),
.B1(n_153),
.B2(n_17),
.Y(n_197)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_197),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_120),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_206),
.C(n_182),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_200),
.A2(n_204),
.B(n_208),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_160),
.B(n_110),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_203),
.Y(n_219)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_171),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_167),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_161),
.C(n_168),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_169),
.B(n_33),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_210),
.Y(n_221)
);

AND2x6_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_16),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_178),
.Y(n_210)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_212),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_206),
.C(n_199),
.Y(n_240)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_217),
.B(n_218),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_193),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_189),
.B(n_161),
.Y(n_222)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_222),
.Y(n_248)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_211),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_223),
.B(n_233),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_172),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_225),
.C(n_186),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_164),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_180),
.Y(n_226)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_205),
.Y(n_227)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_227),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_228),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_229),
.A2(n_231),
.B1(n_200),
.B2(n_207),
.Y(n_246)
);

INVx8_ASAP7_75t_L g231 ( 
.A(n_209),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_181),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_185),
.Y(n_234)
);

OA22x2_ASAP7_75t_L g247 ( 
.A1(n_234),
.A2(n_239),
.B1(n_36),
.B2(n_34),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_198),
.B(n_210),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_236),
.B(n_238),
.Y(n_258)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_190),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_202),
.B(n_0),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_242),
.C(n_243),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_244),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_186),
.C(n_195),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_225),
.C(n_236),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_226),
.B(n_195),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_197),
.C(n_203),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_259),
.C(n_261),
.Y(n_269)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_246),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_247),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_212),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_252),
.Y(n_279)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_234),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_231),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_204),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_237),
.A2(n_208),
.B1(n_209),
.B2(n_66),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_253),
.A2(n_221),
.B1(n_215),
.B2(n_217),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_36),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_220),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_22),
.C(n_65),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_222),
.B(n_65),
.C(n_61),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_61),
.C(n_59),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_219),
.C(n_216),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_254),
.A2(n_237),
.B1(n_229),
.B2(n_230),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_263),
.A2(n_280),
.B1(n_260),
.B2(n_26),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_219),
.Y(n_265)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_265),
.Y(n_285)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_266),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_255),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_271),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_244),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_257),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_277),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_215),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_275),
.B(n_276),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_227),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_258),
.Y(n_277)
);

OAI321xp33_ASAP7_75t_L g284 ( 
.A1(n_278),
.A2(n_247),
.A3(n_274),
.B1(n_239),
.B2(n_263),
.C(n_265),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_245),
.A2(n_216),
.B1(n_213),
.B2(n_239),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_270),
.C(n_243),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_289),
.C(n_269),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_272),
.A2(n_248),
.B1(n_242),
.B2(n_213),
.Y(n_282)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_282),
.Y(n_298)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_283),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_284),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_279),
.B(n_241),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_293),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_247),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_269),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_291),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_264),
.B(n_57),
.Y(n_293)
);

A2O1A1Ixp33_ASAP7_75t_L g294 ( 
.A1(n_265),
.A2(n_9),
.B(n_14),
.C(n_13),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_294),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_296),
.B(n_304),
.C(n_309),
.Y(n_317)
);

OAI21xp33_ASAP7_75t_L g299 ( 
.A1(n_285),
.A2(n_264),
.B(n_278),
.Y(n_299)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_299),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_294),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_301),
.B(n_307),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_303),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_295),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_293),
.C(n_287),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_292),
.A2(n_123),
.B1(n_57),
.B2(n_6),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_305),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_288),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_286),
.C(n_1),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_308),
.A2(n_5),
.B1(n_11),
.B2(n_10),
.Y(n_310)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_310),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_4),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_316),
.Y(n_323)
);

BUFx12f_ASAP7_75t_SL g313 ( 
.A(n_296),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_313),
.B(n_304),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_297),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_300),
.B(n_4),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_318),
.B(n_300),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_321),
.B(n_322),
.C(n_327),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_313),
.A2(n_298),
.B(n_306),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_324),
.A2(n_325),
.B(n_326),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_305),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_317),
.A2(n_3),
.B(n_6),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_311),
.B(n_319),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_325),
.A2(n_312),
.B(n_315),
.Y(n_328)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_328),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_323),
.A2(n_315),
.B(n_3),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_331),
.A2(n_332),
.B(n_7),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_323),
.A2(n_320),
.B(n_7),
.Y(n_332)
);

AOI31xp33_ASAP7_75t_L g335 ( 
.A1(n_333),
.A2(n_330),
.A3(n_329),
.B(n_7),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_334),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_0),
.C(n_1),
.Y(n_337)
);

AOI221xp5_ASAP7_75t_SL g338 ( 
.A1(n_337),
.A2(n_1),
.B1(n_2),
.B2(n_43),
.C(n_313),
.Y(n_338)
);

BUFx24_ASAP7_75t_SL g339 ( 
.A(n_338),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_339),
.A2(n_2),
.B(n_336),
.Y(n_340)
);


endmodule