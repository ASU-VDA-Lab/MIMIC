module real_aes_7046_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_756;
wire n_404;
wire n_288;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g258 ( .A1(n_0), .A2(n_259), .B(n_260), .C(n_263), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_1), .B(n_247), .Y(n_264) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_2), .B(n_109), .C(n_110), .Y(n_108) );
INVx1_ASAP7_75t_L g460 ( .A(n_2), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_3), .B(n_175), .Y(n_174) );
A2O1A1Ixp33_ASAP7_75t_L g551 ( .A1(n_4), .A2(n_136), .B(n_139), .C(n_552), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_5), .A2(n_131), .B(n_576), .Y(n_575) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_6), .A2(n_131), .B(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_7), .B(n_247), .Y(n_582) );
AO21x2_ASAP7_75t_L g202 ( .A1(n_8), .A2(n_166), .B(n_203), .Y(n_202) );
AND2x6_ASAP7_75t_L g136 ( .A(n_9), .B(n_137), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_10), .A2(n_136), .B(n_139), .C(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g520 ( .A(n_11), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_12), .B(n_40), .Y(n_114) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_13), .A2(n_468), .B1(n_469), .B2(n_470), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_13), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_14), .B(n_223), .Y(n_554) );
INVx1_ASAP7_75t_L g157 ( .A(n_15), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_16), .B(n_175), .Y(n_209) );
A2O1A1Ixp33_ASAP7_75t_L g537 ( .A1(n_17), .A2(n_176), .B(n_538), .C(n_540), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_18), .B(n_247), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_19), .B(n_151), .Y(n_511) );
A2O1A1Ixp33_ASAP7_75t_L g138 ( .A1(n_20), .A2(n_139), .B(n_142), .C(n_150), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_21), .A2(n_211), .B(n_262), .C(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_22), .B(n_223), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_23), .A2(n_56), .B1(n_450), .B2(n_451), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_23), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_24), .B(n_223), .Y(n_493) );
CKINVDCx16_ASAP7_75t_R g567 ( .A(n_25), .Y(n_567) );
INVx1_ASAP7_75t_L g492 ( .A(n_26), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_27), .A2(n_139), .B(n_150), .C(n_206), .Y(n_205) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_28), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_29), .Y(n_550) );
INVx1_ASAP7_75t_L g508 ( .A(n_30), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_31), .A2(n_131), .B(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g134 ( .A(n_32), .Y(n_134) );
A2O1A1Ixp33_ASAP7_75t_L g187 ( .A1(n_33), .A2(n_179), .B(n_188), .C(n_190), .Y(n_187) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_34), .Y(n_557) );
A2O1A1Ixp33_ASAP7_75t_L g578 ( .A1(n_35), .A2(n_262), .B(n_579), .C(n_581), .Y(n_578) );
INVxp67_ASAP7_75t_L g509 ( .A(n_36), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_37), .B(n_208), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_38), .A2(n_139), .B(n_150), .C(n_491), .Y(n_490) );
CKINVDCx14_ASAP7_75t_R g577 ( .A(n_39), .Y(n_577) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_41), .A2(n_263), .B(n_518), .C(n_519), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_42), .B(n_130), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_43), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_44), .B(n_175), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_45), .B(n_131), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_46), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_47), .Y(n_505) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_48), .A2(n_179), .B(n_188), .C(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_49), .B(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g261 ( .A(n_50), .Y(n_261) );
OAI22xp5_ASAP7_75t_SL g447 ( .A1(n_51), .A2(n_448), .B1(n_449), .B2(n_452), .Y(n_447) );
CKINVDCx16_ASAP7_75t_R g452 ( .A(n_51), .Y(n_452) );
AOI222xp33_ASAP7_75t_L g465 ( .A1(n_52), .A2(n_466), .B1(n_467), .B2(n_476), .C1(n_755), .C2(n_759), .Y(n_465) );
INVx1_ASAP7_75t_L g233 ( .A(n_53), .Y(n_233) );
INVx1_ASAP7_75t_L g526 ( .A(n_54), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_55), .B(n_131), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_56), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_57), .Y(n_159) );
CKINVDCx14_ASAP7_75t_R g516 ( .A(n_58), .Y(n_516) );
INVx1_ASAP7_75t_L g137 ( .A(n_59), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_60), .B(n_131), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_61), .B(n_247), .Y(n_246) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_62), .A2(n_149), .B(n_172), .C(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g156 ( .A(n_63), .Y(n_156) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_64), .A2(n_103), .B1(n_472), .B2(n_473), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_64), .Y(n_473) );
INVx1_ASAP7_75t_SL g580 ( .A(n_65), .Y(n_580) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_66), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_67), .B(n_175), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_68), .B(n_247), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_69), .B(n_176), .Y(n_221) );
INVx1_ASAP7_75t_L g570 ( .A(n_70), .Y(n_570) );
CKINVDCx16_ASAP7_75t_R g257 ( .A(n_71), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_72), .B(n_144), .Y(n_143) );
A2O1A1Ixp33_ASAP7_75t_L g169 ( .A1(n_73), .A2(n_139), .B(n_170), .C(n_179), .Y(n_169) );
CKINVDCx16_ASAP7_75t_R g242 ( .A(n_74), .Y(n_242) );
INVx1_ASAP7_75t_L g112 ( .A(n_75), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_76), .A2(n_131), .B(n_515), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g573 ( .A(n_77), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_78), .A2(n_131), .B(n_535), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_79), .A2(n_105), .B1(n_115), .B2(n_765), .Y(n_104) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_80), .A2(n_130), .B(n_504), .Y(n_503) );
CKINVDCx16_ASAP7_75t_R g489 ( .A(n_81), .Y(n_489) );
INVx1_ASAP7_75t_L g536 ( .A(n_82), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_83), .B(n_147), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_84), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_85), .A2(n_131), .B(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g539 ( .A(n_86), .Y(n_539) );
INVx2_ASAP7_75t_L g154 ( .A(n_87), .Y(n_154) );
INVx1_ASAP7_75t_L g553 ( .A(n_88), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_89), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_90), .B(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g109 ( .A(n_91), .Y(n_109) );
OR2x2_ASAP7_75t_L g457 ( .A(n_91), .B(n_458), .Y(n_457) );
OR2x2_ASAP7_75t_L g479 ( .A(n_91), .B(n_459), .Y(n_479) );
OAI22xp5_ASAP7_75t_SL g470 ( .A1(n_92), .A2(n_471), .B1(n_474), .B2(n_475), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_92), .Y(n_475) );
A2O1A1Ixp33_ASAP7_75t_L g568 ( .A1(n_93), .A2(n_139), .B(n_179), .C(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_94), .B(n_131), .Y(n_186) );
INVx1_ASAP7_75t_L g191 ( .A(n_95), .Y(n_191) );
INVxp67_ASAP7_75t_L g245 ( .A(n_96), .Y(n_245) );
XNOR2xp5_ASAP7_75t_L g119 ( .A(n_97), .B(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_97), .B(n_166), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_98), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g171 ( .A(n_99), .Y(n_171) );
INVx1_ASAP7_75t_L g217 ( .A(n_100), .Y(n_217) );
INVx2_ASAP7_75t_L g529 ( .A(n_101), .Y(n_529) );
AND2x2_ASAP7_75t_L g235 ( .A(n_102), .B(n_153), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_103), .Y(n_472) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_107), .Y(n_767) );
OR2x2_ASAP7_75t_SL g107 ( .A(n_108), .B(n_113), .Y(n_107) );
OR2x2_ASAP7_75t_L g480 ( .A(n_109), .B(n_459), .Y(n_480) );
NOR2x2_ASAP7_75t_L g761 ( .A(n_109), .B(n_458), .Y(n_761) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
INVxp67_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x2_ASAP7_75t_L g459 ( .A(n_114), .B(n_460), .Y(n_459) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_118), .B(n_464), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g764 ( .A(n_117), .Y(n_764) );
OAI21xp5_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_454), .B(n_461), .Y(n_118) );
OAI22xp5_ASAP7_75t_SL g120 ( .A1(n_121), .A2(n_446), .B1(n_447), .B2(n_453), .Y(n_120) );
OAI22xp5_ASAP7_75t_SL g755 ( .A1(n_121), .A2(n_482), .B1(n_756), .B2(n_757), .Y(n_755) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx2_ASAP7_75t_L g453 ( .A(n_122), .Y(n_453) );
AND3x1_ASAP7_75t_L g122 ( .A(n_123), .B(n_350), .C(n_407), .Y(n_122) );
NOR3xp33_ASAP7_75t_L g123 ( .A(n_124), .B(n_295), .C(n_331), .Y(n_123) );
OAI211xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_197), .B(n_249), .C(n_282), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_161), .Y(n_125) );
HB1xp67_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x4_ASAP7_75t_L g252 ( .A(n_127), .B(n_253), .Y(n_252) );
INVx5_ASAP7_75t_L g281 ( .A(n_127), .Y(n_281) );
AND2x2_ASAP7_75t_L g354 ( .A(n_127), .B(n_270), .Y(n_354) );
AND2x2_ASAP7_75t_L g392 ( .A(n_127), .B(n_298), .Y(n_392) );
AND2x2_ASAP7_75t_L g412 ( .A(n_127), .B(n_254), .Y(n_412) );
OR2x6_ASAP7_75t_L g127 ( .A(n_128), .B(n_158), .Y(n_127) );
AOI21xp5_ASAP7_75t_SL g128 ( .A1(n_129), .A2(n_138), .B(n_151), .Y(n_128) );
BUFx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_136), .Y(n_131) );
NAND2x1p5_ASAP7_75t_L g218 ( .A(n_132), .B(n_136), .Y(n_218) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_135), .Y(n_132) );
INVx1_ASAP7_75t_L g149 ( .A(n_133), .Y(n_149) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g140 ( .A(n_134), .Y(n_140) );
INVx1_ASAP7_75t_L g212 ( .A(n_134), .Y(n_212) );
INVx1_ASAP7_75t_L g141 ( .A(n_135), .Y(n_141) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_135), .Y(n_145) );
INVx3_ASAP7_75t_L g176 ( .A(n_135), .Y(n_176) );
INVx1_ASAP7_75t_L g208 ( .A(n_135), .Y(n_208) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_135), .Y(n_223) );
BUFx3_ASAP7_75t_L g150 ( .A(n_136), .Y(n_150) );
INVx4_ASAP7_75t_SL g180 ( .A(n_136), .Y(n_180) );
INVx5_ASAP7_75t_L g189 ( .A(n_139), .Y(n_189) );
AND2x6_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_140), .Y(n_178) );
BUFx3_ASAP7_75t_L g194 ( .A(n_140), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_146), .B(n_148), .Y(n_142) );
INVx2_ASAP7_75t_L g147 ( .A(n_144), .Y(n_147) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx4_ASAP7_75t_L g173 ( .A(n_145), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_L g190 ( .A1(n_147), .A2(n_191), .B(n_192), .C(n_193), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_L g232 ( .A1(n_147), .A2(n_193), .B(n_233), .C(n_234), .Y(n_232) );
O2A1O1Ixp5_ASAP7_75t_L g552 ( .A1(n_147), .A2(n_553), .B(n_554), .C(n_555), .Y(n_552) );
O2A1O1Ixp33_ASAP7_75t_L g569 ( .A1(n_147), .A2(n_555), .B(n_570), .C(n_571), .Y(n_569) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_148), .A2(n_175), .B(n_492), .C(n_493), .Y(n_491) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_149), .B(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_152), .B(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g160 ( .A(n_153), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_153), .A2(n_186), .B(n_187), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_153), .A2(n_230), .B(n_231), .Y(n_229) );
O2A1O1Ixp33_ASAP7_75t_L g488 ( .A1(n_153), .A2(n_218), .B(n_489), .C(n_490), .Y(n_488) );
OA21x2_ASAP7_75t_L g513 ( .A1(n_153), .A2(n_514), .B(n_521), .Y(n_513) );
AND2x2_ASAP7_75t_SL g153 ( .A(n_154), .B(n_155), .Y(n_153) );
AND2x2_ASAP7_75t_L g167 ( .A(n_154), .B(n_155), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
AO21x2_ASAP7_75t_L g548 ( .A1(n_160), .A2(n_549), .B(n_556), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_161), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g161 ( .A(n_162), .B(n_184), .Y(n_161) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_162), .Y(n_293) );
AND2x2_ASAP7_75t_L g307 ( .A(n_162), .B(n_253), .Y(n_307) );
INVx1_ASAP7_75t_L g330 ( .A(n_162), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_162), .B(n_281), .Y(n_369) );
OR2x2_ASAP7_75t_L g406 ( .A(n_162), .B(n_251), .Y(n_406) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_163), .Y(n_342) );
AND2x2_ASAP7_75t_L g349 ( .A(n_163), .B(n_254), .Y(n_349) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AND2x2_ASAP7_75t_L g270 ( .A(n_164), .B(n_254), .Y(n_270) );
BUFx2_ASAP7_75t_L g298 ( .A(n_164), .Y(n_298) );
AO21x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_168), .B(n_182), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_165), .B(n_183), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_165), .B(n_196), .Y(n_195) );
AO21x2_ASAP7_75t_L g215 ( .A1(n_165), .A2(n_216), .B(n_224), .Y(n_215) );
INVx3_ASAP7_75t_L g247 ( .A(n_165), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_165), .B(n_495), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_165), .B(n_557), .Y(n_556) );
AO21x2_ASAP7_75t_L g565 ( .A1(n_165), .A2(n_566), .B(n_572), .Y(n_565) );
INVx4_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_166), .A2(n_204), .B(n_205), .Y(n_203) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_166), .Y(n_239) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g226 ( .A(n_167), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_169), .B(n_181), .Y(n_168) );
O2A1O1Ixp33_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_174), .C(n_177), .Y(n_170) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
OAI22xp33_ASAP7_75t_L g507 ( .A1(n_173), .A2(n_175), .B1(n_508), .B2(n_509), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_173), .B(n_529), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_173), .B(n_539), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_175), .B(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g259 ( .A(n_175), .Y(n_259) );
INVx5_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_176), .B(n_520), .Y(n_519) );
HB1xp67_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx3_ASAP7_75t_L g581 ( .A(n_178), .Y(n_581) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
O2A1O1Ixp33_ASAP7_75t_L g241 ( .A1(n_180), .A2(n_189), .B(n_242), .C(n_243), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_SL g256 ( .A1(n_180), .A2(n_189), .B(n_257), .C(n_258), .Y(n_256) );
O2A1O1Ixp33_ASAP7_75t_SL g504 ( .A1(n_180), .A2(n_189), .B(n_505), .C(n_506), .Y(n_504) );
O2A1O1Ixp33_ASAP7_75t_SL g515 ( .A1(n_180), .A2(n_189), .B(n_516), .C(n_517), .Y(n_515) );
O2A1O1Ixp33_ASAP7_75t_SL g525 ( .A1(n_180), .A2(n_189), .B(n_526), .C(n_527), .Y(n_525) );
O2A1O1Ixp33_ASAP7_75t_SL g535 ( .A1(n_180), .A2(n_189), .B(n_536), .C(n_537), .Y(n_535) );
O2A1O1Ixp33_ASAP7_75t_L g576 ( .A1(n_180), .A2(n_189), .B(n_577), .C(n_578), .Y(n_576) );
INVx5_ASAP7_75t_L g251 ( .A(n_184), .Y(n_251) );
BUFx2_ASAP7_75t_L g274 ( .A(n_184), .Y(n_274) );
AND2x2_ASAP7_75t_L g431 ( .A(n_184), .B(n_285), .Y(n_431) );
OR2x6_ASAP7_75t_L g184 ( .A(n_185), .B(n_195), .Y(n_184) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g263 ( .A(n_194), .Y(n_263) );
INVx1_ASAP7_75t_L g540 ( .A(n_194), .Y(n_540) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NAND2xp33_ASAP7_75t_L g198 ( .A(n_199), .B(n_236), .Y(n_198) );
OAI221xp5_ASAP7_75t_L g331 ( .A1(n_199), .A2(n_332), .B1(n_339), .B2(n_340), .C(n_343), .Y(n_331) );
OR2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_213), .Y(n_199) );
AND2x2_ASAP7_75t_L g237 ( .A(n_200), .B(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_200), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_SL g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g266 ( .A(n_201), .B(n_214), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_201), .B(n_215), .Y(n_276) );
OR2x2_ASAP7_75t_L g287 ( .A(n_201), .B(n_238), .Y(n_287) );
AND2x2_ASAP7_75t_L g290 ( .A(n_201), .B(n_278), .Y(n_290) );
AND2x2_ASAP7_75t_L g306 ( .A(n_201), .B(n_227), .Y(n_306) );
OR2x2_ASAP7_75t_L g322 ( .A(n_201), .B(n_215), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_201), .B(n_238), .Y(n_384) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_202), .B(n_227), .Y(n_376) );
AND2x2_ASAP7_75t_L g379 ( .A(n_202), .B(n_215), .Y(n_379) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_209), .B(n_210), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_210), .A2(n_221), .B(n_222), .Y(n_220) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx3_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
OR2x2_ASAP7_75t_L g300 ( .A(n_213), .B(n_287), .Y(n_300) );
INVx2_ASAP7_75t_L g326 ( .A(n_213), .Y(n_326) );
OR2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_227), .Y(n_213) );
AND2x2_ASAP7_75t_L g248 ( .A(n_214), .B(n_228), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_214), .B(n_238), .Y(n_305) );
OR2x2_ASAP7_75t_L g316 ( .A(n_214), .B(n_228), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_214), .B(n_278), .Y(n_375) );
OAI221xp5_ASAP7_75t_L g408 ( .A1(n_214), .A2(n_409), .B1(n_411), .B2(n_413), .C(n_416), .Y(n_408) );
INVx5_ASAP7_75t_SL g214 ( .A(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_215), .B(n_238), .Y(n_347) );
OAI21xp5_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_218), .B(n_219), .Y(n_216) );
OAI21xp5_ASAP7_75t_L g549 ( .A1(n_218), .A2(n_550), .B(n_551), .Y(n_549) );
OAI21xp5_ASAP7_75t_L g566 ( .A1(n_218), .A2(n_567), .B(n_568), .Y(n_566) );
INVx4_ASAP7_75t_L g262 ( .A(n_223), .Y(n_262) );
INVx2_ASAP7_75t_L g518 ( .A(n_223), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_225), .B(n_226), .Y(n_224) );
INVx2_ASAP7_75t_L g501 ( .A(n_226), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_227), .B(n_278), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_227), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g294 ( .A(n_227), .B(n_266), .Y(n_294) );
OR2x2_ASAP7_75t_L g338 ( .A(n_227), .B(n_238), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_227), .B(n_290), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_227), .B(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g403 ( .A(n_227), .B(n_404), .Y(n_403) );
INVx5_ASAP7_75t_SL g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_SL g267 ( .A(n_228), .B(n_237), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_SL g271 ( .A1(n_228), .A2(n_272), .B(n_275), .C(n_279), .Y(n_271) );
OR2x2_ASAP7_75t_L g309 ( .A(n_228), .B(n_305), .Y(n_309) );
OR2x2_ASAP7_75t_L g345 ( .A(n_228), .B(n_287), .Y(n_345) );
OAI311xp33_ASAP7_75t_L g351 ( .A1(n_228), .A2(n_290), .A3(n_352), .B1(n_355), .C1(n_362), .Y(n_351) );
AND2x2_ASAP7_75t_L g402 ( .A(n_228), .B(n_238), .Y(n_402) );
AND2x2_ASAP7_75t_L g410 ( .A(n_228), .B(n_265), .Y(n_410) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_228), .Y(n_428) );
AND2x2_ASAP7_75t_L g445 ( .A(n_228), .B(n_266), .Y(n_445) );
OR2x6_ASAP7_75t_L g228 ( .A(n_229), .B(n_235), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_237), .B(n_248), .Y(n_236) );
AND2x2_ASAP7_75t_L g273 ( .A(n_237), .B(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g429 ( .A(n_237), .Y(n_429) );
AND2x2_ASAP7_75t_L g265 ( .A(n_238), .B(n_266), .Y(n_265) );
INVx3_ASAP7_75t_L g278 ( .A(n_238), .Y(n_278) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_238), .Y(n_321) );
INVxp67_ASAP7_75t_L g360 ( .A(n_238), .Y(n_360) );
OA21x2_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_240), .B(n_246), .Y(n_238) );
OA21x2_ASAP7_75t_L g523 ( .A1(n_239), .A2(n_524), .B(n_530), .Y(n_523) );
OA21x2_ASAP7_75t_L g533 ( .A1(n_239), .A2(n_534), .B(n_541), .Y(n_533) );
OA21x2_ASAP7_75t_L g574 ( .A1(n_239), .A2(n_575), .B(n_582), .Y(n_574) );
OA21x2_ASAP7_75t_L g254 ( .A1(n_247), .A2(n_255), .B(n_264), .Y(n_254) );
AND2x2_ASAP7_75t_L g438 ( .A(n_248), .B(n_286), .Y(n_438) );
AOI221xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_265), .B1(n_267), .B2(n_268), .C(n_271), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_251), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g291 ( .A(n_251), .B(n_281), .Y(n_291) );
AND2x2_ASAP7_75t_L g299 ( .A(n_251), .B(n_253), .Y(n_299) );
OR2x2_ASAP7_75t_L g311 ( .A(n_251), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g329 ( .A(n_251), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g353 ( .A(n_251), .B(n_354), .Y(n_353) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_251), .Y(n_373) );
AND2x2_ASAP7_75t_L g425 ( .A(n_251), .B(n_349), .Y(n_425) );
OAI31xp33_ASAP7_75t_L g433 ( .A1(n_251), .A2(n_302), .A3(n_401), .B(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_252), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_SL g397 ( .A(n_252), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_252), .B(n_406), .Y(n_405) );
AND2x4_ASAP7_75t_L g285 ( .A(n_253), .B(n_281), .Y(n_285) );
INVx1_ASAP7_75t_L g372 ( .A(n_253), .Y(n_372) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g422 ( .A(n_254), .B(n_281), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_262), .B(n_580), .Y(n_579) );
INVx2_ASAP7_75t_L g555 ( .A(n_263), .Y(n_555) );
INVx1_ASAP7_75t_SL g432 ( .A(n_265), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_266), .B(n_337), .Y(n_336) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_267), .A2(n_379), .B1(n_417), .B2(n_420), .Y(n_416) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g280 ( .A(n_270), .B(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g339 ( .A(n_270), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_270), .B(n_291), .Y(n_444) );
INVx1_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g414 ( .A(n_273), .B(n_415), .Y(n_414) );
AOI21xp5_ASAP7_75t_L g332 ( .A1(n_274), .A2(n_333), .B(n_335), .Y(n_332) );
OR2x2_ASAP7_75t_L g340 ( .A(n_274), .B(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g361 ( .A(n_274), .B(n_349), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_274), .B(n_372), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_274), .B(n_412), .Y(n_411) );
OAI221xp5_ASAP7_75t_SL g388 ( .A1(n_275), .A2(n_389), .B1(n_394), .B2(n_397), .C(n_398), .Y(n_388) );
OR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
OR2x2_ASAP7_75t_L g365 ( .A(n_276), .B(n_338), .Y(n_365) );
INVx1_ASAP7_75t_L g404 ( .A(n_276), .Y(n_404) );
INVx2_ASAP7_75t_L g380 ( .A(n_277), .Y(n_380) );
INVx1_ASAP7_75t_L g314 ( .A(n_278), .Y(n_314) );
INVx1_ASAP7_75t_SL g279 ( .A(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g319 ( .A(n_281), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_281), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g348 ( .A(n_281), .B(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g436 ( .A(n_281), .B(n_406), .Y(n_436) );
AOI222xp33_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_286), .B1(n_288), .B2(n_291), .C1(n_292), .C2(n_294), .Y(n_282) );
INVxp67_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g292 ( .A(n_285), .B(n_293), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_285), .A2(n_335), .B1(n_363), .B2(n_364), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_285), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
OAI21xp33_ASAP7_75t_SL g323 ( .A1(n_294), .A2(n_324), .B(n_327), .Y(n_323) );
OAI211xp5_ASAP7_75t_SL g295 ( .A1(n_296), .A2(n_300), .B(n_301), .C(n_323), .Y(n_295) );
INVxp67_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
AOI221xp5_ASAP7_75t_L g301 ( .A1(n_299), .A2(n_302), .B1(n_307), .B2(n_308), .C(n_310), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_299), .B(n_387), .Y(n_386) );
INVxp67_ASAP7_75t_L g393 ( .A(n_299), .Y(n_393) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
AND2x2_ASAP7_75t_L g395 ( .A(n_304), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g312 ( .A(n_307), .Y(n_312) );
AND2x2_ASAP7_75t_L g318 ( .A(n_307), .B(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OAI22xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_313), .B1(n_317), .B2(n_320), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_314), .B(n_326), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_315), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g415 ( .A(n_319), .Y(n_415) );
AND2x2_ASAP7_75t_L g434 ( .A(n_319), .B(n_349), .Y(n_434) );
OR2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_326), .B(n_383), .Y(n_442) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_329), .B(n_397), .Y(n_440) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g363 ( .A(n_341), .Y(n_363) );
BUFx2_ASAP7_75t_L g387 ( .A(n_342), .Y(n_387) );
OAI21xp5_ASAP7_75t_SL g343 ( .A1(n_344), .A2(n_346), .B(n_348), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NOR3xp33_ASAP7_75t_L g350 ( .A(n_351), .B(n_366), .C(n_388), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OAI21xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_358), .B(n_361), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
A2O1A1Ixp33_ASAP7_75t_SL g366 ( .A1(n_367), .A2(n_370), .B(n_374), .C(n_377), .Y(n_366) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_367), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NOR2xp67_ASAP7_75t_SL g371 ( .A(n_372), .B(n_373), .Y(n_371) );
OR2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
INVx1_ASAP7_75t_SL g396 ( .A(n_376), .Y(n_396) );
OAI21xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_381), .B(n_385), .Y(n_377) );
AND2x4_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
AND2x2_ASAP7_75t_L g401 ( .A(n_379), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_391), .B(n_393), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_401), .B1(n_403), .B2(n_405), .Y(n_398) );
INVx2_ASAP7_75t_SL g419 ( .A(n_406), .Y(n_419) );
NOR3xp33_ASAP7_75t_L g407 ( .A(n_408), .B(n_423), .C(n_435), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVxp67_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVxp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_419), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
OAI221xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_426), .B1(n_430), .B2(n_432), .C(n_433), .Y(n_423) );
A2O1A1Ixp33_ASAP7_75t_L g435 ( .A1(n_424), .A2(n_436), .B(n_437), .C(n_439), .Y(n_435) );
INVx1_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
INVxp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_441), .B1(n_443), .B2(n_445), .Y(n_439) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_453), .A2(n_477), .B1(n_480), .B2(n_481), .Y(n_476) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_457), .Y(n_463) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
NAND3xp33_ASAP7_75t_L g464 ( .A(n_461), .B(n_465), .C(n_762), .Y(n_464) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g474 ( .A(n_471), .Y(n_474) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g756 ( .A(n_478), .Y(n_756) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g758 ( .A(n_480), .Y(n_758) );
INVx1_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
OR5x1_ASAP7_75t_L g482 ( .A(n_483), .B(n_649), .C(n_713), .D(n_729), .E(n_744), .Y(n_482) );
NAND4xp25_ASAP7_75t_L g483 ( .A(n_484), .B(n_583), .C(n_610), .D(n_633), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_531), .B(n_542), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_486), .B(n_496), .Y(n_485) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx3_ASAP7_75t_SL g562 ( .A(n_487), .Y(n_562) );
AND2x4_ASAP7_75t_L g596 ( .A(n_487), .B(n_585), .Y(n_596) );
OR2x2_ASAP7_75t_L g606 ( .A(n_487), .B(n_564), .Y(n_606) );
OR2x2_ASAP7_75t_L g652 ( .A(n_487), .B(n_499), .Y(n_652) );
AND2x2_ASAP7_75t_L g666 ( .A(n_487), .B(n_563), .Y(n_666) );
AND2x2_ASAP7_75t_L g709 ( .A(n_487), .B(n_599), .Y(n_709) );
AND2x2_ASAP7_75t_L g716 ( .A(n_487), .B(n_574), .Y(n_716) );
AND2x2_ASAP7_75t_L g735 ( .A(n_487), .B(n_625), .Y(n_735) );
AND2x2_ASAP7_75t_L g753 ( .A(n_487), .B(n_595), .Y(n_753) );
OR2x6_ASAP7_75t_L g487 ( .A(n_488), .B(n_494), .Y(n_487) );
INVx1_ASAP7_75t_L g718 ( .A(n_496), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_497), .B(n_512), .Y(n_496) );
AND2x2_ASAP7_75t_L g628 ( .A(n_497), .B(n_563), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_497), .B(n_648), .Y(n_647) );
AOI32xp33_ASAP7_75t_L g661 ( .A1(n_497), .A2(n_662), .A3(n_665), .B1(n_667), .B2(n_671), .Y(n_661) );
AND2x2_ASAP7_75t_L g731 ( .A(n_497), .B(n_625), .Y(n_731) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g595 ( .A(n_499), .B(n_564), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_499), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g637 ( .A(n_499), .B(n_584), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_499), .B(n_716), .Y(n_715) );
AO21x2_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_502), .B(n_510), .Y(n_499) );
INVx1_ASAP7_75t_L g600 ( .A(n_500), .Y(n_600) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
OA21x2_ASAP7_75t_L g599 ( .A1(n_503), .A2(n_511), .B(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g602 ( .A(n_512), .B(n_546), .Y(n_602) );
AND2x2_ASAP7_75t_L g678 ( .A(n_512), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_SL g750 ( .A(n_512), .Y(n_750) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_522), .Y(n_512) );
OR2x2_ASAP7_75t_L g545 ( .A(n_513), .B(n_523), .Y(n_545) );
AND2x2_ASAP7_75t_L g559 ( .A(n_513), .B(n_560), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_513), .B(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g609 ( .A(n_513), .Y(n_609) );
AND2x2_ASAP7_75t_L g636 ( .A(n_513), .B(n_523), .Y(n_636) );
BUFx3_ASAP7_75t_L g639 ( .A(n_513), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_513), .B(n_614), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_513), .B(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g590 ( .A(n_522), .Y(n_590) );
AND2x2_ASAP7_75t_L g608 ( .A(n_522), .B(n_588), .Y(n_608) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g619 ( .A(n_523), .B(n_533), .Y(n_619) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_523), .Y(n_632) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_532), .B(n_639), .Y(n_689) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_SL g560 ( .A(n_533), .Y(n_560) );
NAND3xp33_ASAP7_75t_L g607 ( .A(n_533), .B(n_608), .C(n_609), .Y(n_607) );
OR2x2_ASAP7_75t_L g615 ( .A(n_533), .B(n_588), .Y(n_615) );
AND2x2_ASAP7_75t_L g635 ( .A(n_533), .B(n_588), .Y(n_635) );
AND2x2_ASAP7_75t_L g679 ( .A(n_533), .B(n_548), .Y(n_679) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_558), .B(n_561), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_544), .B(n_546), .Y(n_543) );
AND2x2_ASAP7_75t_L g754 ( .A(n_544), .B(n_679), .Y(n_754) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_545), .A2(n_652), .B1(n_694), .B2(n_696), .Y(n_693) );
OR2x2_ASAP7_75t_L g700 ( .A(n_545), .B(n_615), .Y(n_700) );
OR2x2_ASAP7_75t_L g724 ( .A(n_545), .B(n_725), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_545), .B(n_644), .Y(n_737) );
AND2x2_ASAP7_75t_L g630 ( .A(n_546), .B(n_631), .Y(n_630) );
AOI21xp5_ASAP7_75t_L g717 ( .A1(n_546), .A2(n_703), .B(n_718), .Y(n_717) );
AOI32xp33_ASAP7_75t_L g738 ( .A1(n_546), .A2(n_628), .A3(n_739), .B1(n_741), .B2(n_742), .Y(n_738) );
OR2x2_ASAP7_75t_L g749 ( .A(n_546), .B(n_750), .Y(n_749) );
CKINVDCx16_ASAP7_75t_R g546 ( .A(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g617 ( .A(n_547), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_547), .B(n_631), .Y(n_696) );
BUFx3_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx4_ASAP7_75t_L g588 ( .A(n_548), .Y(n_588) );
AND2x2_ASAP7_75t_L g654 ( .A(n_548), .B(n_619), .Y(n_654) );
AND3x2_ASAP7_75t_L g663 ( .A(n_548), .B(n_559), .C(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g589 ( .A(n_560), .B(n_590), .Y(n_589) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_560), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_560), .B(n_588), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
AND2x2_ASAP7_75t_L g584 ( .A(n_562), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g624 ( .A(n_562), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g642 ( .A(n_562), .B(n_574), .Y(n_642) );
AND2x2_ASAP7_75t_L g660 ( .A(n_562), .B(n_564), .Y(n_660) );
OR2x2_ASAP7_75t_L g674 ( .A(n_562), .B(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g720 ( .A(n_562), .B(n_648), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_563), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_574), .Y(n_563) );
AND2x2_ASAP7_75t_L g621 ( .A(n_564), .B(n_599), .Y(n_621) );
OR2x2_ASAP7_75t_L g675 ( .A(n_564), .B(n_599), .Y(n_675) );
AND2x2_ASAP7_75t_L g728 ( .A(n_564), .B(n_585), .Y(n_728) );
INVx2_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
BUFx2_ASAP7_75t_L g626 ( .A(n_565), .Y(n_626) );
AND2x2_ASAP7_75t_L g648 ( .A(n_565), .B(n_574), .Y(n_648) );
INVx2_ASAP7_75t_L g585 ( .A(n_574), .Y(n_585) );
INVx1_ASAP7_75t_L g605 ( .A(n_574), .Y(n_605) );
AOI211xp5_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_586), .B(n_591), .C(n_603), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_584), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g747 ( .A(n_584), .Y(n_747) );
AND2x2_ASAP7_75t_L g625 ( .A(n_585), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_588), .B(n_589), .Y(n_597) );
INVx1_ASAP7_75t_L g682 ( .A(n_588), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_588), .B(n_609), .Y(n_706) );
AND2x2_ASAP7_75t_L g722 ( .A(n_588), .B(n_636), .Y(n_722) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_589), .B(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g613 ( .A(n_590), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_597), .B1(n_598), .B2(n_601), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_594), .B(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_595), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g620 ( .A(n_596), .B(n_621), .Y(n_620) );
AOI221xp5_ASAP7_75t_SL g685 ( .A1(n_596), .A2(n_638), .B1(n_686), .B2(n_691), .C(n_693), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_596), .B(n_659), .Y(n_692) );
INVx1_ASAP7_75t_L g752 ( .A(n_598), .Y(n_752) );
BUFx3_ASAP7_75t_L g659 ( .A(n_599), .Y(n_659) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AOI21xp33_ASAP7_75t_SL g603 ( .A1(n_604), .A2(n_606), .B(n_607), .Y(n_603) );
INVx1_ASAP7_75t_L g668 ( .A(n_605), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_605), .B(n_659), .Y(n_712) );
INVx1_ASAP7_75t_L g669 ( .A(n_606), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_606), .B(n_659), .Y(n_670) );
INVxp67_ASAP7_75t_L g690 ( .A(n_608), .Y(n_690) );
AND2x2_ASAP7_75t_L g631 ( .A(n_609), .B(n_632), .Y(n_631) );
O2A1O1Ixp33_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_616), .B(n_620), .C(n_622), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
INVx1_ASAP7_75t_SL g645 ( .A(n_613), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_614), .B(n_645), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_614), .B(n_636), .Y(n_687) );
INVx2_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_617), .A2(n_623), .B1(n_627), .B2(n_629), .Y(n_622) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g638 ( .A(n_619), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g683 ( .A(n_619), .B(n_684), .Y(n_683) );
OAI21xp33_ASAP7_75t_L g686 ( .A1(n_621), .A2(n_687), .B(n_688), .Y(n_686) );
INVx1_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
AOI221xp5_ASAP7_75t_L g633 ( .A1(n_625), .A2(n_634), .B1(n_637), .B2(n_638), .C(n_640), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_625), .B(n_659), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_625), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g741 ( .A(n_631), .Y(n_741) );
INVxp67_ASAP7_75t_L g664 ( .A(n_632), .Y(n_664) );
INVx1_ASAP7_75t_L g671 ( .A(n_634), .Y(n_671) );
AND2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
AND2x2_ASAP7_75t_L g710 ( .A(n_635), .B(n_639), .Y(n_710) );
INVx1_ASAP7_75t_L g684 ( .A(n_639), .Y(n_684) );
NAND2xp5_ASAP7_75t_SL g714 ( .A(n_639), .B(n_654), .Y(n_714) );
OAI32xp33_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_643), .A3(n_645), .B1(n_646), .B2(n_647), .Y(n_640) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_SL g653 ( .A(n_648), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_648), .B(n_680), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_648), .B(n_709), .Y(n_740) );
NAND2x1p5_ASAP7_75t_L g748 ( .A(n_648), .B(n_659), .Y(n_748) );
NAND5xp2_ASAP7_75t_L g649 ( .A(n_650), .B(n_672), .C(n_685), .D(n_697), .E(n_698), .Y(n_649) );
AOI221xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_654), .B1(n_655), .B2(n_657), .C(n_661), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NAND2xp33_ASAP7_75t_SL g676 ( .A(n_656), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_659), .B(n_728), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_660), .A2(n_673), .B1(n_676), .B2(n_680), .Y(n_672) );
INVx2_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
OAI211xp5_ASAP7_75t_SL g667 ( .A1(n_663), .A2(n_668), .B(n_669), .C(n_670), .Y(n_667) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_SL g695 ( .A(n_675), .Y(n_695) );
INVx1_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_684), .B(n_733), .Y(n_743) );
OR2x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AOI222xp33_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_701), .B1(n_703), .B2(n_707), .C1(n_710), .C2(n_711), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
OAI221xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_715), .B1(n_717), .B2(n_719), .C(n_721), .Y(n_713) );
INVx1_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
OAI21xp33_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .B(n_726), .Y(n_721) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g733 ( .A(n_725), .Y(n_733) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
OAI221xp5_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_732), .B1(n_734), .B2(n_736), .C(n_738), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
INVxp67_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
A2O1A1Ixp33_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_748), .B(n_749), .C(n_751), .Y(n_744) );
INVxp67_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
OAI21xp33_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_753), .B(n_754), .Y(n_751) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_SL g759 ( .A(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_SL g763 ( .A(n_764), .Y(n_763) );
BUFx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
endmodule