module fake_jpeg_17107_n_146 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_146);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_L g30 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_30),
.A2(n_28),
.B1(n_27),
.B2(n_14),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_32),
.B(n_33),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_13),
.B(n_2),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_28),
.Y(n_48)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_21),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_41),
.B(n_48),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_53),
.B1(n_2),
.B2(n_3),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_35),
.A2(n_23),
.B1(n_14),
.B2(n_13),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_51),
.A2(n_39),
.B1(n_24),
.B2(n_22),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_21),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_56),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_32),
.A2(n_23),
.B1(n_27),
.B2(n_20),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_15),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_31),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_59),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_31),
.Y(n_59)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_66),
.Y(n_86)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_65),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_39),
.B1(n_20),
.B2(n_26),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_64),
.A2(n_68),
.B1(n_72),
.B2(n_74),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_50),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_25),
.Y(n_66)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_25),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_73),
.Y(n_93)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_50),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_25),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_44),
.A2(n_17),
.B1(n_3),
.B2(n_25),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_40),
.B(n_37),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_76),
.B(n_77),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_40),
.B(n_37),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_67),
.B(n_9),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_79),
.B(n_88),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_81),
.Y(n_105)
);

NOR3xp33_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_47),
.C(n_40),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_71),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_29),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_89),
.C(n_77),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_3),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_76),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_16),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_47),
.C(n_29),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_16),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_91),
.B(n_69),
.Y(n_103)
);

NAND3xp33_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_106),
.C(n_69),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_102),
.C(n_80),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_92),
.A2(n_74),
.B1(n_58),
.B2(n_62),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_107),
.B1(n_90),
.B2(n_88),
.Y(n_109)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_99),
.A2(n_100),
.B(n_102),
.Y(n_116)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_101),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_60),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_58),
.C(n_47),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_104),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_82),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_82),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_114),
.C(n_115),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_109),
.A2(n_99),
.B1(n_98),
.B2(n_106),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_112),
.B(n_105),
.Y(n_119)
);

OAI22x1_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_90),
.B1(n_84),
.B2(n_87),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_113),
.A2(n_116),
.B1(n_117),
.B2(n_16),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_87),
.C(n_45),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_65),
.C(n_61),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_125),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_99),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_124),
.C(n_16),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_123),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_113),
.A2(n_63),
.B1(n_54),
.B2(n_68),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_17),
.C(n_54),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_112),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_118),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_127),
.A2(n_128),
.B(n_125),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_111),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_122),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_130),
.A2(n_124),
.B(n_120),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_133),
.B(n_135),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_134),
.A2(n_136),
.B(n_137),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_132),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_131),
.A2(n_6),
.B(n_7),
.Y(n_137)
);

XOR2x2_ASAP7_75t_SL g139 ( 
.A(n_133),
.B(n_127),
.Y(n_139)
);

AO21x1_ASAP7_75t_L g143 ( 
.A1(n_139),
.A2(n_141),
.B(n_8),
.Y(n_143)
);

NOR2xp67_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_128),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_140),
.B(n_8),
.Y(n_142)
);

BUFx24_ASAP7_75t_SL g144 ( 
.A(n_142),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_138),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_143),
.Y(n_146)
);


endmodule