module fake_jpeg_21794_n_102 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_102);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_102;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx5p33_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_25),
.B(n_12),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_26),
.A2(n_28),
.B1(n_34),
.B2(n_24),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_13),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_31),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_28)
);

AND2x2_ASAP7_75t_SL g29 ( 
.A(n_13),
.B(n_23),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_13),
.C(n_22),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_1),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_33),
.Y(n_43)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

AOI21xp33_ASAP7_75t_L g32 ( 
.A1(n_14),
.A2(n_3),
.B(n_4),
.Y(n_32)
);

AND2x4_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_18),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_24),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_23),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_36),
.A2(n_14),
.B(n_9),
.Y(n_63)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_41),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_49),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g40 ( 
.A1(n_32),
.A2(n_23),
.B1(n_19),
.B2(n_18),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_28),
.B1(n_31),
.B2(n_29),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_12),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_19),
.B(n_16),
.Y(n_59)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_45),
.Y(n_54)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_15),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_48),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_25),
.B(n_17),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_26),
.B(n_14),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

OAI32xp33_ASAP7_75t_L g76 ( 
.A1(n_51),
.A2(n_61),
.A3(n_64),
.B1(n_40),
.B2(n_45),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_27),
.B(n_31),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_52),
.A2(n_63),
.B(n_49),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_15),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_60),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_40),
.B(n_37),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_43),
.B(n_17),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_50),
.A2(n_16),
.B1(n_18),
.B2(n_14),
.Y(n_61)
);

AO21x2_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_14),
.B(n_7),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_35),
.Y(n_66)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_42),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_68),
.A2(n_58),
.B1(n_54),
.B2(n_52),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_38),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_75),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_39),
.C(n_44),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_74),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_72),
.A2(n_76),
.B1(n_63),
.B2(n_62),
.Y(n_83)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_73),
.A2(n_51),
.B1(n_62),
.B2(n_64),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_82),
.B1(n_83),
.B2(n_61),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_69),
.Y(n_85)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_86),
.A2(n_89),
.B1(n_76),
.B2(n_82),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_71),
.C(n_74),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_88),
.C(n_90),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_55),
.C(n_59),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_84),
.C(n_78),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_85),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_60),
.C(n_65),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_68),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_96),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_55),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_94),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_93),
.C(n_96),
.Y(n_100)
);

AOI322xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_10),
.A3(n_40),
.B1(n_55),
.B2(n_57),
.C1(n_98),
.C2(n_99),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);


endmodule