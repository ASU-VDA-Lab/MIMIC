module fake_jpeg_7602_n_205 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_205);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_205;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_33),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_39),
.Y(n_53)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_35),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_1),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_17),
.Y(n_50)
);

HAxp5_ASAP7_75t_SL g37 ( 
.A(n_23),
.B(n_2),
.CON(n_37),
.SN(n_37)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_20),
.B1(n_28),
.B2(n_25),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_29),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_36),
.A2(n_29),
.B1(n_26),
.B2(n_27),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_43),
.B1(n_49),
.B2(n_58),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_26),
.B1(n_17),
.B2(n_21),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_26),
.B1(n_18),
.B2(n_28),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_44),
.A2(n_47),
.B(n_55),
.Y(n_72)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_52),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_18),
.B1(n_27),
.B2(n_25),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_21),
.B1(n_17),
.B2(n_24),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_34),
.Y(n_59)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_30),
.B(n_21),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_15),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_57),
.Y(n_74)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_24),
.B1(n_20),
.B2(n_22),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_67),
.Y(n_82)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_62),
.Y(n_80)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_66),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_35),
.B1(n_15),
.B2(n_19),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_68),
.B1(n_49),
.B2(n_44),
.Y(n_79)
);

OR2x2_ASAP7_75t_SL g65 ( 
.A(n_58),
.B(n_34),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_65),
.A2(n_47),
.B(n_41),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_32),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_33),
.C(n_30),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_43),
.A2(n_35),
.B1(n_19),
.B2(n_22),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_69),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_32),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_75),
.Y(n_89)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_76),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_42),
.B(n_30),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_77),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_79),
.B(n_61),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_92),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_51),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_85),
.B(n_87),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_48),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_91),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_51),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_65),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_32),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_80),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_45),
.B1(n_52),
.B2(n_40),
.Y(n_94)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_72),
.A2(n_51),
.B1(n_57),
.B2(n_40),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_41),
.B(n_32),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_98),
.B(n_106),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_67),
.C(n_72),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_87),
.C(n_85),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_101),
.A2(n_95),
.B1(n_89),
.B2(n_91),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_92),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_107),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_77),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_59),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_79),
.A2(n_61),
.B(n_76),
.C(n_62),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_108),
.A2(n_114),
.B(n_115),
.Y(n_118)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_111),
.B(n_112),
.Y(n_122)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_77),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_113),
.B(n_96),
.Y(n_131)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_116),
.B(n_123),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_119),
.A2(n_121),
.B1(n_132),
.B2(n_109),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_101),
.A2(n_93),
.B1(n_94),
.B2(n_90),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_82),
.Y(n_124)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_108),
.A2(n_84),
.B1(n_82),
.B2(n_86),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_125),
.A2(n_133),
.B(n_100),
.Y(n_136)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_128),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_82),
.Y(n_127)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_130),
.C(n_100),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_80),
.C(n_96),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_131),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_103),
.A2(n_40),
.B1(n_57),
.B2(n_86),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_115),
.A2(n_32),
.B(n_41),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_118),
.A2(n_108),
.B1(n_103),
.B2(n_114),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_134),
.A2(n_113),
.B(n_128),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_136),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_130),
.C(n_129),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_110),
.Y(n_140)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_106),
.Y(n_142)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_119),
.A2(n_114),
.B(n_104),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_143),
.A2(n_127),
.B(n_124),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_110),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_144),
.B(n_147),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_126),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_125),
.A2(n_109),
.B1(n_112),
.B2(n_111),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_148),
.A2(n_122),
.B1(n_117),
.B2(n_133),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_116),
.B(n_98),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_149),
.B(n_69),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_148),
.A2(n_121),
.B1(n_123),
.B2(n_118),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_154),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_157),
.C(n_161),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_137),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_159),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_158),
.A2(n_160),
.B(n_145),
.Y(n_170)
);

AO22x1_ASAP7_75t_L g160 ( 
.A1(n_134),
.A2(n_51),
.B1(n_38),
.B2(n_31),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_32),
.C(n_38),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_38),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_141),
.C(n_143),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_161),
.B(n_135),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_167),
.Y(n_175)
);

BUFx24_ASAP7_75t_SL g168 ( 
.A(n_153),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_174),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_146),
.C(n_139),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_171),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_170),
.A2(n_173),
.B(n_2),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_139),
.C(n_144),
.Y(n_171)
);

OAI21x1_ASAP7_75t_L g173 ( 
.A1(n_155),
.A2(n_140),
.B(n_145),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_38),
.C(n_19),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_SL g176 ( 
.A1(n_172),
.A2(n_158),
.B(n_156),
.C(n_160),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_176),
.A2(n_180),
.B1(n_3),
.B2(n_4),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_172),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_182),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_166),
.A2(n_162),
.B1(n_163),
.B2(n_13),
.Y(n_178)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_165),
.A2(n_73),
.B1(n_3),
.B2(n_4),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_13),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_181),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_176),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_190),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_11),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_10),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_3),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_189),
.A2(n_6),
.B(n_7),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_186),
.A2(n_176),
.B(n_183),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_193),
.C(n_194),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_186),
.A2(n_179),
.B1(n_5),
.B2(n_6),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_4),
.C(n_5),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_196),
.Y(n_198)
);

FAx1_ASAP7_75t_SL g199 ( 
.A(n_191),
.B(n_185),
.CI(n_7),
.CON(n_199),
.SN(n_199)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_199),
.B(n_200),
.Y(n_202)
);

OAI221xp5_ASAP7_75t_L g200 ( 
.A1(n_191),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_8),
.C(n_9),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_201),
.B(n_10),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_198),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_204),
.Y(n_205)
);


endmodule