module fake_jpeg_12599_n_191 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_191);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_191;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_11),
.B(n_33),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_7),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx4f_ASAP7_75t_SL g59 ( 
.A(n_38),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_46),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_5),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_37),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_1),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_13),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_14),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_9),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

BUFx16f_ASAP7_75t_L g78 ( 
.A(n_3),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_0),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_82),
.B(n_83),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_64),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_0),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_84),
.B(n_50),
.Y(n_96)
);

INVx4_ASAP7_75t_SL g85 ( 
.A(n_64),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_55),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_58),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_56),
.B1(n_73),
.B2(n_68),
.Y(n_101)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_89),
.A2(n_71),
.B1(n_61),
.B2(n_52),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_85),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_90),
.A2(n_56),
.B1(n_70),
.B2(n_77),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_92),
.A2(n_101),
.B1(n_105),
.B2(n_80),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_96),
.B(n_103),
.Y(n_106)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_81),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_67),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_104),
.B(n_66),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_77),
.B1(n_69),
.B2(n_76),
.Y(n_105)
);

OAI32xp33_ASAP7_75t_L g107 ( 
.A1(n_95),
.A2(n_50),
.A3(n_51),
.B1(n_79),
.B2(n_54),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_117),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_108),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_141)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g135 ( 
.A(n_109),
.Y(n_135)
);

OAI21xp33_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_91),
.B(n_94),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_114),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_101),
.A2(n_55),
.B1(n_74),
.B2(n_75),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_111),
.A2(n_18),
.B(n_19),
.Y(n_149)
);

BUFx8_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_72),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_115),
.B(n_2),
.Y(n_133)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

AO22x1_ASAP7_75t_SL g118 ( 
.A1(n_92),
.A2(n_78),
.B1(n_59),
.B2(n_62),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_59),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_119),
.B(n_6),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_51),
.B1(n_63),
.B2(n_60),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_120),
.A2(n_121),
.B1(n_106),
.B2(n_116),
.Y(n_129)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_124),
.Y(n_132)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

INVx3_ASAP7_75t_SL g126 ( 
.A(n_100),
.Y(n_126)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_31),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_136),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_115),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_123),
.B(n_112),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_138),
.B(n_143),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_141),
.B1(n_144),
.B2(n_147),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_32),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_36),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_108),
.A2(n_10),
.B1(n_16),
.B2(n_17),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_20),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_162),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_132),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_153),
.B(n_160),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_157),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_128),
.B(n_29),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_159),
.B(n_164),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_35),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_166),
.Y(n_168)
);

AND2x6_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_39),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_41),
.Y(n_165)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_145),
.A2(n_42),
.B(n_44),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_45),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_167),
.B(n_134),
.Y(n_169)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_151),
.A2(n_130),
.B1(n_149),
.B2(n_139),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_171),
.A2(n_161),
.B1(n_156),
.B2(n_150),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_177),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_173),
.A2(n_166),
.B(n_158),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_178),
.A2(n_179),
.B(n_181),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_170),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_174),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_182),
.B(n_169),
.Y(n_184)
);

NAND4xp25_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_183),
.C(n_180),
.D(n_178),
.Y(n_185)
);

AOI322xp5_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_164),
.A3(n_175),
.B1(n_176),
.B2(n_168),
.C1(n_172),
.C2(n_154),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_168),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_187),
.Y(n_188)
);

BUFx24_ASAP7_75t_SL g189 ( 
.A(n_188),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_163),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_140),
.Y(n_191)
);


endmodule