module fake_jpeg_1855_n_191 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_191);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_191;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_15),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_27),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_13),
.B(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_8),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_30),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_69),
.Y(n_77)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_70),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_56),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_71),
.A2(n_59),
.B1(n_50),
.B2(n_48),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_65),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_69),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_59),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_81),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_79),
.B1(n_71),
.B2(n_69),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_66),
.A2(n_56),
.B1(n_48),
.B2(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_47),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_52),
.C(n_54),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_63),
.Y(n_88)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_86),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_88),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_52),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_94),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_66),
.B1(n_70),
.B2(n_67),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_90),
.A2(n_91),
.B1(n_100),
.B2(n_21),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_80),
.A2(n_66),
.B1(n_70),
.B2(n_61),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_54),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_51),
.B(n_62),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_95),
.A2(n_0),
.B(n_4),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_77),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_65),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_51),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_72),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_75),
.A2(n_65),
.B1(n_64),
.B2(n_49),
.Y(n_100)
);

AO21x1_ASAP7_75t_L g101 ( 
.A1(n_95),
.A2(n_62),
.B(n_55),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_101),
.A2(n_110),
.B(n_7),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_73),
.C(n_83),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_107),
.C(n_102),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_73),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_115),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_106),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_72),
.B(n_70),
.C(n_57),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_60),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_112),
.B(n_116),
.Y(n_121)
);

BUFx8_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_113),
.Y(n_131)
);

AOI32xp33_ASAP7_75t_L g115 ( 
.A1(n_88),
.A2(n_57),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_118),
.Y(n_137)
);

NAND2xp33_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_4),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_119),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_113),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_124),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_97),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

OAI32xp33_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_90),
.A3(n_91),
.B1(n_92),
.B2(n_85),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_23),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_135),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_128),
.A2(n_113),
.B1(n_9),
.B2(n_10),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_104),
.B(n_5),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_129),
.B(n_132),
.Y(n_150)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_119),
.A2(n_22),
.B1(n_42),
.B2(n_39),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_133),
.A2(n_24),
.B(n_35),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_101),
.B(n_6),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_134),
.B(n_117),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_45),
.C(n_37),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_8),
.Y(n_145)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_138),
.B(n_109),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_139),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_143),
.Y(n_158)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_124),
.A2(n_105),
.B1(n_110),
.B2(n_120),
.Y(n_142)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_148),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_128),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_147),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_127),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_151),
.A2(n_154),
.B(n_152),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_153),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_139),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_126),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_130),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_17),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_29),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_131),
.C(n_25),
.Y(n_164)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_160),
.Y(n_172)
);

OAI322xp33_ASAP7_75t_L g161 ( 
.A1(n_156),
.A2(n_122),
.A3(n_137),
.B1(n_133),
.B2(n_136),
.C1(n_131),
.C2(n_32),
.Y(n_161)
);

OAI322xp33_ASAP7_75t_L g170 ( 
.A1(n_161),
.A2(n_164),
.A3(n_168),
.B1(n_146),
.B2(n_157),
.C1(n_151),
.C2(n_18),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_167),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_175)
);

NOR3xp33_ASAP7_75t_SL g169 ( 
.A(n_158),
.B(n_154),
.C(n_144),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_165),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_170),
.A2(n_159),
.B(n_162),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_149),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_173),
.C(n_163),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_149),
.C(n_142),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_167),
.A2(n_150),
.B1(n_19),
.B2(n_20),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_174),
.A2(n_175),
.B1(n_176),
.B2(n_160),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_165),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_178),
.Y(n_183)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_172),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_179),
.A2(n_180),
.B1(n_174),
.B2(n_163),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_181),
.A2(n_171),
.B1(n_173),
.B2(n_164),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_182),
.A2(n_184),
.B1(n_181),
.B2(n_161),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_184),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_183),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_187),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_169),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_189),
.A2(n_20),
.B(n_18),
.Y(n_190)
);

NOR2xp67_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_19),
.Y(n_191)
);


endmodule