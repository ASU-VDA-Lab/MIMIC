module fake_ariane_2431_n_1961 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1961);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1961;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_279;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_967;
wire n_274;
wire n_337;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1860;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_1211;
wire n_996;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

BUFx2_ASAP7_75t_L g207 ( 
.A(n_114),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_71),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_70),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_161),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_41),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_117),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_181),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_183),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_67),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_154),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_2),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_52),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_11),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_155),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_136),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_113),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_33),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_24),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_6),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_50),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_25),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_61),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_30),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_200),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_56),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_0),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_74),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_73),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_140),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_59),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_39),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_76),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_44),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_112),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_118),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_66),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_93),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_100),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_197),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_116),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_25),
.Y(n_248)
);

INVxp33_ASAP7_75t_L g249 ( 
.A(n_106),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_92),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_195),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_31),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_88),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_4),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_50),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_110),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_158),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_127),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_153),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_35),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_83),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_105),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_16),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_194),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_86),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_91),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_119),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_63),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_125),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_188),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_142),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_196),
.Y(n_272)
);

BUFx5_ASAP7_75t_L g273 ( 
.A(n_148),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_206),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_169),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_190),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_203),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_202),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_144),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_168),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_132),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_33),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_73),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_71),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_184),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_174),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_35),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_74),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_21),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_177),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_53),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_179),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_59),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_95),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_7),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_162),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_69),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_126),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_27),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_47),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_107),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_98),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_157),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_52),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_147),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_69),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_63),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_78),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_156),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_2),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_152),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_31),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_115),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_3),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_57),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_186),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_23),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_159),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_101),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_137),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_55),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_70),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_24),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_84),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_173),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_187),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_139),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_131),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_90),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_151),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_96),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_180),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_145),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_10),
.Y(n_334)
);

INVxp33_ASAP7_75t_L g335 ( 
.A(n_182),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_72),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_143),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_128),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_146),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_133),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_176),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_89),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_49),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_138),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_164),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_9),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_167),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_41),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_166),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_32),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_10),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_62),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_109),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_51),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_26),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_12),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_193),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_189),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_16),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_121),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_171),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_11),
.Y(n_362)
);

BUFx10_ASAP7_75t_L g363 ( 
.A(n_8),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_14),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_97),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_18),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_163),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_102),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_22),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_64),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_201),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_130),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_87),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_170),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_29),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_72),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_0),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_149),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_18),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_58),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_124),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_61),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_46),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_123),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_129),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_12),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_37),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_82),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_204),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_85),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_64),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_67),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_15),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_54),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_75),
.Y(n_395)
);

INVx2_ASAP7_75t_SL g396 ( 
.A(n_39),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_134),
.Y(n_397)
);

INVx2_ASAP7_75t_SL g398 ( 
.A(n_13),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_27),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_6),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_111),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_150),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_32),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_3),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_7),
.Y(n_405)
);

CKINVDCx14_ASAP7_75t_R g406 ( 
.A(n_34),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_224),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_210),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_284),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_406),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_241),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_207),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g413 ( 
.A(n_383),
.B(n_1),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_284),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_267),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_245),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_210),
.Y(n_417)
);

NOR2xp67_ASAP7_75t_L g418 ( 
.A(n_396),
.B(n_1),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_383),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_224),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_267),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_284),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_251),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_258),
.Y(n_424)
);

NOR2xp67_ASAP7_75t_L g425 ( 
.A(n_396),
.B(n_4),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_207),
.B(n_5),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_212),
.B(n_5),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g428 ( 
.A(n_310),
.B(n_8),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_213),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_213),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_220),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_272),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_331),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_220),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_211),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_221),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_280),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_224),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_212),
.B(n_9),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_331),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_295),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_295),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_397),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_397),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_361),
.Y(n_445)
);

CKINVDCx14_ASAP7_75t_R g446 ( 
.A(n_231),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_295),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_361),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_285),
.Y(n_449)
);

INVxp67_ASAP7_75t_SL g450 ( 
.A(n_304),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_286),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_303),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_342),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_357),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_360),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_304),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_209),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_304),
.Y(n_458)
);

INVxp33_ASAP7_75t_SL g459 ( 
.A(n_217),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_218),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_365),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_221),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_346),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_225),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_208),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_346),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_366),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_211),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_394),
.Y(n_469)
);

INVxp67_ASAP7_75t_SL g470 ( 
.A(n_346),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_227),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_215),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_230),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_398),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_257),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_222),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_232),
.Y(n_477)
);

INVxp67_ASAP7_75t_SL g478 ( 
.A(n_224),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_363),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_257),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_215),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_363),
.B(n_13),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_405),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_405),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_257),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_265),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_233),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_265),
.Y(n_488)
);

OR2x2_ASAP7_75t_L g489 ( 
.A(n_219),
.B(n_14),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_219),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_234),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_226),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_226),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_229),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_229),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_238),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_235),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_222),
.B(n_15),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_237),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_265),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_243),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_246),
.Y(n_502)
);

NOR2xp67_ASAP7_75t_L g503 ( 
.A(n_398),
.B(n_17),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_246),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_238),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_250),
.B(n_19),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_252),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_363),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_255),
.Y(n_509)
);

CKINVDCx14_ASAP7_75t_R g510 ( 
.A(n_363),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_260),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_407),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_407),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_445),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_420),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_420),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_438),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_438),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_463),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_408),
.B(n_224),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_457),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_466),
.Y(n_522)
);

INVx5_ASAP7_75t_L g523 ( 
.A(n_482),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_408),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_417),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_417),
.B(n_224),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_429),
.Y(n_527)
);

NAND2x1_ASAP7_75t_L g528 ( 
.A(n_482),
.B(n_256),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_478),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_429),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_430),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_430),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_431),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_431),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_434),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_434),
.Y(n_536)
);

OA21x2_ASAP7_75t_L g537 ( 
.A1(n_436),
.A2(n_259),
.B(n_250),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_436),
.B(n_240),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_462),
.Y(n_539)
);

OAI21x1_ASAP7_75t_L g540 ( 
.A1(n_506),
.A2(n_374),
.B(n_256),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_462),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_476),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_427),
.B(n_249),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_476),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_443),
.B(n_335),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_502),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_450),
.B(n_259),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_502),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_465),
.A2(n_254),
.B1(n_282),
.B2(n_228),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_504),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_504),
.B(n_240),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_470),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_472),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_481),
.Y(n_554)
);

NOR2x1_ASAP7_75t_L g555 ( 
.A(n_412),
.B(n_239),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_483),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_409),
.B(n_278),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_484),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_490),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_492),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_414),
.B(n_278),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_494),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_495),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_496),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_505),
.Y(n_565)
);

CKINVDCx16_ASAP7_75t_R g566 ( 
.A(n_479),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_422),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_511),
.Y(n_568)
);

OA21x2_ASAP7_75t_L g569 ( 
.A1(n_498),
.A2(n_313),
.B(n_308),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_441),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_442),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_447),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_456),
.B(n_308),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_458),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_435),
.B(n_313),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_489),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_489),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_474),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_418),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_468),
.B(n_318),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_493),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_425),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_415),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_474),
.B(n_318),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_503),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_412),
.B(n_325),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_413),
.Y(n_587)
);

INVx5_ASAP7_75t_L g588 ( 
.A(n_446),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_428),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_445),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_428),
.Y(n_591)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_448),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_413),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_426),
.Y(n_594)
);

BUFx10_ASAP7_75t_L g595 ( 
.A(n_547),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_529),
.B(n_552),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_529),
.B(n_552),
.Y(n_597)
);

INVx4_ASAP7_75t_L g598 ( 
.A(n_588),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_531),
.Y(n_599)
);

OR2x2_ASAP7_75t_L g600 ( 
.A(n_578),
.B(n_469),
.Y(n_600)
);

HB1xp67_ASAP7_75t_L g601 ( 
.A(n_514),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_531),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_512),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_588),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_552),
.B(n_459),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_524),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_512),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_594),
.B(n_421),
.Y(n_608)
);

NAND3xp33_ASAP7_75t_L g609 ( 
.A(n_594),
.B(n_448),
.C(n_439),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_531),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_588),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_531),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_531),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_531),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_531),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_513),
.Y(n_616)
);

BUFx10_ASAP7_75t_L g617 ( 
.A(n_547),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_531),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_591),
.B(n_510),
.Y(n_619)
);

INVx1_ASAP7_75t_SL g620 ( 
.A(n_568),
.Y(n_620)
);

AO22x2_ASAP7_75t_L g621 ( 
.A1(n_528),
.A2(n_419),
.B1(n_352),
.B2(n_399),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_L g622 ( 
.A1(n_594),
.A2(n_421),
.B1(n_440),
.B2(n_433),
.Y(n_622)
);

AND2x2_ASAP7_75t_SL g623 ( 
.A(n_545),
.B(n_256),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_591),
.B(n_440),
.Y(n_624)
);

AND2x6_ASAP7_75t_L g625 ( 
.A(n_576),
.B(n_374),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_578),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_532),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_523),
.B(n_444),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g629 ( 
.A(n_578),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_513),
.Y(n_630)
);

NOR2x1p5_ASAP7_75t_L g631 ( 
.A(n_578),
.B(n_444),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_588),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_522),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_532),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_588),
.Y(n_635)
);

AOI21x1_ASAP7_75t_L g636 ( 
.A1(n_528),
.A2(n_326),
.B(n_325),
.Y(n_636)
);

XOR2xp5_ASAP7_75t_R g637 ( 
.A(n_566),
.B(n_467),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_513),
.Y(n_638)
);

INVx8_ASAP7_75t_L g639 ( 
.A(n_588),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_523),
.Y(n_640)
);

OR2x2_ASAP7_75t_L g641 ( 
.A(n_566),
.B(n_452),
.Y(n_641)
);

AND2x2_ASAP7_75t_SL g642 ( 
.A(n_545),
.B(n_374),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_523),
.B(n_475),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_513),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_515),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_515),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_592),
.B(n_464),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_591),
.B(n_464),
.Y(n_648)
);

CKINVDCx6p67_ASAP7_75t_R g649 ( 
.A(n_583),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_532),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_532),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_532),
.Y(n_652)
);

INVxp33_ASAP7_75t_L g653 ( 
.A(n_514),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_515),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_515),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_592),
.B(n_471),
.Y(n_656)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_590),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_532),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_568),
.Y(n_659)
);

NAND2xp33_ASAP7_75t_R g660 ( 
.A(n_583),
.B(n_452),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_569),
.A2(n_485),
.B1(n_486),
.B2(n_480),
.Y(n_661)
);

INVxp67_ASAP7_75t_SL g662 ( 
.A(n_534),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_523),
.B(n_488),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_569),
.A2(n_500),
.B1(n_248),
.B2(n_299),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_523),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_532),
.Y(n_666)
);

INVx5_ASAP7_75t_L g667 ( 
.A(n_532),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_536),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_523),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_588),
.Y(n_670)
);

INVx8_ASAP7_75t_L g671 ( 
.A(n_588),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_516),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_592),
.B(n_471),
.Y(n_673)
);

INVxp33_ASAP7_75t_SL g674 ( 
.A(n_590),
.Y(n_674)
);

OAI22xp5_ASAP7_75t_L g675 ( 
.A1(n_591),
.A2(n_355),
.B1(n_477),
.B2(n_473),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_536),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_524),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_516),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_523),
.B(n_473),
.Y(n_679)
);

BUFx2_ASAP7_75t_L g680 ( 
.A(n_583),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_527),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_569),
.A2(n_248),
.B1(n_299),
.B2(n_293),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_581),
.B(n_293),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_523),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_576),
.B(n_477),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_576),
.B(n_487),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_523),
.B(n_576),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_516),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_591),
.B(n_487),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_522),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_576),
.B(n_491),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_576),
.B(n_491),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_527),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_587),
.B(n_454),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_543),
.B(n_499),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_543),
.B(n_499),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_536),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_576),
.B(n_501),
.Y(n_698)
);

OR2x6_ASAP7_75t_L g699 ( 
.A(n_528),
.B(n_576),
.Y(n_699)
);

BUFx4f_ASAP7_75t_L g700 ( 
.A(n_569),
.Y(n_700)
);

OAI22xp33_ASAP7_75t_L g701 ( 
.A1(n_584),
.A2(n_507),
.B1(n_501),
.B2(n_497),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_569),
.A2(n_300),
.B1(n_321),
.B2(n_315),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_581),
.B(n_300),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_516),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_517),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_588),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_568),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_581),
.B(n_315),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_517),
.Y(n_709)
);

INVx5_ASAP7_75t_L g710 ( 
.A(n_536),
.Y(n_710)
);

AND2x6_ASAP7_75t_L g711 ( 
.A(n_520),
.B(n_326),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_536),
.Y(n_712)
);

INVx1_ASAP7_75t_SL g713 ( 
.A(n_581),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_521),
.A2(n_507),
.B1(n_509),
.B2(n_460),
.Y(n_714)
);

INVxp33_ASAP7_75t_L g715 ( 
.A(n_549),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_517),
.Y(n_716)
);

INVxp67_ASAP7_75t_SL g717 ( 
.A(n_534),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_521),
.A2(n_351),
.B1(n_268),
.B2(n_404),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_549),
.Y(n_719)
);

AND2x6_ASAP7_75t_L g720 ( 
.A(n_520),
.B(n_344),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_555),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_589),
.B(n_410),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_589),
.A2(n_297),
.B1(n_403),
.B2(n_400),
.Y(n_723)
);

OR2x6_ASAP7_75t_L g724 ( 
.A(n_577),
.B(n_321),
.Y(n_724)
);

OAI22xp33_ASAP7_75t_L g725 ( 
.A1(n_584),
.A2(n_575),
.B1(n_580),
.B2(n_589),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_536),
.Y(n_726)
);

AND3x2_ASAP7_75t_L g727 ( 
.A(n_579),
.B(n_585),
.C(n_582),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_517),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_536),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_536),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_527),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_589),
.B(n_508),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_577),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_535),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_569),
.A2(n_343),
.B1(n_375),
.B2(n_386),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_522),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_522),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_555),
.B(n_577),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_535),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_535),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_522),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_522),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_713),
.B(n_725),
.Y(n_743)
);

INVxp67_ASAP7_75t_L g744 ( 
.A(n_600),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_626),
.B(n_577),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_626),
.B(n_579),
.Y(n_746)
);

O2A1O1Ixp33_ASAP7_75t_L g747 ( 
.A1(n_698),
.A2(n_575),
.B(n_580),
.C(n_534),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_682),
.A2(n_537),
.B1(n_525),
.B2(n_530),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_733),
.A2(n_579),
.B1(n_585),
.B2(n_582),
.Y(n_749)
);

NOR2xp67_ASAP7_75t_L g750 ( 
.A(n_657),
.B(n_454),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_600),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_595),
.B(n_617),
.Y(n_752)
);

INVx8_ASAP7_75t_L g753 ( 
.A(n_699),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_733),
.B(n_533),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_731),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_605),
.B(n_533),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_595),
.B(n_587),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_608),
.B(n_533),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_734),
.Y(n_759)
);

INVxp67_ASAP7_75t_SL g760 ( 
.A(n_629),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_647),
.B(n_533),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_633),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_606),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_677),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_656),
.B(n_533),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_673),
.B(n_587),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_680),
.B(n_593),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_700),
.B(n_534),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_695),
.A2(n_582),
.B1(n_585),
.B2(n_593),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_648),
.B(n_593),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_680),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_629),
.B(n_586),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_595),
.B(n_586),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_687),
.A2(n_717),
.B(n_662),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_732),
.B(n_461),
.Y(n_775)
);

NAND3xp33_ASAP7_75t_L g776 ( 
.A(n_722),
.B(n_567),
.C(n_570),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_603),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_601),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_648),
.B(n_534),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_607),
.Y(n_780)
);

NAND3xp33_ASAP7_75t_L g781 ( 
.A(n_696),
.B(n_567),
.C(n_570),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_637),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_689),
.B(n_542),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_624),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_616),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_689),
.B(n_542),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_633),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_681),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_693),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_619),
.B(n_542),
.Y(n_790)
);

INVxp67_ASAP7_75t_L g791 ( 
.A(n_660),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_617),
.B(n_574),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_700),
.B(n_617),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_739),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_619),
.B(n_544),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_624),
.B(n_544),
.Y(n_796)
);

OR2x6_ASAP7_75t_L g797 ( 
.A(n_641),
.B(n_556),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_721),
.B(n_574),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_721),
.B(n_574),
.Y(n_799)
);

OR2x6_ASAP7_75t_L g800 ( 
.A(n_641),
.B(n_556),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_738),
.B(n_544),
.Y(n_801)
);

OAI21xp33_ASAP7_75t_L g802 ( 
.A1(n_723),
.A2(n_550),
.B(n_559),
.Y(n_802)
);

NAND2xp33_ASAP7_75t_L g803 ( 
.A(n_679),
.B(n_550),
.Y(n_803)
);

INVxp33_ASAP7_75t_SL g804 ( 
.A(n_707),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_701),
.B(n_550),
.Y(n_805)
);

NAND3xp33_ASAP7_75t_L g806 ( 
.A(n_622),
.B(n_570),
.C(n_461),
.Y(n_806)
);

AO221x1_ASAP7_75t_L g807 ( 
.A1(n_621),
.A2(n_240),
.B1(n_336),
.B2(n_343),
.C(n_350),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_623),
.B(n_553),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_623),
.B(n_553),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_699),
.A2(n_563),
.B1(n_559),
.B2(n_554),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_740),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_596),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_642),
.B(n_553),
.Y(n_813)
);

INVx4_ASAP7_75t_L g814 ( 
.A(n_699),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_642),
.B(n_572),
.Y(n_815)
);

A2O1A1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_700),
.A2(n_540),
.B(n_554),
.C(n_553),
.Y(n_816)
);

INVx4_ASAP7_75t_L g817 ( 
.A(n_699),
.Y(n_817)
);

INVxp67_ASAP7_75t_L g818 ( 
.A(n_620),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_609),
.B(n_572),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_597),
.Y(n_820)
);

NOR3xp33_ASAP7_75t_L g821 ( 
.A(n_675),
.B(n_554),
.C(n_553),
.Y(n_821)
);

NOR2xp67_ASAP7_75t_SL g822 ( 
.A(n_685),
.B(n_336),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_683),
.B(n_554),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_686),
.B(n_691),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_630),
.Y(n_825)
);

OR2x6_ASAP7_75t_L g826 ( 
.A(n_631),
.B(n_563),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_683),
.B(n_554),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_630),
.Y(n_828)
);

NAND2xp33_ASAP7_75t_L g829 ( 
.A(n_639),
.B(n_525),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_683),
.B(n_572),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_692),
.A2(n_574),
.B1(n_572),
.B2(n_560),
.Y(n_831)
);

HB1xp67_ASAP7_75t_L g832 ( 
.A(n_724),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_639),
.A2(n_540),
.B(n_530),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_703),
.B(n_572),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_638),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_703),
.B(n_574),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_674),
.B(n_558),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_674),
.B(n_558),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_703),
.B(n_525),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_714),
.B(n_558),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_708),
.B(n_525),
.Y(n_841)
);

INVx1_ASAP7_75t_SL g842 ( 
.A(n_659),
.Y(n_842)
);

O2A1O1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_724),
.A2(n_539),
.B(n_541),
.C(n_530),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_640),
.B(n_558),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_L g845 ( 
.A1(n_724),
.A2(n_560),
.B1(n_565),
.B2(n_562),
.Y(n_845)
);

NAND2x1p5_ASAP7_75t_L g846 ( 
.A(n_640),
.B(n_537),
.Y(n_846)
);

NOR2xp67_ASAP7_75t_L g847 ( 
.A(n_694),
.B(n_560),
.Y(n_847)
);

INVx2_ASAP7_75t_SL g848 ( 
.A(n_727),
.Y(n_848)
);

BUFx10_ASAP7_75t_L g849 ( 
.A(n_707),
.Y(n_849)
);

INVxp67_ASAP7_75t_L g850 ( 
.A(n_694),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_665),
.B(n_558),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_665),
.B(n_558),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_643),
.B(n_571),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_638),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_644),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_663),
.B(n_571),
.Y(n_856)
);

HB1xp67_ASAP7_75t_L g857 ( 
.A(n_724),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_628),
.B(n_571),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_708),
.B(n_530),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_708),
.B(n_539),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_644),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_664),
.B(n_539),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_653),
.B(n_558),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_645),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_718),
.B(n_558),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_711),
.B(n_539),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_711),
.B(n_541),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_669),
.B(n_571),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_669),
.B(n_564),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_711),
.B(n_541),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_684),
.B(n_564),
.Y(n_871)
);

NAND2xp33_ASAP7_75t_L g872 ( 
.A(n_639),
.B(n_541),
.Y(n_872)
);

OR2x6_ASAP7_75t_L g873 ( 
.A(n_621),
.B(n_557),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_684),
.B(n_564),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_599),
.B(n_627),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_702),
.B(n_564),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_633),
.B(n_564),
.Y(n_877)
);

NOR2xp67_ASAP7_75t_L g878 ( 
.A(n_645),
.B(n_560),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_711),
.B(n_546),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_711),
.B(n_546),
.Y(n_880)
);

BUFx6f_ASAP7_75t_L g881 ( 
.A(n_633),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_711),
.B(n_546),
.Y(n_882)
);

AOI22xp5_ASAP7_75t_L g883 ( 
.A1(n_720),
.A2(n_565),
.B1(n_562),
.B2(n_564),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_720),
.B(n_416),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_742),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_599),
.B(n_564),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_599),
.B(n_564),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_735),
.A2(n_537),
.B1(n_548),
.B2(n_546),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_633),
.B(n_548),
.Y(n_889)
);

NAND3xp33_ASAP7_75t_L g890 ( 
.A(n_661),
.B(n_561),
.C(n_557),
.Y(n_890)
);

AND2x6_ASAP7_75t_SL g891 ( 
.A(n_637),
.B(n_350),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_690),
.B(n_548),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_L g893 ( 
.A1(n_621),
.A2(n_537),
.B1(n_548),
.B2(n_562),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_720),
.B(n_562),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_646),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_720),
.B(n_565),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_SL g897 ( 
.A(n_649),
.B(n_423),
.Y(n_897)
);

AO22x2_ASAP7_75t_L g898 ( 
.A1(n_715),
.A2(n_395),
.B1(n_362),
.B2(n_364),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_654),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_627),
.B(n_666),
.Y(n_900)
);

AO21x1_ASAP7_75t_L g901 ( 
.A1(n_793),
.A2(n_540),
.B(n_636),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_803),
.A2(n_671),
.B(n_639),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_766),
.B(n_720),
.Y(n_903)
);

INVxp67_ASAP7_75t_L g904 ( 
.A(n_751),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_751),
.B(n_744),
.Y(n_905)
);

INVx8_ASAP7_75t_L g906 ( 
.A(n_753),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_768),
.A2(n_671),
.B(n_632),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_812),
.B(n_720),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_768),
.A2(n_671),
.B(n_632),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_755),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_850),
.B(n_424),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_767),
.B(n_432),
.Y(n_912)
);

O2A1O1Ixp5_ASAP7_75t_L g913 ( 
.A1(n_819),
.A2(n_636),
.B(n_730),
.C(n_729),
.Y(n_913)
);

AOI21x1_ASAP7_75t_L g914 ( 
.A1(n_793),
.A2(n_610),
.B(n_602),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_757),
.A2(n_449),
.B1(n_451),
.B2(n_437),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_820),
.B(n_625),
.Y(n_916)
);

OR2x6_ASAP7_75t_L g917 ( 
.A(n_753),
.B(n_565),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_760),
.A2(n_671),
.B(n_632),
.Y(n_918)
);

INVx2_ASAP7_75t_SL g919 ( 
.A(n_849),
.Y(n_919)
);

INVx1_ASAP7_75t_SL g920 ( 
.A(n_842),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_743),
.A2(n_666),
.B1(n_668),
.B2(n_627),
.Y(n_921)
);

O2A1O1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_757),
.A2(n_364),
.B(n_375),
.C(n_362),
.Y(n_922)
);

INVx4_ASAP7_75t_L g923 ( 
.A(n_753),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_791),
.B(n_719),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_752),
.B(n_719),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_832),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_770),
.B(n_625),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_875),
.A2(n_598),
.B(n_604),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_784),
.B(n_625),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_875),
.A2(n_598),
.B(n_604),
.Y(n_930)
);

O2A1O1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_779),
.A2(n_756),
.B(n_745),
.C(n_773),
.Y(n_931)
);

NOR2x2_ASAP7_75t_L g932 ( 
.A(n_797),
.B(n_659),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_900),
.A2(n_598),
.B(n_611),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_900),
.A2(n_635),
.B(n_611),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_847),
.B(n_752),
.Y(n_935)
);

OAI21xp5_ASAP7_75t_L g936 ( 
.A1(n_816),
.A2(n_610),
.B(n_602),
.Y(n_936)
);

A2O1A1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_815),
.A2(n_819),
.B(n_824),
.C(n_792),
.Y(n_937)
);

INVx1_ASAP7_75t_SL g938 ( 
.A(n_771),
.Y(n_938)
);

BUFx4f_ASAP7_75t_L g939 ( 
.A(n_797),
.Y(n_939)
);

NOR2xp67_ASAP7_75t_L g940 ( 
.A(n_818),
.B(n_778),
.Y(n_940)
);

INVx4_ASAP7_75t_L g941 ( 
.A(n_814),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_SL g942 ( 
.A1(n_804),
.A2(n_455),
.B1(n_453),
.B2(n_263),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_814),
.B(n_690),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_774),
.A2(n_833),
.B(n_858),
.Y(n_944)
);

BUFx12f_ASAP7_75t_L g945 ( 
.A(n_849),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_783),
.B(n_625),
.Y(n_946)
);

O2A1O1Ixp5_ASAP7_75t_L g947 ( 
.A1(n_865),
.A2(n_730),
.B(n_729),
.C(n_612),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_817),
.Y(n_948)
);

O2A1O1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_790),
.A2(n_386),
.B(n_393),
.C(n_379),
.Y(n_949)
);

A2O1A1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_815),
.A2(n_668),
.B(n_666),
.C(n_613),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_759),
.Y(n_951)
);

BUFx4f_ASAP7_75t_L g952 ( 
.A(n_797),
.Y(n_952)
);

INVxp67_ASAP7_75t_L g953 ( 
.A(n_832),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_786),
.B(n_625),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_858),
.A2(n_670),
.B(n_635),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_763),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_795),
.B(n_625),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_817),
.B(n_690),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_775),
.B(n_668),
.Y(n_959)
);

O2A1O1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_796),
.A2(n_393),
.B(n_395),
.C(n_379),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_764),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_824),
.A2(n_792),
.B(n_799),
.C(n_798),
.Y(n_962)
);

INVxp67_ASAP7_75t_SL g963 ( 
.A(n_857),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_769),
.B(n_561),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_749),
.B(n_573),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_747),
.A2(n_613),
.B(n_612),
.Y(n_966)
);

CKINVDCx10_ASAP7_75t_R g967 ( 
.A(n_800),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_857),
.B(n_614),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_761),
.A2(n_706),
.B(n_670),
.Y(n_969)
);

AO21x1_ASAP7_75t_L g970 ( 
.A1(n_853),
.A2(n_615),
.B(n_614),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_762),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_758),
.B(n_573),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_765),
.A2(n_706),
.B(n_618),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_808),
.B(n_690),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_754),
.B(n_520),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_886),
.A2(n_618),
.B(n_615),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_788),
.B(n_520),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_886),
.A2(n_650),
.B(n_634),
.Y(n_978)
);

OR2x2_ASAP7_75t_L g979 ( 
.A(n_800),
.B(n_520),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_789),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_777),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_887),
.A2(n_650),
.B(n_634),
.Y(n_982)
);

O2A1O1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_805),
.A2(n_772),
.B(n_838),
.C(n_837),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_887),
.A2(n_872),
.B(n_829),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_892),
.A2(n_652),
.B(n_651),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_794),
.B(n_811),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_762),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_890),
.B(n_520),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_798),
.B(n_526),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_892),
.A2(n_652),
.B(n_651),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_801),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_839),
.Y(n_992)
);

OAI21xp33_ASAP7_75t_SL g993 ( 
.A1(n_810),
.A2(n_746),
.B(n_799),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_821),
.A2(n_726),
.B(n_676),
.C(n_712),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_844),
.A2(n_676),
.B(n_658),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_844),
.A2(n_697),
.B(n_658),
.Y(n_996)
);

O2A1O1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_802),
.A2(n_726),
.B(n_712),
.C(n_697),
.Y(n_997)
);

INVx4_ASAP7_75t_L g998 ( 
.A(n_762),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_809),
.A2(n_742),
.B(n_741),
.C(n_737),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_823),
.B(n_526),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_851),
.A2(n_737),
.B(n_736),
.Y(n_1001)
);

HB1xp67_ASAP7_75t_L g1002 ( 
.A(n_827),
.Y(n_1002)
);

NOR2x1p5_ASAP7_75t_SL g1003 ( 
.A(n_825),
.B(n_736),
.Y(n_1003)
);

BUFx2_ASAP7_75t_SL g1004 ( 
.A(n_750),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_813),
.A2(n_741),
.B1(n_690),
.B2(n_537),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_884),
.Y(n_1006)
);

INVx4_ASAP7_75t_L g1007 ( 
.A(n_762),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_781),
.A2(n_537),
.B1(n_283),
.B2(n_387),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_841),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_853),
.A2(n_672),
.B(n_655),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_851),
.A2(n_710),
.B(n_667),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_787),
.Y(n_1012)
);

OAI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_856),
.A2(n_672),
.B(n_655),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_787),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_863),
.B(n_678),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_787),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_776),
.B(n_526),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_884),
.B(n_526),
.Y(n_1018)
);

NAND3xp33_ASAP7_75t_L g1019 ( 
.A(n_806),
.B(n_288),
.C(n_287),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_787),
.Y(n_1020)
);

INVx4_ASAP7_75t_L g1021 ( 
.A(n_881),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_881),
.B(n_667),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_852),
.A2(n_710),
.B(n_667),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_830),
.B(n_526),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_840),
.B(n_678),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_852),
.A2(n_710),
.B(n_667),
.Y(n_1026)
);

O2A1O1Ixp5_ASAP7_75t_L g1027 ( 
.A1(n_889),
.A2(n_519),
.B(n_526),
.C(n_538),
.Y(n_1027)
);

OAI21xp33_ASAP7_75t_L g1028 ( 
.A1(n_834),
.A2(n_291),
.B(n_289),
.Y(n_1028)
);

O2A1O1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_843),
.A2(n_836),
.B(n_874),
.C(n_877),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_859),
.B(n_538),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_860),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_845),
.Y(n_1032)
);

AOI22xp33_ASAP7_75t_SL g1033 ( 
.A1(n_898),
.A2(n_317),
.B1(n_356),
.B2(n_359),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_846),
.A2(n_728),
.B(n_704),
.Y(n_1034)
);

AOI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_826),
.A2(n_274),
.B1(n_344),
.B2(n_345),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_826),
.B(n_688),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_780),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_785),
.Y(n_1038)
);

O2A1O1Ixp5_ASAP7_75t_L g1039 ( 
.A1(n_877),
.A2(n_519),
.B(n_551),
.C(n_538),
.Y(n_1039)
);

OAI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_846),
.A2(n_705),
.B(n_688),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_881),
.B(n_667),
.Y(n_1041)
);

AOI21xp33_ASAP7_75t_L g1042 ( 
.A1(n_894),
.A2(n_709),
.B(n_705),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_874),
.A2(n_710),
.B(n_709),
.Y(n_1043)
);

NAND3xp33_ASAP7_75t_L g1044 ( 
.A(n_822),
.B(n_307),
.C(n_306),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_881),
.B(n_710),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_826),
.B(n_716),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_869),
.A2(n_716),
.B(n_551),
.Y(n_1047)
);

INVx11_ASAP7_75t_L g1048 ( 
.A(n_897),
.Y(n_1048)
);

BUFx3_ASAP7_75t_L g1049 ( 
.A(n_782),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_868),
.B(n_538),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_869),
.A2(n_551),
.B(n_538),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_868),
.B(n_538),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_893),
.B(n_551),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_871),
.A2(n_551),
.B(n_216),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_835),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_893),
.B(n_551),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_828),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_871),
.A2(n_223),
.B(n_214),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_885),
.A2(n_242),
.B(n_236),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_854),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_866),
.B(n_522),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_885),
.A2(n_247),
.B(n_244),
.Y(n_1062)
);

BUFx2_ASAP7_75t_L g1063 ( 
.A(n_891),
.Y(n_1063)
);

O2A1O1Ixp33_ASAP7_75t_SL g1064 ( 
.A1(n_867),
.A2(n_345),
.B(n_384),
.C(n_373),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_873),
.B(n_312),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_870),
.B(n_349),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_848),
.B(n_314),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_899),
.A2(n_261),
.B(n_253),
.Y(n_1068)
);

BUFx2_ASAP7_75t_L g1069 ( 
.A(n_873),
.Y(n_1069)
);

AOI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_896),
.A2(n_274),
.B1(n_367),
.B2(n_349),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_855),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_861),
.A2(n_264),
.B(n_262),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_864),
.A2(n_269),
.B(n_266),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_879),
.A2(n_373),
.B(n_367),
.C(n_384),
.Y(n_1074)
);

O2A1O1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_880),
.A2(n_316),
.B(n_301),
.C(n_281),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_984),
.A2(n_882),
.B(n_876),
.Y(n_1076)
);

O2A1O1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_937),
.A2(n_895),
.B(n_862),
.C(n_316),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_923),
.B(n_883),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_962),
.A2(n_831),
.B1(n_748),
.B2(n_888),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_944),
.A2(n_888),
.B(n_748),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_911),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_906),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_923),
.B(n_878),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_945),
.Y(n_1084)
);

INVx4_ASAP7_75t_L g1085 ( 
.A(n_906),
.Y(n_1085)
);

AO21x1_ASAP7_75t_L g1086 ( 
.A1(n_974),
.A2(n_518),
.B(n_807),
.Y(n_1086)
);

AOI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_1033),
.A2(n_334),
.B1(n_370),
.B2(n_369),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_956),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_925),
.B(n_322),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_961),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_972),
.A2(n_319),
.B(n_332),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_906),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_903),
.A2(n_330),
.B(n_402),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_939),
.B(n_323),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_913),
.A2(n_518),
.B(n_348),
.Y(n_1095)
);

O2A1O1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_922),
.A2(n_904),
.B(n_959),
.C(n_925),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_980),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_915),
.B(n_354),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_910),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_R g1100 ( 
.A(n_967),
.B(n_376),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_963),
.B(n_377),
.Y(n_1101)
);

OAI21xp33_ASAP7_75t_SL g1102 ( 
.A1(n_964),
.A2(n_518),
.B(n_20),
.Y(n_1102)
);

BUFx12f_ASAP7_75t_L g1103 ( 
.A(n_919),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_952),
.B(n_380),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_963),
.B(n_382),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_936),
.A2(n_401),
.B(n_270),
.Y(n_1106)
);

INVx3_ASAP7_75t_L g1107 ( 
.A(n_941),
.Y(n_1107)
);

AND2x4_ASAP7_75t_L g1108 ( 
.A(n_917),
.B(n_19),
.Y(n_1108)
);

O2A1O1Ixp5_ASAP7_75t_L g1109 ( 
.A1(n_970),
.A2(n_240),
.B(n_21),
.C(n_22),
.Y(n_1109)
);

INVx2_ASAP7_75t_SL g1110 ( 
.A(n_1048),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_971),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_905),
.B(n_904),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_938),
.B(n_391),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_924),
.B(n_392),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_951),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_902),
.A2(n_390),
.B(n_389),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_993),
.A2(n_240),
.B(n_385),
.C(n_381),
.Y(n_1117)
);

INVx5_ASAP7_75t_L g1118 ( 
.A(n_917),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_924),
.B(n_20),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_965),
.A2(n_240),
.B1(n_378),
.B2(n_372),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_920),
.B(n_271),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_986),
.A2(n_388),
.B1(n_371),
.B2(n_368),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1002),
.B(n_23),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_1033),
.A2(n_358),
.B1(n_353),
.B2(n_347),
.Y(n_1124)
);

AOI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_942),
.A2(n_305),
.B1(n_340),
.B2(n_339),
.Y(n_1125)
);

A2O1A1Ixp33_ASAP7_75t_SL g1126 ( 
.A1(n_959),
.A2(n_966),
.B(n_931),
.C(n_994),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1057),
.Y(n_1127)
);

INVx2_ASAP7_75t_SL g1128 ( 
.A(n_1049),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_917),
.B(n_26),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_1004),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_913),
.A2(n_950),
.B(n_999),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_935),
.A2(n_341),
.B(n_338),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_973),
.A2(n_337),
.B(n_333),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_940),
.B(n_275),
.Y(n_1134)
);

OAI21xp33_ASAP7_75t_L g1135 ( 
.A1(n_1028),
.A2(n_329),
.B(n_328),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_971),
.Y(n_1136)
);

BUFx5_ASAP7_75t_L g1137 ( 
.A(n_1032),
.Y(n_1137)
);

AND2x4_ASAP7_75t_L g1138 ( 
.A(n_941),
.B(n_28),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_928),
.A2(n_327),
.B(n_324),
.Y(n_1139)
);

INVx5_ASAP7_75t_L g1140 ( 
.A(n_971),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_953),
.B(n_276),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1050),
.A2(n_320),
.B1(n_311),
.B2(n_309),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_SL g1143 ( 
.A1(n_1063),
.A2(n_302),
.B1(n_298),
.B2(n_296),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_926),
.B(n_28),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_930),
.A2(n_294),
.B(n_292),
.Y(n_1145)
);

NAND3xp33_ASAP7_75t_SL g1146 ( 
.A(n_1035),
.B(n_290),
.C(n_279),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_983),
.A2(n_277),
.B(n_273),
.C(n_34),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_971),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_1006),
.B(n_29),
.Y(n_1149)
);

OAI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1052),
.A2(n_30),
.B1(n_36),
.B2(n_37),
.Y(n_1150)
);

INVxp67_ASAP7_75t_L g1151 ( 
.A(n_926),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1002),
.B(n_991),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_953),
.B(n_36),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_992),
.B(n_38),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1009),
.B(n_38),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_SL g1156 ( 
.A(n_1006),
.B(n_273),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_968),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_1157)
);

AO21x2_ASAP7_75t_L g1158 ( 
.A1(n_1034),
.A2(n_273),
.B(n_80),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_933),
.A2(n_81),
.B(n_205),
.Y(n_1159)
);

NAND2xp33_ASAP7_75t_L g1160 ( 
.A(n_987),
.B(n_273),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_989),
.A2(n_40),
.B1(n_42),
.B2(n_44),
.Y(n_1161)
);

O2A1O1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_960),
.A2(n_45),
.B(n_46),
.C(n_47),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1065),
.A2(n_273),
.B1(n_51),
.B2(n_53),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_969),
.A2(n_104),
.B(n_199),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_979),
.B(n_48),
.Y(n_1165)
);

O2A1O1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_949),
.A2(n_48),
.B(n_54),
.C(n_55),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_977),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1047),
.A2(n_122),
.B(n_192),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1036),
.B(n_60),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_L g1170 ( 
.A1(n_1018),
.A2(n_273),
.B1(n_62),
.B2(n_65),
.Y(n_1170)
);

A2O1A1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1029),
.A2(n_273),
.B(n_66),
.C(n_68),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_976),
.A2(n_141),
.B(n_191),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_1036),
.B(n_60),
.Y(n_1173)
);

BUFx4f_ASAP7_75t_L g1174 ( 
.A(n_948),
.Y(n_1174)
);

INVx1_ASAP7_75t_SL g1175 ( 
.A(n_932),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1031),
.B(n_75),
.Y(n_1176)
);

OR2x2_ASAP7_75t_L g1177 ( 
.A(n_1067),
.B(n_77),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_978),
.A2(n_79),
.B(n_94),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_948),
.B(n_99),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1046),
.B(n_273),
.Y(n_1180)
);

INVx2_ASAP7_75t_SL g1181 ( 
.A(n_987),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_982),
.A2(n_103),
.B(n_108),
.Y(n_1182)
);

A2O1A1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_908),
.A2(n_968),
.B(n_916),
.C(n_997),
.Y(n_1183)
);

INVx3_ASAP7_75t_L g1184 ( 
.A(n_998),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1040),
.A2(n_120),
.B(n_135),
.Y(n_1185)
);

O2A1O1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1008),
.A2(n_160),
.B(n_165),
.C(n_172),
.Y(n_1186)
);

NOR2x1_ASAP7_75t_R g1187 ( 
.A(n_998),
.B(n_175),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1030),
.B(n_178),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_975),
.A2(n_1024),
.B1(n_1000),
.B2(n_927),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_1019),
.B(n_185),
.Y(n_1190)
);

BUFx8_ASAP7_75t_L g1191 ( 
.A(n_1014),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_946),
.A2(n_954),
.B(n_1001),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1017),
.A2(n_957),
.B1(n_1070),
.B2(n_988),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_SL g1194 ( 
.A(n_1007),
.B(n_1021),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1071),
.B(n_1012),
.Y(n_1195)
);

O2A1O1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_921),
.A2(n_1074),
.B(n_1064),
.C(n_1039),
.Y(n_1196)
);

BUFx3_ASAP7_75t_L g1197 ( 
.A(n_1071),
.Y(n_1197)
);

INVx3_ASAP7_75t_L g1198 ( 
.A(n_1007),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1069),
.A2(n_1060),
.B1(n_1038),
.B2(n_1055),
.Y(n_1199)
);

INVx4_ASAP7_75t_L g1200 ( 
.A(n_1014),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1051),
.A2(n_1053),
.B1(n_1056),
.B2(n_929),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_981),
.Y(n_1202)
);

INVx4_ASAP7_75t_L g1203 ( 
.A(n_1014),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_1012),
.B(n_1016),
.Y(n_1204)
);

CKINVDCx12_ASAP7_75t_R g1205 ( 
.A(n_1037),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_1020),
.B(n_1021),
.Y(n_1206)
);

O2A1O1Ixp33_ASAP7_75t_SL g1207 ( 
.A1(n_1022),
.A2(n_1041),
.B(n_1045),
.C(n_974),
.Y(n_1207)
);

NOR3xp33_ASAP7_75t_L g1208 ( 
.A(n_1044),
.B(n_1039),
.C(n_1027),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1066),
.A2(n_1015),
.B1(n_1061),
.B2(n_1025),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1020),
.B(n_1066),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_934),
.A2(n_990),
.B(n_985),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1025),
.B(n_1058),
.Y(n_1212)
);

O2A1O1Ixp33_ASAP7_75t_L g1213 ( 
.A1(n_1068),
.A2(n_1027),
.B(n_1073),
.C(n_1072),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_943),
.B(n_958),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_1075),
.B(n_1062),
.Y(n_1215)
);

INVx3_ASAP7_75t_SL g1216 ( 
.A(n_1022),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_1059),
.B(n_1010),
.Y(n_1217)
);

INVx3_ASAP7_75t_L g1218 ( 
.A(n_1191),
.Y(n_1218)
);

OAI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1080),
.A2(n_1005),
.B(n_947),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_1118),
.B(n_1041),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1189),
.A2(n_1045),
.B(n_1013),
.Y(n_1221)
);

AO31x2_ASAP7_75t_L g1222 ( 
.A1(n_1086),
.A2(n_901),
.A3(n_1043),
.B(n_1054),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_SL g1223 ( 
.A(n_1118),
.B(n_1042),
.Y(n_1223)
);

INVx5_ASAP7_75t_L g1224 ( 
.A(n_1092),
.Y(n_1224)
);

BUFx2_ASAP7_75t_L g1225 ( 
.A(n_1081),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1118),
.B(n_1003),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1088),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1114),
.A2(n_947),
.B(n_955),
.C(n_1061),
.Y(n_1228)
);

BUFx12f_ASAP7_75t_L g1229 ( 
.A(n_1084),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1192),
.A2(n_914),
.B(n_995),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1211),
.A2(n_996),
.B(n_909),
.Y(n_1231)
);

OA21x2_ASAP7_75t_L g1232 ( 
.A1(n_1095),
.A2(n_1011),
.B(n_1023),
.Y(n_1232)
);

OAI22x1_ASAP7_75t_L g1233 ( 
.A1(n_1175),
.A2(n_1026),
.B1(n_907),
.B2(n_918),
.Y(n_1233)
);

OAI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1095),
.A2(n_1183),
.B(n_1189),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1152),
.B(n_1151),
.Y(n_1235)
);

AO31x2_ASAP7_75t_L g1236 ( 
.A1(n_1201),
.A2(n_1079),
.A3(n_1117),
.B(n_1193),
.Y(n_1236)
);

INVx3_ASAP7_75t_L g1237 ( 
.A(n_1191),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1126),
.A2(n_1188),
.B(n_1212),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_1100),
.Y(n_1239)
);

CKINVDCx20_ASAP7_75t_R g1240 ( 
.A(n_1130),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1217),
.A2(n_1131),
.B(n_1076),
.Y(n_1241)
);

O2A1O1Ixp33_ASAP7_75t_SL g1242 ( 
.A1(n_1171),
.A2(n_1119),
.B(n_1147),
.C(n_1089),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1090),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_SL g1244 ( 
.A(n_1137),
.B(n_1096),
.Y(n_1244)
);

INVx4_ASAP7_75t_L g1245 ( 
.A(n_1092),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1201),
.A2(n_1193),
.B(n_1131),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1215),
.A2(n_1196),
.B(n_1185),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1164),
.A2(n_1159),
.B(n_1077),
.Y(n_1248)
);

OR2x6_ASAP7_75t_L g1249 ( 
.A(n_1108),
.B(n_1129),
.Y(n_1249)
);

AOI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1169),
.A2(n_1173),
.B1(n_1165),
.B2(n_1087),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1168),
.A2(n_1207),
.B(n_1178),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1113),
.B(n_1121),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1172),
.A2(n_1182),
.B(n_1213),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1144),
.B(n_1149),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_SL g1255 ( 
.A1(n_1154),
.A2(n_1155),
.B(n_1176),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_1137),
.B(n_1174),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_SL g1257 ( 
.A(n_1118),
.B(n_1175),
.Y(n_1257)
);

AOI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1157),
.A2(n_1153),
.B1(n_1124),
.B2(n_1120),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1106),
.A2(n_1158),
.B(n_1174),
.Y(n_1259)
);

INVx3_ASAP7_75t_L g1260 ( 
.A(n_1085),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_SL g1261 ( 
.A1(n_1123),
.A2(n_1186),
.B(n_1210),
.Y(n_1261)
);

AOI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1120),
.A2(n_1150),
.B1(n_1146),
.B2(n_1149),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1097),
.Y(n_1263)
);

AOI222xp33_ASAP7_75t_L g1264 ( 
.A1(n_1150),
.A2(n_1161),
.B1(n_1167),
.B2(n_1108),
.C1(n_1129),
.C2(n_1099),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1209),
.A2(n_1109),
.B(n_1180),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1110),
.B(n_1141),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_1103),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1115),
.B(n_1101),
.Y(n_1268)
);

OR2x2_ASAP7_75t_L g1269 ( 
.A(n_1105),
.B(n_1127),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_SL g1270 ( 
.A(n_1187),
.B(n_1156),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1158),
.A2(n_1194),
.B(n_1208),
.Y(n_1271)
);

BUFx10_ASAP7_75t_L g1272 ( 
.A(n_1138),
.Y(n_1272)
);

BUFx10_ASAP7_75t_L g1273 ( 
.A(n_1128),
.Y(n_1273)
);

INVx4_ASAP7_75t_L g1274 ( 
.A(n_1092),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1194),
.A2(n_1093),
.B(n_1204),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1202),
.Y(n_1276)
);

NOR2xp67_ASAP7_75t_L g1277 ( 
.A(n_1107),
.B(n_1085),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1216),
.B(n_1197),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1137),
.Y(n_1279)
);

INVx2_ASAP7_75t_SL g1280 ( 
.A(n_1082),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1161),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1214),
.A2(n_1179),
.B(n_1140),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1177),
.B(n_1125),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1167),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1205),
.Y(n_1285)
);

O2A1O1Ixp33_ASAP7_75t_SL g1286 ( 
.A1(n_1206),
.A2(n_1190),
.B(n_1166),
.C(n_1162),
.Y(n_1286)
);

OAI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1102),
.A2(n_1091),
.B(n_1163),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_SL g1288 ( 
.A(n_1137),
.B(n_1078),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1184),
.A2(n_1198),
.B(n_1107),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_1143),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1137),
.Y(n_1291)
);

AND2x4_ASAP7_75t_L g1292 ( 
.A(n_1082),
.B(n_1083),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1179),
.A2(n_1140),
.B(n_1160),
.Y(n_1293)
);

AOI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1078),
.A2(n_1170),
.B1(n_1156),
.B2(n_1104),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1140),
.A2(n_1116),
.B(n_1135),
.Y(n_1295)
);

OA22x2_ASAP7_75t_L g1296 ( 
.A1(n_1094),
.A2(n_1134),
.B1(n_1083),
.B2(n_1181),
.Y(n_1296)
);

A2O1A1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1195),
.A2(n_1132),
.B(n_1145),
.C(n_1139),
.Y(n_1297)
);

AO31x2_ASAP7_75t_L g1298 ( 
.A1(n_1133),
.A2(n_1142),
.A3(n_1122),
.B(n_1203),
.Y(n_1298)
);

OAI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1200),
.A2(n_1203),
.B(n_1140),
.Y(n_1299)
);

BUFx4f_ASAP7_75t_L g1300 ( 
.A(n_1111),
.Y(n_1300)
);

CKINVDCx6p67_ASAP7_75t_R g1301 ( 
.A(n_1111),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1199),
.B(n_1184),
.Y(n_1302)
);

AO32x2_ASAP7_75t_L g1303 ( 
.A1(n_1200),
.A2(n_1111),
.A3(n_1136),
.B1(n_1148),
.B2(n_1198),
.Y(n_1303)
);

OA21x2_ASAP7_75t_L g1304 ( 
.A1(n_1136),
.A2(n_1095),
.B(n_1131),
.Y(n_1304)
);

CKINVDCx20_ASAP7_75t_R g1305 ( 
.A(n_1136),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_1148),
.B(n_939),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1148),
.A2(n_1192),
.B(n_1211),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1080),
.A2(n_944),
.B(n_984),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1080),
.A2(n_944),
.B(n_984),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1080),
.A2(n_944),
.B(n_984),
.Y(n_1310)
);

OAI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1080),
.A2(n_937),
.B(n_962),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_1081),
.Y(n_1312)
);

O2A1O1Ixp33_ASAP7_75t_SL g1313 ( 
.A1(n_1126),
.A2(n_962),
.B(n_793),
.C(n_937),
.Y(n_1313)
);

INVx1_ASAP7_75t_SL g1314 ( 
.A(n_1216),
.Y(n_1314)
);

BUFx4_ASAP7_75t_SL g1315 ( 
.A(n_1084),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1080),
.A2(n_944),
.B(n_984),
.Y(n_1316)
);

O2A1O1Ixp33_ASAP7_75t_SL g1317 ( 
.A1(n_1126),
.A2(n_962),
.B(n_793),
.C(n_937),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1088),
.Y(n_1318)
);

AO31x2_ASAP7_75t_L g1319 ( 
.A1(n_1086),
.A2(n_970),
.A3(n_901),
.B(n_1080),
.Y(n_1319)
);

OAI22x1_ASAP7_75t_L g1320 ( 
.A1(n_1175),
.A2(n_915),
.B1(n_925),
.B2(n_1114),
.Y(n_1320)
);

NAND3xp33_ASAP7_75t_L g1321 ( 
.A(n_1114),
.B(n_1171),
.C(n_1119),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1088),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1080),
.A2(n_944),
.B(n_984),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1098),
.A2(n_715),
.B1(n_642),
.B2(n_623),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1080),
.A2(n_944),
.B(n_984),
.Y(n_1325)
);

AOI221xp5_ASAP7_75t_L g1326 ( 
.A1(n_1114),
.A2(n_701),
.B1(n_1098),
.B2(n_732),
.C(n_775),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1112),
.B(n_744),
.Y(n_1327)
);

NOR2xp67_ASAP7_75t_SL g1328 ( 
.A(n_1084),
.B(n_945),
.Y(n_1328)
);

HB1xp67_ASAP7_75t_L g1329 ( 
.A(n_1081),
.Y(n_1329)
);

INVx4_ASAP7_75t_L g1330 ( 
.A(n_1092),
.Y(n_1330)
);

BUFx2_ASAP7_75t_L g1331 ( 
.A(n_1081),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1080),
.A2(n_944),
.B(n_984),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1081),
.B(n_912),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1112),
.B(n_744),
.Y(n_1334)
);

XOR2xp5_ASAP7_75t_L g1335 ( 
.A(n_1084),
.B(n_782),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1192),
.A2(n_1211),
.B(n_944),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1080),
.A2(n_944),
.B(n_984),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1114),
.B(n_804),
.Y(n_1338)
);

OA21x2_ASAP7_75t_L g1339 ( 
.A1(n_1095),
.A2(n_1131),
.B(n_944),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1089),
.A2(n_1114),
.B1(n_757),
.B2(n_752),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1080),
.A2(n_944),
.B(n_984),
.Y(n_1341)
);

O2A1O1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1114),
.A2(n_1089),
.B(n_1119),
.C(n_1096),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1098),
.A2(n_715),
.B1(n_642),
.B2(n_623),
.Y(n_1343)
);

O2A1O1Ixp33_ASAP7_75t_L g1344 ( 
.A1(n_1114),
.A2(n_1089),
.B(n_1119),
.C(n_1096),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1088),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1080),
.A2(n_944),
.B(n_984),
.Y(n_1346)
);

AOI31xp67_ASAP7_75t_L g1347 ( 
.A1(n_1217),
.A2(n_1215),
.A3(n_974),
.B(n_1212),
.Y(n_1347)
);

AOI22x1_ASAP7_75t_SL g1348 ( 
.A1(n_1175),
.A2(n_659),
.B1(n_782),
.B2(n_707),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_1100),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_1092),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1080),
.A2(n_944),
.B(n_984),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1080),
.A2(n_944),
.B(n_984),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1112),
.B(n_744),
.Y(n_1353)
);

OAI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1114),
.A2(n_757),
.B(n_937),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1080),
.A2(n_937),
.B(n_962),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1088),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1088),
.Y(n_1357)
);

AOI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1114),
.A2(n_925),
.B1(n_732),
.B2(n_1098),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1192),
.A2(n_1211),
.B(n_944),
.Y(n_1359)
);

OAI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1080),
.A2(n_937),
.B(n_962),
.Y(n_1360)
);

AND2x6_ASAP7_75t_L g1361 ( 
.A(n_1108),
.B(n_1129),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1088),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1080),
.A2(n_944),
.B(n_984),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1080),
.A2(n_944),
.B(n_984),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1081),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1112),
.B(n_744),
.Y(n_1366)
);

AOI221x1_ASAP7_75t_L g1367 ( 
.A1(n_1171),
.A2(n_1150),
.B1(n_1161),
.B2(n_1147),
.C(n_1117),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1080),
.A2(n_944),
.B(n_984),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1080),
.A2(n_944),
.B(n_984),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1080),
.A2(n_944),
.B(n_984),
.Y(n_1370)
);

CKINVDCx20_ASAP7_75t_R g1371 ( 
.A(n_1239),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1358),
.A2(n_1326),
.B1(n_1250),
.B2(n_1324),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1250),
.A2(n_1343),
.B1(n_1320),
.B2(n_1264),
.Y(n_1373)
);

INVx1_ASAP7_75t_SL g1374 ( 
.A(n_1314),
.Y(n_1374)
);

INVx2_ASAP7_75t_SL g1375 ( 
.A(n_1273),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_SL g1376 ( 
.A1(n_1283),
.A2(n_1270),
.B1(n_1361),
.B2(n_1354),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1264),
.A2(n_1321),
.B1(n_1258),
.B2(n_1284),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1319),
.Y(n_1378)
);

INVx6_ASAP7_75t_L g1379 ( 
.A(n_1224),
.Y(n_1379)
);

INVx1_ASAP7_75t_SL g1380 ( 
.A(n_1314),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1243),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1319),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1258),
.A2(n_1281),
.B1(n_1262),
.B2(n_1234),
.Y(n_1383)
);

CKINVDCx11_ASAP7_75t_R g1384 ( 
.A(n_1229),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1262),
.A2(n_1234),
.B1(n_1246),
.B2(n_1340),
.Y(n_1385)
);

AOI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1252),
.A2(n_1338),
.B1(n_1290),
.B2(n_1361),
.Y(n_1386)
);

OAI22xp33_ASAP7_75t_R g1387 ( 
.A1(n_1266),
.A2(n_1269),
.B1(n_1329),
.B2(n_1365),
.Y(n_1387)
);

CKINVDCx16_ASAP7_75t_R g1388 ( 
.A(n_1335),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1305),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1263),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1246),
.A2(n_1361),
.B1(n_1333),
.B2(n_1294),
.Y(n_1391)
);

INVx6_ASAP7_75t_L g1392 ( 
.A(n_1224),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1294),
.A2(n_1287),
.B1(n_1355),
.B2(n_1360),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1287),
.A2(n_1355),
.B1(n_1360),
.B2(n_1311),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1318),
.Y(n_1395)
);

INVx8_ASAP7_75t_L g1396 ( 
.A(n_1249),
.Y(n_1396)
);

BUFx4_ASAP7_75t_SL g1397 ( 
.A(n_1349),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1342),
.A2(n_1344),
.B1(n_1249),
.B2(n_1311),
.Y(n_1398)
);

OAI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1367),
.A2(n_1268),
.B1(n_1366),
.B2(n_1327),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1244),
.A2(n_1331),
.B1(n_1225),
.B2(n_1334),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1296),
.A2(n_1339),
.B1(n_1254),
.B2(n_1255),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1353),
.B(n_1312),
.Y(n_1402)
);

CKINVDCx20_ASAP7_75t_R g1403 ( 
.A(n_1267),
.Y(n_1403)
);

INVx5_ASAP7_75t_L g1404 ( 
.A(n_1218),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_1348),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1322),
.B(n_1345),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1356),
.A2(n_1357),
.B1(n_1362),
.B2(n_1276),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_1285),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1292),
.B(n_1278),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1347),
.Y(n_1410)
);

INVx1_ASAP7_75t_SL g1411 ( 
.A(n_1272),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1257),
.B(n_1272),
.Y(n_1412)
);

INVx6_ASAP7_75t_L g1413 ( 
.A(n_1245),
.Y(n_1413)
);

INVx1_ASAP7_75t_SL g1414 ( 
.A(n_1350),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_SL g1415 ( 
.A1(n_1257),
.A2(n_1223),
.B1(n_1261),
.B2(n_1271),
.Y(n_1415)
);

OAI21xp33_ASAP7_75t_SL g1416 ( 
.A1(n_1256),
.A2(n_1289),
.B(n_1288),
.Y(n_1416)
);

INVx2_ASAP7_75t_SL g1417 ( 
.A(n_1218),
.Y(n_1417)
);

CKINVDCx8_ASAP7_75t_R g1418 ( 
.A(n_1350),
.Y(n_1418)
);

BUFx3_ASAP7_75t_L g1419 ( 
.A(n_1237),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1303),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1302),
.A2(n_1304),
.B1(n_1219),
.B2(n_1259),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1219),
.A2(n_1221),
.B1(n_1238),
.B2(n_1306),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1303),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_1237),
.Y(n_1424)
);

OAI22x1_ASAP7_75t_L g1425 ( 
.A1(n_1220),
.A2(n_1226),
.B1(n_1279),
.B2(n_1291),
.Y(n_1425)
);

OAI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1282),
.A2(n_1247),
.B1(n_1369),
.B2(n_1316),
.Y(n_1426)
);

CKINVDCx11_ASAP7_75t_R g1427 ( 
.A(n_1301),
.Y(n_1427)
);

OAI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1308),
.A2(n_1370),
.B1(n_1368),
.B2(n_1309),
.Y(n_1428)
);

BUFx12f_ASAP7_75t_L g1429 ( 
.A(n_1245),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_1274),
.Y(n_1430)
);

BUFx8_ASAP7_75t_L g1431 ( 
.A(n_1280),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1223),
.A2(n_1265),
.B1(n_1220),
.B2(n_1364),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1330),
.B(n_1260),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1310),
.A2(n_1363),
.B1(n_1346),
.B2(n_1352),
.Y(n_1434)
);

INVx4_ASAP7_75t_L g1435 ( 
.A(n_1300),
.Y(n_1435)
);

AOI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1242),
.A2(n_1328),
.B1(n_1286),
.B2(n_1226),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_SL g1437 ( 
.A1(n_1293),
.A2(n_1251),
.B1(n_1295),
.B2(n_1275),
.Y(n_1437)
);

INVx3_ASAP7_75t_SL g1438 ( 
.A(n_1260),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1323),
.A2(n_1341),
.B1(n_1337),
.B2(n_1332),
.Y(n_1439)
);

OAI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1325),
.A2(n_1351),
.B1(n_1241),
.B2(n_1277),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_SL g1441 ( 
.A(n_1299),
.Y(n_1441)
);

AOI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1313),
.A2(n_1317),
.B1(n_1233),
.B2(n_1228),
.Y(n_1442)
);

OAI22xp33_ASAP7_75t_R g1443 ( 
.A1(n_1236),
.A2(n_1297),
.B1(n_1253),
.B2(n_1298),
.Y(n_1443)
);

CKINVDCx20_ASAP7_75t_R g1444 ( 
.A(n_1299),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_SL g1445 ( 
.A1(n_1236),
.A2(n_1232),
.B1(n_1248),
.B2(n_1359),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1232),
.A2(n_1236),
.B1(n_1336),
.B2(n_1230),
.Y(n_1446)
);

BUFx4f_ASAP7_75t_SL g1447 ( 
.A(n_1298),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1307),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1231),
.A2(n_1033),
.B1(n_1358),
.B2(n_1326),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_SL g1450 ( 
.A1(n_1298),
.A2(n_898),
.B1(n_1283),
.B2(n_411),
.Y(n_1450)
);

INVx3_ASAP7_75t_L g1451 ( 
.A(n_1222),
.Y(n_1451)
);

INVx4_ASAP7_75t_L g1452 ( 
.A(n_1222),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1315),
.Y(n_1453)
);

INVxp67_ASAP7_75t_SL g1454 ( 
.A(n_1235),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1227),
.Y(n_1455)
);

BUFx10_ASAP7_75t_L g1456 ( 
.A(n_1239),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1227),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1227),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1358),
.B(n_1235),
.Y(n_1459)
);

BUFx6f_ASAP7_75t_L g1460 ( 
.A(n_1303),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1358),
.A2(n_1033),
.B1(n_1326),
.B2(n_1250),
.Y(n_1461)
);

INVx1_ASAP7_75t_SL g1462 ( 
.A(n_1314),
.Y(n_1462)
);

BUFx12f_ASAP7_75t_L g1463 ( 
.A(n_1239),
.Y(n_1463)
);

CKINVDCx20_ASAP7_75t_R g1464 ( 
.A(n_1239),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1227),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_SL g1466 ( 
.A1(n_1283),
.A2(n_898),
.B1(n_411),
.B2(n_423),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1227),
.Y(n_1467)
);

BUFx2_ASAP7_75t_SL g1468 ( 
.A(n_1240),
.Y(n_1468)
);

BUFx8_ASAP7_75t_L g1469 ( 
.A(n_1229),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1358),
.A2(n_1033),
.B1(n_1326),
.B2(n_1250),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1254),
.B(n_1333),
.Y(n_1471)
);

CKINVDCx11_ASAP7_75t_R g1472 ( 
.A(n_1229),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1358),
.A2(n_1033),
.B1(n_1326),
.B2(n_1250),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1227),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1227),
.Y(n_1475)
);

BUFx2_ASAP7_75t_L g1476 ( 
.A(n_1305),
.Y(n_1476)
);

BUFx3_ASAP7_75t_L g1477 ( 
.A(n_1305),
.Y(n_1477)
);

CKINVDCx20_ASAP7_75t_R g1478 ( 
.A(n_1239),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1312),
.Y(n_1479)
);

BUFx2_ASAP7_75t_SL g1480 ( 
.A(n_1240),
.Y(n_1480)
);

BUFx10_ASAP7_75t_L g1481 ( 
.A(n_1239),
.Y(n_1481)
);

CKINVDCx11_ASAP7_75t_R g1482 ( 
.A(n_1229),
.Y(n_1482)
);

CKINVDCx6p67_ASAP7_75t_R g1483 ( 
.A(n_1229),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1358),
.A2(n_1033),
.B1(n_1326),
.B2(n_1250),
.Y(n_1484)
);

CKINVDCx20_ASAP7_75t_R g1485 ( 
.A(n_1239),
.Y(n_1485)
);

BUFx6f_ASAP7_75t_L g1486 ( 
.A(n_1303),
.Y(n_1486)
);

OAI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1358),
.A2(n_1250),
.B1(n_1258),
.B2(n_1249),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1358),
.A2(n_1033),
.B1(n_1326),
.B2(n_1250),
.Y(n_1488)
);

CKINVDCx11_ASAP7_75t_R g1489 ( 
.A(n_1229),
.Y(n_1489)
);

BUFx3_ASAP7_75t_L g1490 ( 
.A(n_1305),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1358),
.A2(n_1033),
.B1(n_1326),
.B2(n_1250),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1358),
.A2(n_1033),
.B1(n_1326),
.B2(n_1250),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_SL g1493 ( 
.A1(n_1283),
.A2(n_898),
.B1(n_411),
.B2(n_423),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1358),
.A2(n_1033),
.B1(n_1326),
.B2(n_1250),
.Y(n_1494)
);

BUFx4f_ASAP7_75t_SL g1495 ( 
.A(n_1229),
.Y(n_1495)
);

INVx4_ASAP7_75t_L g1496 ( 
.A(n_1224),
.Y(n_1496)
);

INVx4_ASAP7_75t_L g1497 ( 
.A(n_1224),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_SL g1498 ( 
.A1(n_1283),
.A2(n_898),
.B1(n_411),
.B2(n_423),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1358),
.A2(n_1033),
.B1(n_1326),
.B2(n_1250),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1358),
.A2(n_1250),
.B1(n_1326),
.B2(n_1258),
.Y(n_1500)
);

OAI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1358),
.A2(n_1250),
.B1(n_1258),
.B2(n_1249),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1227),
.Y(n_1502)
);

BUFx12f_ASAP7_75t_L g1503 ( 
.A(n_1239),
.Y(n_1503)
);

INVx1_ASAP7_75t_SL g1504 ( 
.A(n_1314),
.Y(n_1504)
);

CKINVDCx11_ASAP7_75t_R g1505 ( 
.A(n_1229),
.Y(n_1505)
);

BUFx12f_ASAP7_75t_L g1506 ( 
.A(n_1239),
.Y(n_1506)
);

A2O1A1Ixp33_ASAP7_75t_L g1507 ( 
.A1(n_1461),
.A2(n_1470),
.B(n_1494),
.C(n_1492),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1420),
.Y(n_1508)
);

AO21x2_ASAP7_75t_L g1509 ( 
.A1(n_1428),
.A2(n_1382),
.B(n_1378),
.Y(n_1509)
);

INVx2_ASAP7_75t_SL g1510 ( 
.A(n_1460),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1479),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1454),
.Y(n_1512)
);

CKINVDCx20_ASAP7_75t_R g1513 ( 
.A(n_1371),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1466),
.A2(n_1498),
.B1(n_1493),
.B2(n_1470),
.Y(n_1514)
);

BUFx6f_ASAP7_75t_L g1515 ( 
.A(n_1486),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1400),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1459),
.B(n_1402),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1399),
.B(n_1377),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1434),
.A2(n_1439),
.B(n_1446),
.Y(n_1519)
);

INVx2_ASAP7_75t_SL g1520 ( 
.A(n_1404),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1406),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1423),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1381),
.Y(n_1523)
);

INVx3_ASAP7_75t_L g1524 ( 
.A(n_1410),
.Y(n_1524)
);

OR2x6_ASAP7_75t_L g1525 ( 
.A(n_1396),
.B(n_1425),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1390),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1394),
.B(n_1383),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1383),
.B(n_1385),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1395),
.Y(n_1529)
);

BUFx2_ASAP7_75t_L g1530 ( 
.A(n_1416),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1455),
.Y(n_1531)
);

BUFx2_ASAP7_75t_L g1532 ( 
.A(n_1451),
.Y(n_1532)
);

AO31x2_ASAP7_75t_L g1533 ( 
.A1(n_1500),
.A2(n_1452),
.A3(n_1398),
.B(n_1448),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1457),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1458),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1399),
.B(n_1377),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1465),
.Y(n_1537)
);

BUFx2_ASAP7_75t_L g1538 ( 
.A(n_1447),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1467),
.Y(n_1539)
);

NAND2x1_ASAP7_75t_L g1540 ( 
.A(n_1422),
.B(n_1442),
.Y(n_1540)
);

CKINVDCx6p67_ASAP7_75t_R g1541 ( 
.A(n_1388),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1474),
.Y(n_1542)
);

OAI21x1_ASAP7_75t_L g1543 ( 
.A1(n_1434),
.A2(n_1439),
.B(n_1446),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1475),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1502),
.Y(n_1545)
);

OAI21x1_ASAP7_75t_L g1546 ( 
.A1(n_1432),
.A2(n_1422),
.B(n_1421),
.Y(n_1546)
);

AO21x1_ASAP7_75t_SL g1547 ( 
.A1(n_1385),
.A2(n_1393),
.B(n_1449),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1393),
.B(n_1421),
.Y(n_1548)
);

BUFx2_ASAP7_75t_L g1549 ( 
.A(n_1447),
.Y(n_1549)
);

INVx3_ASAP7_75t_L g1550 ( 
.A(n_1441),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1443),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1407),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_1444),
.Y(n_1553)
);

AO21x2_ASAP7_75t_L g1554 ( 
.A1(n_1426),
.A2(n_1440),
.B(n_1501),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1440),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1426),
.Y(n_1556)
);

OAI21xp5_ASAP7_75t_L g1557 ( 
.A1(n_1461),
.A2(n_1488),
.B(n_1473),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1445),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1432),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1473),
.A2(n_1488),
.B1(n_1484),
.B2(n_1491),
.Y(n_1560)
);

AOI21x1_ASAP7_75t_L g1561 ( 
.A1(n_1412),
.A2(n_1433),
.B(n_1409),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1415),
.Y(n_1562)
);

INVxp33_ASAP7_75t_L g1563 ( 
.A(n_1471),
.Y(n_1563)
);

AO21x2_ASAP7_75t_L g1564 ( 
.A1(n_1487),
.A2(n_1501),
.B(n_1436),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1487),
.B(n_1373),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1437),
.Y(n_1566)
);

INVx2_ASAP7_75t_SL g1567 ( 
.A(n_1396),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1401),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1401),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1449),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1391),
.B(n_1372),
.Y(n_1571)
);

INVx3_ASAP7_75t_L g1572 ( 
.A(n_1419),
.Y(n_1572)
);

BUFx2_ASAP7_75t_L g1573 ( 
.A(n_1419),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1391),
.B(n_1373),
.Y(n_1574)
);

OA21x2_ASAP7_75t_L g1575 ( 
.A1(n_1484),
.A2(n_1491),
.B(n_1492),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1376),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1494),
.B(n_1499),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1499),
.B(n_1386),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1387),
.Y(n_1579)
);

OA21x2_ASAP7_75t_L g1580 ( 
.A1(n_1414),
.A2(n_1450),
.B(n_1374),
.Y(n_1580)
);

OAI322xp33_ASAP7_75t_L g1581 ( 
.A1(n_1380),
.A2(n_1462),
.A3(n_1504),
.B1(n_1417),
.B2(n_1405),
.C1(n_1411),
.C2(n_1375),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1477),
.B(n_1490),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1490),
.B(n_1389),
.Y(n_1583)
);

AO21x2_ASAP7_75t_L g1584 ( 
.A1(n_1379),
.A2(n_1392),
.B(n_1438),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1438),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1476),
.B(n_1480),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1418),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1496),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1413),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1497),
.B(n_1435),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1468),
.B(n_1424),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1431),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1431),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1430),
.Y(n_1594)
);

NAND2x1p5_ASAP7_75t_L g1595 ( 
.A(n_1429),
.B(n_1427),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1408),
.Y(n_1596)
);

NOR2x1_ASAP7_75t_SL g1597 ( 
.A(n_1584),
.B(n_1525),
.Y(n_1597)
);

AOI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1560),
.A2(n_1483),
.B1(n_1495),
.B2(n_1403),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1551),
.B(n_1469),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1582),
.B(n_1481),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1582),
.B(n_1481),
.Y(n_1601)
);

INVx3_ASAP7_75t_L g1602 ( 
.A(n_1572),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1563),
.B(n_1456),
.Y(n_1603)
);

O2A1O1Ixp33_ASAP7_75t_L g1604 ( 
.A1(n_1507),
.A2(n_1478),
.B(n_1485),
.C(n_1464),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1526),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_1513),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1583),
.B(n_1456),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1528),
.A2(n_1495),
.B1(n_1453),
.B2(n_1463),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1551),
.B(n_1469),
.Y(n_1609)
);

AO32x2_ASAP7_75t_L g1610 ( 
.A1(n_1510),
.A2(n_1384),
.A3(n_1505),
.B1(n_1472),
.B2(n_1482),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1512),
.B(n_1503),
.Y(n_1611)
);

BUFx2_ASAP7_75t_L g1612 ( 
.A(n_1573),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1557),
.A2(n_1489),
.B1(n_1506),
.B2(n_1397),
.Y(n_1613)
);

INVxp67_ASAP7_75t_L g1614 ( 
.A(n_1530),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1511),
.B(n_1521),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_1541),
.Y(n_1616)
);

OAI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1518),
.A2(n_1536),
.B(n_1528),
.Y(n_1617)
);

OAI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1540),
.A2(n_1527),
.B(n_1566),
.Y(n_1618)
);

O2A1O1Ixp33_ASAP7_75t_SL g1619 ( 
.A1(n_1540),
.A2(n_1592),
.B(n_1593),
.C(n_1516),
.Y(n_1619)
);

AO32x2_ASAP7_75t_L g1620 ( 
.A1(n_1510),
.A2(n_1520),
.A3(n_1567),
.B1(n_1531),
.B2(n_1561),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_SL g1621 ( 
.A(n_1579),
.B(n_1550),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1553),
.B(n_1586),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1517),
.B(n_1548),
.Y(n_1623)
);

OA21x2_ASAP7_75t_L g1624 ( 
.A1(n_1519),
.A2(n_1543),
.B(n_1546),
.Y(n_1624)
);

OAI22xp5_ASAP7_75t_SL g1625 ( 
.A1(n_1579),
.A2(n_1595),
.B1(n_1514),
.B2(n_1575),
.Y(n_1625)
);

OAI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1527),
.A2(n_1565),
.B1(n_1577),
.B2(n_1575),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1548),
.B(n_1556),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1556),
.B(n_1555),
.Y(n_1628)
);

OAI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1566),
.A2(n_1575),
.B(n_1578),
.Y(n_1629)
);

AND2x2_ASAP7_75t_SL g1630 ( 
.A(n_1530),
.B(n_1538),
.Y(n_1630)
);

A2O1A1Ixp33_ASAP7_75t_L g1631 ( 
.A1(n_1578),
.A2(n_1574),
.B(n_1571),
.C(n_1562),
.Y(n_1631)
);

A2O1A1Ixp33_ASAP7_75t_L g1632 ( 
.A1(n_1574),
.A2(n_1571),
.B(n_1562),
.C(n_1576),
.Y(n_1632)
);

OAI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1555),
.A2(n_1570),
.B(n_1543),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1581),
.B(n_1564),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1524),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1523),
.Y(n_1636)
);

AOI221xp5_ASAP7_75t_L g1637 ( 
.A1(n_1581),
.A2(n_1558),
.B1(n_1552),
.B2(n_1568),
.C(n_1569),
.Y(n_1637)
);

AOI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1554),
.A2(n_1564),
.B(n_1509),
.Y(n_1638)
);

INVx1_ASAP7_75t_SL g1639 ( 
.A(n_1541),
.Y(n_1639)
);

AO32x2_ASAP7_75t_L g1640 ( 
.A1(n_1520),
.A2(n_1567),
.A3(n_1561),
.B1(n_1552),
.B2(n_1533),
.Y(n_1640)
);

BUFx3_ASAP7_75t_L g1641 ( 
.A(n_1595),
.Y(n_1641)
);

INVxp67_ASAP7_75t_L g1642 ( 
.A(n_1532),
.Y(n_1642)
);

OR2x6_ASAP7_75t_L g1643 ( 
.A(n_1538),
.B(n_1549),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1572),
.B(n_1591),
.Y(n_1644)
);

NAND3xp33_ASAP7_75t_L g1645 ( 
.A(n_1585),
.B(n_1559),
.C(n_1588),
.Y(n_1645)
);

NOR2xp33_ASAP7_75t_L g1646 ( 
.A(n_1596),
.B(n_1594),
.Y(n_1646)
);

O2A1O1Ixp33_ASAP7_75t_SL g1647 ( 
.A1(n_1592),
.A2(n_1593),
.B(n_1594),
.C(n_1585),
.Y(n_1647)
);

AO21x1_ASAP7_75t_L g1648 ( 
.A1(n_1529),
.A2(n_1535),
.B(n_1534),
.Y(n_1648)
);

BUFx3_ASAP7_75t_L g1649 ( 
.A(n_1595),
.Y(n_1649)
);

HB1xp67_ASAP7_75t_L g1650 ( 
.A(n_1524),
.Y(n_1650)
);

INVxp33_ASAP7_75t_L g1651 ( 
.A(n_1587),
.Y(n_1651)
);

OAI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1559),
.A2(n_1580),
.B(n_1547),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1614),
.B(n_1515),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1614),
.B(n_1515),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1648),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1615),
.B(n_1533),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1636),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1627),
.B(n_1533),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1623),
.B(n_1533),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1630),
.B(n_1515),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1630),
.B(n_1515),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1635),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1639),
.B(n_1589),
.Y(n_1663)
);

AOI22xp33_ASAP7_75t_L g1664 ( 
.A1(n_1625),
.A2(n_1547),
.B1(n_1564),
.B2(n_1580),
.Y(n_1664)
);

INVxp67_ASAP7_75t_SL g1665 ( 
.A(n_1642),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1623),
.B(n_1533),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1628),
.B(n_1554),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1605),
.B(n_1522),
.Y(n_1668)
);

OAI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1634),
.A2(n_1580),
.B1(n_1539),
.B2(n_1537),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1612),
.B(n_1522),
.Y(n_1670)
);

INVx2_ASAP7_75t_SL g1671 ( 
.A(n_1643),
.Y(n_1671)
);

NOR2x1_ASAP7_75t_L g1672 ( 
.A(n_1645),
.B(n_1554),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1624),
.Y(n_1673)
);

INVx2_ASAP7_75t_SL g1674 ( 
.A(n_1643),
.Y(n_1674)
);

INVx4_ASAP7_75t_L g1675 ( 
.A(n_1641),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1628),
.B(n_1508),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1624),
.Y(n_1677)
);

NAND4xp25_ASAP7_75t_L g1678 ( 
.A(n_1604),
.B(n_1544),
.C(n_1542),
.D(n_1537),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1640),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1640),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1640),
.Y(n_1681)
);

INVx1_ASAP7_75t_SL g1682 ( 
.A(n_1644),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1650),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1650),
.Y(n_1684)
);

INVxp67_ASAP7_75t_L g1685 ( 
.A(n_1621),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1620),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1622),
.B(n_1545),
.Y(n_1687)
);

INVxp67_ASAP7_75t_SL g1688 ( 
.A(n_1638),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1663),
.B(n_1616),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1673),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1682),
.B(n_1620),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1682),
.B(n_1620),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1657),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1660),
.B(n_1643),
.Y(n_1694)
);

INVx2_ASAP7_75t_SL g1695 ( 
.A(n_1683),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1687),
.B(n_1620),
.Y(n_1696)
);

INVx4_ASAP7_75t_L g1697 ( 
.A(n_1675),
.Y(n_1697)
);

OAI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1664),
.A2(n_1634),
.B1(n_1631),
.B2(n_1632),
.Y(n_1698)
);

BUFx2_ASAP7_75t_L g1699 ( 
.A(n_1665),
.Y(n_1699)
);

BUFx6f_ASAP7_75t_L g1700 ( 
.A(n_1673),
.Y(n_1700)
);

BUFx3_ASAP7_75t_L g1701 ( 
.A(n_1671),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1660),
.B(n_1661),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1659),
.B(n_1633),
.Y(n_1703)
);

HB1xp67_ASAP7_75t_L g1704 ( 
.A(n_1662),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1657),
.Y(n_1705)
);

AOI31xp67_ASAP7_75t_L g1706 ( 
.A1(n_1673),
.A2(n_1677),
.A3(n_1679),
.B(n_1683),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1667),
.B(n_1626),
.Y(n_1707)
);

INVxp67_ASAP7_75t_SL g1708 ( 
.A(n_1655),
.Y(n_1708)
);

OAI21xp5_ASAP7_75t_SL g1709 ( 
.A1(n_1678),
.A2(n_1604),
.B(n_1613),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1668),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1677),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1687),
.B(n_1602),
.Y(n_1712)
);

INVxp67_ASAP7_75t_L g1713 ( 
.A(n_1655),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1659),
.B(n_1626),
.Y(n_1714)
);

AND2x4_ASAP7_75t_L g1715 ( 
.A(n_1674),
.B(n_1597),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1666),
.B(n_1638),
.Y(n_1716)
);

AND2x2_ASAP7_75t_SL g1717 ( 
.A(n_1664),
.B(n_1658),
.Y(n_1717)
);

INVx1_ASAP7_75t_SL g1718 ( 
.A(n_1670),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1668),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1685),
.B(n_1606),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1670),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1679),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1679),
.Y(n_1723)
);

OR3x1_ASAP7_75t_L g1724 ( 
.A(n_1678),
.B(n_1646),
.C(n_1610),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1676),
.Y(n_1725)
);

AOI221xp5_ASAP7_75t_L g1726 ( 
.A1(n_1669),
.A2(n_1617),
.B1(n_1637),
.B2(n_1629),
.C(n_1618),
.Y(n_1726)
);

OAI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1672),
.A2(n_1637),
.B1(n_1618),
.B2(n_1617),
.Y(n_1727)
);

INVx3_ASAP7_75t_L g1728 ( 
.A(n_1700),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1722),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1722),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1722),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1696),
.B(n_1686),
.Y(n_1732)
);

INVx4_ASAP7_75t_L g1733 ( 
.A(n_1697),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1723),
.Y(n_1734)
);

INVx1_ASAP7_75t_SL g1735 ( 
.A(n_1724),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1696),
.B(n_1686),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1723),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1696),
.B(n_1653),
.Y(n_1738)
);

NOR2xp67_ASAP7_75t_L g1739 ( 
.A(n_1713),
.B(n_1680),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1691),
.B(n_1685),
.Y(n_1740)
);

INVxp67_ASAP7_75t_SL g1741 ( 
.A(n_1708),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1715),
.B(n_1688),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1706),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1706),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1693),
.Y(n_1745)
);

BUFx2_ASAP7_75t_L g1746 ( 
.A(n_1699),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1691),
.B(n_1692),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1714),
.B(n_1680),
.Y(n_1748)
);

HB1xp67_ASAP7_75t_L g1749 ( 
.A(n_1704),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1693),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1705),
.Y(n_1751)
);

INVx3_ASAP7_75t_L g1752 ( 
.A(n_1700),
.Y(n_1752)
);

CKINVDCx20_ASAP7_75t_R g1753 ( 
.A(n_1689),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1714),
.B(n_1681),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1691),
.B(n_1665),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1700),
.Y(n_1756)
);

HB1xp67_ASAP7_75t_L g1757 ( 
.A(n_1704),
.Y(n_1757)
);

NOR2x1p5_ASAP7_75t_L g1758 ( 
.A(n_1697),
.B(n_1649),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1692),
.B(n_1712),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1700),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1725),
.B(n_1681),
.Y(n_1761)
);

HB1xp67_ASAP7_75t_L g1762 ( 
.A(n_1699),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1700),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1692),
.B(n_1684),
.Y(n_1764)
);

NOR2xp33_ASAP7_75t_R g1765 ( 
.A(n_1720),
.B(n_1613),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1700),
.Y(n_1766)
);

AND2x4_ASAP7_75t_L g1767 ( 
.A(n_1715),
.B(n_1688),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1695),
.B(n_1654),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1735),
.B(n_1694),
.Y(n_1769)
);

AOI221xp5_ASAP7_75t_SL g1770 ( 
.A1(n_1735),
.A2(n_1713),
.B1(n_1724),
.B2(n_1727),
.C(n_1698),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1745),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1740),
.B(n_1759),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1740),
.B(n_1759),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1748),
.B(n_1725),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1743),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1745),
.Y(n_1776)
);

INVx2_ASAP7_75t_SL g1777 ( 
.A(n_1758),
.Y(n_1777)
);

OR2x2_ASAP7_75t_L g1778 ( 
.A(n_1748),
.B(n_1707),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1740),
.B(n_1694),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1745),
.Y(n_1780)
);

INVx1_ASAP7_75t_SL g1781 ( 
.A(n_1753),
.Y(n_1781)
);

AND2x4_ASAP7_75t_L g1782 ( 
.A(n_1758),
.B(n_1708),
.Y(n_1782)
);

NAND2x1p5_ASAP7_75t_L g1783 ( 
.A(n_1758),
.B(n_1672),
.Y(n_1783)
);

OAI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1741),
.A2(n_1709),
.B(n_1727),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1741),
.B(n_1718),
.Y(n_1785)
);

OAI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1739),
.A2(n_1709),
.B(n_1717),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1759),
.B(n_1702),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1762),
.B(n_1718),
.Y(n_1788)
);

AOI21xp33_ASAP7_75t_L g1789 ( 
.A1(n_1743),
.A2(n_1698),
.B(n_1717),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1743),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1750),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1762),
.B(n_1724),
.Y(n_1792)
);

HB1xp67_ASAP7_75t_L g1793 ( 
.A(n_1739),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1746),
.B(n_1710),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1750),
.Y(n_1795)
);

NOR2x1p5_ASAP7_75t_L g1796 ( 
.A(n_1748),
.B(n_1599),
.Y(n_1796)
);

OR2x2_ASAP7_75t_L g1797 ( 
.A(n_1754),
.B(n_1707),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1750),
.Y(n_1798)
);

AO22x1_ASAP7_75t_L g1799 ( 
.A1(n_1743),
.A2(n_1651),
.B1(n_1608),
.B2(n_1599),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1746),
.B(n_1710),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1746),
.B(n_1719),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1755),
.B(n_1719),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1739),
.Y(n_1803)
);

INVxp67_ASAP7_75t_L g1804 ( 
.A(n_1749),
.Y(n_1804)
);

AOI222xp33_ASAP7_75t_L g1805 ( 
.A1(n_1747),
.A2(n_1726),
.B1(n_1717),
.B2(n_1669),
.C1(n_1629),
.C2(n_1716),
.Y(n_1805)
);

OR2x2_ASAP7_75t_L g1806 ( 
.A(n_1754),
.B(n_1721),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1755),
.B(n_1721),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1751),
.Y(n_1808)
);

NAND2x1p5_ASAP7_75t_L g1809 ( 
.A(n_1733),
.B(n_1697),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1755),
.B(n_1656),
.Y(n_1810)
);

BUFx2_ASAP7_75t_L g1811 ( 
.A(n_1733),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1751),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1754),
.B(n_1656),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1744),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1759),
.B(n_1702),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1772),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1771),
.Y(n_1817)
);

INVxp67_ASAP7_75t_L g1818 ( 
.A(n_1781),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1784),
.B(n_1747),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1772),
.Y(n_1820)
);

AND2x4_ASAP7_75t_L g1821 ( 
.A(n_1769),
.B(n_1733),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1771),
.Y(n_1822)
);

NAND2x1_ASAP7_75t_L g1823 ( 
.A(n_1782),
.B(n_1773),
.Y(n_1823)
);

INVx1_ASAP7_75t_SL g1824 ( 
.A(n_1769),
.Y(n_1824)
);

OAI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1786),
.A2(n_1726),
.B1(n_1744),
.B2(n_1703),
.Y(n_1825)
);

INVx2_ASAP7_75t_SL g1826 ( 
.A(n_1782),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1805),
.B(n_1747),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1778),
.B(n_1761),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1776),
.Y(n_1829)
);

INVxp67_ASAP7_75t_SL g1830 ( 
.A(n_1775),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1778),
.B(n_1747),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1770),
.B(n_1738),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1773),
.B(n_1732),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1776),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1779),
.B(n_1732),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1798),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1796),
.B(n_1738),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1797),
.B(n_1732),
.Y(n_1838)
);

OR2x2_ASAP7_75t_L g1839 ( 
.A(n_1797),
.B(n_1732),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1774),
.B(n_1736),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1774),
.B(n_1736),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1798),
.Y(n_1842)
);

AOI22xp5_ASAP7_75t_L g1843 ( 
.A1(n_1789),
.A2(n_1744),
.B1(n_1736),
.B2(n_1716),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1804),
.B(n_1738),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1787),
.B(n_1736),
.Y(n_1845)
);

NAND2x1p5_ASAP7_75t_L g1846 ( 
.A(n_1782),
.B(n_1733),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1787),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1779),
.B(n_1733),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1815),
.Y(n_1849)
);

OR2x2_ASAP7_75t_L g1850 ( 
.A(n_1806),
.B(n_1802),
.Y(n_1850)
);

AOI22xp33_ASAP7_75t_L g1851 ( 
.A1(n_1775),
.A2(n_1744),
.B1(n_1652),
.B2(n_1580),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1806),
.B(n_1761),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1830),
.Y(n_1853)
);

HB1xp67_ASAP7_75t_L g1854 ( 
.A(n_1818),
.Y(n_1854)
);

AOI21xp5_ASAP7_75t_L g1855 ( 
.A1(n_1825),
.A2(n_1799),
.B(n_1792),
.Y(n_1855)
);

AND2x2_ASAP7_75t_SL g1856 ( 
.A(n_1827),
.B(n_1811),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1824),
.B(n_1815),
.Y(n_1857)
);

NOR3xp33_ASAP7_75t_L g1858 ( 
.A(n_1825),
.B(n_1799),
.C(n_1790),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1817),
.Y(n_1859)
);

AOI221x1_ASAP7_75t_SL g1860 ( 
.A1(n_1819),
.A2(n_1814),
.B1(n_1790),
.B2(n_1785),
.C(n_1788),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1822),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1829),
.Y(n_1862)
);

AOI21xp5_ASAP7_75t_L g1863 ( 
.A1(n_1832),
.A2(n_1803),
.B(n_1793),
.Y(n_1863)
);

OAI21xp33_ASAP7_75t_L g1864 ( 
.A1(n_1843),
.A2(n_1800),
.B(n_1794),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1834),
.Y(n_1865)
);

OAI221xp5_ASAP7_75t_SL g1866 ( 
.A1(n_1831),
.A2(n_1814),
.B1(n_1813),
.B2(n_1810),
.C(n_1598),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1836),
.Y(n_1867)
);

NAND3xp33_ASAP7_75t_L g1868 ( 
.A(n_1851),
.B(n_1811),
.C(n_1733),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1835),
.B(n_1777),
.Y(n_1869)
);

AOI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1823),
.A2(n_1777),
.B(n_1753),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1842),
.Y(n_1871)
);

OAI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1838),
.A2(n_1783),
.B1(n_1767),
.B2(n_1742),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1816),
.B(n_1801),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1830),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1816),
.B(n_1807),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1820),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1820),
.B(n_1749),
.Y(n_1877)
);

OAI22xp5_ASAP7_75t_L g1878 ( 
.A1(n_1839),
.A2(n_1783),
.B1(n_1742),
.B2(n_1767),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1847),
.Y(n_1879)
);

AOI221xp5_ASAP7_75t_L g1880 ( 
.A1(n_1860),
.A2(n_1851),
.B1(n_1828),
.B2(n_1844),
.C(n_1826),
.Y(n_1880)
);

A2O1A1Ixp33_ASAP7_75t_L g1881 ( 
.A1(n_1855),
.A2(n_1828),
.B(n_1841),
.C(n_1840),
.Y(n_1881)
);

NOR2xp33_ASAP7_75t_L g1882 ( 
.A(n_1854),
.B(n_1856),
.Y(n_1882)
);

INVx1_ASAP7_75t_SL g1883 ( 
.A(n_1854),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1853),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1853),
.Y(n_1885)
);

AOI221xp5_ASAP7_75t_L g1886 ( 
.A1(n_1858),
.A2(n_1826),
.B1(n_1835),
.B2(n_1852),
.C(n_1833),
.Y(n_1886)
);

OAI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1856),
.A2(n_1845),
.B1(n_1849),
.B2(n_1847),
.Y(n_1887)
);

AOI21xp5_ASAP7_75t_L g1888 ( 
.A1(n_1863),
.A2(n_1821),
.B(n_1848),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1869),
.B(n_1821),
.Y(n_1889)
);

AOI221xp5_ASAP7_75t_L g1890 ( 
.A1(n_1866),
.A2(n_1833),
.B1(n_1837),
.B2(n_1849),
.C(n_1850),
.Y(n_1890)
);

OAI22xp5_ASAP7_75t_L g1891 ( 
.A1(n_1868),
.A2(n_1821),
.B1(n_1846),
.B2(n_1783),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1869),
.Y(n_1892)
);

AOI22xp5_ASAP7_75t_L g1893 ( 
.A1(n_1874),
.A2(n_1864),
.B1(n_1879),
.B2(n_1857),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1879),
.Y(n_1894)
);

AOI22xp5_ASAP7_75t_L g1895 ( 
.A1(n_1872),
.A2(n_1767),
.B1(n_1742),
.B2(n_1848),
.Y(n_1895)
);

NOR3xp33_ASAP7_75t_L g1896 ( 
.A(n_1870),
.B(n_1608),
.C(n_1609),
.Y(n_1896)
);

OAI221xp5_ASAP7_75t_L g1897 ( 
.A1(n_1878),
.A2(n_1875),
.B1(n_1876),
.B2(n_1873),
.C(n_1846),
.Y(n_1897)
);

AOI32xp33_ASAP7_75t_L g1898 ( 
.A1(n_1876),
.A2(n_1742),
.A3(n_1767),
.B1(n_1764),
.B2(n_1728),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1877),
.B(n_1757),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1859),
.Y(n_1900)
);

AOI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1861),
.A2(n_1742),
.B1(n_1767),
.B2(n_1734),
.Y(n_1901)
);

INVx1_ASAP7_75t_SL g1902 ( 
.A(n_1883),
.Y(n_1902)
);

INVx1_ASAP7_75t_SL g1903 ( 
.A(n_1883),
.Y(n_1903)
);

OAI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1881),
.A2(n_1767),
.B1(n_1742),
.B2(n_1809),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_SL g1905 ( 
.A(n_1882),
.B(n_1765),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1894),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1892),
.B(n_1862),
.Y(n_1907)
);

NOR2x1_ASAP7_75t_L g1908 ( 
.A(n_1884),
.B(n_1865),
.Y(n_1908)
);

XNOR2x1_ASAP7_75t_L g1909 ( 
.A(n_1893),
.B(n_1609),
.Y(n_1909)
);

INVx1_ASAP7_75t_SL g1910 ( 
.A(n_1889),
.Y(n_1910)
);

INVx1_ASAP7_75t_SL g1911 ( 
.A(n_1899),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1885),
.Y(n_1912)
);

OAI22xp5_ASAP7_75t_SL g1913 ( 
.A1(n_1887),
.A2(n_1871),
.B1(n_1867),
.B2(n_1809),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_SL g1914 ( 
.A(n_1886),
.B(n_1809),
.Y(n_1914)
);

AOI31xp33_ASAP7_75t_L g1915 ( 
.A1(n_1902),
.A2(n_1900),
.A3(n_1880),
.B(n_1888),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1903),
.B(n_1890),
.Y(n_1916)
);

OAI22xp33_ASAP7_75t_L g1917 ( 
.A1(n_1911),
.A2(n_1895),
.B1(n_1901),
.B2(n_1897),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1908),
.Y(n_1918)
);

O2A1O1Ixp33_ASAP7_75t_L g1919 ( 
.A1(n_1905),
.A2(n_1891),
.B(n_1896),
.C(n_1812),
.Y(n_1919)
);

NAND3xp33_ASAP7_75t_SL g1920 ( 
.A(n_1910),
.B(n_1898),
.C(n_1765),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1914),
.B(n_1768),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1907),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1906),
.B(n_1757),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1909),
.Y(n_1924)
);

AND4x1_ASAP7_75t_L g1925 ( 
.A(n_1912),
.B(n_1913),
.C(n_1610),
.D(n_1914),
.Y(n_1925)
);

AOI31xp33_ASAP7_75t_L g1926 ( 
.A1(n_1916),
.A2(n_1904),
.A3(n_1611),
.B(n_1607),
.Y(n_1926)
);

AND4x2_ASAP7_75t_L g1927 ( 
.A(n_1915),
.B(n_1610),
.C(n_1808),
.D(n_1812),
.Y(n_1927)
);

OAI221xp5_ASAP7_75t_SL g1928 ( 
.A1(n_1925),
.A2(n_1763),
.B1(n_1756),
.B2(n_1760),
.C(n_1766),
.Y(n_1928)
);

A2O1A1Ixp33_ASAP7_75t_L g1929 ( 
.A1(n_1915),
.A2(n_1763),
.B(n_1756),
.C(n_1760),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1918),
.B(n_1780),
.Y(n_1930)
);

AOI222xp33_ASAP7_75t_L g1931 ( 
.A1(n_1924),
.A2(n_1729),
.B1(n_1730),
.B2(n_1731),
.C1(n_1734),
.C2(n_1737),
.Y(n_1931)
);

OAI211xp5_ASAP7_75t_L g1932 ( 
.A1(n_1929),
.A2(n_1922),
.B(n_1923),
.C(n_1919),
.Y(n_1932)
);

AOI221xp5_ASAP7_75t_L g1933 ( 
.A1(n_1928),
.A2(n_1917),
.B1(n_1920),
.B2(n_1921),
.C(n_1808),
.Y(n_1933)
);

AOI222xp33_ASAP7_75t_L g1934 ( 
.A1(n_1927),
.A2(n_1730),
.B1(n_1729),
.B2(n_1731),
.C1(n_1734),
.C2(n_1737),
.Y(n_1934)
);

A2O1A1Ixp33_ASAP7_75t_L g1935 ( 
.A1(n_1926),
.A2(n_1756),
.B(n_1766),
.C(n_1760),
.Y(n_1935)
);

OAI211xp5_ASAP7_75t_L g1936 ( 
.A1(n_1930),
.A2(n_1752),
.B(n_1728),
.C(n_1795),
.Y(n_1936)
);

AOI221xp5_ASAP7_75t_L g1937 ( 
.A1(n_1931),
.A2(n_1791),
.B1(n_1756),
.B2(n_1760),
.C(n_1763),
.Y(n_1937)
);

AOI221xp5_ASAP7_75t_L g1938 ( 
.A1(n_1928),
.A2(n_1763),
.B1(n_1766),
.B2(n_1711),
.C(n_1690),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1932),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1934),
.Y(n_1940)
);

NAND4xp75_ASAP7_75t_L g1941 ( 
.A(n_1933),
.B(n_1610),
.C(n_1611),
.D(n_1766),
.Y(n_1941)
);

OAI211xp5_ASAP7_75t_L g1942 ( 
.A1(n_1936),
.A2(n_1728),
.B(n_1752),
.C(n_1697),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1935),
.B(n_1751),
.Y(n_1943)
);

NOR2xp67_ASAP7_75t_L g1944 ( 
.A(n_1937),
.B(n_1728),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1939),
.B(n_1938),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1940),
.B(n_1728),
.Y(n_1946)
);

HB1xp67_ASAP7_75t_L g1947 ( 
.A(n_1941),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1946),
.Y(n_1948)
);

AOI22xp33_ASAP7_75t_SL g1949 ( 
.A1(n_1948),
.A2(n_1947),
.B1(n_1945),
.B2(n_1943),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1949),
.Y(n_1950)
);

XOR2x2_ASAP7_75t_L g1951 ( 
.A(n_1949),
.B(n_1944),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1950),
.Y(n_1952)
);

INVx1_ASAP7_75t_SL g1953 ( 
.A(n_1951),
.Y(n_1953)
);

NOR2xp33_ASAP7_75t_L g1954 ( 
.A(n_1952),
.B(n_1942),
.Y(n_1954)
);

OAI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1953),
.A2(n_1752),
.B1(n_1728),
.B2(n_1764),
.Y(n_1955)
);

OAI21x1_ASAP7_75t_L g1956 ( 
.A1(n_1954),
.A2(n_1752),
.B(n_1601),
.Y(n_1956)
);

AND3x4_ASAP7_75t_L g1957 ( 
.A(n_1955),
.B(n_1701),
.C(n_1590),
.Y(n_1957)
);

NOR2xp33_ASAP7_75t_L g1958 ( 
.A(n_1957),
.B(n_1729),
.Y(n_1958)
);

XNOR2xp5_ASAP7_75t_L g1959 ( 
.A(n_1958),
.B(n_1956),
.Y(n_1959)
);

OAI221xp5_ASAP7_75t_R g1960 ( 
.A1(n_1959),
.A2(n_1752),
.B1(n_1647),
.B2(n_1764),
.C(n_1600),
.Y(n_1960)
);

AOI211xp5_ASAP7_75t_L g1961 ( 
.A1(n_1960),
.A2(n_1603),
.B(n_1619),
.C(n_1752),
.Y(n_1961)
);


endmodule