module fake_ariane_298_n_5534 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_646, n_197, n_640, n_463, n_176, n_691, n_34, n_404, n_172, n_678, n_651, n_347, n_423, n_183, n_469, n_479, n_603, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_610, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_20, n_690, n_416, n_283, n_50, n_187, n_525, n_367, n_649, n_598, n_345, n_374, n_318, n_103, n_244, n_643, n_679, n_226, n_220, n_261, n_682, n_36, n_663, n_370, n_189, n_72, n_286, n_443, n_586, n_57, n_686, n_605, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_607, n_670, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_631, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_665, n_59, n_336, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_668, n_339, n_672, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_648, n_269, n_597, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_645, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_600, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_677, n_222, n_478, n_510, n_256, n_326, n_681, n_227, n_48, n_188, n_323, n_550, n_635, n_330, n_400, n_689, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_644, n_293, n_620, n_228, n_325, n_276, n_93, n_688, n_636, n_427, n_108, n_587, n_497, n_303, n_671, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_611, n_238, n_365, n_429, n_455, n_654, n_588, n_638, n_136, n_334, n_192, n_661, n_488, n_667, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_684, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_579, n_459, n_685, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_616, n_617, n_658, n_630, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_601, n_683, n_565, n_281, n_24, n_7, n_628, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_660, n_464, n_575, n_546, n_297, n_662, n_641, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_639, n_217, n_452, n_673, n_676, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_680, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_148, n_652, n_451, n_613, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_674, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_656, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_629, n_664, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_655, n_99, n_540, n_216, n_544, n_5, n_599, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_657, n_513, n_288, n_179, n_395, n_621, n_195, n_606, n_213, n_110, n_304, n_659, n_67, n_509, n_583, n_306, n_666, n_313, n_92, n_430, n_626, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_669, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_615, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_425, n_431, n_508, n_624, n_118, n_121, n_618, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_687, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_642, n_97, n_408, n_595, n_322, n_251, n_506, n_602, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_653, n_359, n_155, n_573, n_127, n_531, n_675, n_5534);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_646;
input n_197;
input n_640;
input n_463;
input n_176;
input n_691;
input n_34;
input n_404;
input n_172;
input n_678;
input n_651;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_603;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_20;
input n_690;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_643;
input n_679;
input n_226;
input n_220;
input n_261;
input n_682;
input n_36;
input n_663;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_686;
input n_605;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_670;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_665;
input n_59;
input n_336;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_668;
input n_339;
input n_672;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_648;
input n_269;
input n_597;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_645;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_600;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_677;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_681;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_635;
input n_330;
input n_400;
input n_689;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_644;
input n_293;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_688;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_303;
input n_671;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_654;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_661;
input n_488;
input n_667;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_684;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_685;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_616;
input n_617;
input n_658;
input n_630;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_601;
input n_683;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_660;
input n_464;
input n_575;
input n_546;
input n_297;
input n_662;
input n_641;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_639;
input n_217;
input n_452;
input n_673;
input n_676;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_680;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_652;
input n_451;
input n_613;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_674;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_656;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_629;
input n_664;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_655;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_599;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_657;
input n_513;
input n_288;
input n_179;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_659;
input n_67;
input n_509;
input n_583;
input n_306;
input n_666;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_669;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_615;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_425;
input n_431;
input n_508;
input n_624;
input n_118;
input n_121;
input n_618;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_687;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_653;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;
input n_675;

output n_5534;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_4030;
wire n_4770;
wire n_5093;
wire n_3152;
wire n_4586;
wire n_3056;
wire n_3500;
wire n_2679;
wire n_5402;
wire n_2182;
wire n_2680;
wire n_3264;
wire n_1250;
wire n_2993;
wire n_4283;
wire n_2879;
wire n_4403;
wire n_4962;
wire n_1430;
wire n_2002;
wire n_1238;
wire n_2729;
wire n_4302;
wire n_4547;
wire n_5090;
wire n_3765;
wire n_864;
wire n_5302;
wire n_1096;
wire n_1379;
wire n_2376;
wire n_2790;
wire n_2207;
wire n_3954;
wire n_4982;
wire n_2042;
wire n_1131;
wire n_5479;
wire n_2646;
wire n_737;
wire n_2653;
wire n_4610;
wire n_3115;
wire n_4028;
wire n_5263;
wire n_2482;
wire n_1682;
wire n_958;
wire n_2554;
wire n_4321;
wire n_1985;
wire n_2621;
wire n_4853;
wire n_1909;
wire n_5229;
wire n_4260;
wire n_903;
wire n_3348;
wire n_3261;
wire n_1761;
wire n_1690;
wire n_2807;
wire n_1018;
wire n_4512;
wire n_4132;
wire n_1364;
wire n_2390;
wire n_4500;
wire n_2322;
wire n_1107;
wire n_2663;
wire n_5481;
wire n_4824;
wire n_5340;
wire n_3545;
wire n_1428;
wire n_1284;
wire n_4741;
wire n_1241;
wire n_4143;
wire n_4273;
wire n_901;
wire n_4136;
wire n_3144;
wire n_2359;
wire n_1519;
wire n_4567;
wire n_786;
wire n_3552;
wire n_2950;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_2301;
wire n_3121;
wire n_2847;
wire n_3015;
wire n_3870;
wire n_3749;
wire n_1676;
wire n_1085;
wire n_3482;
wire n_5403;
wire n_823;
wire n_1900;
wire n_4268;
wire n_863;
wire n_3960;
wire n_2433;
wire n_3975;
wire n_899;
wire n_2004;
wire n_4018;
wire n_1495;
wire n_3325;
wire n_4227;
wire n_5158;
wire n_5152;
wire n_1917;
wire n_2456;
wire n_5092;
wire n_1924;
wire n_1811;
wire n_3612;
wire n_4505;
wire n_1840;
wire n_5247;
wire n_5464;
wire n_4476;
wire n_844;
wire n_1267;
wire n_2956;
wire n_5210;
wire n_1213;
wire n_2382;
wire n_780;
wire n_5292;
wire n_1918;
wire n_4119;
wire n_4443;
wire n_4000;
wire n_2686;
wire n_5086;
wire n_1949;
wire n_1140;
wire n_3458;
wire n_3511;
wire n_2077;
wire n_1121;
wire n_3012;
wire n_1947;
wire n_4529;
wire n_3850;
wire n_1216;
wire n_4908;
wire n_3754;
wire n_5060;
wire n_4432;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2116;
wire n_4530;
wire n_1432;
wire n_2245;
wire n_5391;
wire n_5452;
wire n_3359;
wire n_3841;
wire n_5249;
wire n_851;
wire n_3900;
wire n_3413;
wire n_5076;
wire n_3539;
wire n_5062;
wire n_2134;
wire n_3862;
wire n_930;
wire n_4912;
wire n_4226;
wire n_4311;
wire n_3284;
wire n_5046;
wire n_1386;
wire n_3506;
wire n_4827;
wire n_1842;
wire n_4993;
wire n_3678;
wire n_2791;
wire n_1661;
wire n_3212;
wire n_4871;
wire n_3529;
wire n_4405;
wire n_966;
wire n_992;
wire n_3549;
wire n_3914;
wire n_1692;
wire n_2611;
wire n_5468;
wire n_3029;
wire n_4745;
wire n_2398;
wire n_4233;
wire n_4791;
wire n_5056;
wire n_1178;
wire n_2015;
wire n_5204;
wire n_2877;
wire n_4951;
wire n_4959;
wire n_3000;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_2161;
wire n_746;
wire n_1357;
wire n_1787;
wire n_1389;
wire n_3172;
wire n_2659;
wire n_4033;
wire n_3747;
wire n_4905;
wire n_4508;
wire n_4045;
wire n_4894;
wire n_3651;
wire n_1812;
wire n_3614;
wire n_959;
wire n_2257;
wire n_1101;
wire n_1343;
wire n_3116;
wire n_4141;
wire n_3784;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_1623;
wire n_3559;
wire n_5179;
wire n_2435;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_1087;
wire n_2388;
wire n_2273;
wire n_1911;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_3700;
wire n_4307;
wire n_2795;
wire n_1841;
wire n_1680;
wire n_2954;
wire n_4438;
wire n_974;
wire n_3814;
wire n_4367;
wire n_5134;
wire n_2467;
wire n_4195;
wire n_5091;
wire n_4866;
wire n_1447;
wire n_1220;
wire n_2019;
wire n_698;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_5454;
wire n_1209;
wire n_4254;
wire n_3438;
wire n_2625;
wire n_5373;
wire n_1578;
wire n_3147;
wire n_3661;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_1568;
wire n_2919;
wire n_3108;
wire n_2632;
wire n_4314;
wire n_2980;
wire n_1728;
wire n_4315;
wire n_3239;
wire n_2631;
wire n_3311;
wire n_3516;
wire n_4442;
wire n_4857;
wire n_1651;
wire n_3087;
wire n_4637;
wire n_5523;
wire n_2697;
wire n_1263;
wire n_1817;
wire n_3704;
wire n_4296;
wire n_2677;
wire n_2483;
wire n_5088;
wire n_1032;
wire n_1592;
wire n_5392;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_3589;
wire n_1743;
wire n_720;
wire n_1943;
wire n_5138;
wire n_4588;
wire n_5149;
wire n_1163;
wire n_3054;
wire n_4970;
wire n_5280;
wire n_4153;
wire n_1868;
wire n_5052;
wire n_3601;
wire n_5137;
wire n_2373;
wire n_3881;
wire n_5089;
wire n_2099;
wire n_3759;
wire n_3323;
wire n_4643;
wire n_2617;
wire n_808;
wire n_2476;
wire n_2814;
wire n_4133;
wire n_2636;
wire n_1439;
wire n_3466;
wire n_2074;
wire n_5031;
wire n_1665;
wire n_2122;
wire n_4543;
wire n_4337;
wire n_5082;
wire n_4788;
wire n_1414;
wire n_2067;
wire n_4555;
wire n_5230;
wire n_1901;
wire n_4486;
wire n_3465;
wire n_2117;
wire n_1053;
wire n_5296;
wire n_5398;
wire n_1906;
wire n_2194;
wire n_4780;
wire n_4640;
wire n_1828;
wire n_1304;
wire n_3335;
wire n_3007;
wire n_2267;
wire n_1349;
wire n_1061;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_3370;
wire n_874;
wire n_3949;
wire n_2286;
wire n_5192;
wire n_4247;
wire n_707;
wire n_5051;
wire n_5336;
wire n_3036;
wire n_2783;
wire n_4583;
wire n_1015;
wire n_1162;
wire n_4292;
wire n_2118;
wire n_1490;
wire n_3764;
wire n_1553;
wire n_4773;
wire n_1760;
wire n_5028;
wire n_1086;
wire n_3025;
wire n_3051;
wire n_986;
wire n_1104;
wire n_2802;
wire n_887;
wire n_2125;
wire n_1156;
wire n_4974;
wire n_5123;
wire n_2861;
wire n_4344;
wire n_5242;
wire n_3130;
wire n_1188;
wire n_1498;
wire n_4856;
wire n_2618;
wire n_4216;
wire n_957;
wire n_1242;
wire n_2707;
wire n_2849;
wire n_1489;
wire n_2756;
wire n_3781;
wire n_2217;
wire n_4864;
wire n_2226;
wire n_5127;
wire n_4313;
wire n_5255;
wire n_4460;
wire n_4670;
wire n_1119;
wire n_3713;
wire n_1863;
wire n_4798;
wire n_1500;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_4229;
wire n_5071;
wire n_3337;
wire n_1189;
wire n_3750;
wire n_3424;
wire n_3356;
wire n_1523;
wire n_2190;
wire n_3931;
wire n_2516;
wire n_4991;
wire n_3070;
wire n_1005;
wire n_3275;
wire n_5198;
wire n_3245;
wire n_2894;
wire n_2452;
wire n_4182;
wire n_2827;
wire n_3214;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_5009;
wire n_3710;
wire n_1844;
wire n_1957;
wire n_1953;
wire n_1219;
wire n_710;
wire n_3944;
wire n_4729;
wire n_1793;
wire n_4446;
wire n_4662;
wire n_4800;
wire n_1373;
wire n_1540;
wire n_5427;
wire n_4440;
wire n_1797;
wire n_4425;
wire n_5450;
wire n_832;
wire n_744;
wire n_2821;
wire n_3696;
wire n_1331;
wire n_4781;
wire n_1529;
wire n_3531;
wire n_5124;
wire n_4237;
wire n_5297;
wire n_4828;
wire n_3333;
wire n_4652;
wire n_4114;
wire n_1007;
wire n_1580;
wire n_3135;
wire n_4925;
wire n_2448;
wire n_2211;
wire n_951;
wire n_5318;
wire n_5374;
wire n_2424;
wire n_4697;
wire n_4765;
wire n_5108;
wire n_722;
wire n_3277;
wire n_4863;
wire n_1766;
wire n_5463;
wire n_1338;
wire n_2978;
wire n_4859;
wire n_4568;
wire n_3617;
wire n_704;
wire n_2958;
wire n_1044;
wire n_1714;
wire n_4429;
wire n_5435;
wire n_3340;
wire n_5053;
wire n_5476;
wire n_5483;
wire n_1243;
wire n_5511;
wire n_3486;
wire n_2457;
wire n_2992;
wire n_3197;
wire n_3256;
wire n_1878;
wire n_3646;
wire n_2520;
wire n_811;
wire n_791;
wire n_3864;
wire n_4694;
wire n_1025;
wire n_4664;
wire n_3450;
wire n_4633;
wire n_2026;
wire n_4050;
wire n_3173;
wire n_1406;
wire n_5073;
wire n_4306;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_3266;
wire n_3102;
wire n_1499;
wire n_4288;
wire n_3452;
wire n_4098;
wire n_2691;
wire n_4511;
wire n_3422;
wire n_4675;
wire n_695;
wire n_2991;
wire n_5419;
wire n_1596;
wire n_4289;
wire n_4972;
wire n_2723;
wire n_1476;
wire n_2016;
wire n_3925;
wire n_4689;
wire n_5165;
wire n_2850;
wire n_1874;
wire n_5077;
wire n_3780;
wire n_1657;
wire n_3753;
wire n_1488;
wire n_4846;
wire n_1330;
wire n_906;
wire n_2295;
wire n_5225;
wire n_4076;
wire n_3142;
wire n_3129;
wire n_3495;
wire n_3843;
wire n_4805;
wire n_2606;
wire n_2386;
wire n_4822;
wire n_1829;
wire n_4635;
wire n_1450;
wire n_5532;
wire n_3740;
wire n_5441;
wire n_2417;
wire n_1815;
wire n_1493;
wire n_2911;
wire n_3313;
wire n_2354;
wire n_4281;
wire n_3945;
wire n_3726;
wire n_4419;
wire n_5405;
wire n_1256;
wire n_5365;
wire n_3560;
wire n_3345;
wire n_3421;
wire n_1448;
wire n_1009;
wire n_3548;
wire n_4906;
wire n_4630;
wire n_4829;
wire n_2612;
wire n_5259;
wire n_3236;
wire n_1995;
wire n_1397;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_4966;
wire n_2250;
wire n_1117;
wire n_3321;
wire n_1303;
wire n_4188;
wire n_2001;
wire n_2506;
wire n_2413;
wire n_4825;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_2626;
wire n_2892;
wire n_2605;
wire n_2804;
wire n_5006;
wire n_4882;
wire n_3206;
wire n_1035;
wire n_3475;
wire n_4878;
wire n_2070;
wire n_3842;
wire n_1367;
wire n_4202;
wire n_2044;
wire n_3886;
wire n_825;
wire n_732;
wire n_2619;
wire n_1192;
wire n_5141;
wire n_3098;
wire n_4503;
wire n_1291;
wire n_5208;
wire n_5113;
wire n_3987;
wire n_5205;
wire n_4249;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_2711;
wire n_3223;
wire n_3386;
wire n_3921;
wire n_2177;
wire n_2766;
wire n_4196;
wire n_1197;
wire n_2613;
wire n_1517;
wire n_2647;
wire n_5508;
wire n_5105;
wire n_3920;
wire n_3444;
wire n_3851;
wire n_1671;
wire n_5027;
wire n_1048;
wire n_2343;
wire n_775;
wire n_3380;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2411;
wire n_4631;
wire n_1504;
wire n_2110;
wire n_5377;
wire n_3822;
wire n_889;
wire n_4355;
wire n_3818;
wire n_3587;
wire n_2608;
wire n_1948;
wire n_4155;
wire n_810;
wire n_4278;
wire n_4710;
wire n_1959;
wire n_3497;
wire n_4542;
wire n_5451;
wire n_3243;
wire n_4326;
wire n_2121;
wire n_3865;
wire n_5460;
wire n_4685;
wire n_3927;
wire n_2068;
wire n_3595;
wire n_1194;
wire n_4060;
wire n_1647;
wire n_1454;
wire n_2459;
wire n_941;
wire n_3396;
wire n_5517;
wire n_5426;
wire n_4093;
wire n_4123;
wire n_4294;
wire n_1521;
wire n_1940;
wire n_3683;
wire n_4452;
wire n_3887;
wire n_3195;
wire n_4722;
wire n_3048;
wire n_3339;
wire n_4164;
wire n_4126;
wire n_5030;
wire n_2963;
wire n_2561;
wire n_1056;
wire n_3168;
wire n_5320;
wire n_4079;
wire n_1749;
wire n_1653;
wire n_4088;
wire n_2669;
wire n_3911;
wire n_3802;
wire n_4366;
wire n_1584;
wire n_848;
wire n_5125;
wire n_4922;
wire n_4733;
wire n_1814;
wire n_2441;
wire n_4041;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_4935;
wire n_4509;
wire n_2073;
wire n_4004;
wire n_5238;
wire n_750;
wire n_834;
wire n_3630;
wire n_1612;
wire n_800;
wire n_1910;
wire n_2189;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_2602;
wire n_724;
wire n_2931;
wire n_3433;
wire n_3597;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_3786;
wire n_875;
wire n_2828;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_4204;
wire n_3553;
wire n_5323;
wire n_3645;
wire n_793;
wire n_4996;
wire n_1485;
wire n_2883;
wire n_4411;
wire n_4317;
wire n_3550;
wire n_5510;
wire n_4785;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_1805;
wire n_4068;
wire n_5440;
wire n_2270;
wire n_4163;
wire n_3294;
wire n_2443;
wire n_3610;
wire n_5011;
wire n_1554;
wire n_3279;
wire n_5513;
wire n_972;
wire n_4262;
wire n_2923;
wire n_2843;
wire n_3714;
wire n_4832;
wire n_3676;
wire n_2010;
wire n_5197;
wire n_1679;
wire n_3109;
wire n_1952;
wire n_2394;
wire n_3125;
wire n_5128;
wire n_2356;
wire n_4672;
wire n_2564;
wire n_3558;
wire n_3034;
wire n_3502;
wire n_783;
wire n_4053;
wire n_1127;
wire n_1008;
wire n_3963;
wire n_3091;
wire n_1024;
wire n_5157;
wire n_4496;
wire n_2518;
wire n_936;
wire n_4596;
wire n_5178;
wire n_3105;
wire n_1525;
wire n_4628;
wire n_1775;
wire n_908;
wire n_1036;
wire n_4083;
wire n_1270;
wire n_1272;
wire n_2794;
wire n_2901;
wire n_3940;
wire n_3225;
wire n_3621;
wire n_5529;
wire n_3473;
wire n_3680;
wire n_3565;
wire n_5388;
wire n_5354;
wire n_2453;
wire n_3331;
wire n_1788;
wire n_2138;
wire n_3040;
wire n_4230;
wire n_3360;
wire n_1930;
wire n_1809;
wire n_3585;
wire n_1843;
wire n_2000;
wire n_5276;
wire n_4037;
wire n_3804;
wire n_4659;
wire n_3211;
wire n_917;
wire n_5196;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2215;
wire n_3847;
wire n_4073;
wire n_1261;
wire n_3633;
wire n_857;
wire n_1235;
wire n_2584;
wire n_4001;
wire n_1462;
wire n_1064;
wire n_1446;
wire n_1701;
wire n_3111;
wire n_731;
wire n_1813;
wire n_2997;
wire n_1573;
wire n_3258;
wire n_758;
wire n_3691;
wire n_2252;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_4339;
wire n_4690;
wire n_2987;
wire n_1473;
wire n_1076;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2733;
wire n_2445;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_3316;
wire n_4023;
wire n_4253;
wire n_2522;
wire n_3632;
wire n_1344;
wire n_4064;
wire n_3351;
wire n_5478;
wire n_1141;
wire n_3457;
wire n_5384;
wire n_840;
wire n_2324;
wire n_5283;
wire n_3454;
wire n_2139;
wire n_2521;
wire n_2740;
wire n_1991;
wire n_4066;
wire n_4681;
wire n_3303;
wire n_4414;
wire n_2541;
wire n_5094;
wire n_3232;
wire n_1113;
wire n_3768;
wire n_4295;
wire n_1615;
wire n_4100;
wire n_1265;
wire n_2372;
wire n_2105;
wire n_3445;
wire n_1806;
wire n_4087;
wire n_1409;
wire n_1684;
wire n_1588;
wire n_1148;
wire n_1673;
wire n_4473;
wire n_4619;
wire n_5371;
wire n_2290;
wire n_4398;
wire n_5026;
wire n_2856;
wire n_3235;
wire n_5350;
wire n_3265;
wire n_3018;
wire n_1875;
wire n_2429;
wire n_5286;
wire n_4449;
wire n_3285;
wire n_4607;
wire n_1039;
wire n_5040;
wire n_1150;
wire n_4266;
wire n_1628;
wire n_2971;
wire n_4407;
wire n_4695;
wire n_1136;
wire n_1190;
wire n_3628;
wire n_4777;
wire n_5243;
wire n_3941;
wire n_1915;
wire n_5399;
wire n_2846;
wire n_3371;
wire n_4918;
wire n_3872;
wire n_4415;
wire n_5110;
wire n_1964;
wire n_3659;
wire n_3928;
wire n_1777;
wire n_3366;
wire n_3441;
wire n_3020;
wire n_4146;
wire n_4947;
wire n_708;
wire n_2545;
wire n_2513;
wire n_4408;
wire n_2115;
wire n_2017;
wire n_1810;
wire n_1347;
wire n_4976;
wire n_860;
wire n_3555;
wire n_3534;
wire n_4548;
wire n_2670;
wire n_3556;
wire n_896;
wire n_4574;
wire n_2644;
wire n_4557;
wire n_3071;
wire n_1698;
wire n_1337;
wire n_774;
wire n_2148;
wire n_1168;
wire n_4663;
wire n_3296;
wire n_3794;
wire n_3762;
wire n_4624;
wire n_4963;
wire n_5136;
wire n_4205;
wire n_3293;
wire n_4902;
wire n_1683;
wire n_4686;
wire n_2384;
wire n_1705;
wire n_768;
wire n_3707;
wire n_1091;
wire n_3895;
wire n_3149;
wire n_3934;
wire n_4338;
wire n_2058;
wire n_3231;
wire n_1846;
wire n_4161;
wire n_5304;
wire n_5437;
wire n_1581;
wire n_946;
wire n_757;
wire n_2047;
wire n_3058;
wire n_1655;
wire n_3398;
wire n_3709;
wire n_1146;
wire n_5355;
wire n_998;
wire n_3592;
wire n_5321;
wire n_2536;
wire n_1604;
wire n_3399;
wire n_4772;
wire n_1368;
wire n_963;
wire n_4120;
wire n_925;
wire n_2880;
wire n_1313;
wire n_3722;
wire n_1001;
wire n_4716;
wire n_1115;
wire n_4654;
wire n_1339;
wire n_1051;
wire n_5116;
wire n_3771;
wire n_719;
wire n_3158;
wire n_3221;
wire n_2316;
wire n_1010;
wire n_2830;
wire n_5500;
wire n_4622;
wire n_4757;
wire n_803;
wire n_1871;
wire n_4016;
wire n_3334;
wire n_2940;
wire n_3427;
wire n_3162;
wire n_4591;
wire n_5515;
wire n_3083;
wire n_4570;
wire n_2491;
wire n_1931;
wire n_2259;
wire n_5337;
wire n_849;
wire n_5059;
wire n_4655;
wire n_1820;
wire n_1233;
wire n_4493;
wire n_1808;
wire n_1635;
wire n_1704;
wire n_4896;
wire n_4851;
wire n_2479;
wire n_886;
wire n_1308;
wire n_1451;
wire n_1487;
wire n_5528;
wire n_3432;
wire n_2163;
wire n_1938;
wire n_2484;
wire n_5358;
wire n_1469;
wire n_4901;
wire n_3480;
wire n_1355;
wire n_4213;
wire n_4127;
wire n_2500;
wire n_2334;
wire n_5467;
wire n_1169;
wire n_789;
wire n_3181;
wire n_5493;
wire n_1916;
wire n_4602;
wire n_1713;
wire n_1436;
wire n_2818;
wire n_4900;
wire n_3578;
wire n_1109;
wire n_2537;
wire n_3745;
wire n_3487;
wire n_3668;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1566;
wire n_2837;
wire n_717;
wire n_952;
wire n_2446;
wire n_4116;
wire n_5360;
wire n_2671;
wire n_2702;
wire n_4363;
wire n_3561;
wire n_1839;
wire n_1138;
wire n_4103;
wire n_2529;
wire n_2374;
wire n_5439;
wire n_1225;
wire n_3154;
wire n_1366;
wire n_3938;
wire n_2278;
wire n_1424;
wire n_4736;
wire n_2976;
wire n_4842;
wire n_5250;
wire n_4416;
wire n_4439;
wire n_870;
wire n_4985;
wire n_3382;
wire n_3930;
wire n_3808;
wire n_5471;
wire n_2248;
wire n_813;
wire n_4660;
wire n_3081;
wire n_5497;
wire n_5519;
wire n_995;
wire n_2579;
wire n_1961;
wire n_1535;
wire n_2960;
wire n_3270;
wire n_871;
wire n_2844;
wire n_1979;
wire n_829;
wire n_4814;
wire n_2221;
wire n_5502;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1736;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_3657;
wire n_2634;
wire n_2746;
wire n_5098;
wire n_721;
wire n_1084;
wire n_1276;
wire n_5145;
wire n_2878;
wire n_3830;
wire n_3252;
wire n_5466;
wire n_1528;
wire n_3315;
wire n_3523;
wire n_3999;
wire n_3420;
wire n_3859;
wire n_868;
wire n_5213;
wire n_3474;
wire n_2458;
wire n_3150;
wire n_5491;
wire n_1542;
wire n_4831;
wire n_4782;
wire n_1539;
wire n_2859;
wire n_5216;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1636;
wire n_4597;
wire n_4546;
wire n_5187;
wire n_4031;
wire n_5119;
wire n_1254;
wire n_4147;
wire n_1703;
wire n_3073;
wire n_3571;
wire n_4576;
wire n_3297;
wire n_5148;
wire n_3003;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_5330;
wire n_1560;
wire n_2899;
wire n_4284;
wire n_3274;
wire n_3877;
wire n_5526;
wire n_5202;
wire n_3817;
wire n_2722;
wire n_3728;
wire n_5107;
wire n_4680;
wire n_5067;
wire n_1012;
wire n_2061;
wire n_2685;
wire n_2512;
wire n_1790;
wire n_2788;
wire n_1443;
wire n_5264;
wire n_2595;
wire n_1465;
wire n_3084;
wire n_705;
wire n_4593;
wire n_4562;
wire n_3860;
wire n_2909;
wire n_3554;
wire n_2717;
wire n_1391;
wire n_2981;
wire n_1006;
wire n_4995;
wire n_1159;
wire n_4498;
wire n_772;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_1675;
wire n_2466;
wire n_3758;
wire n_5423;
wire n_2568;
wire n_2271;
wire n_2326;
wire n_3485;
wire n_1594;
wire n_4109;
wire n_1935;
wire n_3777;
wire n_1872;
wire n_1585;
wire n_3767;
wire n_3692;
wire n_1351;
wire n_3234;
wire n_2216;
wire n_2426;
wire n_4850;
wire n_1260;
wire n_3716;
wire n_2926;
wire n_4937;
wire n_798;
wire n_3391;
wire n_912;
wire n_4786;
wire n_5203;
wire n_4354;
wire n_4235;
wire n_3159;
wire n_2855;
wire n_794;
wire n_2848;
wire n_3306;
wire n_2185;
wire n_4345;
wire n_1292;
wire n_1026;
wire n_3460;
wire n_1610;
wire n_5155;
wire n_2202;
wire n_2952;
wire n_3530;
wire n_2693;
wire n_5408;
wire n_3240;
wire n_5066;
wire n_931;
wire n_3362;
wire n_4992;
wire n_4130;
wire n_967;
wire n_5130;
wire n_4175;
wire n_1079;
wire n_5200;
wire n_3393;
wire n_2836;
wire n_2864;
wire n_4456;
wire n_1717;
wire n_2172;
wire n_2601;
wire n_1880;
wire n_2365;
wire n_1399;
wire n_1855;
wire n_2333;
wire n_3629;
wire n_4948;
wire n_5413;
wire n_1903;
wire n_2147;
wire n_4020;
wire n_5150;
wire n_5111;
wire n_1226;
wire n_2224;
wire n_1970;
wire n_3724;
wire n_3287;
wire n_2167;
wire n_2293;
wire n_3046;
wire n_2921;
wire n_1240;
wire n_4984;
wire n_4055;
wire n_4410;
wire n_3980;
wire n_5444;
wire n_3257;
wire n_3730;
wire n_3979;
wire n_5097;
wire n_2695;
wire n_2598;
wire n_3727;
wire n_976;
wire n_4003;
wire n_1832;
wire n_767;
wire n_2302;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_3342;
wire n_2895;
wire n_3796;
wire n_3884;
wire n_4492;
wire n_3625;
wire n_3375;
wire n_2768;
wire n_3760;
wire n_4975;
wire n_3515;
wire n_2363;
wire n_5306;
wire n_2728;
wire n_2025;
wire n_3744;
wire n_5457;
wire n_5159;
wire n_4022;
wire n_1020;
wire n_2495;
wire n_1058;
wire n_4336;
wire n_5314;
wire n_5231;
wire n_5064;
wire n_2223;
wire n_1279;
wire n_2511;
wire n_3981;
wire n_2681;
wire n_1689;
wire n_2535;
wire n_1255;
wire n_3031;
wire n_2335;
wire n_5482;
wire n_3215;
wire n_1401;
wire n_3138;
wire n_776;
wire n_2860;
wire n_2041;
wire n_1933;
wire n_4494;
wire n_4201;
wire n_5287;
wire n_4719;
wire n_3577;
wire n_4074;
wire n_3994;
wire n_4636;
wire n_4983;
wire n_3185;
wire n_1217;
wire n_2662;
wire n_4386;
wire n_3917;
wire n_1231;
wire n_5041;
wire n_4275;
wire n_3774;
wire n_5023;
wire n_5524;
wire n_926;
wire n_2296;
wire n_2178;
wire n_4243;
wire n_2765;
wire n_4225;
wire n_4658;
wire n_4186;
wire n_1501;
wire n_2241;
wire n_4699;
wire n_5139;
wire n_4096;
wire n_2531;
wire n_1570;
wire n_3377;
wire n_1518;
wire n_4907;
wire n_3961;
wire n_5153;
wire n_855;
wire n_2059;
wire n_4713;
wire n_1287;
wire n_1611;
wire n_3374;
wire n_4870;
wire n_4818;
wire n_4916;
wire n_4323;
wire n_1899;
wire n_5376;
wire n_3508;
wire n_4129;
wire n_5488;
wire n_1105;
wire n_3599;
wire n_4480;
wire n_3734;
wire n_3401;
wire n_983;
wire n_699;
wire n_3542;
wire n_3263;
wire n_2523;
wire n_1945;
wire n_2418;
wire n_1377;
wire n_1614;
wire n_5328;
wire n_3819;
wire n_3222;
wire n_1740;
wire n_4616;
wire n_5016;
wire n_5470;
wire n_1092;
wire n_3205;
wire n_4374;
wire n_2225;
wire n_1963;
wire n_3868;
wire n_729;
wire n_2218;
wire n_1122;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_5362;
wire n_2754;
wire n_4580;
wire n_1218;
wire n_3611;
wire n_5147;
wire n_4826;
wire n_3959;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_877;
wire n_3995;
wire n_3908;
wire n_1055;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_1089;
wire n_1502;
wire n_3501;
wire n_1478;
wire n_2555;
wire n_3216;
wire n_3568;
wire n_2708;
wire n_735;
wire n_4844;
wire n_1294;
wire n_4049;
wire n_2661;
wire n_845;
wire n_1649;
wire n_2470;
wire n_1297;
wire n_3551;
wire n_1708;
wire n_5037;
wire n_4677;
wire n_5189;
wire n_4525;
wire n_3364;
wire n_2643;
wire n_755;
wire n_3766;
wire n_3985;
wire n_5055;
wire n_4369;
wire n_3826;
wire n_2266;
wire n_4324;
wire n_842;
wire n_1898;
wire n_1741;
wire n_1907;
wire n_742;
wire n_5160;
wire n_1719;
wire n_2742;
wire n_769;
wire n_3671;
wire n_2366;
wire n_1753;
wire n_5484;
wire n_1372;
wire n_1895;
wire n_4104;
wire n_982;
wire n_3791;
wire n_915;
wire n_2008;
wire n_4989;
wire n_3064;
wire n_3199;
wire n_2127;
wire n_3151;
wire n_3016;
wire n_2460;
wire n_1319;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_4898;
wire n_4081;
wire n_2292;
wire n_2480;
wire n_4528;
wire n_2772;
wire n_1700;
wire n_1332;
wire n_5385;
wire n_1747;
wire n_3990;
wire n_1171;
wire n_4069;
wire n_3582;
wire n_4280;
wire n_1867;
wire n_3993;
wire n_2576;
wire n_3459;
wire n_4811;
wire n_2696;
wire n_5256;
wire n_4779;
wire n_2140;
wire n_2157;
wire n_1966;
wire n_5380;
wire n_1400;
wire n_3735;
wire n_1527;
wire n_1513;
wire n_3656;
wire n_4524;
wire n_2831;
wire n_3069;
wire n_4657;
wire n_4891;
wire n_2629;
wire n_3369;
wire n_1257;
wire n_1954;
wire n_3964;
wire n_5364;
wire n_3302;
wire n_2486;
wire n_1897;
wire n_5469;
wire n_2137;
wire n_3685;
wire n_4977;
wire n_2492;
wire n_2939;
wire n_3425;
wire n_4876;
wire n_5021;
wire n_1449;
wire n_2900;
wire n_797;
wire n_2912;
wire n_1405;
wire n_3813;
wire n_5312;
wire n_2622;
wire n_3447;
wire n_1757;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_3124;
wire n_3811;
wire n_4200;
wire n_2249;
wire n_3411;
wire n_5222;
wire n_3463;
wire n_2785;
wire n_730;
wire n_4938;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_1856;
wire n_1524;
wire n_2928;
wire n_5505;
wire n_1118;
wire n_4604;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_1293;
wire n_961;
wire n_726;
wire n_5504;
wire n_878;
wire n_4118;
wire n_3857;
wire n_3110;
wire n_4239;
wire n_3157;
wire n_1180;
wire n_1697;
wire n_2730;
wire n_5129;
wire n_806;
wire n_1350;
wire n_4704;
wire n_2720;
wire n_1561;
wire n_5494;
wire n_2405;
wire n_2700;
wire n_1616;
wire n_2416;
wire n_2064;
wire n_3640;
wire n_5161;
wire n_1557;
wire n_4744;
wire n_5378;
wire n_4706;
wire n_3879;
wire n_2022;
wire n_4343;
wire n_1505;
wire n_2408;
wire n_4764;
wire n_5389;
wire n_4990;
wire n_2986;
wire n_949;
wire n_2454;
wire n_3591;
wire n_2760;
wire n_4919;
wire n_1208;
wire n_3317;
wire n_4835;
wire n_1151;
wire n_4420;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_5266;
wire n_4559;
wire n_4742;
wire n_5038;
wire n_3566;
wire n_1133;
wire n_883;
wire n_4372;
wire n_5396;
wire n_4097;
wire n_4162;
wire n_5293;
wire n_779;
wire n_4790;
wire n_4173;
wire n_5309;
wire n_3573;
wire n_2943;
wire n_3319;
wire n_2247;
wire n_2230;
wire n_1269;
wire n_4727;
wire n_1547;
wire n_1438;
wire n_3654;
wire n_1047;
wire n_3783;
wire n_4008;
wire n_2158;
wire n_3643;
wire n_2285;
wire n_3184;
wire n_1288;
wire n_2173;
wire n_3982;
wire n_3647;
wire n_1143;
wire n_3973;
wire n_4799;
wire n_4534;
wire n_4960;
wire n_1153;
wire n_1103;
wire n_3738;
wire n_894;
wire n_1380;
wire n_2020;
wire n_2310;
wire n_3600;
wire n_1023;
wire n_914;
wire n_5382;
wire n_4327;
wire n_3190;
wire n_3027;
wire n_4011;
wire n_3695;
wire n_3800;
wire n_3462;
wire n_3906;
wire n_3395;
wire n_3011;
wire n_2820;
wire n_3733;
wire n_1165;
wire n_3967;
wire n_4370;
wire n_4816;
wire n_4091;
wire n_5058;
wire n_1417;
wire n_3096;
wire n_4166;
wire n_2777;
wire n_5356;
wire n_2234;
wire n_1341;
wire n_3233;
wire n_2431;
wire n_3322;
wire n_1603;
wire n_4478;
wire n_2935;
wire n_4246;
wire n_715;
wire n_1066;
wire n_2863;
wire n_2331;
wire n_4632;
wire n_4061;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_4754;
wire n_1534;
wire n_1290;
wire n_4375;
wire n_2396;
wire n_3368;
wire n_1559;
wire n_3117;
wire n_4684;
wire n_743;
wire n_1546;
wire n_3384;
wire n_5279;
wire n_2592;
wire n_3490;
wire n_962;
wire n_5043;
wire n_4241;
wire n_1622;
wire n_2751;
wire n_3113;
wire n_4183;
wire n_918;
wire n_1968;
wire n_5020;
wire n_2842;
wire n_2196;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_3720;
wire n_5232;
wire n_2560;
wire n_4256;
wire n_1164;
wire n_1193;
wire n_1345;
wire n_5035;
wire n_3037;
wire n_1336;
wire n_1033;
wire n_5453;
wire n_4333;
wire n_5339;
wire n_5443;
wire n_1166;
wire n_2007;
wire n_3363;
wire n_1158;
wire n_1803;
wire n_872;
wire n_3522;
wire n_4455;
wire n_3241;
wire n_3899;
wire n_3481;
wire n_5101;
wire n_2236;
wire n_692;
wire n_4457;
wire n_2150;
wire n_1816;
wire n_2803;
wire n_2887;
wire n_2648;
wire n_4735;
wire n_3305;
wire n_3810;
wire n_5170;
wire n_4062;
wire n_2093;
wire n_3354;
wire n_2204;
wire n_1481;
wire n_2040;
wire n_2151;
wire n_2455;
wire n_827;
wire n_3437;
wire n_2231;
wire n_4212;
wire n_4584;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_4477;
wire n_4110;
wire n_5182;
wire n_1221;
wire n_4217;
wire n_5277;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_1579;
wire n_4949;
wire n_2181;
wire n_2014;
wire n_2974;
wire n_923;
wire n_1124;
wire n_1326;
wire n_3969;
wire n_2282;
wire n_4605;
wire n_981;
wire n_3873;
wire n_4649;
wire n_1204;
wire n_994;
wire n_2428;
wire n_1360;
wire n_2858;
wire n_3076;
wire n_3410;
wire n_5415;
wire n_856;
wire n_4592;
wire n_4999;
wire n_1564;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_1361;
wire n_4656;
wire n_1520;
wire n_4862;
wire n_1411;
wire n_1359;
wire n_3536;
wire n_1721;
wire n_3782;
wire n_1317;
wire n_3594;
wire n_5383;
wire n_2385;
wire n_1980;
wire n_4177;
wire n_2501;
wire n_1385;
wire n_1998;
wire n_5029;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_3855;
wire n_2985;
wire n_5218;
wire n_2630;
wire n_2028;
wire n_919;
wire n_3114;
wire n_2092;
wire n_3622;
wire n_2817;
wire n_2773;
wire n_2402;
wire n_1458;
wire n_3047;
wire n_3163;
wire n_5361;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_5512;
wire n_2808;
wire n_2344;
wire n_3520;
wire n_2392;
wire n_3272;
wire n_3122;
wire n_3687;
wire n_2787;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2770;
wire n_4550;
wire n_4347;
wire n_702;
wire n_5193;
wire n_4933;
wire n_968;
wire n_4144;
wire n_5514;
wire n_2375;
wire n_3278;
wire n_4167;
wire n_3608;
wire n_4895;
wire n_1282;
wire n_4726;
wire n_5143;
wire n_1755;
wire n_5188;
wire n_5049;
wire n_2212;
wire n_5308;
wire n_4434;
wire n_5068;
wire n_2569;
wire n_4019;
wire n_4199;
wire n_816;
wire n_1322;
wire n_3829;
wire n_4510;
wire n_5057;
wire n_5425;
wire n_5273;
wire n_2469;
wire n_1125;
wire n_2358;
wire n_1710;
wire n_3546;
wire n_2355;
wire n_1390;
wire n_3068;
wire n_1629;
wire n_1094;
wire n_1510;
wire n_3002;
wire n_1099;
wire n_5248;
wire n_4899;
wire n_3146;
wire n_3038;
wire n_759;
wire n_4156;
wire n_1727;
wire n_3693;
wire n_3132;
wire n_5002;
wire n_5487;
wire n_5531;
wire n_831;
wire n_3681;
wire n_3970;
wire n_778;
wire n_2351;
wire n_1619;
wire n_3188;
wire n_4448;
wire n_3218;
wire n_1152;
wire n_2447;
wire n_2101;
wire n_4193;
wire n_1236;
wire n_4579;
wire n_4776;
wire n_2704;
wire n_1334;
wire n_3729;
wire n_4471;
wire n_4392;
wire n_3103;
wire n_2048;
wire n_3028;
wire n_4691;
wire n_3148;
wire n_3775;
wire n_5461;
wire n_3966;
wire n_4397;
wire n_3616;
wire n_4753;
wire n_4803;
wire n_1289;
wire n_1831;
wire n_3874;
wire n_2191;
wire n_4165;
wire n_2056;
wire n_2852;
wire n_2515;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1941;
wire n_3637;
wire n_1017;
wire n_734;
wire n_4893;
wire n_2240;
wire n_4258;
wire n_709;
wire n_2917;
wire n_3194;
wire n_2085;
wire n_2432;
wire n_5033;
wire n_1686;
wire n_4232;
wire n_5075;
wire n_2097;
wire n_3461;
wire n_1410;
wire n_939;
wire n_2297;
wire n_4203;
wire n_5400;
wire n_1325;
wire n_1223;
wire n_5347;
wire n_2957;
wire n_1983;
wire n_4767;
wire n_4569;
wire n_948;
wire n_3820;
wire n_5144;
wire n_3072;
wire n_2961;
wire n_4468;
wire n_5509;
wire n_1923;
wire n_3848;
wire n_3631;
wire n_5169;
wire n_4885;
wire n_1479;
wire n_4698;
wire n_1031;
wire n_3674;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_5349;
wire n_3763;
wire n_933;
wire n_3499;
wire n_1821;
wire n_3947;
wire n_3910;
wire n_2585;
wire n_5183;
wire n_3361;
wire n_2995;
wire n_4533;
wire n_4287;
wire n_3228;
wire n_2164;
wire n_1732;
wire n_2678;
wire n_1186;
wire n_2052;
wire n_4761;
wire n_4627;
wire n_4556;
wire n_2205;
wire n_2183;
wire n_1724;
wire n_3088;
wire n_1707;
wire n_2080;
wire n_5254;
wire n_3590;
wire n_1126;
wire n_5079;
wire n_2761;
wire n_2357;
wire n_4520;
wire n_895;
wire n_1639;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_3849;
wire n_4263;
wire n_4444;
wire n_5039;
wire n_1818;
wire n_4265;
wire n_3557;
wire n_1598;
wire n_2269;
wire n_1583;
wire n_4612;
wire n_5375;
wire n_5438;
wire n_1264;
wire n_4149;
wire n_1827;
wire n_4958;
wire n_1752;
wire n_2361;
wire n_4538;
wire n_3030;
wire n_3505;
wire n_3075;
wire n_1102;
wire n_2239;
wire n_1296;
wire n_4730;
wire n_4421;
wire n_2464;
wire n_3697;
wire n_882;
wire n_2304;
wire n_2514;
wire n_1299;
wire n_3430;
wire n_2063;
wire n_3489;
wire n_5012;
wire n_2079;
wire n_2152;
wire n_4967;
wire n_2517;
wire n_4696;
wire n_3484;
wire n_4971;
wire n_2095;
wire n_2738;
wire n_2590;
wire n_4661;
wire n_2797;
wire n_3041;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_5422;
wire n_5246;
wire n_4376;
wire n_3832;
wire n_3525;
wire n_3712;
wire n_1069;
wire n_4305;
wire n_2037;
wire n_2953;
wire n_2823;
wire n_3684;
wire n_5404;
wire n_913;
wire n_1681;
wire n_4834;
wire n_1507;
wire n_5332;
wire n_2866;
wire n_3153;
wire n_1174;
wire n_2346;
wire n_4692;
wire n_1353;
wire n_3268;
wire n_2559;
wire n_1383;
wire n_4259;
wire n_2030;
wire n_850;
wire n_4299;
wire n_2407;
wire n_5367;
wire n_2243;
wire n_5288;
wire n_2694;
wire n_3742;
wire n_4965;
wire n_1837;
wire n_4178;
wire n_2006;
wire n_4953;
wire n_4813;
wire n_3352;
wire n_2367;
wire n_5294;
wire n_2731;
wire n_3703;
wire n_5411;
wire n_1246;
wire n_5265;
wire n_2123;
wire n_2238;
wire n_4793;
wire n_4802;
wire n_1196;
wire n_3435;
wire n_2380;
wire n_1187;
wire n_4897;
wire n_1298;
wire n_1745;
wire n_4674;
wire n_4796;
wire n_1088;
wire n_766;
wire n_5184;
wire n_2750;
wire n_2547;
wire n_945;
wire n_4575;
wire n_3665;
wire n_3063;
wire n_3281;
wire n_3535;
wire n_5061;
wire n_2288;
wire n_3858;
wire n_4653;
wire n_4589;
wire n_3220;
wire n_4581;
wire n_4625;
wire n_2107;
wire n_5070;
wire n_4845;
wire n_4148;
wire n_3679;
wire n_738;
wire n_4968;
wire n_2342;
wire n_4590;
wire n_5177;
wire n_3856;
wire n_4038;
wire n_5316;
wire n_2735;
wire n_953;
wire n_4214;
wire n_1888;
wire n_5290;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_3419;
wire n_989;
wire n_5048;
wire n_2233;
wire n_5363;
wire n_795;
wire n_4892;
wire n_1936;
wire n_3890;
wire n_821;
wire n_770;
wire n_1514;
wire n_2782;
wire n_3929;
wire n_971;
wire n_4353;
wire n_2201;
wire n_4950;
wire n_1650;
wire n_4176;
wire n_4124;
wire n_4431;
wire n_1404;
wire n_3347;
wire n_4797;
wire n_4823;
wire n_5462;
wire n_4488;
wire n_5278;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_5214;
wire n_3756;
wire n_4077;
wire n_3209;
wire n_5220;
wire n_4608;
wire n_3948;
wire n_4839;
wire n_1074;
wire n_1765;
wire n_1977;
wire n_2650;
wire n_4454;
wire n_4184;
wire n_2332;
wire n_2391;
wire n_1295;
wire n_2060;
wire n_3883;
wire n_1013;
wire n_4032;
wire n_2571;
wire n_4929;
wire n_2874;
wire n_4117;
wire n_3049;
wire n_3634;
wire n_5436;
wire n_2341;
wire n_1654;
wire n_3066;
wire n_2045;
wire n_3913;
wire n_5341;
wire n_2575;
wire n_3739;
wire n_1230;
wire n_5140;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_4541;
wire n_3271;
wire n_3164;
wire n_3861;
wire n_5096;
wire n_2043;
wire n_4171;
wire n_4815;
wire n_4665;
wire n_4884;
wire n_3580;
wire n_1437;
wire n_4276;
wire n_1378;
wire n_5268;
wire n_5050;
wire n_5240;
wire n_5503;
wire n_1461;
wire n_1876;
wire n_1830;
wire n_5001;
wire n_1112;
wire n_700;
wire n_4174;
wire n_5131;
wire n_5174;
wire n_2145;
wire n_4801;
wire n_4582;
wire n_4774;
wire n_4108;
wire n_5289;
wire n_3119;
wire n_4740;
wire n_1108;
wire n_1274;
wire n_4394;
wire n_4920;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_5069;
wire n_916;
wire n_2810;
wire n_1884;
wire n_1555;
wire n_762;
wire n_1253;
wire n_1468;
wire n_4378;
wire n_5166;
wire n_2683;
wire n_4180;
wire n_4459;
wire n_3624;
wire n_1182;
wire n_4594;
wire n_2748;
wire n_4642;
wire n_1376;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1506;
wire n_3544;
wire n_5300;
wire n_2072;
wire n_3852;
wire n_5233;
wire n_5381;
wire n_1491;
wire n_2628;
wire n_3219;
wire n_1083;
wire n_5333;
wire n_4914;
wire n_3510;
wire n_4587;
wire n_1139;
wire n_3688;
wire n_5008;
wire n_1312;
wire n_3871;
wire n_892;
wire n_3757;
wire n_1567;
wire n_2219;
wire n_2100;
wire n_3666;
wire n_990;
wire n_867;
wire n_3479;
wire n_944;
wire n_5499;
wire n_749;
wire n_2888;
wire n_3998;
wire n_4150;
wire n_1920;
wire n_4285;
wire n_2668;
wire n_2701;
wire n_2400;
wire n_3741;
wire n_2567;
wire n_2557;
wire n_1908;
wire n_1155;
wire n_2755;
wire n_1071;
wire n_5109;
wire n_712;
wire n_909;
wire n_1392;
wire n_2066;
wire n_5281;
wire n_2762;
wire n_964;
wire n_2220;
wire n_4433;
wire n_2829;
wire n_1914;
wire n_2253;
wire n_2130;
wire n_4861;
wire n_2021;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_1633;
wire n_4621;
wire n_3187;
wire n_4451;
wire n_5285;
wire n_2328;
wire n_2434;
wire n_1234;
wire n_3936;
wire n_2261;
wire n_3082;
wire n_5162;
wire n_5442;
wire n_2473;
wire n_4784;
wire n_2438;
wire n_3210;
wire n_3867;
wire n_3397;
wire n_1646;
wire n_2262;
wire n_4613;
wire n_2565;
wire n_1237;
wire n_1095;
wire n_3078;
wire n_3971;
wire n_5117;
wire n_4979;
wire n_3869;
wire n_1531;
wire n_2113;
wire n_1387;
wire n_3711;
wire n_5054;
wire n_3171;
wire n_5394;
wire n_4751;
wire n_4242;
wire n_1951;
wire n_2490;
wire n_2558;
wire n_1496;
wire n_2812;
wire n_3300;
wire n_5496;
wire n_3104;
wire n_4122;
wire n_2132;
wire n_4522;
wire n_4952;
wire n_4426;
wire n_4362;
wire n_3267;
wire n_3946;
wire n_2112;
wire n_2640;
wire n_5000;
wire n_4634;
wire n_4932;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2983;
wire n_5211;
wire n_4089;
wire n_3513;
wire n_1173;
wire n_3498;
wire n_5132;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_4506;
wire n_4728;
wire n_1886;
wire n_4346;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2481;
wire n_3863;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_1365;
wire n_3968;
wire n_3675;
wire n_2437;
wire n_2841;
wire n_3332;
wire n_2055;
wire n_2998;
wire n_1423;
wire n_4359;
wire n_1609;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_4447;
wire n_2937;
wire n_4293;
wire n_5176;
wire n_4039;
wire n_1798;
wire n_3057;
wire n_1608;
wire n_3983;
wire n_703;
wire n_3318;
wire n_3385;
wire n_3773;
wire n_3494;
wire n_1278;
wire n_5074;
wire n_3788;
wire n_3939;
wire n_727;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_3260;
wire n_2496;
wire n_3349;
wire n_4348;
wire n_1602;
wire n_3139;
wire n_3801;
wire n_2338;
wire n_5261;
wire n_1080;
wire n_3636;
wire n_3653;
wire n_3823;
wire n_3403;
wire n_2057;
wire n_1205;
wire n_2716;
wire n_2944;
wire n_2780;
wire n_3439;
wire n_1120;
wire n_1202;
wire n_4084;
wire n_1371;
wire n_4240;
wire n_2033;
wire n_4121;
wire n_3602;
wire n_2774;
wire n_2799;
wire n_4393;
wire n_3984;
wire n_1586;
wire n_1431;
wire n_4389;
wire n_1763;
wire n_4461;
wire n_2763;
wire n_3156;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_4615;
wire n_3044;
wire n_3492;
wire n_3737;
wire n_2379;
wire n_3579;
wire n_1667;
wire n_888;
wire n_3896;
wire n_2300;
wire n_4067;
wire n_1677;
wire n_5244;
wire n_5114;
wire n_4551;
wire n_4521;
wire n_2284;
wire n_3005;
wire n_5420;
wire n_2283;
wire n_5206;
wire n_2526;
wire n_1097;
wire n_1711;
wire n_4387;
wire n_3186;
wire n_2508;
wire n_2594;
wire n_1239;
wire n_5298;
wire n_3417;
wire n_890;
wire n_3626;
wire n_4598;
wire n_4464;
wire n_5106;
wire n_4789;
wire n_3180;
wire n_3423;
wire n_1081;
wire n_2119;
wire n_2493;
wire n_5080;
wire n_4565;
wire n_3392;
wire n_1800;
wire n_5081;
wire n_2904;
wire n_3353;
wire n_2946;
wire n_3512;
wire n_1860;
wire n_1734;
wire n_4552;
wire n_2840;
wire n_4482;
wire n_837;
wire n_812;
wire n_4172;
wire n_4040;
wire n_3024;
wire n_5406;
wire n_4328;
wire n_1854;
wire n_5191;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_2893;
wire n_4940;
wire n_785;
wire n_3161;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1394;
wire n_5085;
wire n_3365;
wire n_4113;
wire n_873;
wire n_3977;
wire n_2468;
wire n_2171;
wire n_4112;
wire n_2035;
wire n_4928;
wire n_2614;
wire n_5428;
wire n_2494;
wire n_1538;
wire n_4865;
wire n_2128;
wire n_4071;
wire n_4436;
wire n_3586;
wire n_4160;
wire n_1668;
wire n_4137;
wire n_1078;
wire n_5417;
wire n_4545;
wire n_4758;
wire n_1161;
wire n_4840;
wire n_3097;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_1191;
wire n_4535;
wire n_4385;
wire n_1215;
wire n_3748;
wire n_4731;
wire n_2337;
wire n_1786;
wire n_3732;
wire n_1804;
wire n_4671;
wire n_2272;
wire n_4766;
wire n_4558;
wire n_1318;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_4319;
wire n_2929;
wire n_4358;
wire n_1526;
wire n_4874;
wire n_2656;
wire n_4904;
wire n_1997;
wire n_1137;
wire n_1258;
wire n_1733;
wire n_4651;
wire n_943;
wire n_3167;
wire n_4748;
wire n_1807;
wire n_1123;
wire n_2857;
wire n_1784;
wire n_4618;
wire n_3787;
wire n_4025;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_752;
wire n_985;
wire n_5506;
wire n_5475;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_1352;
wire n_5431;
wire n_5100;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_5315;
wire n_2633;
wire n_3708;
wire n_2907;
wire n_1429;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1154;
wire n_4910;
wire n_1759;
wire n_2325;
wire n_4724;
wire n_1130;
wire n_3718;
wire n_756;
wire n_3390;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_4666;
wire n_4082;
wire n_3140;
wire n_2320;
wire n_979;
wire n_3976;
wire n_3381;
wire n_897;
wire n_2546;
wire n_2813;
wire n_3736;
wire n_4466;
wire n_891;
wire n_885;
wire n_1659;
wire n_3955;
wire n_5366;
wire n_5322;
wire n_1864;
wire n_5414;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_3336;
wire n_3635;
wire n_3541;
wire n_2502;
wire n_5151;
wire n_714;
wire n_3605;
wire n_5307;
wire n_2170;
wire n_4721;
wire n_725;
wire n_1577;
wire n_5003;
wire n_3840;
wire n_2198;
wire n_5369;
wire n_3067;
wire n_3809;
wire n_4921;
wire n_1852;
wire n_801;
wire n_4377;
wire n_818;
wire n_2410;
wire n_2314;
wire n_5156;
wire n_5270;
wire n_3468;
wire n_1877;
wire n_4301;
wire n_5313;
wire n_2133;
wire n_2497;
wire n_879;
wire n_5446;
wire n_4561;
wire n_1541;
wire n_3291;
wire n_1472;
wire n_1050;
wire n_2578;
wire n_1201;
wire n_1185;
wire n_2475;
wire n_4715;
wire n_2715;
wire n_2665;
wire n_4879;
wire n_5044;
wire n_3755;
wire n_1090;
wire n_4536;
wire n_4304;
wire n_4927;
wire n_4078;
wire n_5459;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_4418;
wire n_3341;
wire n_4125;
wire n_5390;
wire n_5351;
wire n_5267;
wire n_1116;
wire n_5024;
wire n_3043;
wire n_2747;
wire n_1511;
wire n_5275;
wire n_3226;
wire n_3378;
wire n_1641;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_2845;
wire n_4151;
wire n_4412;
wire n_2036;
wire n_843;
wire n_3358;
wire n_2003;
wire n_2533;
wire n_1307;
wire n_4682;
wire n_1128;
wire n_2419;
wire n_2330;
wire n_5078;
wire n_4810;
wire n_3189;
wire n_2309;
wire n_4957;
wire n_4855;
wire n_1955;
wire n_3289;
wire n_1440;
wire n_1370;
wire n_5005;
wire n_1549;
wire n_5207;
wire n_2658;
wire n_3620;
wire n_4601;
wire n_1065;
wire n_4518;
wire n_2767;
wire n_5474;
wire n_3376;
wire n_1362;
wire n_3123;
wire n_5447;
wire n_2692;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_4308;
wire n_2862;
wire n_4325;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_4711;
wire n_2749;
wire n_4413;
wire n_1210;
wire n_3307;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2833;
wire n_1038;
wire n_3723;
wire n_4135;
wire n_5223;
wire n_3880;
wire n_3904;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_3405;
wire n_2313;
wire n_1022;
wire n_5465;
wire n_3532;
wire n_5154;
wire n_2609;
wire n_1767;
wire n_4138;
wire n_1040;
wire n_3131;
wire n_1973;
wire n_1444;
wire n_820;
wire n_2882;
wire n_2303;
wire n_4384;
wire n_4639;
wire n_1664;
wire n_4577;
wire n_2154;
wire n_1986;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_3926;
wire n_4481;
wire n_984;
wire n_5087;
wire n_1552;
wire n_2938;
wire n_2498;
wire n_3992;
wire n_1772;
wire n_1311;
wire n_3106;
wire n_2881;
wire n_3092;
wire n_4270;
wire n_697;
wire n_4620;
wire n_5397;
wire n_4924;
wire n_4044;
wire n_2305;
wire n_880;
wire n_3304;
wire n_4388;
wire n_3247;
wire n_739;
wire n_1028;
wire n_4271;
wire n_2180;
wire n_4406;
wire n_2809;
wire n_975;
wire n_1645;
wire n_932;
wire n_2276;
wire n_3301;
wire n_2910;
wire n_2503;
wire n_3785;
wire n_5492;
wire n_2465;
wire n_5501;
wire n_2972;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_3178;
wire n_2251;
wire n_3100;
wire n_3721;
wire n_3389;
wire n_2126;
wire n_2425;
wire n_4973;
wire n_4792;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_2487;
wire n_5473;
wire n_1834;
wire n_1011;
wire n_2534;
wire n_2941;
wire n_4286;
wire n_3638;
wire n_3576;
wire n_4858;
wire n_1445;
wire n_5370;
wire n_4435;
wire n_3248;
wire n_5317;
wire n_5458;
wire n_2387;
wire n_4318;
wire n_5227;
wire n_830;
wire n_987;
wire n_2510;
wire n_3570;
wire n_3227;
wire n_5359;
wire n_4673;
wire n_2793;
wire n_5282;
wire n_2639;
wire n_4738;
wire n_2603;
wire n_5386;
wire n_1167;
wire n_4554;
wire n_4526;
wire n_4105;
wire n_969;
wire n_3663;
wire n_1663;
wire n_2086;
wire n_1926;
wire n_1630;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_3431;
wire n_3355;
wire n_1738;
wire n_3897;
wire n_1735;
wire n_4005;
wire n_4181;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_956;
wire n_765;
wire n_4092;
wire n_4875;
wire n_4255;
wire n_2758;
wire n_5036;
wire n_1271;
wire n_2186;
wire n_4647;
wire n_3575;
wire n_2471;
wire n_3042;
wire n_1067;
wire n_1323;
wire n_1937;
wire n_4142;
wire n_5118;
wire n_900;
wire n_5485;
wire n_5525;
wire n_3004;
wire n_1551;
wire n_4849;
wire n_5271;
wire n_2039;
wire n_1285;
wire n_733;
wire n_761;
wire n_3838;
wire n_4059;
wire n_5194;
wire n_5445;
wire n_2734;
wire n_4499;
wire n_4504;
wire n_3598;
wire n_4917;
wire n_2420;
wire n_3273;
wire n_2918;
wire n_835;
wire n_1865;
wire n_2641;
wire n_2463;
wire n_2580;
wire n_1792;
wire n_5245;
wire n_2062;
wire n_4489;
wire n_822;
wire n_1459;
wire n_2153;
wire n_5329;
wire n_5472;
wire n_839;
wire n_1754;
wire n_4833;
wire n_3394;
wire n_2235;
wire n_1575;
wire n_4564;
wire n_1848;
wire n_1172;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_3581;
wire n_5072;
wire n_3778;
wire n_4322;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_4080;
wire n_2206;
wire n_997;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_3001;
wire n_5260;
wire n_4981;
wire n_2347;
wire n_4676;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_2362;
wire n_5372;
wire n_4507;
wire n_4756;
wire n_1576;
wire n_2422;
wire n_2933;
wire n_3387;
wire n_3952;
wire n_4365;
wire n_3584;
wire n_4349;
wire n_3446;
wire n_1059;
wire n_2736;
wire n_3825;
wire n_4198;
wire n_977;
wire n_2339;
wire n_2532;
wire n_4373;
wire n_1866;
wire n_2664;
wire n_4154;
wire n_4390;
wire n_1782;
wire n_1558;
wire n_4107;
wire n_2519;
wire n_4380;
wire n_4361;
wire n_4609;
wire n_2360;
wire n_4453;
wire n_723;
wire n_1393;
wire n_4571;
wire n_3137;
wire n_2544;
wire n_809;
wire n_3032;
wire n_4886;
wire n_5172;
wire n_881;
wire n_1477;
wire n_1019;
wire n_1982;
wire n_5311;
wire n_910;
wire n_5164;
wire n_4964;
wire n_4700;
wire n_4002;
wire n_1114;
wire n_1742;
wire n_4679;
wire n_3815;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_1273;
wire n_2982;
wire n_5495;
wire n_4483;
wire n_3061;
wire n_3504;
wire n_2587;
wire n_4693;
wire n_1043;
wire n_5121;
wire n_4956;
wire n_2869;
wire n_5379;
wire n_4487;
wire n_2674;
wire n_1737;
wire n_1613;
wire n_3026;
wire n_2979;
wire n_4329;
wire n_5291;
wire n_4010;
wire n_4501;
wire n_4808;
wire n_3902;
wire n_3244;
wire n_1779;
wire n_2562;
wire n_954;
wire n_3112;
wire n_2051;
wire n_3196;
wire n_2673;
wire n_4678;
wire n_1591;
wire n_5301;
wire n_5126;
wire n_2548;
wire n_3488;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_3779;
wire n_1063;
wire n_991;
wire n_2275;
wire n_4606;
wire n_3834;
wire n_4303;
wire n_2029;
wire n_1912;
wire n_3923;
wire n_938;
wire n_1891;
wire n_5348;
wire n_1000;
wire n_4868;
wire n_4072;
wire n_2792;
wire n_4465;
wire n_2596;
wire n_5217;
wire n_3986;
wire n_3725;
wire n_4026;
wire n_4245;
wire n_5520;
wire n_2524;
wire n_3894;
wire n_1702;
wire n_4852;
wire n_3202;
wire n_4290;
wire n_4945;
wire n_1232;
wire n_1211;
wire n_996;
wire n_1082;
wire n_1725;
wire n_2318;
wire n_866;
wire n_2819;
wire n_1722;
wire n_2229;
wire n_1644;
wire n_3547;
wire n_4014;
wire n_2551;
wire n_2255;
wire n_1252;
wire n_3045;
wire n_773;
wire n_5135;
wire n_4599;
wire n_2706;
wire n_4222;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_5448;
wire n_2573;
wire n_2336;
wire n_5412;
wire n_1662;
wire n_3249;
wire n_3483;
wire n_4046;
wire n_4701;
wire n_1925;
wire n_782;
wire n_2915;
wire n_4869;
wire n_3213;
wire n_5533;
wire n_4047;
wire n_1244;
wire n_1796;
wire n_2719;
wire n_2876;
wire n_4063;
wire n_5224;
wire n_2778;
wire n_1574;
wire n_3033;
wire n_893;
wire n_1582;
wire n_1981;
wire n_2824;
wire n_5327;
wire n_4417;
wire n_796;
wire n_1374;
wire n_2089;
wire n_4688;
wire n_4939;
wire n_1486;
wire n_3619;
wire n_4013;
wire n_3434;
wire n_4342;
wire n_4903;
wire n_2131;
wire n_3853;
wire n_4382;
wire n_2509;
wire n_4085;
wire n_5486;
wire n_2135;
wire n_4475;
wire n_5432;
wire n_1463;
wire n_4626;
wire n_4997;
wire n_5065;
wire n_924;
wire n_781;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_2436;
wire n_3517;
wire n_1706;
wire n_2461;
wire n_3719;
wire n_1214;
wire n_3526;
wire n_3888;
wire n_3198;
wire n_1853;
wire n_764;
wire n_1503;
wire n_5295;
wire n_1181;
wire n_1999;
wire n_4841;
wire n_4683;
wire n_5173;
wire n_2873;
wire n_2084;
wire n_3330;
wire n_3514;
wire n_3383;
wire n_1835;
wire n_3965;
wire n_1457;
wire n_3905;
wire n_3797;
wire n_1836;
wire n_3416;
wire n_4600;
wire n_1453;
wire n_3943;
wire n_3145;
wire n_2908;
wire n_4106;
wire n_2156;
wire n_1184;
wire n_754;
wire n_2323;
wire n_1073;
wire n_4549;
wire n_1277;
wire n_1746;
wire n_1062;
wire n_4702;
wire n_5102;
wire n_4954;
wire n_740;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_3283;
wire n_4331;
wire n_4159;
wire n_3451;
wire n_4734;
wire n_2832;
wire n_1688;
wire n_2370;
wire n_1944;
wire n_2914;
wire n_1988;
wire n_1718;
wire n_4515;
wire n_2149;
wire n_2277;
wire n_2539;
wire n_2078;
wire n_1145;
wire n_4809;
wire n_787;
wire n_4012;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_5212;
wire n_4760;
wire n_1207;
wire n_3606;
wire n_2232;
wire n_1847;
wire n_4320;
wire n_5084;
wire n_5251;
wire n_1314;
wire n_1512;
wire n_884;
wire n_4980;
wire n_3324;
wire n_2192;
wire n_5407;
wire n_2988;
wire n_4560;
wire n_3230;
wire n_3793;
wire n_859;
wire n_5042;
wire n_4768;
wire n_1889;
wire n_693;
wire n_5368;
wire n_929;
wire n_3207;
wire n_3641;
wire n_3828;
wire n_1850;
wire n_3183;
wire n_3607;
wire n_1637;
wire n_2427;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_5310;
wire n_2769;
wire n_1548;
wire n_4987;
wire n_3013;
wire n_4572;
wire n_1396;
wire n_2739;
wire n_3962;
wire n_4988;
wire n_2902;
wire n_4360;
wire n_1544;
wire n_4540;
wire n_2094;
wire n_3854;
wire n_1354;
wire n_2349;
wire n_3652;
wire n_3449;
wire n_1021;
wire n_3089;
wire n_4854;
wire n_1595;
wire n_1142;
wire n_5477;
wire n_2727;
wire n_942;
wire n_5234;
wire n_1416;
wire n_1599;
wire n_4747;
wire n_3472;
wire n_2527;
wire n_3126;
wire n_2759;
wire n_5007;
wire n_4881;
wire n_2038;
wire n_3958;
wire n_4495;
wire n_4737;
wire n_1838;
wire n_4357;
wire n_2806;
wire n_4502;
wire n_3191;
wire n_1716;
wire n_5334;
wire n_3562;
wire n_2281;
wire n_5253;
wire n_3588;
wire n_1590;
wire n_3280;
wire n_4115;
wire n_5274;
wire n_5418;
wire n_5019;
wire n_1819;
wire n_3095;
wire n_947;
wire n_3698;
wire n_4513;
wire n_1179;
wire n_696;
wire n_1442;
wire n_4775;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_2499;
wire n_2549;
wire n_804;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_3885;
wire n_955;
wire n_4264;
wire n_2166;
wire n_3192;
wire n_4709;
wire n_1562;
wire n_3250;
wire n_4223;
wire n_3538;
wire n_3915;
wire n_3839;
wire n_5490;
wire n_1972;
wire n_4718;
wire n_3717;
wire n_5489;
wire n_3407;
wire n_3875;
wire n_4029;
wire n_4206;
wire n_2415;
wire n_4099;
wire n_3120;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_5342;
wire n_4794;
wire n_4843;
wire n_5215;
wire n_3937;
wire n_4763;
wire n_1418;
wire n_4170;
wire n_2462;
wire n_2155;
wire n_2439;
wire n_4838;
wire n_4795;
wire n_3604;
wire n_5430;
wire n_824;
wire n_4272;
wire n_5195;
wire n_3176;
wire n_3792;
wire n_4267;
wire n_2083;
wire n_815;
wire n_2753;
wire n_1340;
wire n_3021;
wire n_4352;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_3912;
wire n_3950;
wire n_2898;
wire n_1825;
wire n_3567;
wire n_2682;
wire n_5112;
wire n_5326;
wire n_1627;
wire n_2903;
wire n_5303;
wire n_3812;
wire n_3127;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_5530;
wire n_965;
wire n_934;
wire n_2213;
wire n_4056;
wire n_4806;
wire n_1674;
wire n_4015;
wire n_2924;
wire n_4445;
wire n_4462;
wire n_5299;
wire n_4219;
wire n_4484;
wire n_4723;
wire n_2142;
wire n_4517;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_4043;
wire n_1042;
wire n_3170;
wire n_2311;
wire n_1455;
wire n_2287;
wire n_836;
wire n_3415;
wire n_3464;
wire n_3414;
wire n_4234;
wire n_760;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_3467;
wire n_713;
wire n_3179;
wire n_5522;
wire n_4836;
wire n_3889;
wire n_5262;
wire n_3262;
wire n_5319;
wire n_927;
wire n_3699;
wire n_706;
wire n_2120;
wire n_1419;
wire n_3816;
wire n_3528;
wire n_4207;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_4725;
wire n_2312;
wire n_1826;
wire n_4880;
wire n_2834;
wire n_4051;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_5335;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_4334;
wire n_5284;
wire n_4978;
wire n_3246;
wire n_3299;
wire n_980;
wire n_1618;
wire n_1869;
wire n_3623;
wire n_905;
wire n_2718;
wire n_4707;
wire n_2687;
wire n_4923;
wire n_4911;
wire n_3876;
wire n_5516;
wire n_3615;
wire n_1802;
wire n_2811;
wire n_3019;
wire n_5168;
wire n_3200;
wire n_3642;
wire n_2146;
wire n_4274;
wire n_3276;
wire n_5433;
wire n_3682;
wire n_5429;
wire n_4007;
wire n_1456;
wire n_1879;
wire n_2129;
wire n_814;
wire n_5120;
wire n_3572;
wire n_2975;
wire n_2399;
wire n_1134;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_2027;
wire n_2932;
wire n_3118;
wire n_4441;
wire n_3039;
wire n_3922;
wire n_2195;
wire n_5455;
wire n_1467;
wire n_5209;
wire n_4458;
wire n_2159;
wire n_4889;
wire n_3831;
wire n_1744;
wire n_4523;
wire n_3618;
wire n_3705;
wire n_3022;
wire n_1709;
wire n_5099;
wire n_3286;
wire n_2023;
wire n_3974;
wire n_3443;
wire n_2599;
wire n_3988;
wire n_5022;
wire n_2075;
wire n_1726;
wire n_2031;
wire n_3761;
wire n_3996;
wire n_5353;
wire n_4771;
wire n_2853;
wire n_3350;
wire n_1098;
wire n_3009;
wire n_777;
wire n_5219;
wire n_920;
wire n_3951;
wire n_5518;
wire n_3035;
wire n_4261;
wire n_1132;
wire n_1823;
wire n_5236;
wire n_4236;
wire n_3942;
wire n_3023;
wire n_2254;
wire n_3290;
wire n_1402;
wire n_3957;
wire n_3418;
wire n_1607;
wire n_861;
wire n_1666;
wire n_5103;
wire n_4648;
wire n_2214;
wire n_2256;
wire n_3326;
wire n_2732;
wire n_1883;
wire n_4094;
wire n_2776;
wire n_3224;
wire n_1969;
wire n_2949;
wire n_4269;
wire n_1927;
wire n_1222;
wire n_3803;
wire n_5239;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_4913;
wire n_2449;
wire n_4428;
wire n_745;
wire n_1572;
wire n_4463;
wire n_5357;
wire n_3648;
wire n_1975;
wire n_5421;
wire n_1388;
wire n_1266;
wire n_4396;
wire n_1990;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_1075;
wire n_1890;
wire n_4034;
wire n_4228;
wire n_1227;
wire n_3166;
wire n_3649;
wire n_3065;
wire n_5045;
wire n_5237;
wire n_3924;
wire n_3997;
wire n_3564;
wire n_862;
wire n_2637;
wire n_3795;
wire n_4931;
wire n_2306;
wire n_2071;
wire n_3953;
wire n_4400;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_5434;
wire n_1532;
wire n_1030;
wire n_5181;
wire n_3208;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_852;
wire n_2916;
wire n_1060;
wire n_4424;
wire n_4351;
wire n_4192;
wire n_1748;
wire n_1301;
wire n_3400;
wire n_1466;
wire n_2581;
wire n_1783;
wire n_5146;
wire n_4646;
wire n_4221;
wire n_1037;
wire n_3650;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_4035;
wire n_1480;
wire n_3670;
wire n_2540;
wire n_4190;
wire n_1605;
wire n_3060;
wire n_2984;
wire n_4009;
wire n_2489;
wire n_5013;
wire n_4145;
wire n_876;
wire n_5017;
wire n_736;
wire n_2265;
wire n_3524;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_2106;
wire n_4717;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_854;
wire n_2091;
wire n_4312;
wire n_5424;
wire n_3789;
wire n_1658;
wire n_1072;
wire n_1305;
wire n_4750;
wire n_2348;
wire n_1873;
wire n_2667;
wire n_2725;
wire n_3746;
wire n_4537;
wire n_1046;
wire n_3694;
wire n_771;
wire n_5456;
wire n_3893;
wire n_4847;
wire n_2307;
wire n_3702;
wire n_1984;
wire n_3453;
wire n_1556;
wire n_5345;
wire n_2815;
wire n_4427;
wire n_1824;
wire n_1492;
wire n_4065;
wire n_4705;
wire n_819;
wire n_1971;
wire n_2945;
wire n_1324;
wire n_3543;
wire n_1776;
wire n_3448;
wire n_4279;
wire n_2936;
wire n_3609;
wire n_4330;
wire n_4152;
wire n_2698;
wire n_4783;
wire n_3017;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2789;
wire n_5409;
wire n_2525;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_807;
wire n_5142;
wire n_3907;
wire n_4603;
wire n_5010;
wire n_4332;
wire n_1987;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_802;
wire n_5401;
wire n_4595;
wire n_960;
wire n_2352;
wire n_5201;
wire n_790;
wire n_5416;
wire n_4404;
wire n_2377;
wire n_2652;
wire n_5498;
wire n_4054;
wire n_1286;
wire n_4617;
wire n_1685;
wire n_2477;
wire n_4611;
wire n_2279;
wire n_3169;
wire n_2222;
wire n_1052;
wire n_4732;
wire n_2076;
wire n_2203;
wire n_1426;
wire n_4969;
wire n_5252;
wire n_5063;
wire n_4641;
wire n_4399;
wire n_4140;
wire n_5171;
wire n_2607;
wire n_3343;
wire n_4712;
wire n_3309;
wire n_2796;
wire n_858;
wire n_5393;
wire n_4817;
wire n_2136;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_2771;
wire n_2403;
wire n_2947;
wire n_928;
wire n_3769;
wire n_1565;
wire n_4437;
wire n_3055;
wire n_4070;
wire n_5346;
wire n_748;
wire n_1045;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_4139;
wire n_4769;
wire n_1958;
wire n_4867;
wire n_3667;
wire n_2713;
wire n_1422;
wire n_1965;
wire n_5167;
wire n_5257;
wire n_4450;
wire n_2934;
wire n_5104;
wire n_2210;
wire n_4368;
wire n_3141;
wire n_2053;
wire n_5272;
wire n_3476;
wire n_1049;
wire n_4430;
wire n_3238;
wire n_2450;
wire n_5338;
wire n_1356;
wire n_1773;
wire n_3175;
wire n_4544;
wire n_2666;
wire n_728;
wire n_4191;
wire n_4409;
wire n_2401;
wire n_3255;
wire n_2588;
wire n_935;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_2478;
wire n_911;
wire n_3509;
wire n_1403;
wire n_5395;
wire n_3006;
wire n_4531;
wire n_3770;
wire n_3456;
wire n_4532;
wire n_3790;
wire n_907;
wire n_847;
wire n_747;
wire n_1135;
wire n_2566;
wire n_5095;
wire n_3101;
wire n_3662;
wire n_5199;
wire n_4257;
wire n_4282;
wire n_4341;
wire n_1694;
wire n_1695;
wire n_4027;
wire n_4309;
wire n_4650;
wire n_5480;
wire n_3077;
wire n_4944;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_4994;
wire n_3533;
wire n_5175;
wire n_1994;
wire n_3978;
wire n_3836;
wire n_3409;
wire n_4381;
wire n_3583;
wire n_4316;
wire n_4860;
wire n_4469;
wire n_3540;
wire n_4930;
wire n_5352;
wire n_1157;
wire n_3563;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_3689;
wire n_1789;
wire n_763;
wire n_2174;
wire n_3442;
wire n_3972;
wire n_2315;
wire n_4209;
wire n_1687;
wire n_4703;
wire n_4934;
wire n_2638;
wire n_2046;
wire n_1756;
wire n_4350;
wire n_1606;
wire n_1587;
wire n_2340;
wire n_4804;
wire n_2444;
wire n_4888;
wire n_1014;
wire n_1427;
wire n_2977;
wire n_3991;
wire n_4936;
wire n_2199;
wire n_4669;
wire n_5228;
wire n_1100;
wire n_1617;
wire n_2600;
wire n_3436;
wire n_1962;
wire n_3806;
wire n_4759;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3833;
wire n_1175;
wire n_4887;
wire n_3751;
wire n_3402;
wire n_1621;
wire n_5186;
wire n_4585;
wire n_1785;
wire n_3406;
wire n_3664;
wire n_4218;
wire n_4687;
wire n_1381;
wire n_3686;
wire n_1183;
wire n_4720;
wire n_2889;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_3470;
wire n_5221;
wire n_1407;
wire n_2865;
wire n_973;
wire n_4762;
wire n_3844;
wire n_3259;
wire n_2572;
wire n_4490;
wire n_1248;
wire n_1176;
wire n_3677;
wire n_1054;
wire n_5387;
wire n_3292;
wire n_3989;
wire n_4644;
wire n_4752;
wire n_4746;
wire n_1057;
wire n_4131;
wire n_5449;
wire n_4215;
wire n_978;
wire n_2488;
wire n_1509;
wire n_828;
wire n_4158;
wire n_3079;
wire n_5190;
wire n_3269;
wire n_5325;
wire n_4231;
wire n_5047;
wire n_2591;
wire n_5004;
wire n_4926;
wire n_2050;
wire n_2197;
wire n_4872;
wire n_4778;
wire n_5344;
wire n_2550;
wire n_1536;
wire n_3177;
wire n_4667;
wire n_1471;
wire n_3440;
wire n_3658;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1620;
wire n_2542;
wire n_2165;
wire n_4837;
wire n_4210;
wire n_788;
wire n_2169;
wire n_5133;
wire n_5305;
wire n_2175;
wire n_1625;
wire n_4578;
wire n_3644;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_1922;
wire n_940;
wire n_1537;
wire n_4877;
wire n_2065;
wire n_4470;
wire n_4187;
wire n_1904;
wire n_4998;
wire n_2395;
wire n_2868;
wire n_1530;
wire n_4057;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_898;
wire n_3328;
wire n_2012;
wire n_3182;
wire n_2967;
wire n_5343;
wire n_1093;
wire n_4021;
wire n_3379;
wire n_4379;
wire n_2268;
wire n_3469;
wire n_1452;
wire n_2835;
wire n_2111;
wire n_3743;
wire n_2948;
wire n_5015;
wire n_3099;
wire n_5527;
wire n_2897;
wire n_4812;
wire n_4497;
wire n_2583;
wire n_3155;
wire n_4300;
wire n_2024;
wire n_1770;
wire n_701;
wire n_1003;
wire n_4472;
wire n_2699;
wire n_3901;
wire n_5180;
wire n_1640;
wire n_2973;
wire n_2710;
wire n_2505;
wire n_4519;
wire n_5025;
wire n_2397;
wire n_3878;
wire n_4197;
wire n_2721;
wire n_1892;
wire n_2615;
wire n_4787;
wire n_1212;
wire n_4310;
wire n_4566;
wire n_3933;
wire n_4371;
wire n_1902;
wire n_2784;
wire n_3898;
wire n_694;
wire n_4749;
wire n_1845;
wire n_921;
wire n_2104;
wire n_2552;
wire n_1470;
wire n_1533;
wire n_5083;
wire n_3253;
wire n_2088;
wire n_1275;
wire n_4238;
wire n_904;
wire n_2005;
wire n_1696;
wire n_2108;
wire n_3824;
wire n_2246;
wire n_3846;
wire n_5122;
wire n_1497;
wire n_4189;
wire n_2472;
wire n_2705;
wire n_4479;
wire n_3845;
wire n_3203;
wire n_4986;
wire n_1316;
wire n_4668;
wire n_950;
wire n_711;
wire n_4168;
wire n_1369;
wire n_4298;
wire n_4743;
wire n_1781;
wire n_4250;
wire n_3143;
wire n_3690;
wire n_3229;
wire n_2188;
wire n_2430;
wire n_2504;
wire n_4211;
wire n_3094;
wire n_741;
wire n_5185;
wire n_2964;
wire n_5032;
wire n_865;
wire n_5034;
wire n_3312;
wire n_1041;
wire n_2451;
wire n_2913;
wire n_993;
wire n_1862;
wire n_3752;
wire n_3672;
wire n_922;
wire n_1004;
wire n_2839;
wire n_3237;
wire n_4128;
wire n_4036;
wire n_5269;
wire n_3655;
wire n_2955;
wire n_1764;
wire n_4807;
wire n_5115;
wire n_902;
wire n_1723;
wire n_3918;
wire n_5324;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_1946;
wire n_4383;
wire n_4830;
wire n_4391;
wire n_4095;
wire n_1310;
wire n_4485;
wire n_3593;
wire n_5163;
wire n_1229;
wire n_2582;
wire n_3327;
wire n_4356;
wire n_1896;
wire n_1516;
wire n_4890;
wire n_2485;
wire n_2563;
wire n_4224;
wire n_1670;
wire n_1799;
wire n_5507;
wire n_4573;
wire n_1328;
wire n_4943;
wire n_2875;
wire n_3519;
wire n_2209;
wire n_4042;
wire n_4244;
wire n_1928;
wire n_4708;
wire n_4883;
wire n_4553;
wire n_1634;
wire n_1203;
wire n_1699;
wire n_5226;
wire n_2081;
wire n_937;
wire n_1474;
wire n_1631;
wire n_1794;
wire n_1375;
wire n_3053;
wire n_5014;
wire n_3772;
wire n_2891;
wire n_4335;
wire n_3128;
wire n_4277;
wire n_4614;
wire n_4629;
wire n_1002;
wire n_4516;
wire n_5235;
wire n_1129;
wire n_1464;
wire n_2798;
wire n_3217;
wire n_1249;
wire n_3821;
wire n_3201;
wire n_3503;
wire n_1870;
wire n_4467;
wire n_5521;
wire n_2654;
wire n_3935;
wire n_1861;
wire n_1228;
wire n_2319;
wire n_2965;
wire n_4955;
wire n_5410;
wire n_1251;
wire n_1989;
wire n_2689;
wire n_1762;
wire n_3798;
wire n_3080;
wire n_5241;
wire n_4248;
wire n_1672;
wire n_2228;
wire n_4645;
wire n_5331;
wire n_3308;
wire n_841;
wire n_3204;
wire n_4134;
wire n_5018;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_2345;
wire n_1730;
wire n_5258;

INVx1_ASAP7_75t_L g692 ( 
.A(n_679),
.Y(n_692)
);

CKINVDCx20_ASAP7_75t_R g693 ( 
.A(n_9),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_95),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_664),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_94),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_399),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_499),
.Y(n_698)
);

CKINVDCx20_ASAP7_75t_R g699 ( 
.A(n_439),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_363),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_516),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_253),
.Y(n_702)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_94),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_128),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_356),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_90),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_475),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_632),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_45),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_431),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_39),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_539),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_47),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_429),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_431),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_165),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_164),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_486),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_311),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_122),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_276),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_298),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_432),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_466),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_520),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_49),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_635),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_507),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_666),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_86),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_556),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_98),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_576),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_191),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_365),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_271),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_467),
.Y(n_737)
);

BUFx8_ASAP7_75t_SL g738 ( 
.A(n_17),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_538),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_88),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_190),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_453),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_629),
.Y(n_743)
);

CKINVDCx20_ASAP7_75t_R g744 ( 
.A(n_315),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_2),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_590),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_179),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_444),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_476),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_198),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_498),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_325),
.Y(n_752)
);

CKINVDCx14_ASAP7_75t_R g753 ( 
.A(n_241),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_441),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_402),
.Y(n_755)
);

INVx1_ASAP7_75t_SL g756 ( 
.A(n_50),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_225),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_666),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_311),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_547),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_395),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_82),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_302),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_63),
.Y(n_764)
);

INVxp67_ASAP7_75t_SL g765 ( 
.A(n_389),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_47),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_98),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_135),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_399),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_472),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_251),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_154),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_502),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_637),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_101),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_433),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_262),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_602),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_97),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_29),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_555),
.Y(n_781)
);

INVx1_ASAP7_75t_SL g782 ( 
.A(n_496),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_273),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_274),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_689),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_456),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_138),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_208),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_16),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_679),
.Y(n_790)
);

CKINVDCx20_ASAP7_75t_R g791 ( 
.A(n_526),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_505),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_501),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_306),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_591),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_132),
.Y(n_796)
);

BUFx3_ASAP7_75t_L g797 ( 
.A(n_327),
.Y(n_797)
);

INVx1_ASAP7_75t_SL g798 ( 
.A(n_310),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_174),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_677),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_474),
.Y(n_801)
);

CKINVDCx20_ASAP7_75t_R g802 ( 
.A(n_408),
.Y(n_802)
);

CKINVDCx20_ASAP7_75t_R g803 ( 
.A(n_49),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_192),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_211),
.Y(n_805)
);

CKINVDCx20_ASAP7_75t_R g806 ( 
.A(n_686),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_542),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_558),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_214),
.Y(n_809)
);

BUFx5_ASAP7_75t_L g810 ( 
.A(n_415),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_654),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_86),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_218),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_673),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_587),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_183),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_341),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_455),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_482),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_651),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_447),
.Y(n_821)
);

CKINVDCx20_ASAP7_75t_R g822 ( 
.A(n_133),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_197),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_471),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_39),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_119),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_404),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_385),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_196),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_471),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_360),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_392),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_585),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_676),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_446),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_577),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_16),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_680),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_672),
.Y(n_839)
);

BUFx3_ASAP7_75t_L g840 ( 
.A(n_557),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_610),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_147),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_468),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_623),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_224),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_174),
.Y(n_846)
);

INVx1_ASAP7_75t_SL g847 ( 
.A(n_72),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_428),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_187),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_187),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_336),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_682),
.Y(n_852)
);

BUFx10_ASAP7_75t_L g853 ( 
.A(n_59),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_233),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_78),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_516),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_123),
.Y(n_857)
);

BUFx10_ASAP7_75t_L g858 ( 
.A(n_678),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_360),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_572),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_510),
.Y(n_861)
);

BUFx5_ASAP7_75t_L g862 ( 
.A(n_127),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_7),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_281),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_557),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_598),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_290),
.Y(n_867)
);

CKINVDCx20_ASAP7_75t_R g868 ( 
.A(n_248),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_301),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_570),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_19),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_133),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_517),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_435),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_404),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_355),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_222),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_364),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_614),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_185),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_192),
.Y(n_881)
);

CKINVDCx20_ASAP7_75t_R g882 ( 
.A(n_612),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_594),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_549),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_475),
.Y(n_885)
);

CKINVDCx20_ASAP7_75t_R g886 ( 
.A(n_338),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_590),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_220),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_391),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_656),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_316),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_600),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_281),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_175),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_240),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_110),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_416),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_576),
.Y(n_898)
);

CKINVDCx16_ASAP7_75t_R g899 ( 
.A(n_2),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_463),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_318),
.Y(n_901)
);

CKINVDCx20_ASAP7_75t_R g902 ( 
.A(n_97),
.Y(n_902)
);

CKINVDCx20_ASAP7_75t_R g903 ( 
.A(n_132),
.Y(n_903)
);

CKINVDCx20_ASAP7_75t_R g904 ( 
.A(n_596),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_465),
.Y(n_905)
);

BUFx10_ASAP7_75t_L g906 ( 
.A(n_618),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_513),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_422),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_683),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_396),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_44),
.Y(n_911)
);

BUFx10_ASAP7_75t_L g912 ( 
.A(n_374),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_684),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_540),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_676),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_459),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_490),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_568),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_349),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_327),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_4),
.Y(n_921)
);

INVx1_ASAP7_75t_SL g922 ( 
.A(n_363),
.Y(n_922)
);

INVx3_ASAP7_75t_L g923 ( 
.A(n_586),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_535),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_37),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_354),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_522),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_30),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_302),
.Y(n_929)
);

CKINVDCx16_ASAP7_75t_R g930 ( 
.A(n_128),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_686),
.Y(n_931)
);

INVxp67_ASAP7_75t_SL g932 ( 
.A(n_427),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_7),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_401),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_319),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_190),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_610),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_448),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_357),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_553),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_631),
.Y(n_941)
);

INVxp67_ASAP7_75t_SL g942 ( 
.A(n_172),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_681),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_626),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_18),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_287),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_120),
.Y(n_947)
);

INVxp33_ASAP7_75t_SL g948 ( 
.A(n_125),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_27),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_88),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_453),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_296),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_632),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_397),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_226),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_565),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_48),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_51),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_110),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_313),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_112),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_601),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_682),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_602),
.Y(n_964)
);

INVx2_ASAP7_75t_SL g965 ( 
.A(n_371),
.Y(n_965)
);

BUFx10_ASAP7_75t_L g966 ( 
.A(n_477),
.Y(n_966)
);

BUFx3_ASAP7_75t_L g967 ( 
.A(n_161),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_467),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_611),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_344),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_506),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_9),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_197),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_495),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_635),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_527),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_647),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_7),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_135),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_407),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_654),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_138),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_459),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_627),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_0),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_214),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_109),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_675),
.Y(n_988)
);

INVx2_ASAP7_75t_SL g989 ( 
.A(n_649),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_120),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_643),
.Y(n_991)
);

INVx1_ASAP7_75t_SL g992 ( 
.A(n_612),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_162),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_413),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_306),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_198),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_179),
.Y(n_997)
);

CKINVDCx20_ASAP7_75t_R g998 ( 
.A(n_305),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_366),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_190),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_532),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_381),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_186),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_21),
.Y(n_1004)
);

CKINVDCx16_ASAP7_75t_R g1005 ( 
.A(n_674),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_519),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_246),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_208),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_473),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_449),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_276),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_554),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_194),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_50),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_232),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_508),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_0),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_37),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_617),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_67),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_426),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_535),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_318),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_118),
.B(n_109),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_136),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_162),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_553),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_495),
.Y(n_1028)
);

BUFx10_ASAP7_75t_L g1029 ( 
.A(n_740),
.Y(n_1029)
);

INVxp67_ASAP7_75t_L g1030 ( 
.A(n_738),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_753),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_758),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_1005),
.Y(n_1033)
);

CKINVDCx20_ASAP7_75t_R g1034 ( 
.A(n_693),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_874),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_874),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_698),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_700),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_874),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_923),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_923),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_923),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_862),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_862),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_862),
.Y(n_1045)
);

BUFx5_ASAP7_75t_L g1046 ( 
.A(n_694),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_710),
.Y(n_1047)
);

CKINVDCx16_ASAP7_75t_R g1048 ( 
.A(n_899),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_862),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_758),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_862),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_718),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_862),
.Y(n_1053)
);

CKINVDCx20_ASAP7_75t_R g1054 ( 
.A(n_703),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_862),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_719),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_862),
.Y(n_1057)
);

INVx1_ASAP7_75t_SL g1058 ( 
.A(n_699),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_722),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_945),
.Y(n_1060)
);

HB1xp67_ASAP7_75t_L g1061 ( 
.A(n_930),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_945),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_810),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_724),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_967),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_720),
.Y(n_1066)
);

INVx2_ASAP7_75t_SL g1067 ( 
.A(n_853),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_728),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_810),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_810),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_967),
.Y(n_1071)
);

HB1xp67_ASAP7_75t_L g1072 ( 
.A(n_696),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_731),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_810),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_733),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_735),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_982),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_982),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_736),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_810),
.Y(n_1080)
);

CKINVDCx14_ASAP7_75t_R g1081 ( 
.A(n_853),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1008),
.Y(n_1082)
);

INVxp67_ASAP7_75t_SL g1083 ( 
.A(n_740),
.Y(n_1083)
);

INVx2_ASAP7_75t_SL g1084 ( 
.A(n_853),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1008),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_740),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_758),
.Y(n_1087)
);

XOR2xp5_ASAP7_75t_L g1088 ( 
.A(n_803),
.B(n_822),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_739),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_740),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_742),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_740),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_775),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_775),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_775),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_775),
.Y(n_1096)
);

CKINVDCx20_ASAP7_75t_R g1097 ( 
.A(n_902),
.Y(n_1097)
);

INVx2_ASAP7_75t_SL g1098 ( 
.A(n_743),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_775),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_871),
.Y(n_1100)
);

CKINVDCx14_ASAP7_75t_R g1101 ( 
.A(n_858),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_871),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_748),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_751),
.Y(n_1104)
);

CKINVDCx20_ASAP7_75t_R g1105 ( 
.A(n_903),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_810),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_755),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_871),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_871),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_948),
.B(n_0),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_757),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_871),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_704),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_872),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_810),
.Y(n_1115)
);

CKINVDCx14_ASAP7_75t_R g1116 ( 
.A(n_858),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_758),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_810),
.Y(n_1118)
);

INVx3_ASAP7_75t_L g1119 ( 
.A(n_758),
.Y(n_1119)
);

HB1xp67_ASAP7_75t_L g1120 ( 
.A(n_713),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_872),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_872),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_759),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_872),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_761),
.Y(n_1125)
);

HB1xp67_ASAP7_75t_L g1126 ( 
.A(n_716),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_872),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_959),
.Y(n_1128)
);

INVxp67_ASAP7_75t_L g1129 ( 
.A(n_779),
.Y(n_1129)
);

INVxp67_ASAP7_75t_L g1130 ( 
.A(n_787),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_771),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_959),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_773),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_774),
.Y(n_1134)
);

BUFx10_ASAP7_75t_L g1135 ( 
.A(n_959),
.Y(n_1135)
);

BUFx8_ASAP7_75t_SL g1136 ( 
.A(n_744),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_959),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_959),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_743),
.Y(n_1139)
);

CKINVDCx20_ASAP7_75t_R g1140 ( 
.A(n_754),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_749),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_776),
.Y(n_1142)
);

INVxp67_ASAP7_75t_SL g1143 ( 
.A(n_812),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_749),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_769),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_777),
.Y(n_1146)
);

BUFx5_ASAP7_75t_L g1147 ( 
.A(n_694),
.Y(n_1147)
);

NOR2xp67_ASAP7_75t_L g1148 ( 
.A(n_1024),
.B(n_1),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_781),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_778),
.Y(n_1150)
);

CKINVDCx20_ASAP7_75t_R g1151 ( 
.A(n_791),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_769),
.Y(n_1152)
);

INVx1_ASAP7_75t_SL g1153 ( 
.A(n_802),
.Y(n_1153)
);

INVxp67_ASAP7_75t_SL g1154 ( 
.A(n_812),
.Y(n_1154)
);

INVx1_ASAP7_75t_SL g1155 ( 
.A(n_806),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_783),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_797),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_797),
.Y(n_1158)
);

CKINVDCx14_ASAP7_75t_R g1159 ( 
.A(n_858),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_785),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_790),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_794),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_840),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_840),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_988),
.Y(n_1165)
);

INVxp67_ASAP7_75t_SL g1166 ( 
.A(n_842),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_778),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_800),
.Y(n_1168)
);

BUFx2_ASAP7_75t_L g1169 ( 
.A(n_717),
.Y(n_1169)
);

BUFx5_ASAP7_75t_L g1170 ( 
.A(n_706),
.Y(n_1170)
);

CKINVDCx16_ASAP7_75t_R g1171 ( 
.A(n_906),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_988),
.Y(n_1172)
);

CKINVDCx14_ASAP7_75t_R g1173 ( 
.A(n_906),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_778),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_778),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_706),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_801),
.Y(n_1177)
);

CKINVDCx14_ASAP7_75t_R g1178 ( 
.A(n_906),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_709),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_778),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_811),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_867),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_709),
.Y(n_1183)
);

CKINVDCx20_ASAP7_75t_R g1184 ( 
.A(n_868),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_711),
.Y(n_1185)
);

CKINVDCx20_ASAP7_75t_R g1186 ( 
.A(n_882),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_711),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_734),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_734),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_813),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_741),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_741),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_745),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_745),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_767),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_767),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_815),
.Y(n_1197)
);

CKINVDCx16_ASAP7_75t_R g1198 ( 
.A(n_912),
.Y(n_1198)
);

INVxp67_ASAP7_75t_L g1199 ( 
.A(n_692),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_821),
.Y(n_1200)
);

BUFx2_ASAP7_75t_L g1201 ( 
.A(n_726),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_805),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_730),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_827),
.Y(n_1204)
);

CKINVDCx16_ASAP7_75t_R g1205 ( 
.A(n_912),
.Y(n_1205)
);

HB1xp67_ASAP7_75t_L g1206 ( 
.A(n_732),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_805),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_809),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_809),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_867),
.Y(n_1210)
);

CKINVDCx20_ASAP7_75t_R g1211 ( 
.A(n_886),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_823),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_823),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_837),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_828),
.Y(n_1215)
);

CKINVDCx14_ASAP7_75t_R g1216 ( 
.A(n_912),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_831),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_837),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_849),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_832),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_849),
.Y(n_1221)
);

BUFx2_ASAP7_75t_L g1222 ( 
.A(n_747),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_833),
.Y(n_1223)
);

BUFx6f_ASAP7_75t_L g1224 ( 
.A(n_867),
.Y(n_1224)
);

CKINVDCx20_ASAP7_75t_R g1225 ( 
.A(n_904),
.Y(n_1225)
);

CKINVDCx14_ASAP7_75t_R g1226 ( 
.A(n_966),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_880),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_880),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_838),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_839),
.Y(n_1230)
);

CKINVDCx20_ASAP7_75t_R g1231 ( 
.A(n_998),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_841),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_896),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_844),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_896),
.Y(n_1235)
);

CKINVDCx16_ASAP7_75t_R g1236 ( 
.A(n_966),
.Y(n_1236)
);

NOR2xp67_ASAP7_75t_L g1237 ( 
.A(n_965),
.B(n_1),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_845),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_848),
.Y(n_1239)
);

NOR2xp67_ASAP7_75t_L g1240 ( 
.A(n_965),
.B(n_1),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_851),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_925),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_856),
.Y(n_1243)
);

INVx1_ASAP7_75t_SL g1244 ( 
.A(n_756),
.Y(n_1244)
);

CKINVDCx16_ASAP7_75t_R g1245 ( 
.A(n_966),
.Y(n_1245)
);

INVxp67_ASAP7_75t_L g1246 ( 
.A(n_692),
.Y(n_1246)
);

INVxp67_ASAP7_75t_SL g1247 ( 
.A(n_842),
.Y(n_1247)
);

CKINVDCx16_ASAP7_75t_R g1248 ( 
.A(n_989),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_989),
.B(n_2),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_859),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_861),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_925),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_933),
.Y(n_1253)
);

OR2x2_ASAP7_75t_L g1254 ( 
.A(n_933),
.B(n_972),
.Y(n_1254)
);

INVxp67_ASAP7_75t_SL g1255 ( 
.A(n_846),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_869),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_949),
.Y(n_1257)
);

INVxp67_ASAP7_75t_SL g1258 ( 
.A(n_846),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_949),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_958),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_870),
.Y(n_1261)
);

INVx1_ASAP7_75t_SL g1262 ( 
.A(n_847),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_873),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_876),
.Y(n_1264)
);

INVxp67_ASAP7_75t_SL g1265 ( 
.A(n_958),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_877),
.Y(n_1266)
);

BUFx10_ASAP7_75t_L g1267 ( 
.A(n_867),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_972),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_883),
.Y(n_1269)
);

INVxp67_ASAP7_75t_L g1270 ( 
.A(n_695),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_884),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_973),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_885),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_973),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_990),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_990),
.Y(n_1276)
);

CKINVDCx20_ASAP7_75t_R g1277 ( 
.A(n_750),
.Y(n_1277)
);

CKINVDCx20_ASAP7_75t_R g1278 ( 
.A(n_762),
.Y(n_1278)
);

CKINVDCx20_ASAP7_75t_R g1279 ( 
.A(n_764),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_888),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1025),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_889),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_766),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1025),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_867),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_890),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_695),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_892),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_895),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_701),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_701),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_705),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_897),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_705),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_898),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1022),
.Y(n_1296)
);

INVxp33_ASAP7_75t_SL g1297 ( 
.A(n_768),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_707),
.Y(n_1298)
);

INVx1_ASAP7_75t_SL g1299 ( 
.A(n_702),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_707),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_708),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_901),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_907),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_908),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1022),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_708),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_909),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_712),
.Y(n_1308)
);

BUFx2_ASAP7_75t_SL g1309 ( 
.A(n_1022),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_913),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_712),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_715),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_715),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_914),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_915),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1022),
.Y(n_1316)
);

BUFx3_ASAP7_75t_L g1317 ( 
.A(n_1022),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_721),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_721),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_723),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_916),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_919),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_723),
.Y(n_1323)
);

NOR2xp67_ASAP7_75t_L g1324 ( 
.A(n_697),
.B(n_3),
.Y(n_1324)
);

INVx1_ASAP7_75t_SL g1325 ( 
.A(n_737),
.Y(n_1325)
);

INVxp67_ASAP7_75t_L g1326 ( 
.A(n_725),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_920),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_927),
.Y(n_1328)
);

CKINVDCx20_ASAP7_75t_R g1329 ( 
.A(n_772),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_929),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_931),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_937),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_939),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_725),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_727),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_L g1336 ( 
.A(n_697),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_727),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_780),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_940),
.Y(n_1339)
);

CKINVDCx20_ASAP7_75t_R g1340 ( 
.A(n_788),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_746),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_746),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_752),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_752),
.Y(n_1344)
);

BUFx5_ASAP7_75t_L g1345 ( 
.A(n_760),
.Y(n_1345)
);

INVx1_ASAP7_75t_SL g1346 ( 
.A(n_782),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_941),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_943),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_944),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_714),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_714),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_951),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_952),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_760),
.Y(n_1354)
);

BUFx3_ASAP7_75t_L g1355 ( 
.A(n_784),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_763),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_763),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_729),
.Y(n_1358)
);

BUFx3_ASAP7_75t_L g1359 ( 
.A(n_792),
.Y(n_1359)
);

BUFx3_ASAP7_75t_L g1360 ( 
.A(n_793),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_729),
.Y(n_1361)
);

INVxp67_ASAP7_75t_L g1362 ( 
.A(n_770),
.Y(n_1362)
);

CKINVDCx20_ASAP7_75t_R g1363 ( 
.A(n_789),
.Y(n_1363)
);

CKINVDCx20_ASAP7_75t_R g1364 ( 
.A(n_796),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_953),
.Y(n_1365)
);

BUFx2_ASAP7_75t_L g1366 ( 
.A(n_799),
.Y(n_1366)
);

INVxp67_ASAP7_75t_L g1367 ( 
.A(n_770),
.Y(n_1367)
);

CKINVDCx20_ASAP7_75t_R g1368 ( 
.A(n_804),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_960),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_807),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_786),
.Y(n_1371)
);

INVx2_ASAP7_75t_SL g1372 ( 
.A(n_786),
.Y(n_1372)
);

INVx1_ASAP7_75t_SL g1373 ( 
.A(n_798),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_807),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_808),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_808),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_962),
.Y(n_1377)
);

CKINVDCx16_ASAP7_75t_R g1378 ( 
.A(n_922),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_963),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_964),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_878),
.B(n_3),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_814),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_814),
.Y(n_1383)
);

INVxp67_ASAP7_75t_L g1384 ( 
.A(n_817),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_817),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_818),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_968),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_969),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_818),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_819),
.Y(n_1390)
);

BUFx3_ASAP7_75t_L g1391 ( 
.A(n_795),
.Y(n_1391)
);

CKINVDCx20_ASAP7_75t_R g1392 ( 
.A(n_816),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1083),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1035),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1036),
.Y(n_1395)
);

INVxp67_ASAP7_75t_SL g1396 ( 
.A(n_1063),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1031),
.B(n_825),
.Y(n_1397)
);

CKINVDCx20_ASAP7_75t_R g1398 ( 
.A(n_1034),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1039),
.Y(n_1399)
);

NOR2xp67_ASAP7_75t_L g1400 ( 
.A(n_1125),
.B(n_970),
.Y(n_1400)
);

INVxp67_ASAP7_75t_SL g1401 ( 
.A(n_1063),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1244),
.B(n_878),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_1031),
.B(n_826),
.Y(n_1403)
);

NOR2xp67_ASAP7_75t_L g1404 ( 
.A(n_1131),
.B(n_971),
.Y(n_1404)
);

CKINVDCx20_ASAP7_75t_R g1405 ( 
.A(n_1034),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_1136),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1058),
.Y(n_1407)
);

CKINVDCx20_ASAP7_75t_R g1408 ( 
.A(n_1054),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1040),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_1153),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1041),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1042),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_1155),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1143),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_1133),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1154),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1166),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_1134),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1247),
.Y(n_1419)
);

OR2x2_ASAP7_75t_L g1420 ( 
.A(n_1262),
.B(n_819),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_1142),
.Y(n_1421)
);

CKINVDCx20_ASAP7_75t_R g1422 ( 
.A(n_1054),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1255),
.Y(n_1423)
);

INVxp67_ASAP7_75t_SL g1424 ( 
.A(n_1174),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1258),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1265),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_1146),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1060),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1062),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1065),
.Y(n_1430)
);

INVxp67_ASAP7_75t_L g1431 ( 
.A(n_1299),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1071),
.Y(n_1432)
);

INVxp67_ASAP7_75t_L g1433 ( 
.A(n_1325),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1077),
.Y(n_1434)
);

CKINVDCx20_ASAP7_75t_R g1435 ( 
.A(n_1066),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1078),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1082),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1085),
.Y(n_1438)
);

INVxp67_ASAP7_75t_SL g1439 ( 
.A(n_1174),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1149),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_1156),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1287),
.Y(n_1442)
);

INVxp67_ASAP7_75t_L g1443 ( 
.A(n_1346),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1290),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1291),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_1160),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_1161),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_1197),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1292),
.Y(n_1449)
);

NOR2xp67_ASAP7_75t_L g1450 ( 
.A(n_1204),
.B(n_976),
.Y(n_1450)
);

CKINVDCx20_ASAP7_75t_R g1451 ( 
.A(n_1066),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_1215),
.Y(n_1452)
);

INVxp67_ASAP7_75t_SL g1453 ( 
.A(n_1182),
.Y(n_1453)
);

INVxp67_ASAP7_75t_SL g1454 ( 
.A(n_1182),
.Y(n_1454)
);

INVxp67_ASAP7_75t_SL g1455 ( 
.A(n_1317),
.Y(n_1455)
);

CKINVDCx20_ASAP7_75t_R g1456 ( 
.A(n_1097),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_1248),
.B(n_829),
.Y(n_1457)
);

CKINVDCx16_ASAP7_75t_R g1458 ( 
.A(n_1048),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_1217),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_1220),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1294),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1298),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_1223),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1373),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1300),
.Y(n_1465)
);

CKINVDCx20_ASAP7_75t_R g1466 ( 
.A(n_1097),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_1229),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1301),
.Y(n_1468)
);

CKINVDCx16_ASAP7_75t_R g1469 ( 
.A(n_1171),
.Y(n_1469)
);

CKINVDCx20_ASAP7_75t_R g1470 ( 
.A(n_1105),
.Y(n_1470)
);

CKINVDCx20_ASAP7_75t_R g1471 ( 
.A(n_1105),
.Y(n_1471)
);

CKINVDCx20_ASAP7_75t_R g1472 ( 
.A(n_1140),
.Y(n_1472)
);

CKINVDCx16_ASAP7_75t_R g1473 ( 
.A(n_1198),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1230),
.Y(n_1474)
);

CKINVDCx20_ASAP7_75t_R g1475 ( 
.A(n_1140),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1306),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_1232),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1308),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1311),
.Y(n_1479)
);

CKINVDCx20_ASAP7_75t_R g1480 ( 
.A(n_1151),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1312),
.Y(n_1481)
);

CKINVDCx20_ASAP7_75t_R g1482 ( 
.A(n_1151),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1313),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_1234),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1081),
.B(n_1101),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_1238),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1318),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_1239),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_1241),
.Y(n_1489)
);

CKINVDCx20_ASAP7_75t_R g1490 ( 
.A(n_1184),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1319),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1320),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_1243),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1323),
.Y(n_1494)
);

INVxp67_ASAP7_75t_SL g1495 ( 
.A(n_1317),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1297),
.B(n_850),
.Y(n_1496)
);

CKINVDCx20_ASAP7_75t_R g1497 ( 
.A(n_1184),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1334),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1061),
.Y(n_1499)
);

INVxp67_ASAP7_75t_L g1500 ( 
.A(n_1113),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1335),
.Y(n_1501)
);

INVxp67_ASAP7_75t_L g1502 ( 
.A(n_1169),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1337),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1341),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1342),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_1250),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1297),
.B(n_855),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1343),
.Y(n_1508)
);

INVxp67_ASAP7_75t_L g1509 ( 
.A(n_1201),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1344),
.Y(n_1510)
);

CKINVDCx20_ASAP7_75t_R g1511 ( 
.A(n_1186),
.Y(n_1511)
);

CKINVDCx16_ASAP7_75t_R g1512 ( 
.A(n_1205),
.Y(n_1512)
);

CKINVDCx20_ASAP7_75t_R g1513 ( 
.A(n_1186),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_1251),
.Y(n_1514)
);

CKINVDCx16_ASAP7_75t_R g1515 ( 
.A(n_1236),
.Y(n_1515)
);

CKINVDCx20_ASAP7_75t_R g1516 ( 
.A(n_1211),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1354),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1356),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_1256),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1357),
.Y(n_1520)
);

CKINVDCx20_ASAP7_75t_R g1521 ( 
.A(n_1211),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1370),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1374),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1098),
.B(n_1014),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_1261),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1375),
.Y(n_1526)
);

NOR2xp67_ASAP7_75t_L g1527 ( 
.A(n_1263),
.B(n_977),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1033),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1376),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1382),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_1264),
.Y(n_1531)
);

CKINVDCx20_ASAP7_75t_R g1532 ( 
.A(n_1225),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1383),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1385),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_1387),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_1037),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_1037),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1386),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_1038),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1389),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1067),
.B(n_857),
.Y(n_1541)
);

NOR2xp67_ASAP7_75t_L g1542 ( 
.A(n_1030),
.B(n_980),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1390),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_1038),
.Y(n_1544)
);

CKINVDCx20_ASAP7_75t_R g1545 ( 
.A(n_1225),
.Y(n_1545)
);

NOR2xp67_ASAP7_75t_L g1546 ( 
.A(n_1047),
.B(n_1052),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_1047),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1029),
.Y(n_1548)
);

BUFx3_ASAP7_75t_L g1549 ( 
.A(n_1267),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1029),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1029),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_1052),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_1056),
.Y(n_1553)
);

CKINVDCx20_ASAP7_75t_R g1554 ( 
.A(n_1231),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1135),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1135),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1135),
.Y(n_1557)
);

BUFx3_ASAP7_75t_L g1558 ( 
.A(n_1267),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_1056),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1043),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1044),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1049),
.Y(n_1562)
);

BUFx2_ASAP7_75t_SL g1563 ( 
.A(n_1277),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_1059),
.Y(n_1564)
);

CKINVDCx20_ASAP7_75t_R g1565 ( 
.A(n_1231),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1051),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_1059),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1067),
.B(n_863),
.Y(n_1568)
);

CKINVDCx20_ASAP7_75t_R g1569 ( 
.A(n_1277),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_1064),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1053),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1055),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_1064),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_1068),
.Y(n_1574)
);

BUFx2_ASAP7_75t_L g1575 ( 
.A(n_1278),
.Y(n_1575)
);

CKINVDCx20_ASAP7_75t_R g1576 ( 
.A(n_1278),
.Y(n_1576)
);

INVxp33_ASAP7_75t_SL g1577 ( 
.A(n_1033),
.Y(n_1577)
);

INVxp67_ASAP7_75t_L g1578 ( 
.A(n_1203),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1057),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1176),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1179),
.Y(n_1581)
);

CKINVDCx20_ASAP7_75t_R g1582 ( 
.A(n_1279),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1032),
.Y(n_1583)
);

BUFx6f_ASAP7_75t_L g1584 ( 
.A(n_1032),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1183),
.Y(n_1585)
);

INVxp67_ASAP7_75t_SL g1586 ( 
.A(n_1119),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_1116),
.Y(n_1587)
);

INVxp33_ASAP7_75t_L g1588 ( 
.A(n_1088),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1032),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1185),
.Y(n_1590)
);

CKINVDCx20_ASAP7_75t_R g1591 ( 
.A(n_1279),
.Y(n_1591)
);

CKINVDCx20_ASAP7_75t_R g1592 ( 
.A(n_1329),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1159),
.Y(n_1593)
);

HB1xp67_ASAP7_75t_L g1594 ( 
.A(n_1329),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_1173),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_1178),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1187),
.Y(n_1597)
);

HB1xp67_ASAP7_75t_L g1598 ( 
.A(n_1340),
.Y(n_1598)
);

CKINVDCx20_ASAP7_75t_R g1599 ( 
.A(n_1340),
.Y(n_1599)
);

INVxp67_ASAP7_75t_SL g1600 ( 
.A(n_1119),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_1216),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_1226),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1188),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1189),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1191),
.Y(n_1605)
);

CKINVDCx20_ASAP7_75t_R g1606 ( 
.A(n_1363),
.Y(n_1606)
);

CKINVDCx20_ASAP7_75t_R g1607 ( 
.A(n_1363),
.Y(n_1607)
);

BUFx6f_ASAP7_75t_L g1608 ( 
.A(n_1032),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_1378),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_1068),
.Y(n_1610)
);

CKINVDCx20_ASAP7_75t_R g1611 ( 
.A(n_1364),
.Y(n_1611)
);

NOR2xp67_ASAP7_75t_L g1612 ( 
.A(n_1073),
.B(n_983),
.Y(n_1612)
);

INVxp67_ASAP7_75t_SL g1613 ( 
.A(n_1119),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1192),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1364),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1193),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1194),
.Y(n_1617)
);

CKINVDCx20_ASAP7_75t_R g1618 ( 
.A(n_1368),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1195),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_1073),
.Y(n_1620)
);

BUFx2_ASAP7_75t_SL g1621 ( 
.A(n_1368),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1196),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1084),
.B(n_881),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1098),
.B(n_1026),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1084),
.B(n_1139),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_1075),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_1075),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1202),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_1076),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1207),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1208),
.Y(n_1631)
);

CKINVDCx16_ASAP7_75t_R g1632 ( 
.A(n_1245),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_1076),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1209),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1032),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_1079),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_1079),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1089),
.Y(n_1638)
);

INVxp67_ASAP7_75t_L g1639 ( 
.A(n_1222),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1212),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1213),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1214),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1218),
.Y(n_1643)
);

CKINVDCx20_ASAP7_75t_R g1644 ( 
.A(n_1392),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1219),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1221),
.Y(n_1646)
);

BUFx2_ASAP7_75t_L g1647 ( 
.A(n_1392),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1089),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1227),
.Y(n_1649)
);

CKINVDCx16_ASAP7_75t_R g1650 ( 
.A(n_1072),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1228),
.Y(n_1651)
);

CKINVDCx20_ASAP7_75t_R g1652 ( 
.A(n_1091),
.Y(n_1652)
);

CKINVDCx20_ASAP7_75t_R g1653 ( 
.A(n_1091),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_1103),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_1103),
.Y(n_1655)
);

INVxp33_ASAP7_75t_L g1656 ( 
.A(n_1120),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1233),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1283),
.B(n_900),
.Y(n_1658)
);

HB1xp67_ASAP7_75t_L g1659 ( 
.A(n_1104),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1235),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1104),
.B(n_894),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1242),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_1107),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1252),
.Y(n_1664)
);

INVxp67_ASAP7_75t_SL g1665 ( 
.A(n_1050),
.Y(n_1665)
);

BUFx2_ASAP7_75t_SL g1666 ( 
.A(n_1267),
.Y(n_1666)
);

CKINVDCx20_ASAP7_75t_R g1667 ( 
.A(n_1107),
.Y(n_1667)
);

INVxp67_ASAP7_75t_L g1668 ( 
.A(n_1366),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_1111),
.Y(n_1669)
);

NAND2xp33_ASAP7_75t_R g1670 ( 
.A(n_1111),
.B(n_911),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1253),
.Y(n_1671)
);

INVxp67_ASAP7_75t_L g1672 ( 
.A(n_1126),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1257),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1259),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1260),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_L g1676 ( 
.A(n_1123),
.B(n_921),
.Y(n_1676)
);

CKINVDCx20_ASAP7_75t_R g1677 ( 
.A(n_1123),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_1162),
.Y(n_1678)
);

INVxp67_ASAP7_75t_L g1679 ( 
.A(n_1206),
.Y(n_1679)
);

CKINVDCx20_ASAP7_75t_R g1680 ( 
.A(n_1162),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1268),
.Y(n_1681)
);

CKINVDCx20_ASAP7_75t_R g1682 ( 
.A(n_1168),
.Y(n_1682)
);

INVxp67_ASAP7_75t_SL g1683 ( 
.A(n_1050),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1272),
.Y(n_1684)
);

INVxp67_ASAP7_75t_SL g1685 ( 
.A(n_1050),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1274),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1168),
.B(n_928),
.Y(n_1687)
);

CKINVDCx20_ASAP7_75t_R g1688 ( 
.A(n_1177),
.Y(n_1688)
);

INVxp67_ASAP7_75t_SL g1689 ( 
.A(n_1050),
.Y(n_1689)
);

NOR2xp67_ASAP7_75t_L g1690 ( 
.A(n_1177),
.B(n_984),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_1181),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_1181),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1275),
.Y(n_1693)
);

INVxp67_ASAP7_75t_L g1694 ( 
.A(n_1338),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1141),
.B(n_1010),
.Y(n_1695)
);

CKINVDCx16_ASAP7_75t_R g1696 ( 
.A(n_1355),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1050),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1276),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1281),
.Y(n_1699)
);

INVx3_ASAP7_75t_L g1700 ( 
.A(n_1584),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1666),
.B(n_1046),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1426),
.B(n_1355),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1428),
.Y(n_1703)
);

HB1xp67_ASAP7_75t_L g1704 ( 
.A(n_1464),
.Y(n_1704)
);

OA21x2_ASAP7_75t_L g1705 ( 
.A1(n_1560),
.A2(n_1045),
.B(n_1069),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1561),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1429),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1430),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1432),
.Y(n_1709)
);

OAI22x1_ASAP7_75t_R g1710 ( 
.A1(n_1569),
.A2(n_1377),
.B1(n_1379),
.B2(n_1369),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1402),
.B(n_1359),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1562),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1434),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1436),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1586),
.B(n_1046),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1696),
.B(n_1658),
.Y(n_1716)
);

BUFx6f_ASAP7_75t_L g1717 ( 
.A(n_1584),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1566),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1437),
.Y(n_1719)
);

CKINVDCx5p33_ASAP7_75t_R g1720 ( 
.A(n_1427),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1431),
.B(n_1359),
.Y(n_1721)
);

OA21x2_ASAP7_75t_L g1722 ( 
.A1(n_1571),
.A2(n_1045),
.B(n_1069),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1438),
.Y(n_1723)
);

BUFx6f_ASAP7_75t_L g1724 ( 
.A(n_1584),
.Y(n_1724)
);

NAND2xp33_ASAP7_75t_L g1725 ( 
.A(n_1427),
.B(n_1046),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1433),
.B(n_1360),
.Y(n_1726)
);

AND2x4_ASAP7_75t_L g1727 ( 
.A(n_1414),
.B(n_1360),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1572),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1548),
.B(n_1190),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1416),
.B(n_1391),
.Y(n_1730)
);

INVx6_ASAP7_75t_L g1731 ( 
.A(n_1549),
.Y(n_1731)
);

AOI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1496),
.A2(n_1110),
.B1(n_1200),
.B2(n_1190),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1579),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1394),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1583),
.Y(n_1735)
);

CKINVDCx20_ASAP7_75t_R g1736 ( 
.A(n_1398),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1395),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1443),
.B(n_1391),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1420),
.B(n_1442),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1499),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1399),
.Y(n_1741)
);

BUFx6f_ASAP7_75t_L g1742 ( 
.A(n_1584),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1409),
.Y(n_1743)
);

CKINVDCx20_ASAP7_75t_R g1744 ( 
.A(n_1398),
.Y(n_1744)
);

BUFx8_ASAP7_75t_L g1745 ( 
.A(n_1575),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_SL g1746 ( 
.A(n_1507),
.B(n_1046),
.Y(n_1746)
);

INVx5_ASAP7_75t_L g1747 ( 
.A(n_1584),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1600),
.B(n_1046),
.Y(n_1748)
);

CKINVDCx8_ASAP7_75t_R g1749 ( 
.A(n_1563),
.Y(n_1749)
);

AND2x4_ASAP7_75t_L g1750 ( 
.A(n_1417),
.B(n_1237),
.Y(n_1750)
);

BUFx6f_ASAP7_75t_L g1751 ( 
.A(n_1608),
.Y(n_1751)
);

BUFx2_ASAP7_75t_L g1752 ( 
.A(n_1609),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1613),
.B(n_1046),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1650),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_1440),
.Y(n_1755)
);

BUFx6f_ASAP7_75t_L g1756 ( 
.A(n_1608),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1583),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1393),
.B(n_1046),
.Y(n_1758)
);

INVx3_ASAP7_75t_L g1759 ( 
.A(n_1608),
.Y(n_1759)
);

INVxp33_ASAP7_75t_SL g1760 ( 
.A(n_1440),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1589),
.Y(n_1761)
);

AOI22x1_ASAP7_75t_SL g1762 ( 
.A1(n_1569),
.A2(n_947),
.B1(n_950),
.B2(n_936),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_1441),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1550),
.B(n_1147),
.Y(n_1764)
);

BUFx6f_ASAP7_75t_L g1765 ( 
.A(n_1608),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1411),
.Y(n_1766)
);

INVx6_ASAP7_75t_L g1767 ( 
.A(n_1549),
.Y(n_1767)
);

INVx3_ASAP7_75t_L g1768 ( 
.A(n_1608),
.Y(n_1768)
);

CKINVDCx5p33_ASAP7_75t_R g1769 ( 
.A(n_1441),
.Y(n_1769)
);

BUFx2_ASAP7_75t_L g1770 ( 
.A(n_1609),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1551),
.B(n_1147),
.Y(n_1771)
);

BUFx2_ASAP7_75t_L g1772 ( 
.A(n_1652),
.Y(n_1772)
);

OA21x2_ASAP7_75t_L g1773 ( 
.A1(n_1665),
.A2(n_1074),
.B(n_1070),
.Y(n_1773)
);

BUFx6f_ASAP7_75t_L g1774 ( 
.A(n_1589),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1635),
.Y(n_1775)
);

AND2x4_ASAP7_75t_L g1776 ( 
.A(n_1419),
.B(n_1240),
.Y(n_1776)
);

XNOR2x1_ASAP7_75t_L g1777 ( 
.A(n_1407),
.B(n_1200),
.Y(n_1777)
);

AOI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1541),
.A2(n_1266),
.B1(n_1271),
.B2(n_1269),
.Y(n_1778)
);

OA21x2_ASAP7_75t_L g1779 ( 
.A1(n_1683),
.A2(n_1074),
.B(n_1070),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1412),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1635),
.Y(n_1781)
);

CKINVDCx5p33_ASAP7_75t_R g1782 ( 
.A(n_1446),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1444),
.Y(n_1783)
);

BUFx2_ASAP7_75t_L g1784 ( 
.A(n_1500),
.Y(n_1784)
);

INVx3_ASAP7_75t_L g1785 ( 
.A(n_1697),
.Y(n_1785)
);

AND2x4_ASAP7_75t_L g1786 ( 
.A(n_1423),
.B(n_1367),
.Y(n_1786)
);

AND2x4_ASAP7_75t_L g1787 ( 
.A(n_1425),
.B(n_1384),
.Y(n_1787)
);

AND2x4_ASAP7_75t_L g1788 ( 
.A(n_1625),
.B(n_1199),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1555),
.B(n_1266),
.Y(n_1789)
);

BUFx6f_ASAP7_75t_L g1790 ( 
.A(n_1697),
.Y(n_1790)
);

BUFx2_ASAP7_75t_L g1791 ( 
.A(n_1502),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1556),
.B(n_1147),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1557),
.B(n_1568),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1623),
.B(n_1147),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1558),
.B(n_1147),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1445),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1449),
.B(n_1144),
.Y(n_1797)
);

INVx3_ASAP7_75t_L g1798 ( 
.A(n_1558),
.Y(n_1798)
);

OAI21x1_ASAP7_75t_L g1799 ( 
.A1(n_1685),
.A2(n_1106),
.B(n_1080),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1424),
.B(n_1147),
.Y(n_1800)
);

BUFx6f_ASAP7_75t_L g1801 ( 
.A(n_1699),
.Y(n_1801)
);

INVx3_ASAP7_75t_L g1802 ( 
.A(n_1580),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1461),
.Y(n_1803)
);

OAI22xp5_ASAP7_75t_L g1804 ( 
.A1(n_1457),
.A2(n_1148),
.B1(n_961),
.B2(n_978),
.Y(n_1804)
);

AND2x4_ASAP7_75t_L g1805 ( 
.A(n_1462),
.B(n_1246),
.Y(n_1805)
);

AND2x4_ASAP7_75t_L g1806 ( 
.A(n_1465),
.B(n_1270),
.Y(n_1806)
);

INVx3_ASAP7_75t_L g1807 ( 
.A(n_1581),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_1446),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1468),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1585),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1476),
.B(n_1145),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1478),
.Y(n_1812)
);

AND2x4_ASAP7_75t_L g1813 ( 
.A(n_1479),
.B(n_1326),
.Y(n_1813)
);

NOR2x1_ASAP7_75t_L g1814 ( 
.A(n_1546),
.B(n_1254),
.Y(n_1814)
);

AND2x4_ASAP7_75t_L g1815 ( 
.A(n_1481),
.B(n_1362),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1483),
.Y(n_1816)
);

BUFx2_ASAP7_75t_L g1817 ( 
.A(n_1652),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1487),
.Y(n_1818)
);

CKINVDCx20_ASAP7_75t_R g1819 ( 
.A(n_1405),
.Y(n_1819)
);

AND2x4_ASAP7_75t_L g1820 ( 
.A(n_1491),
.B(n_1381),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1590),
.Y(n_1821)
);

AOI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1661),
.A2(n_1269),
.B1(n_1273),
.B2(n_1271),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1492),
.Y(n_1823)
);

AND2x4_ASAP7_75t_L g1824 ( 
.A(n_1494),
.B(n_1129),
.Y(n_1824)
);

AND2x4_ASAP7_75t_L g1825 ( 
.A(n_1498),
.B(n_1130),
.Y(n_1825)
);

INVx4_ASAP7_75t_L g1826 ( 
.A(n_1415),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1439),
.B(n_1147),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1501),
.Y(n_1828)
);

BUFx12f_ASAP7_75t_L g1829 ( 
.A(n_1406),
.Y(n_1829)
);

CKINVDCx20_ASAP7_75t_R g1830 ( 
.A(n_1405),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_SL g1831 ( 
.A(n_1587),
.B(n_1273),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1503),
.Y(n_1832)
);

AND2x6_ASAP7_75t_L g1833 ( 
.A(n_1485),
.B(n_1249),
.Y(n_1833)
);

OAI22xp5_ASAP7_75t_SL g1834 ( 
.A1(n_1576),
.A2(n_1280),
.B1(n_1286),
.B2(n_1282),
.Y(n_1834)
);

INVx4_ASAP7_75t_L g1835 ( 
.A(n_1418),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1597),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_SL g1837 ( 
.A(n_1676),
.B(n_1170),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1603),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1604),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1504),
.Y(n_1840)
);

BUFx2_ASAP7_75t_L g1841 ( 
.A(n_1653),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1505),
.Y(n_1842)
);

CKINVDCx5p33_ASAP7_75t_R g1843 ( 
.A(n_1447),
.Y(n_1843)
);

BUFx6f_ASAP7_75t_L g1844 ( 
.A(n_1698),
.Y(n_1844)
);

AND2x4_ASAP7_75t_L g1845 ( 
.A(n_1508),
.B(n_1152),
.Y(n_1845)
);

INVx3_ASAP7_75t_L g1846 ( 
.A(n_1605),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1614),
.Y(n_1847)
);

INVx3_ASAP7_75t_L g1848 ( 
.A(n_1616),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_L g1849 ( 
.A(n_1397),
.B(n_1280),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1617),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1619),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1510),
.B(n_1157),
.Y(n_1852)
);

HB1xp67_ASAP7_75t_L g1853 ( 
.A(n_1458),
.Y(n_1853)
);

HB1xp67_ASAP7_75t_L g1854 ( 
.A(n_1509),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_SL g1855 ( 
.A(n_1687),
.B(n_1170),
.Y(n_1855)
);

BUFx6f_ASAP7_75t_L g1856 ( 
.A(n_1622),
.Y(n_1856)
);

BUFx6f_ASAP7_75t_L g1857 ( 
.A(n_1628),
.Y(n_1857)
);

INVxp67_ASAP7_75t_L g1858 ( 
.A(n_1670),
.Y(n_1858)
);

INVx3_ASAP7_75t_L g1859 ( 
.A(n_1630),
.Y(n_1859)
);

BUFx2_ASAP7_75t_L g1860 ( 
.A(n_1653),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1631),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1453),
.B(n_1170),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_SL g1863 ( 
.A(n_1447),
.B(n_1448),
.Y(n_1863)
);

OAI22xp5_ASAP7_75t_SL g1864 ( 
.A1(n_1576),
.A2(n_1282),
.B1(n_1288),
.B2(n_1286),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1634),
.Y(n_1865)
);

BUFx6f_ASAP7_75t_L g1866 ( 
.A(n_1640),
.Y(n_1866)
);

BUFx3_ASAP7_75t_L g1867 ( 
.A(n_1421),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_SL g1868 ( 
.A(n_1448),
.B(n_1452),
.Y(n_1868)
);

OAI22xp5_ASAP7_75t_SL g1869 ( 
.A1(n_1582),
.A2(n_1288),
.B1(n_1293),
.B2(n_1289),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1454),
.B(n_1170),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1517),
.Y(n_1871)
);

AND2x4_ASAP7_75t_L g1872 ( 
.A(n_1518),
.B(n_1158),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1455),
.B(n_1170),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1641),
.Y(n_1874)
);

OAI21x1_ASAP7_75t_L g1875 ( 
.A1(n_1689),
.A2(n_1106),
.B(n_1080),
.Y(n_1875)
);

NOR2x1_ASAP7_75t_L g1876 ( 
.A(n_1400),
.B(n_1163),
.Y(n_1876)
);

BUFx8_ASAP7_75t_L g1877 ( 
.A(n_1647),
.Y(n_1877)
);

XNOR2xp5_ASAP7_75t_L g1878 ( 
.A(n_1582),
.B(n_1289),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1642),
.Y(n_1879)
);

INVx3_ASAP7_75t_L g1880 ( 
.A(n_1643),
.Y(n_1880)
);

BUFx12f_ASAP7_75t_L g1881 ( 
.A(n_1587),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1495),
.B(n_1170),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1520),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1522),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1396),
.B(n_1170),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1645),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1523),
.Y(n_1887)
);

INVx4_ASAP7_75t_L g1888 ( 
.A(n_1474),
.Y(n_1888)
);

NOR2xp67_ASAP7_75t_L g1889 ( 
.A(n_1593),
.B(n_1293),
.Y(n_1889)
);

OAI22xp5_ASAP7_75t_SL g1890 ( 
.A1(n_1591),
.A2(n_1295),
.B1(n_1303),
.B2(n_1302),
.Y(n_1890)
);

BUFx6f_ASAP7_75t_L g1891 ( 
.A(n_1646),
.Y(n_1891)
);

AND2x4_ASAP7_75t_L g1892 ( 
.A(n_1526),
.B(n_1529),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1401),
.B(n_1649),
.Y(n_1893)
);

HB1xp67_ASAP7_75t_L g1894 ( 
.A(n_1578),
.Y(n_1894)
);

BUFx2_ASAP7_75t_L g1895 ( 
.A(n_1639),
.Y(n_1895)
);

BUFx6f_ASAP7_75t_L g1896 ( 
.A(n_1651),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1657),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1530),
.B(n_1164),
.Y(n_1898)
);

OAI22xp5_ASAP7_75t_R g1899 ( 
.A1(n_1577),
.A2(n_1302),
.B1(n_1303),
.B2(n_1295),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1533),
.B(n_1165),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1660),
.Y(n_1901)
);

OAI22xp5_ASAP7_75t_SL g1902 ( 
.A1(n_1591),
.A2(n_1304),
.B1(n_1310),
.B2(n_1307),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1662),
.B(n_1309),
.Y(n_1903)
);

BUFx6f_ASAP7_75t_L g1904 ( 
.A(n_1664),
.Y(n_1904)
);

CKINVDCx5p33_ASAP7_75t_R g1905 ( 
.A(n_1452),
.Y(n_1905)
);

BUFx3_ASAP7_75t_L g1906 ( 
.A(n_1477),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1534),
.Y(n_1907)
);

AOI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1672),
.A2(n_1307),
.B1(n_1310),
.B2(n_1304),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1671),
.B(n_1345),
.Y(n_1909)
);

BUFx3_ASAP7_75t_L g1910 ( 
.A(n_1484),
.Y(n_1910)
);

INVx2_ASAP7_75t_SL g1911 ( 
.A(n_1524),
.Y(n_1911)
);

BUFx6f_ASAP7_75t_L g1912 ( 
.A(n_1673),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1674),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1538),
.Y(n_1914)
);

CKINVDCx16_ASAP7_75t_R g1915 ( 
.A(n_1469),
.Y(n_1915)
);

INVx5_ASAP7_75t_L g1916 ( 
.A(n_1473),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1675),
.B(n_1345),
.Y(n_1917)
);

HB1xp67_ASAP7_75t_L g1918 ( 
.A(n_1668),
.Y(n_1918)
);

INVx5_ASAP7_75t_L g1919 ( 
.A(n_1512),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1540),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1681),
.B(n_1345),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1543),
.B(n_1172),
.Y(n_1922)
);

INVx5_ASAP7_75t_L g1923 ( 
.A(n_1515),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1684),
.Y(n_1924)
);

AOI22xp5_ASAP7_75t_L g1925 ( 
.A1(n_1679),
.A2(n_1315),
.B1(n_1321),
.B2(n_1314),
.Y(n_1925)
);

BUFx6f_ASAP7_75t_L g1926 ( 
.A(n_1686),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1693),
.B(n_1350),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1656),
.B(n_1350),
.Y(n_1928)
);

NOR2xp33_ASAP7_75t_L g1929 ( 
.A(n_1403),
.B(n_1314),
.Y(n_1929)
);

BUFx6f_ASAP7_75t_L g1930 ( 
.A(n_1695),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1624),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1612),
.Y(n_1932)
);

BUFx3_ASAP7_75t_L g1933 ( 
.A(n_1486),
.Y(n_1933)
);

INVx3_ASAP7_75t_L g1934 ( 
.A(n_1488),
.Y(n_1934)
);

AND2x4_ASAP7_75t_L g1935 ( 
.A(n_1690),
.B(n_1324),
.Y(n_1935)
);

INVxp67_ASAP7_75t_L g1936 ( 
.A(n_1410),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1404),
.Y(n_1937)
);

BUFx12f_ASAP7_75t_L g1938 ( 
.A(n_1593),
.Y(n_1938)
);

BUFx6f_ASAP7_75t_L g1939 ( 
.A(n_1489),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1694),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1659),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1493),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1450),
.Y(n_1943)
);

BUFx6f_ASAP7_75t_L g1944 ( 
.A(n_1506),
.Y(n_1944)
);

BUFx6f_ASAP7_75t_L g1945 ( 
.A(n_1519),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1525),
.Y(n_1946)
);

BUFx6f_ASAP7_75t_L g1947 ( 
.A(n_1531),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1527),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1535),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1542),
.Y(n_1950)
);

INVx2_ASAP7_75t_SL g1951 ( 
.A(n_1459),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1459),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1460),
.B(n_1345),
.Y(n_1953)
);

BUFx2_ASAP7_75t_L g1954 ( 
.A(n_1667),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1460),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1463),
.Y(n_1956)
);

OAI22xp5_ASAP7_75t_L g1957 ( 
.A1(n_1610),
.A2(n_979),
.B1(n_985),
.B2(n_957),
.Y(n_1957)
);

OA21x2_ASAP7_75t_L g1958 ( 
.A1(n_1610),
.A2(n_1118),
.B(n_1115),
.Y(n_1958)
);

AOI22xp5_ASAP7_75t_L g1959 ( 
.A1(n_1463),
.A2(n_1321),
.B1(n_1322),
.B2(n_1315),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1467),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_SL g1961 ( 
.A(n_1467),
.B(n_1345),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1514),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1514),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1536),
.B(n_1345),
.Y(n_1964)
);

BUFx6f_ASAP7_75t_L g1965 ( 
.A(n_1537),
.Y(n_1965)
);

OAI21x1_ASAP7_75t_L g1966 ( 
.A1(n_1528),
.A2(n_1118),
.B(n_1115),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1539),
.Y(n_1967)
);

BUFx6f_ASAP7_75t_L g1968 ( 
.A(n_1544),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1547),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1552),
.Y(n_1970)
);

HB1xp67_ASAP7_75t_L g1971 ( 
.A(n_1594),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1553),
.Y(n_1972)
);

OA21x2_ASAP7_75t_L g1973 ( 
.A1(n_1620),
.A2(n_1090),
.B(n_1086),
.Y(n_1973)
);

INVx2_ASAP7_75t_SL g1974 ( 
.A(n_1559),
.Y(n_1974)
);

INVx3_ASAP7_75t_L g1975 ( 
.A(n_1564),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1567),
.Y(n_1976)
);

OA21x2_ASAP7_75t_L g1977 ( 
.A1(n_1620),
.A2(n_1093),
.B(n_1092),
.Y(n_1977)
);

BUFx6f_ASAP7_75t_L g1978 ( 
.A(n_1570),
.Y(n_1978)
);

INVx5_ASAP7_75t_L g1979 ( 
.A(n_1632),
.Y(n_1979)
);

BUFx6f_ASAP7_75t_L g1980 ( 
.A(n_1573),
.Y(n_1980)
);

AOI22xp5_ASAP7_75t_L g1981 ( 
.A1(n_1626),
.A2(n_1692),
.B1(n_1627),
.B2(n_1633),
.Y(n_1981)
);

BUFx3_ASAP7_75t_L g1982 ( 
.A(n_1595),
.Y(n_1982)
);

INVx3_ASAP7_75t_L g1983 ( 
.A(n_1574),
.Y(n_1983)
);

BUFx6f_ASAP7_75t_L g1984 ( 
.A(n_1654),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1655),
.B(n_1345),
.Y(n_1985)
);

HB1xp67_ASAP7_75t_L g1986 ( 
.A(n_1598),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1595),
.B(n_1351),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1663),
.Y(n_1988)
);

OAI22xp33_ASAP7_75t_R g1989 ( 
.A1(n_1849),
.A2(n_932),
.B1(n_765),
.B2(n_942),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1721),
.B(n_1626),
.Y(n_1990)
);

NOR2xp33_ASAP7_75t_L g1991 ( 
.A(n_1858),
.B(n_1577),
.Y(n_1991)
);

OAI22xp33_ASAP7_75t_L g1992 ( 
.A1(n_1732),
.A2(n_1981),
.B1(n_1778),
.B2(n_1822),
.Y(n_1992)
);

AND2x4_ASAP7_75t_L g1993 ( 
.A(n_1916),
.B(n_1596),
.Y(n_1993)
);

OAI22xp5_ASAP7_75t_SL g1994 ( 
.A1(n_1736),
.A2(n_1599),
.B1(n_1606),
.B2(n_1592),
.Y(n_1994)
);

XNOR2xp5_ASAP7_75t_L g1995 ( 
.A(n_1777),
.B(n_1472),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1721),
.B(n_1627),
.Y(n_1996)
);

AO22x2_ASAP7_75t_L g1997 ( 
.A1(n_1777),
.A2(n_1621),
.B1(n_1599),
.B2(n_1606),
.Y(n_1997)
);

AOI22xp5_ASAP7_75t_L g1998 ( 
.A1(n_1929),
.A2(n_1633),
.B1(n_1636),
.B2(n_1629),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1801),
.Y(n_1999)
);

AOI22xp5_ASAP7_75t_L g2000 ( 
.A1(n_1725),
.A2(n_1636),
.B1(n_1637),
.B2(n_1629),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1801),
.Y(n_2001)
);

OAI22xp5_ASAP7_75t_SL g2002 ( 
.A1(n_1736),
.A2(n_1607),
.B1(n_1611),
.B2(n_1592),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1726),
.B(n_1637),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1801),
.Y(n_2004)
);

AOI22xp5_ASAP7_75t_L g2005 ( 
.A1(n_1725),
.A2(n_1648),
.B1(n_1692),
.B2(n_1638),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1801),
.Y(n_2006)
);

OAI22xp33_ASAP7_75t_L g2007 ( 
.A1(n_1959),
.A2(n_1648),
.B1(n_1638),
.B2(n_1669),
.Y(n_2007)
);

OA22x2_ASAP7_75t_L g2008 ( 
.A1(n_1754),
.A2(n_1413),
.B1(n_1615),
.B2(n_1678),
.Y(n_2008)
);

OAI22xp5_ASAP7_75t_SL g2009 ( 
.A1(n_1744),
.A2(n_1611),
.B1(n_1618),
.B2(n_1607),
.Y(n_2009)
);

AO22x2_ASAP7_75t_L g2010 ( 
.A1(n_1762),
.A2(n_1644),
.B1(n_1618),
.B2(n_1408),
.Y(n_2010)
);

AOI22xp5_ASAP7_75t_L g2011 ( 
.A1(n_1833),
.A2(n_1931),
.B1(n_1814),
.B2(n_1911),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1726),
.B(n_1691),
.Y(n_2012)
);

OAI22xp33_ASAP7_75t_SL g2013 ( 
.A1(n_1952),
.A2(n_1322),
.B1(n_1328),
.B2(n_1327),
.Y(n_2013)
);

AO22x2_ASAP7_75t_L g2014 ( 
.A1(n_1716),
.A2(n_1644),
.B1(n_1408),
.B2(n_1435),
.Y(n_2014)
);

AOI22xp5_ASAP7_75t_L g2015 ( 
.A1(n_1833),
.A2(n_1327),
.B1(n_1330),
.B2(n_1328),
.Y(n_2015)
);

INVx8_ASAP7_75t_L g2016 ( 
.A(n_1881),
.Y(n_2016)
);

OR2x2_ASAP7_75t_L g2017 ( 
.A(n_1784),
.B(n_1588),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1801),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1927),
.Y(n_2019)
);

OR2x2_ASAP7_75t_L g2020 ( 
.A(n_1784),
.B(n_1602),
.Y(n_2020)
);

OAI22xp33_ASAP7_75t_L g2021 ( 
.A1(n_1831),
.A2(n_1677),
.B1(n_1680),
.B2(n_1667),
.Y(n_2021)
);

OAI22xp5_ASAP7_75t_SL g2022 ( 
.A1(n_1744),
.A2(n_1435),
.B1(n_1451),
.B2(n_1422),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1927),
.Y(n_2023)
);

OAI22xp5_ASAP7_75t_SL g2024 ( 
.A1(n_1819),
.A2(n_1451),
.B1(n_1456),
.B2(n_1422),
.Y(n_2024)
);

OR2x6_ASAP7_75t_L g2025 ( 
.A(n_1829),
.B(n_1472),
.Y(n_2025)
);

AOI22xp5_ASAP7_75t_L g2026 ( 
.A1(n_1833),
.A2(n_1330),
.B1(n_1332),
.B2(n_1331),
.Y(n_2026)
);

AO22x2_ASAP7_75t_L g2027 ( 
.A1(n_1716),
.A2(n_1456),
.B1(n_1470),
.B2(n_1466),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_SL g2028 ( 
.A(n_1939),
.B(n_1347),
.Y(n_2028)
);

OAI22xp33_ASAP7_75t_L g2029 ( 
.A1(n_1951),
.A2(n_1680),
.B1(n_1682),
.B2(n_1677),
.Y(n_2029)
);

AOI22xp5_ASAP7_75t_L g2030 ( 
.A1(n_1833),
.A2(n_1331),
.B1(n_1333),
.B2(n_1332),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_1844),
.Y(n_2031)
);

NOR2xp33_ASAP7_75t_L g2032 ( 
.A(n_1791),
.B(n_1596),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1706),
.Y(n_2033)
);

AND2x2_ASAP7_75t_SL g2034 ( 
.A(n_1915),
.B(n_1682),
.Y(n_2034)
);

INVxp33_ASAP7_75t_L g2035 ( 
.A(n_1704),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1738),
.B(n_1601),
.Y(n_2036)
);

OAI22xp5_ASAP7_75t_SL g2037 ( 
.A1(n_1819),
.A2(n_1470),
.B1(n_1471),
.B2(n_1466),
.Y(n_2037)
);

OA22x2_ASAP7_75t_L g2038 ( 
.A1(n_1834),
.A2(n_1602),
.B1(n_1601),
.B2(n_1333),
.Y(n_2038)
);

INVx2_ASAP7_75t_SL g2039 ( 
.A(n_1738),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1844),
.Y(n_2040)
);

AO22x2_ASAP7_75t_L g2041 ( 
.A1(n_1804),
.A2(n_1471),
.B1(n_1480),
.B2(n_1475),
.Y(n_2041)
);

AOI22xp5_ASAP7_75t_L g2042 ( 
.A1(n_1833),
.A2(n_1339),
.B1(n_1348),
.B2(n_1347),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1791),
.B(n_1339),
.Y(n_2043)
);

INVx2_ASAP7_75t_SL g2044 ( 
.A(n_1895),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1706),
.Y(n_2045)
);

OAI22xp33_ASAP7_75t_L g2046 ( 
.A1(n_1951),
.A2(n_1939),
.B1(n_1945),
.B2(n_1944),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1844),
.Y(n_2047)
);

AO22x2_ASAP7_75t_L g2048 ( 
.A1(n_1957),
.A2(n_1475),
.B1(n_1482),
.B2(n_1480),
.Y(n_2048)
);

OR2x2_ASAP7_75t_L g2049 ( 
.A(n_1895),
.B(n_1752),
.Y(n_2049)
);

OAI22xp33_ASAP7_75t_L g2050 ( 
.A1(n_1939),
.A2(n_1688),
.B1(n_1380),
.B2(n_1388),
.Y(n_2050)
);

OAI22xp33_ASAP7_75t_SL g2051 ( 
.A1(n_1952),
.A2(n_1348),
.B1(n_1352),
.B2(n_1349),
.Y(n_2051)
);

AOI22xp5_ASAP7_75t_L g2052 ( 
.A1(n_1833),
.A2(n_1349),
.B1(n_1353),
.B2(n_1352),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1712),
.Y(n_2053)
);

OAI22xp33_ASAP7_75t_SL g2054 ( 
.A1(n_1955),
.A2(n_1353),
.B1(n_1369),
.B2(n_1365),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_1844),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1844),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1856),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_1928),
.B(n_1365),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1856),
.Y(n_2059)
);

OR2x6_ASAP7_75t_L g2060 ( 
.A(n_1829),
.B(n_1482),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1712),
.Y(n_2061)
);

OAI22xp5_ASAP7_75t_SL g2062 ( 
.A1(n_1830),
.A2(n_1497),
.B1(n_1511),
.B2(n_1490),
.Y(n_2062)
);

AOI22xp5_ASAP7_75t_L g2063 ( 
.A1(n_1911),
.A2(n_1377),
.B1(n_1380),
.B2(n_1379),
.Y(n_2063)
);

AND2x2_ASAP7_75t_SL g2064 ( 
.A(n_1770),
.B(n_1688),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1718),
.Y(n_2065)
);

AOI22xp5_ASAP7_75t_L g2066 ( 
.A1(n_1788),
.A2(n_1388),
.B1(n_992),
.B2(n_987),
.Y(n_2066)
);

INVxp67_ASAP7_75t_SL g2067 ( 
.A(n_1936),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1718),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_SL g2069 ( 
.A(n_1939),
.B(n_994),
.Y(n_2069)
);

OAI22xp33_ASAP7_75t_SL g2070 ( 
.A1(n_1955),
.A2(n_996),
.B1(n_993),
.B2(n_986),
.Y(n_2070)
);

INVx2_ASAP7_75t_SL g2071 ( 
.A(n_1916),
.Y(n_2071)
);

INVxp67_ASAP7_75t_SL g2072 ( 
.A(n_1798),
.Y(n_2072)
);

INVxp67_ASAP7_75t_L g2073 ( 
.A(n_1854),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1728),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_1928),
.B(n_1372),
.Y(n_2075)
);

HB1xp67_ASAP7_75t_L g2076 ( 
.A(n_1740),
.Y(n_2076)
);

AO22x2_ASAP7_75t_L g2077 ( 
.A1(n_1899),
.A2(n_1490),
.B1(n_1511),
.B2(n_1497),
.Y(n_2077)
);

AOI22xp5_ASAP7_75t_L g2078 ( 
.A1(n_1788),
.A2(n_997),
.B1(n_1003),
.B2(n_1000),
.Y(n_2078)
);

NAND2xp33_ASAP7_75t_SL g2079 ( 
.A(n_1826),
.B(n_1835),
.Y(n_2079)
);

OAI22xp33_ASAP7_75t_SL g2080 ( 
.A1(n_1960),
.A2(n_1013),
.B1(n_1017),
.B2(n_1004),
.Y(n_2080)
);

AOI22xp5_ASAP7_75t_L g2081 ( 
.A1(n_1788),
.A2(n_1020),
.B1(n_1018),
.B2(n_999),
.Y(n_2081)
);

AOI22xp5_ASAP7_75t_L g2082 ( 
.A1(n_1961),
.A2(n_1002),
.B1(n_1006),
.B2(n_995),
.Y(n_2082)
);

OAI22xp5_ASAP7_75t_SL g2083 ( 
.A1(n_1830),
.A2(n_1513),
.B1(n_1521),
.B2(n_1516),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_1711),
.B(n_1372),
.Y(n_2084)
);

INVx5_ASAP7_75t_L g2085 ( 
.A(n_1731),
.Y(n_2085)
);

AOI22xp5_ASAP7_75t_L g2086 ( 
.A1(n_1961),
.A2(n_1009),
.B1(n_1011),
.B2(n_1007),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_1711),
.B(n_1351),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1728),
.Y(n_2088)
);

NOR2xp33_ASAP7_75t_SL g2089 ( 
.A(n_1760),
.B(n_1565),
.Y(n_2089)
);

OAI22xp33_ASAP7_75t_L g2090 ( 
.A1(n_1939),
.A2(n_924),
.B1(n_955),
.B2(n_900),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1856),
.Y(n_2091)
);

AO22x2_ASAP7_75t_L g2092 ( 
.A1(n_1899),
.A2(n_1516),
.B1(n_1521),
.B2(n_1513),
.Y(n_2092)
);

AOI22xp5_ASAP7_75t_L g2093 ( 
.A1(n_1930),
.A2(n_1789),
.B1(n_1729),
.B2(n_1892),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_1739),
.B(n_1940),
.Y(n_2094)
);

OAI22xp33_ASAP7_75t_L g2095 ( 
.A1(n_1944),
.A2(n_955),
.B1(n_924),
.B2(n_824),
.Y(n_2095)
);

AOI22xp5_ASAP7_75t_L g2096 ( 
.A1(n_1930),
.A2(n_1892),
.B1(n_1935),
.B2(n_1739),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_1802),
.B(n_1336),
.Y(n_2097)
);

CKINVDCx8_ASAP7_75t_R g2098 ( 
.A(n_1916),
.Y(n_2098)
);

AOI22xp5_ASAP7_75t_L g2099 ( 
.A1(n_1930),
.A2(n_1016),
.B1(n_1019),
.B2(n_1015),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_1940),
.B(n_1358),
.Y(n_2100)
);

OAI22xp33_ASAP7_75t_L g2101 ( 
.A1(n_1944),
.A2(n_824),
.B1(n_830),
.B2(n_820),
.Y(n_2101)
);

AO22x2_ASAP7_75t_L g2102 ( 
.A1(n_1710),
.A2(n_1545),
.B1(n_1554),
.B2(n_1532),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1856),
.Y(n_2103)
);

AND2x2_ASAP7_75t_L g2104 ( 
.A(n_1974),
.B(n_1358),
.Y(n_2104)
);

INVx8_ASAP7_75t_L g2105 ( 
.A(n_1881),
.Y(n_2105)
);

OR2x6_ASAP7_75t_L g2106 ( 
.A(n_1938),
.B(n_1532),
.Y(n_2106)
);

AO22x2_ASAP7_75t_L g2107 ( 
.A1(n_1863),
.A2(n_1554),
.B1(n_1565),
.B2(n_1545),
.Y(n_2107)
);

AO22x2_ASAP7_75t_L g2108 ( 
.A1(n_1863),
.A2(n_830),
.B1(n_834),
.B2(n_820),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_SL g2109 ( 
.A(n_1944),
.B(n_1021),
.Y(n_2109)
);

BUFx10_ASAP7_75t_L g2110 ( 
.A(n_1720),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_1974),
.B(n_1361),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_1894),
.B(n_1918),
.Y(n_2112)
);

AOI22xp5_ASAP7_75t_L g2113 ( 
.A1(n_1930),
.A2(n_1028),
.B1(n_1027),
.B2(n_1284),
.Y(n_2113)
);

INVx2_ASAP7_75t_SL g2114 ( 
.A(n_1916),
.Y(n_2114)
);

OAI22xp33_ASAP7_75t_SL g2115 ( 
.A1(n_1960),
.A2(n_835),
.B1(n_836),
.B2(n_834),
.Y(n_2115)
);

AO22x2_ASAP7_75t_L g2116 ( 
.A1(n_1868),
.A2(n_836),
.B1(n_843),
.B2(n_835),
.Y(n_2116)
);

AOI22xp5_ASAP7_75t_L g2117 ( 
.A1(n_1930),
.A2(n_852),
.B1(n_854),
.B2(n_843),
.Y(n_2117)
);

AOI22xp5_ASAP7_75t_L g2118 ( 
.A1(n_1892),
.A2(n_854),
.B1(n_860),
.B2(n_852),
.Y(n_2118)
);

BUFx3_ASAP7_75t_L g2119 ( 
.A(n_1867),
.Y(n_2119)
);

AOI22xp5_ASAP7_75t_L g2120 ( 
.A1(n_1935),
.A2(n_864),
.B1(n_865),
.B2(n_860),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_1856),
.Y(n_2121)
);

OAI22xp33_ASAP7_75t_SL g2122 ( 
.A1(n_1868),
.A2(n_865),
.B1(n_866),
.B2(n_864),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_SL g2123 ( 
.A(n_1944),
.B(n_1945),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_1857),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_1867),
.B(n_1361),
.Y(n_2125)
);

NAND3x1_ASAP7_75t_L g2126 ( 
.A(n_1934),
.B(n_875),
.C(n_866),
.Y(n_2126)
);

AO22x2_ASAP7_75t_L g2127 ( 
.A1(n_1987),
.A2(n_879),
.B1(n_887),
.B2(n_875),
.Y(n_2127)
);

OAI22xp33_ASAP7_75t_SL g2128 ( 
.A1(n_1942),
.A2(n_887),
.B1(n_891),
.B2(n_879),
.Y(n_2128)
);

AOI22xp5_ASAP7_75t_L g2129 ( 
.A1(n_1935),
.A2(n_893),
.B1(n_905),
.B2(n_891),
.Y(n_2129)
);

INVx4_ASAP7_75t_L g2130 ( 
.A(n_1731),
.Y(n_2130)
);

AOI22xp5_ASAP7_75t_L g2131 ( 
.A1(n_1793),
.A2(n_905),
.B1(n_910),
.B2(n_893),
.Y(n_2131)
);

OAI22xp33_ASAP7_75t_L g2132 ( 
.A1(n_1945),
.A2(n_917),
.B1(n_918),
.B2(n_910),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1733),
.Y(n_2133)
);

AOI22xp5_ASAP7_75t_L g2134 ( 
.A1(n_1953),
.A2(n_918),
.B1(n_926),
.B2(n_917),
.Y(n_2134)
);

OAI22xp5_ASAP7_75t_SL g2135 ( 
.A1(n_1878),
.A2(n_934),
.B1(n_935),
.B2(n_926),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1733),
.Y(n_2136)
);

AOI22xp5_ASAP7_75t_L g2137 ( 
.A1(n_1805),
.A2(n_935),
.B1(n_938),
.B2(n_934),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_1906),
.B(n_1371),
.Y(n_2138)
);

OAI22xp33_ASAP7_75t_L g2139 ( 
.A1(n_1945),
.A2(n_946),
.B1(n_954),
.B2(n_938),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_1857),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_1906),
.B(n_1371),
.Y(n_2141)
);

OR2x6_ASAP7_75t_L g2142 ( 
.A(n_1938),
.B(n_1910),
.Y(n_2142)
);

OA22x2_ASAP7_75t_L g2143 ( 
.A1(n_1864),
.A2(n_954),
.B1(n_956),
.B2(n_946),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_1802),
.B(n_1336),
.Y(n_2144)
);

AOI22xp5_ASAP7_75t_L g2145 ( 
.A1(n_1805),
.A2(n_974),
.B1(n_975),
.B2(n_956),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_1910),
.B(n_1023),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1758),
.Y(n_2147)
);

OAI22xp33_ASAP7_75t_L g2148 ( 
.A1(n_1945),
.A2(n_975),
.B1(n_981),
.B2(n_974),
.Y(n_2148)
);

AOI22xp5_ASAP7_75t_L g2149 ( 
.A1(n_1805),
.A2(n_991),
.B1(n_1001),
.B2(n_981),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1705),
.Y(n_2150)
);

OR2x2_ASAP7_75t_L g2151 ( 
.A(n_1772),
.B(n_991),
.Y(n_2151)
);

AOI22xp5_ASAP7_75t_L g2152 ( 
.A1(n_1806),
.A2(n_1815),
.B1(n_1813),
.B2(n_1802),
.Y(n_2152)
);

BUFx6f_ASAP7_75t_L g2153 ( 
.A(n_1857),
.Y(n_2153)
);

NAND3x1_ASAP7_75t_L g2154 ( 
.A(n_1934),
.B(n_1010),
.C(n_1001),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_1933),
.B(n_1012),
.Y(n_2155)
);

OAI22xp5_ASAP7_75t_SL g2156 ( 
.A1(n_1878),
.A2(n_1023),
.B1(n_1012),
.B2(n_1336),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1705),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_1857),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1705),
.Y(n_2159)
);

AOI22xp5_ASAP7_75t_L g2160 ( 
.A1(n_1806),
.A2(n_1336),
.B1(n_1094),
.B2(n_1096),
.Y(n_2160)
);

OAI22xp5_ASAP7_75t_L g2161 ( 
.A1(n_1807),
.A2(n_1095),
.B1(n_1100),
.B2(n_1099),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_1857),
.Y(n_2162)
);

NOR2xp33_ASAP7_75t_L g2163 ( 
.A(n_1941),
.B(n_218),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_1933),
.B(n_1336),
.Y(n_2164)
);

AO22x2_ASAP7_75t_L g2165 ( 
.A1(n_1987),
.A2(n_1108),
.B1(n_1109),
.B2(n_1102),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_1824),
.B(n_1210),
.Y(n_2166)
);

OAI22xp33_ASAP7_75t_L g2167 ( 
.A1(n_1947),
.A2(n_1180),
.B1(n_1210),
.B2(n_1150),
.Y(n_2167)
);

AO22x2_ASAP7_75t_L g2168 ( 
.A1(n_1941),
.A2(n_1114),
.B1(n_1121),
.B2(n_1112),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_1866),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_1807),
.B(n_1846),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_1824),
.B(n_1305),
.Y(n_2171)
);

OAI22xp33_ASAP7_75t_SL g2172 ( 
.A1(n_1942),
.A2(n_1124),
.B1(n_1127),
.B2(n_1122),
.Y(n_2172)
);

OAI22xp33_ASAP7_75t_L g2173 ( 
.A1(n_1947),
.A2(n_1180),
.B1(n_1285),
.B2(n_1150),
.Y(n_2173)
);

AOI22xp5_ASAP7_75t_L g2174 ( 
.A1(n_1806),
.A2(n_1132),
.B1(n_1137),
.B2(n_1128),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_1866),
.Y(n_2175)
);

INVx3_ASAP7_75t_L g2176 ( 
.A(n_1866),
.Y(n_2176)
);

BUFx6f_ASAP7_75t_SL g2177 ( 
.A(n_1982),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1722),
.Y(n_2178)
);

OAI22xp33_ASAP7_75t_SL g2179 ( 
.A1(n_1946),
.A2(n_1138),
.B1(n_1305),
.B2(n_1285),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_1866),
.Y(n_2180)
);

AOI22xp5_ASAP7_75t_L g2181 ( 
.A1(n_1813),
.A2(n_1316),
.B1(n_1117),
.B2(n_1167),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_1866),
.Y(n_2182)
);

AOI22xp5_ASAP7_75t_L g2183 ( 
.A1(n_1813),
.A2(n_1316),
.B1(n_1117),
.B2(n_1167),
.Y(n_2183)
);

OAI22xp33_ASAP7_75t_SL g2184 ( 
.A1(n_1946),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_2184)
);

AO22x2_ASAP7_75t_L g2185 ( 
.A1(n_1969),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_2185)
);

AOI22xp5_ASAP7_75t_L g2186 ( 
.A1(n_1815),
.A2(n_1117),
.B1(n_1167),
.B2(n_1087),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1722),
.Y(n_2187)
);

AOI22xp5_ASAP7_75t_L g2188 ( 
.A1(n_1815),
.A2(n_1117),
.B1(n_1167),
.B2(n_1087),
.Y(n_2188)
);

NOR2xp33_ASAP7_75t_L g2189 ( 
.A(n_1969),
.B(n_219),
.Y(n_2189)
);

OAI22xp33_ASAP7_75t_SL g2190 ( 
.A1(n_1949),
.A2(n_8),
.B1(n_5),
.B2(n_6),
.Y(n_2190)
);

AOI22xp5_ASAP7_75t_L g2191 ( 
.A1(n_1807),
.A2(n_1117),
.B1(n_1167),
.B2(n_1087),
.Y(n_2191)
);

AO22x2_ASAP7_75t_L g2192 ( 
.A1(n_1970),
.A2(n_9),
.B1(n_6),
.B2(n_8),
.Y(n_2192)
);

OAI22xp5_ASAP7_75t_SL g2193 ( 
.A1(n_1760),
.A2(n_11),
.B1(n_8),
.B2(n_10),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_1891),
.Y(n_2194)
);

OAI22xp5_ASAP7_75t_L g2195 ( 
.A1(n_1846),
.A2(n_1175),
.B1(n_1224),
.B2(n_1087),
.Y(n_2195)
);

OAI22xp5_ASAP7_75t_SL g2196 ( 
.A1(n_1869),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_1824),
.B(n_10),
.Y(n_2197)
);

AOI22xp5_ASAP7_75t_L g2198 ( 
.A1(n_1846),
.A2(n_1175),
.B1(n_1224),
.B2(n_1087),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1722),
.Y(n_2199)
);

OR2x6_ASAP7_75t_L g2200 ( 
.A(n_1947),
.B(n_1853),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_1825),
.B(n_11),
.Y(n_2201)
);

AOI22xp5_ASAP7_75t_L g2202 ( 
.A1(n_1848),
.A2(n_1224),
.B1(n_1296),
.B2(n_1175),
.Y(n_2202)
);

OAI22xp33_ASAP7_75t_L g2203 ( 
.A1(n_1947),
.A2(n_1224),
.B1(n_1296),
.B2(n_1175),
.Y(n_2203)
);

OAI22xp33_ASAP7_75t_L g2204 ( 
.A1(n_1947),
.A2(n_1224),
.B1(n_1296),
.B2(n_1175),
.Y(n_2204)
);

AOI22xp5_ASAP7_75t_L g2205 ( 
.A1(n_1848),
.A2(n_1296),
.B1(n_14),
.B2(n_12),
.Y(n_2205)
);

AOI22xp5_ASAP7_75t_L g2206 ( 
.A1(n_1848),
.A2(n_1859),
.B1(n_1880),
.B2(n_1746),
.Y(n_2206)
);

AOI22xp5_ASAP7_75t_L g2207 ( 
.A1(n_1859),
.A2(n_1296),
.B1(n_14),
.B2(n_12),
.Y(n_2207)
);

AND2x2_ASAP7_75t_L g2208 ( 
.A(n_1825),
.B(n_13),
.Y(n_2208)
);

OA22x2_ASAP7_75t_L g2209 ( 
.A1(n_1890),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_2209)
);

NAND3x1_ASAP7_75t_L g2210 ( 
.A(n_1934),
.B(n_22),
.C(n_13),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_1825),
.B(n_15),
.Y(n_2211)
);

AOI22xp5_ASAP7_75t_L g2212 ( 
.A1(n_1859),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_2212)
);

OAI22xp33_ASAP7_75t_SL g2213 ( 
.A1(n_1949),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_2213)
);

CKINVDCx8_ASAP7_75t_R g2214 ( 
.A(n_1916),
.Y(n_2214)
);

AO22x2_ASAP7_75t_L g2215 ( 
.A1(n_1970),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_2215)
);

OAI22xp33_ASAP7_75t_L g2216 ( 
.A1(n_1720),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_2216)
);

OAI22xp33_ASAP7_75t_L g2217 ( 
.A1(n_1755),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_2217)
);

INVx2_ASAP7_75t_SL g2218 ( 
.A(n_1919),
.Y(n_2218)
);

INVx2_ASAP7_75t_L g2219 ( 
.A(n_1891),
.Y(n_2219)
);

AO22x2_ASAP7_75t_L g2220 ( 
.A1(n_1972),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_2220)
);

OR2x2_ASAP7_75t_L g2221 ( 
.A(n_1817),
.B(n_23),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1909),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1917),
.Y(n_2223)
);

AOI22xp5_ASAP7_75t_L g2224 ( 
.A1(n_1880),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_2224)
);

OR2x6_ASAP7_75t_L g2225 ( 
.A(n_1841),
.B(n_1860),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_1908),
.B(n_24),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_1925),
.B(n_25),
.Y(n_2227)
);

INVx2_ASAP7_75t_SL g2228 ( 
.A(n_1919),
.Y(n_2228)
);

OAI22xp33_ASAP7_75t_L g2229 ( 
.A1(n_1755),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_1826),
.B(n_26),
.Y(n_2230)
);

AO22x2_ASAP7_75t_L g2231 ( 
.A1(n_1972),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_2231)
);

OAI22xp33_ASAP7_75t_L g2232 ( 
.A1(n_1763),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_2232)
);

OAI22xp33_ASAP7_75t_SL g2233 ( 
.A1(n_1956),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_1891),
.Y(n_2234)
);

INVx2_ASAP7_75t_SL g2235 ( 
.A(n_1919),
.Y(n_2235)
);

AOI22xp5_ASAP7_75t_L g2236 ( 
.A1(n_1880),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_2236)
);

AND3x1_ASAP7_75t_L g2237 ( 
.A(n_1962),
.B(n_31),
.C(n_32),
.Y(n_2237)
);

BUFx2_ASAP7_75t_L g2238 ( 
.A(n_1954),
.Y(n_2238)
);

OAI22xp33_ASAP7_75t_L g2239 ( 
.A1(n_1763),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_2239)
);

AND2x2_ASAP7_75t_L g2240 ( 
.A(n_1826),
.B(n_33),
.Y(n_2240)
);

AO22x2_ASAP7_75t_L g2241 ( 
.A1(n_1963),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_1891),
.Y(n_2242)
);

AOI22xp5_ASAP7_75t_L g2243 ( 
.A1(n_1746),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_2243)
);

AND2x2_ASAP7_75t_L g2244 ( 
.A(n_1835),
.B(n_35),
.Y(n_2244)
);

AOI22xp5_ASAP7_75t_L g2245 ( 
.A1(n_1786),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_2245)
);

OAI22xp33_ASAP7_75t_SL g2246 ( 
.A1(n_1769),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_1921),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_1835),
.B(n_38),
.Y(n_2248)
);

AOI22xp5_ASAP7_75t_L g2249 ( 
.A1(n_1786),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_2249)
);

INVx2_ASAP7_75t_SL g2250 ( 
.A(n_1919),
.Y(n_2250)
);

AO22x2_ASAP7_75t_L g2251 ( 
.A1(n_1750),
.A2(n_1776),
.B1(n_1976),
.B2(n_1967),
.Y(n_2251)
);

AOI22xp5_ASAP7_75t_L g2252 ( 
.A1(n_1786),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_SL g2253 ( 
.A(n_1965),
.B(n_219),
.Y(n_2253)
);

AND2x2_ASAP7_75t_L g2254 ( 
.A(n_1888),
.B(n_1787),
.Y(n_2254)
);

AOI22xp5_ASAP7_75t_L g2255 ( 
.A1(n_1787),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_2255)
);

OAI22xp33_ASAP7_75t_SL g2256 ( 
.A1(n_1769),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_2256)
);

AOI22xp5_ASAP7_75t_L g2257 ( 
.A1(n_1787),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1799),
.Y(n_2258)
);

AOI22x1_ASAP7_75t_L g2259 ( 
.A1(n_1932),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_2259)
);

AND2x2_ASAP7_75t_L g2260 ( 
.A(n_1888),
.B(n_46),
.Y(n_2260)
);

AO22x2_ASAP7_75t_L g2261 ( 
.A1(n_1750),
.A2(n_49),
.B1(n_46),
.B2(n_48),
.Y(n_2261)
);

NOR2xp33_ASAP7_75t_L g2262 ( 
.A(n_1988),
.B(n_220),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_1888),
.B(n_50),
.Y(n_2263)
);

AND2x2_ASAP7_75t_L g2264 ( 
.A(n_1975),
.B(n_51),
.Y(n_2264)
);

AOI22xp5_ASAP7_75t_L g2265 ( 
.A1(n_1891),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_2265)
);

INVx2_ASAP7_75t_SL g2266 ( 
.A(n_1919),
.Y(n_2266)
);

OAI22xp33_ASAP7_75t_SL g2267 ( 
.A1(n_1782),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_2267)
);

AO22x2_ASAP7_75t_L g2268 ( 
.A1(n_1750),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_2268)
);

AO22x2_ASAP7_75t_L g2269 ( 
.A1(n_1776),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_1799),
.Y(n_2270)
);

AND2x2_ASAP7_75t_L g2271 ( 
.A(n_1975),
.B(n_1983),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_1896),
.Y(n_2272)
);

OAI22xp33_ASAP7_75t_L g2273 ( 
.A1(n_1782),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_1893),
.B(n_55),
.Y(n_2274)
);

AOI22xp5_ASAP7_75t_L g2275 ( 
.A1(n_1896),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_2275)
);

OR2x2_ASAP7_75t_L g2276 ( 
.A(n_1808),
.B(n_57),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_1964),
.B(n_1985),
.Y(n_2277)
);

BUFx6f_ASAP7_75t_L g2278 ( 
.A(n_1896),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_1875),
.Y(n_2279)
);

OAI22xp33_ASAP7_75t_L g2280 ( 
.A1(n_1808),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_1875),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_SL g2282 ( 
.A(n_1965),
.B(n_221),
.Y(n_2282)
);

AND2x2_ASAP7_75t_L g2283 ( 
.A(n_1975),
.B(n_58),
.Y(n_2283)
);

INVx1_ASAP7_75t_SL g2284 ( 
.A(n_1971),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_1798),
.B(n_59),
.Y(n_2285)
);

AOI22xp5_ASAP7_75t_L g2286 ( 
.A1(n_1896),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_1966),
.Y(n_2287)
);

AOI22xp5_ASAP7_75t_L g2288 ( 
.A1(n_1896),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_2288)
);

OAI22xp5_ASAP7_75t_L g2289 ( 
.A1(n_1798),
.A2(n_222),
.B1(n_223),
.B2(n_221),
.Y(n_2289)
);

OAI22xp33_ASAP7_75t_L g2290 ( 
.A1(n_1843),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_2290)
);

OAI22xp5_ASAP7_75t_SL g2291 ( 
.A1(n_1902),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_2291)
);

AND2x2_ASAP7_75t_L g2292 ( 
.A(n_1983),
.B(n_64),
.Y(n_2292)
);

OAI22xp33_ASAP7_75t_L g2293 ( 
.A1(n_1843),
.A2(n_1905),
.B1(n_1968),
.B2(n_1965),
.Y(n_2293)
);

OAI22xp33_ASAP7_75t_L g2294 ( 
.A1(n_1905),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_1966),
.Y(n_2295)
);

AND2x2_ASAP7_75t_L g2296 ( 
.A(n_1983),
.B(n_65),
.Y(n_2296)
);

OAI22xp33_ASAP7_75t_L g2297 ( 
.A1(n_1965),
.A2(n_1968),
.B1(n_1980),
.B2(n_1978),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_1982),
.B(n_66),
.Y(n_2298)
);

NOR2xp33_ASAP7_75t_L g2299 ( 
.A(n_1937),
.B(n_223),
.Y(n_2299)
);

NAND3x1_ASAP7_75t_L g2300 ( 
.A(n_1745),
.B(n_74),
.C(n_66),
.Y(n_2300)
);

AOI22xp5_ASAP7_75t_L g2301 ( 
.A1(n_1904),
.A2(n_1912),
.B1(n_1926),
.B2(n_1973),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_1965),
.B(n_67),
.Y(n_2302)
);

AO22x2_ASAP7_75t_L g2303 ( 
.A1(n_1776),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_1968),
.B(n_68),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_1715),
.Y(n_2305)
);

OAI22xp5_ASAP7_75t_SL g2306 ( 
.A1(n_1749),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_2306)
);

AOI22xp5_ASAP7_75t_L g2307 ( 
.A1(n_1904),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_1748),
.Y(n_2308)
);

AND2x2_ASAP7_75t_L g2309 ( 
.A(n_1968),
.B(n_70),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_1904),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_2150),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_2150),
.Y(n_2312)
);

NOR2xp33_ASAP7_75t_L g2313 ( 
.A(n_1998),
.B(n_1968),
.Y(n_2313)
);

OR2x2_ASAP7_75t_L g2314 ( 
.A(n_2017),
.B(n_1986),
.Y(n_2314)
);

NOR2xp33_ASAP7_75t_L g2315 ( 
.A(n_1992),
.B(n_1978),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_SL g2316 ( 
.A(n_2293),
.B(n_1978),
.Y(n_2316)
);

INVx8_ASAP7_75t_L g2317 ( 
.A(n_2177),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_SL g2318 ( 
.A(n_2093),
.B(n_1978),
.Y(n_2318)
);

AND2x6_ASAP7_75t_L g2319 ( 
.A(n_2301),
.B(n_1978),
.Y(n_2319)
);

BUFx3_ASAP7_75t_L g2320 ( 
.A(n_2016),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2033),
.Y(n_2321)
);

CKINVDCx16_ASAP7_75t_R g2322 ( 
.A(n_1994),
.Y(n_2322)
);

INVx3_ASAP7_75t_L g2323 ( 
.A(n_2153),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_2271),
.B(n_1980),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_SL g2325 ( 
.A(n_2254),
.B(n_1980),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2033),
.Y(n_2326)
);

INVxp67_ASAP7_75t_L g2327 ( 
.A(n_2044),
.Y(n_2327)
);

BUFx8_ASAP7_75t_SL g2328 ( 
.A(n_2025),
.Y(n_2328)
);

XOR2xp5_ASAP7_75t_L g2329 ( 
.A(n_1995),
.B(n_1980),
.Y(n_2329)
);

NAND2xp33_ASAP7_75t_L g2330 ( 
.A(n_2079),
.B(n_1980),
.Y(n_2330)
);

AND3x2_ASAP7_75t_L g2331 ( 
.A(n_2089),
.B(n_1877),
.C(n_1745),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2045),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2045),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2157),
.Y(n_2334)
);

INVx4_ASAP7_75t_L g2335 ( 
.A(n_2085),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2053),
.Y(n_2336)
);

INVx3_ASAP7_75t_L g2337 ( 
.A(n_2153),
.Y(n_2337)
);

INVx3_ASAP7_75t_L g2338 ( 
.A(n_2153),
.Y(n_2338)
);

INVx3_ASAP7_75t_L g2339 ( 
.A(n_2278),
.Y(n_2339)
);

NOR2xp33_ASAP7_75t_L g2340 ( 
.A(n_1991),
.B(n_1984),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2053),
.Y(n_2341)
);

HB1xp67_ASAP7_75t_L g2342 ( 
.A(n_2284),
.Y(n_2342)
);

INVx2_ASAP7_75t_SL g2343 ( 
.A(n_2085),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2061),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2061),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_2094),
.B(n_1984),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2065),
.Y(n_2347)
);

INVx2_ASAP7_75t_L g2348 ( 
.A(n_2157),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_2087),
.B(n_1984),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_2159),
.Y(n_2350)
);

BUFx10_ASAP7_75t_L g2351 ( 
.A(n_2032),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_SL g2352 ( 
.A(n_2046),
.B(n_1984),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_2152),
.B(n_1984),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2065),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_2019),
.B(n_1702),
.Y(n_2355)
);

AND2x2_ASAP7_75t_L g2356 ( 
.A(n_1990),
.B(n_1820),
.Y(n_2356)
);

BUFx3_ASAP7_75t_L g2357 ( 
.A(n_2016),
.Y(n_2357)
);

INVx3_ASAP7_75t_L g2358 ( 
.A(n_2278),
.Y(n_2358)
);

NAND2xp33_ASAP7_75t_L g2359 ( 
.A(n_2278),
.B(n_1794),
.Y(n_2359)
);

AND3x2_ASAP7_75t_L g2360 ( 
.A(n_2238),
.B(n_1877),
.C(n_1745),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2068),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_2159),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_2023),
.B(n_1702),
.Y(n_2363)
);

CKINVDCx16_ASAP7_75t_R g2364 ( 
.A(n_2002),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_2178),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2068),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2074),
.Y(n_2367)
);

INVx3_ASAP7_75t_L g2368 ( 
.A(n_2130),
.Y(n_2368)
);

AOI22xp33_ASAP7_75t_L g2369 ( 
.A1(n_1989),
.A2(n_1820),
.B1(n_1977),
.B2(n_1973),
.Y(n_2369)
);

AOI21x1_ASAP7_75t_L g2370 ( 
.A1(n_2287),
.A2(n_1855),
.B(n_1837),
.Y(n_2370)
);

BUFx10_ASAP7_75t_L g2371 ( 
.A(n_2177),
.Y(n_2371)
);

BUFx3_ASAP7_75t_L g2372 ( 
.A(n_2105),
.Y(n_2372)
);

OAI22xp33_ASAP7_75t_L g2373 ( 
.A1(n_2000),
.A2(n_1923),
.B1(n_1979),
.B2(n_1749),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_SL g2374 ( 
.A(n_2297),
.B(n_1923),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2178),
.Y(n_2375)
);

INVx2_ASAP7_75t_L g2376 ( 
.A(n_2187),
.Y(n_2376)
);

AND2x6_ASAP7_75t_L g2377 ( 
.A(n_2187),
.B(n_2199),
.Y(n_2377)
);

NOR2xp33_ASAP7_75t_L g2378 ( 
.A(n_2049),
.B(n_1923),
.Y(n_2378)
);

NAND2xp33_ASAP7_75t_L g2379 ( 
.A(n_2170),
.B(n_2206),
.Y(n_2379)
);

AND2x4_ASAP7_75t_L g2380 ( 
.A(n_2119),
.B(n_1923),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2074),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2088),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_2199),
.Y(n_2383)
);

INVx4_ASAP7_75t_L g2384 ( 
.A(n_2085),
.Y(n_2384)
);

INVx2_ASAP7_75t_L g2385 ( 
.A(n_2088),
.Y(n_2385)
);

NOR2x1p5_ASAP7_75t_L g2386 ( 
.A(n_2020),
.B(n_1993),
.Y(n_2386)
);

AND2x6_ASAP7_75t_L g2387 ( 
.A(n_2096),
.B(n_1820),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2133),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2133),
.Y(n_2389)
);

INVx3_ASAP7_75t_L g2390 ( 
.A(n_2130),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2136),
.Y(n_2391)
);

AND2x2_ASAP7_75t_L g2392 ( 
.A(n_1996),
.B(n_1702),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2136),
.Y(n_2393)
);

INVx2_ASAP7_75t_L g2394 ( 
.A(n_2287),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2295),
.Y(n_2395)
);

INVx3_ASAP7_75t_L g2396 ( 
.A(n_2176),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2097),
.Y(n_2397)
);

AND3x2_ASAP7_75t_L g2398 ( 
.A(n_1993),
.B(n_1877),
.C(n_1943),
.Y(n_2398)
);

INVx4_ASAP7_75t_L g2399 ( 
.A(n_2176),
.Y(n_2399)
);

INVx2_ASAP7_75t_SL g2400 ( 
.A(n_2125),
.Y(n_2400)
);

AOI22xp33_ASAP7_75t_L g2401 ( 
.A1(n_1989),
.A2(n_2116),
.B1(n_2108),
.B2(n_2226),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_2295),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2166),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2171),
.Y(n_2404)
);

BUFx3_ASAP7_75t_L g2405 ( 
.A(n_2105),
.Y(n_2405)
);

NOR2xp33_ASAP7_75t_L g2406 ( 
.A(n_2007),
.B(n_1923),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2100),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_SL g2408 ( 
.A(n_2005),
.B(n_1979),
.Y(n_2408)
);

OR2x2_ASAP7_75t_L g2409 ( 
.A(n_2021),
.B(n_1727),
.Y(n_2409)
);

HAxp5_ASAP7_75t_SL g2410 ( 
.A(n_2102),
.B(n_2245),
.CON(n_2410),
.SN(n_2410)
);

AND2x2_ASAP7_75t_L g2411 ( 
.A(n_2003),
.B(n_1727),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2104),
.Y(n_2412)
);

INVx2_ASAP7_75t_SL g2413 ( 
.A(n_2138),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2111),
.Y(n_2414)
);

INVx2_ASAP7_75t_SL g2415 ( 
.A(n_2141),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_SL g2416 ( 
.A(n_2012),
.B(n_1979),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2084),
.Y(n_2417)
);

INVx1_ASAP7_75t_SL g2418 ( 
.A(n_2043),
.Y(n_2418)
);

BUFx3_ASAP7_75t_L g2419 ( 
.A(n_2098),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2258),
.Y(n_2420)
);

BUFx2_ASAP7_75t_L g2421 ( 
.A(n_2225),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_SL g2422 ( 
.A(n_2011),
.B(n_1979),
.Y(n_2422)
);

AND2x2_ASAP7_75t_L g2423 ( 
.A(n_2058),
.B(n_1727),
.Y(n_2423)
);

INVx2_ASAP7_75t_SL g2424 ( 
.A(n_2200),
.Y(n_2424)
);

BUFx6f_ASAP7_75t_L g2425 ( 
.A(n_2214),
.Y(n_2425)
);

AOI22xp33_ASAP7_75t_L g2426 ( 
.A1(n_2108),
.A2(n_1977),
.B1(n_1973),
.B2(n_1912),
.Y(n_2426)
);

NOR2xp33_ASAP7_75t_L g2427 ( 
.A(n_2035),
.B(n_1979),
.Y(n_2427)
);

OAI22xp33_ASAP7_75t_L g2428 ( 
.A1(n_2066),
.A2(n_1889),
.B1(n_1912),
.B2(n_1904),
.Y(n_2428)
);

INVx2_ASAP7_75t_L g2429 ( 
.A(n_2258),
.Y(n_2429)
);

NOR2xp33_ASAP7_75t_L g2430 ( 
.A(n_2073),
.B(n_2050),
.Y(n_2430)
);

INVx2_ASAP7_75t_L g2431 ( 
.A(n_2270),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2270),
.Y(n_2432)
);

INVx3_ASAP7_75t_L g2433 ( 
.A(n_1999),
.Y(n_2433)
);

OR2x2_ASAP7_75t_L g2434 ( 
.A(n_2022),
.B(n_2024),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_2279),
.Y(n_2435)
);

OR2x6_ASAP7_75t_L g2436 ( 
.A(n_2142),
.B(n_1810),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_2279),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2281),
.Y(n_2438)
);

BUFx3_ASAP7_75t_L g2439 ( 
.A(n_2142),
.Y(n_2439)
);

INVx2_ASAP7_75t_L g2440 ( 
.A(n_2281),
.Y(n_2440)
);

INVx3_ASAP7_75t_L g2441 ( 
.A(n_2001),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_SL g2442 ( 
.A(n_2015),
.B(n_1948),
.Y(n_2442)
);

AOI21x1_ASAP7_75t_L g2443 ( 
.A1(n_2144),
.A2(n_1855),
.B(n_1837),
.Y(n_2443)
);

BUFx3_ASAP7_75t_L g2444 ( 
.A(n_2200),
.Y(n_2444)
);

INVx3_ASAP7_75t_L g2445 ( 
.A(n_2004),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2075),
.Y(n_2446)
);

INVx2_ASAP7_75t_SL g2447 ( 
.A(n_2164),
.Y(n_2447)
);

INVx2_ASAP7_75t_L g2448 ( 
.A(n_2006),
.Y(n_2448)
);

CKINVDCx11_ASAP7_75t_R g2449 ( 
.A(n_2110),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_SL g2450 ( 
.A(n_2026),
.B(n_1904),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2039),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_2018),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2168),
.Y(n_2453)
);

BUFx6f_ASAP7_75t_L g2454 ( 
.A(n_2031),
.Y(n_2454)
);

NOR2xp33_ASAP7_75t_L g2455 ( 
.A(n_2063),
.B(n_1950),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2168),
.Y(n_2456)
);

INVx4_ASAP7_75t_L g2457 ( 
.A(n_2040),
.Y(n_2457)
);

INVx3_ASAP7_75t_L g2458 ( 
.A(n_2047),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2274),
.Y(n_2459)
);

BUFx4f_ASAP7_75t_L g2460 ( 
.A(n_2071),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2161),
.Y(n_2461)
);

AND2x6_ASAP7_75t_L g2462 ( 
.A(n_2302),
.B(n_1912),
.Y(n_2462)
);

BUFx6f_ASAP7_75t_L g2463 ( 
.A(n_2055),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2305),
.Y(n_2464)
);

INVx2_ASAP7_75t_L g2465 ( 
.A(n_2056),
.Y(n_2465)
);

INVx2_ASAP7_75t_L g2466 ( 
.A(n_2057),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2305),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2308),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2308),
.Y(n_2469)
);

AND2x6_ASAP7_75t_L g2470 ( 
.A(n_2304),
.B(n_1912),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_SL g2471 ( 
.A(n_2030),
.B(n_2042),
.Y(n_2471)
);

AND2x6_ASAP7_75t_L g2472 ( 
.A(n_2309),
.B(n_1926),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2147),
.Y(n_2473)
);

NOR2xp33_ASAP7_75t_L g2474 ( 
.A(n_2067),
.B(n_1901),
.Y(n_2474)
);

NOR2xp33_ASAP7_75t_L g2475 ( 
.A(n_2052),
.B(n_1901),
.Y(n_2475)
);

NOR2xp33_ASAP7_75t_L g2476 ( 
.A(n_2029),
.B(n_1913),
.Y(n_2476)
);

INVx2_ASAP7_75t_SL g2477 ( 
.A(n_2036),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2147),
.Y(n_2478)
);

NOR2xp33_ASAP7_75t_L g2479 ( 
.A(n_2076),
.B(n_1913),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_SL g2480 ( 
.A(n_2114),
.B(n_1926),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_SL g2481 ( 
.A(n_2218),
.B(n_1926),
.Y(n_2481)
);

INVx3_ASAP7_75t_L g2482 ( 
.A(n_2059),
.Y(n_2482)
);

INVx4_ASAP7_75t_L g2483 ( 
.A(n_2091),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_2103),
.Y(n_2484)
);

INVx2_ASAP7_75t_L g2485 ( 
.A(n_2121),
.Y(n_2485)
);

NAND2x1p5_ASAP7_75t_L g2486 ( 
.A(n_2124),
.B(n_1958),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2140),
.Y(n_2487)
);

AND2x6_ASAP7_75t_L g2488 ( 
.A(n_2243),
.B(n_1926),
.Y(n_2488)
);

BUFx3_ASAP7_75t_L g2489 ( 
.A(n_2110),
.Y(n_2489)
);

AOI22xp33_ASAP7_75t_SL g2490 ( 
.A1(n_2102),
.A2(n_1977),
.B1(n_1845),
.B2(n_1872),
.Y(n_2490)
);

INVx4_ASAP7_75t_L g2491 ( 
.A(n_2158),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_2162),
.Y(n_2492)
);

OR2x2_ASAP7_75t_L g2493 ( 
.A(n_2037),
.B(n_1730),
.Y(n_2493)
);

INVx3_ASAP7_75t_L g2494 ( 
.A(n_2169),
.Y(n_2494)
);

BUFx6f_ASAP7_75t_L g2495 ( 
.A(n_2175),
.Y(n_2495)
);

BUFx6f_ASAP7_75t_L g2496 ( 
.A(n_2180),
.Y(n_2496)
);

INVx2_ASAP7_75t_SL g2497 ( 
.A(n_2146),
.Y(n_2497)
);

AND2x4_ASAP7_75t_L g2498 ( 
.A(n_2228),
.B(n_1845),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2182),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_SL g2500 ( 
.A(n_2235),
.B(n_1701),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_2194),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2219),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2234),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2242),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_SL g2505 ( 
.A(n_2250),
.B(n_1876),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2272),
.Y(n_2506)
);

INVx3_ASAP7_75t_L g2507 ( 
.A(n_2310),
.Y(n_2507)
);

INVx3_ASAP7_75t_L g2508 ( 
.A(n_2266),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_SL g2509 ( 
.A(n_2230),
.B(n_1845),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2222),
.Y(n_2510)
);

INVx4_ASAP7_75t_L g2511 ( 
.A(n_2165),
.Y(n_2511)
);

INVx3_ASAP7_75t_L g2512 ( 
.A(n_2222),
.Y(n_2512)
);

AND2x2_ASAP7_75t_L g2513 ( 
.A(n_2197),
.B(n_1730),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2223),
.Y(n_2514)
);

INVx2_ASAP7_75t_L g2515 ( 
.A(n_2223),
.Y(n_2515)
);

OA22x2_ASAP7_75t_L g2516 ( 
.A1(n_2137),
.A2(n_1872),
.B1(n_1796),
.B2(n_1803),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_SL g2517 ( 
.A(n_2240),
.B(n_1872),
.Y(n_2517)
);

INVx2_ASAP7_75t_L g2518 ( 
.A(n_2247),
.Y(n_2518)
);

AOI22xp5_ASAP7_75t_L g2519 ( 
.A1(n_2227),
.A2(n_1731),
.B1(n_1767),
.B2(n_1797),
.Y(n_2519)
);

OAI22xp5_ASAP7_75t_L g2520 ( 
.A1(n_2072),
.A2(n_1767),
.B1(n_1731),
.B2(n_1764),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2247),
.Y(n_2521)
);

OR2x6_ASAP7_75t_L g2522 ( 
.A(n_2106),
.B(n_1886),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_SL g2523 ( 
.A(n_2244),
.B(n_1903),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2155),
.B(n_1730),
.Y(n_2524)
);

AOI22xp33_ASAP7_75t_L g2525 ( 
.A1(n_2116),
.A2(n_2268),
.B1(n_2269),
.B2(n_2261),
.Y(n_2525)
);

INVx3_ASAP7_75t_L g2526 ( 
.A(n_2264),
.Y(n_2526)
);

BUFx2_ASAP7_75t_L g2527 ( 
.A(n_2225),
.Y(n_2527)
);

BUFx3_ASAP7_75t_L g2528 ( 
.A(n_2025),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_SL g2529 ( 
.A(n_2248),
.B(n_2260),
.Y(n_2529)
);

NOR2xp33_ASAP7_75t_L g2530 ( 
.A(n_2112),
.B(n_1886),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_SL g2531 ( 
.A(n_2263),
.B(n_1810),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_SL g2532 ( 
.A(n_2122),
.B(n_1821),
.Y(n_2532)
);

INVx5_ASAP7_75t_L g2533 ( 
.A(n_2283),
.Y(n_2533)
);

OAI22xp33_ASAP7_75t_L g2534 ( 
.A1(n_2078),
.A2(n_1836),
.B1(n_1838),
.B2(n_1821),
.Y(n_2534)
);

AND2x2_ASAP7_75t_L g2535 ( 
.A(n_2201),
.B(n_1898),
.Y(n_2535)
);

INVx1_ASAP7_75t_SL g2536 ( 
.A(n_2062),
.Y(n_2536)
);

NAND3xp33_ASAP7_75t_L g2537 ( 
.A(n_2189),
.B(n_1707),
.C(n_1703),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2285),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_SL g2539 ( 
.A(n_2298),
.B(n_1836),
.Y(n_2539)
);

NAND3xp33_ASAP7_75t_L g2540 ( 
.A(n_2262),
.B(n_1709),
.C(n_1708),
.Y(n_2540)
);

BUFx8_ASAP7_75t_SL g2541 ( 
.A(n_2060),
.Y(n_2541)
);

AOI22xp5_ASAP7_75t_L g2542 ( 
.A1(n_2208),
.A2(n_2211),
.B1(n_2306),
.B2(n_2291),
.Y(n_2542)
);

INVx2_ASAP7_75t_L g2543 ( 
.A(n_2165),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_2292),
.B(n_1838),
.Y(n_2544)
);

AOI22xp33_ASAP7_75t_L g2545 ( 
.A1(n_2261),
.A2(n_2269),
.B1(n_2268),
.B2(n_2303),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2185),
.Y(n_2546)
);

INVx2_ASAP7_75t_L g2547 ( 
.A(n_2185),
.Y(n_2547)
);

BUFx3_ASAP7_75t_L g2548 ( 
.A(n_2060),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_L g2549 ( 
.A(n_2296),
.B(n_1839),
.Y(n_2549)
);

AND2x2_ASAP7_75t_SL g2550 ( 
.A(n_2237),
.B(n_1958),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2160),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_2134),
.B(n_1839),
.Y(n_2552)
);

INVx2_ASAP7_75t_L g2553 ( 
.A(n_2192),
.Y(n_2553)
);

NOR2xp33_ASAP7_75t_L g2554 ( 
.A(n_2028),
.B(n_1924),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_2192),
.Y(n_2555)
);

INVx3_ASAP7_75t_L g2556 ( 
.A(n_2210),
.Y(n_2556)
);

INVx3_ASAP7_75t_L g2557 ( 
.A(n_2215),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2181),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2183),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2215),
.Y(n_2560)
);

AOI22xp5_ASAP7_75t_L g2561 ( 
.A1(n_2196),
.A2(n_1767),
.B1(n_1811),
.B2(n_1797),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_2220),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2220),
.Y(n_2563)
);

NAND3xp33_ASAP7_75t_L g2564 ( 
.A(n_2299),
.B(n_1714),
.C(n_1713),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2174),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_SL g2566 ( 
.A(n_2064),
.B(n_1847),
.Y(n_2566)
);

INVx2_ASAP7_75t_L g2567 ( 
.A(n_2231),
.Y(n_2567)
);

OAI22xp33_ASAP7_75t_L g2568 ( 
.A1(n_2081),
.A2(n_2249),
.B1(n_2255),
.B2(n_2252),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2186),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2188),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_2231),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2163),
.Y(n_2572)
);

INVx2_ASAP7_75t_L g2573 ( 
.A(n_2191),
.Y(n_2573)
);

INVx3_ASAP7_75t_L g2574 ( 
.A(n_2251),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2251),
.Y(n_2575)
);

BUFx3_ASAP7_75t_L g2576 ( 
.A(n_2106),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_L g2577 ( 
.A(n_2117),
.B(n_1847),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2265),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2275),
.Y(n_2579)
);

NAND2xp5_ASAP7_75t_SL g2580 ( 
.A(n_2034),
.B(n_1850),
.Y(n_2580)
);

NAND3xp33_ASAP7_75t_L g2581 ( 
.A(n_2082),
.B(n_1723),
.C(n_1719),
.Y(n_2581)
);

INVx2_ASAP7_75t_L g2582 ( 
.A(n_2198),
.Y(n_2582)
);

INVx3_ASAP7_75t_L g2583 ( 
.A(n_2126),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_L g2584 ( 
.A(n_2131),
.B(n_1850),
.Y(n_2584)
);

AND2x4_ASAP7_75t_L g2585 ( 
.A(n_2123),
.B(n_1851),
.Y(n_2585)
);

AND2x6_ASAP7_75t_L g2586 ( 
.A(n_2257),
.B(n_1851),
.Y(n_2586)
);

INVx2_ASAP7_75t_L g2587 ( 
.A(n_2202),
.Y(n_2587)
);

INVx4_ASAP7_75t_L g2588 ( 
.A(n_2303),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_L g2589 ( 
.A(n_2145),
.B(n_1861),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_L g2590 ( 
.A(n_2149),
.B(n_1861),
.Y(n_2590)
);

INVx1_ASAP7_75t_SL g2591 ( 
.A(n_2083),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2195),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2286),
.Y(n_2593)
);

INVx3_ASAP7_75t_L g2594 ( 
.A(n_2154),
.Y(n_2594)
);

INVx2_ASAP7_75t_L g2595 ( 
.A(n_2259),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2120),
.B(n_1865),
.Y(n_2596)
);

BUFx6f_ASAP7_75t_SL g2597 ( 
.A(n_2009),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2288),
.Y(n_2598)
);

INVx4_ASAP7_75t_L g2599 ( 
.A(n_2127),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_2129),
.B(n_1865),
.Y(n_2600)
);

INVxp67_ASAP7_75t_L g2601 ( 
.A(n_2151),
.Y(n_2601)
);

AND2x6_ASAP7_75t_L g2602 ( 
.A(n_2212),
.B(n_1874),
.Y(n_2602)
);

CKINVDCx20_ASAP7_75t_R g2603 ( 
.A(n_2135),
.Y(n_2603)
);

AO21x2_ASAP7_75t_L g2604 ( 
.A1(n_2277),
.A2(n_1792),
.B(n_1771),
.Y(n_2604)
);

INVxp33_ASAP7_75t_L g2605 ( 
.A(n_2014),
.Y(n_2605)
);

CKINVDCx5p33_ASAP7_75t_R g2606 ( 
.A(n_2156),
.Y(n_2606)
);

CKINVDCx5p33_ASAP7_75t_R g2607 ( 
.A(n_2013),
.Y(n_2607)
);

NOR2xp33_ASAP7_75t_L g2608 ( 
.A(n_2276),
.B(n_1924),
.Y(n_2608)
);

NOR2xp33_ASAP7_75t_SL g2609 ( 
.A(n_2193),
.B(n_1767),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_2118),
.B(n_1874),
.Y(n_2610)
);

AND2x2_ASAP7_75t_L g2611 ( 
.A(n_2127),
.B(n_1922),
.Y(n_2611)
);

AOI22xp33_ASAP7_75t_L g2612 ( 
.A1(n_2209),
.A2(n_1897),
.B1(n_1879),
.B2(n_1809),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_SL g2613 ( 
.A(n_2101),
.B(n_1879),
.Y(n_2613)
);

INVx4_ASAP7_75t_L g2614 ( 
.A(n_2241),
.Y(n_2614)
);

OR2x6_ASAP7_75t_L g2615 ( 
.A(n_1997),
.B(n_1897),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2307),
.Y(n_2616)
);

NOR2xp33_ASAP7_75t_L g2617 ( 
.A(n_2069),
.B(n_1783),
.Y(n_2617)
);

INVx2_ASAP7_75t_L g2618 ( 
.A(n_2259),
.Y(n_2618)
);

NOR2xp33_ASAP7_75t_L g2619 ( 
.A(n_2109),
.B(n_1812),
.Y(n_2619)
);

OR2x2_ASAP7_75t_L g2620 ( 
.A(n_2221),
.B(n_1811),
.Y(n_2620)
);

INVx2_ASAP7_75t_L g2621 ( 
.A(n_2205),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2207),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2179),
.Y(n_2623)
);

NAND2xp33_ASAP7_75t_R g2624 ( 
.A(n_1997),
.B(n_1958),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2224),
.Y(n_2625)
);

NAND2xp5_ASAP7_75t_L g2626 ( 
.A(n_2113),
.B(n_1816),
.Y(n_2626)
);

NOR2xp33_ASAP7_75t_L g2627 ( 
.A(n_2099),
.B(n_1818),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_L g2628 ( 
.A(n_2132),
.B(n_1823),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2236),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2172),
.Y(n_2630)
);

NOR2xp33_ASAP7_75t_L g2631 ( 
.A(n_2051),
.B(n_1828),
.Y(n_2631)
);

INVx2_ASAP7_75t_L g2632 ( 
.A(n_2241),
.Y(n_2632)
);

INVx2_ASAP7_75t_L g2633 ( 
.A(n_2253),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2289),
.Y(n_2634)
);

INVx3_ASAP7_75t_L g2635 ( 
.A(n_2300),
.Y(n_2635)
);

INVx4_ASAP7_75t_L g2636 ( 
.A(n_2038),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2282),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2115),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2128),
.Y(n_2639)
);

NOR2xp33_ASAP7_75t_L g2640 ( 
.A(n_2054),
.B(n_1832),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2095),
.Y(n_2641)
);

BUFx6f_ASAP7_75t_L g2642 ( 
.A(n_2203),
.Y(n_2642)
);

AND2x6_ASAP7_75t_L g2643 ( 
.A(n_2090),
.B(n_1852),
.Y(n_2643)
);

OAI22xp33_ASAP7_75t_L g2644 ( 
.A1(n_2143),
.A2(n_1842),
.B1(n_1871),
.B2(n_1840),
.Y(n_2644)
);

AND2x2_ASAP7_75t_L g2645 ( 
.A(n_2014),
.B(n_1900),
.Y(n_2645)
);

BUFx3_ASAP7_75t_L g2646 ( 
.A(n_2027),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2167),
.Y(n_2647)
);

AND2x2_ASAP7_75t_L g2648 ( 
.A(n_2027),
.B(n_1900),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_SL g2649 ( 
.A(n_2139),
.B(n_1852),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_2086),
.Y(n_2650)
);

AND2x2_ASAP7_75t_L g2651 ( 
.A(n_2048),
.B(n_1922),
.Y(n_2651)
);

AOI22xp33_ASAP7_75t_L g2652 ( 
.A1(n_2041),
.A2(n_1884),
.B1(n_1887),
.B2(n_1883),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2173),
.Y(n_2653)
);

INVx2_ASAP7_75t_L g2654 ( 
.A(n_2008),
.Y(n_2654)
);

INVx2_ASAP7_75t_L g2655 ( 
.A(n_2107),
.Y(n_2655)
);

BUFx6f_ASAP7_75t_L g2656 ( 
.A(n_2204),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2107),
.Y(n_2657)
);

BUFx6f_ASAP7_75t_L g2658 ( 
.A(n_2184),
.Y(n_2658)
);

AND2x2_ASAP7_75t_L g2659 ( 
.A(n_2048),
.B(n_1898),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2190),
.Y(n_2660)
);

NAND2xp5_ASAP7_75t_SL g2661 ( 
.A(n_2148),
.B(n_1907),
.Y(n_2661)
);

NOR2xp33_ASAP7_75t_L g2662 ( 
.A(n_2070),
.B(n_1914),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2041),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_2213),
.Y(n_2664)
);

BUFx2_ASAP7_75t_L g2665 ( 
.A(n_2077),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2233),
.Y(n_2666)
);

AND2x4_ASAP7_75t_L g2667 ( 
.A(n_2419),
.B(n_1920),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2407),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2412),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2414),
.Y(n_2670)
);

INVx2_ASAP7_75t_L g2671 ( 
.A(n_2385),
.Y(n_2671)
);

INVxp67_ASAP7_75t_L g2672 ( 
.A(n_2342),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_L g2673 ( 
.A(n_2464),
.B(n_1753),
.Y(n_2673)
);

OR2x2_ASAP7_75t_L g2674 ( 
.A(n_2314),
.B(n_2418),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2332),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2333),
.Y(n_2676)
);

BUFx6f_ASAP7_75t_L g2677 ( 
.A(n_2425),
.Y(n_2677)
);

BUFx6f_ASAP7_75t_L g2678 ( 
.A(n_2425),
.Y(n_2678)
);

INVx3_ASAP7_75t_L g2679 ( 
.A(n_2335),
.Y(n_2679)
);

INVxp67_ASAP7_75t_L g2680 ( 
.A(n_2524),
.Y(n_2680)
);

INVxp67_ASAP7_75t_L g2681 ( 
.A(n_2530),
.Y(n_2681)
);

BUFx6f_ASAP7_75t_L g2682 ( 
.A(n_2425),
.Y(n_2682)
);

INVx2_ASAP7_75t_L g2683 ( 
.A(n_2385),
.Y(n_2683)
);

INVx2_ASAP7_75t_L g2684 ( 
.A(n_2321),
.Y(n_2684)
);

NAND3xp33_ASAP7_75t_L g2685 ( 
.A(n_2315),
.B(n_2217),
.C(n_2216),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2336),
.Y(n_2686)
);

INVx6_ASAP7_75t_L g2687 ( 
.A(n_2371),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2464),
.B(n_1734),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_L g2689 ( 
.A(n_2467),
.B(n_1737),
.Y(n_2689)
);

INVx2_ASAP7_75t_SL g2690 ( 
.A(n_2317),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2341),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2344),
.Y(n_2692)
);

NAND2x1p5_ASAP7_75t_L g2693 ( 
.A(n_2425),
.B(n_1773),
.Y(n_2693)
);

OAI22xp5_ASAP7_75t_L g2694 ( 
.A1(n_2467),
.A2(n_2232),
.B1(n_2239),
.B2(n_2229),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2345),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2347),
.Y(n_2696)
);

BUFx6f_ASAP7_75t_L g2697 ( 
.A(n_2425),
.Y(n_2697)
);

AND2x2_ASAP7_75t_L g2698 ( 
.A(n_2611),
.B(n_2077),
.Y(n_2698)
);

AND2x2_ASAP7_75t_L g2699 ( 
.A(n_2611),
.B(n_2092),
.Y(n_2699)
);

HB1xp67_ASAP7_75t_L g2700 ( 
.A(n_2497),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2515),
.Y(n_2701)
);

CKINVDCx5p33_ASAP7_75t_R g2702 ( 
.A(n_2328),
.Y(n_2702)
);

INVxp67_ASAP7_75t_L g2703 ( 
.A(n_2479),
.Y(n_2703)
);

BUFx2_ASAP7_75t_L g2704 ( 
.A(n_2421),
.Y(n_2704)
);

INVx3_ASAP7_75t_L g2705 ( 
.A(n_2335),
.Y(n_2705)
);

INVx2_ASAP7_75t_L g2706 ( 
.A(n_2321),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2515),
.Y(n_2707)
);

INVx4_ASAP7_75t_SL g2708 ( 
.A(n_2387),
.Y(n_2708)
);

INVx4_ASAP7_75t_L g2709 ( 
.A(n_2317),
.Y(n_2709)
);

NAND2x1p5_ASAP7_75t_L g2710 ( 
.A(n_2419),
.B(n_2335),
.Y(n_2710)
);

INVx4_ASAP7_75t_L g2711 ( 
.A(n_2317),
.Y(n_2711)
);

INVx2_ASAP7_75t_L g2712 ( 
.A(n_2326),
.Y(n_2712)
);

AND2x2_ASAP7_75t_L g2713 ( 
.A(n_2356),
.B(n_2092),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2518),
.Y(n_2714)
);

AND2x2_ASAP7_75t_L g2715 ( 
.A(n_2356),
.B(n_2010),
.Y(n_2715)
);

BUFx6f_ASAP7_75t_L g2716 ( 
.A(n_2380),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2518),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2521),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2326),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2521),
.Y(n_2720)
);

INVx2_ASAP7_75t_L g2721 ( 
.A(n_2354),
.Y(n_2721)
);

AND2x4_ASAP7_75t_L g2722 ( 
.A(n_2380),
.B(n_1741),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2354),
.Y(n_2723)
);

NAND2x1p5_ASAP7_75t_L g2724 ( 
.A(n_2384),
.B(n_1773),
.Y(n_2724)
);

NAND2x1p5_ASAP7_75t_L g2725 ( 
.A(n_2384),
.B(n_1773),
.Y(n_2725)
);

AND2x4_ASAP7_75t_L g2726 ( 
.A(n_2380),
.B(n_1743),
.Y(n_2726)
);

INVx2_ASAP7_75t_SL g2727 ( 
.A(n_2317),
.Y(n_2727)
);

AND2x4_ASAP7_75t_L g2728 ( 
.A(n_2386),
.B(n_1766),
.Y(n_2728)
);

AND2x4_ASAP7_75t_L g2729 ( 
.A(n_2436),
.B(n_1780),
.Y(n_2729)
);

BUFx3_ASAP7_75t_L g2730 ( 
.A(n_2320),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2361),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2361),
.Y(n_2732)
);

INVx2_ASAP7_75t_L g2733 ( 
.A(n_2366),
.Y(n_2733)
);

AND2x4_ASAP7_75t_L g2734 ( 
.A(n_2436),
.B(n_1785),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2366),
.Y(n_2735)
);

AND2x2_ASAP7_75t_L g2736 ( 
.A(n_2601),
.B(n_2010),
.Y(n_2736)
);

INVx2_ASAP7_75t_L g2737 ( 
.A(n_2367),
.Y(n_2737)
);

BUFx6f_ASAP7_75t_L g2738 ( 
.A(n_2384),
.Y(n_2738)
);

BUFx6f_ASAP7_75t_L g2739 ( 
.A(n_2444),
.Y(n_2739)
);

AO22x2_ASAP7_75t_L g2740 ( 
.A1(n_2614),
.A2(n_2246),
.B1(n_2267),
.B2(n_2256),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2367),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2381),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_2381),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2468),
.B(n_1885),
.Y(n_2744)
);

BUFx6f_ASAP7_75t_L g2745 ( 
.A(n_2444),
.Y(n_2745)
);

NOR2xp33_ASAP7_75t_L g2746 ( 
.A(n_2409),
.B(n_2080),
.Y(n_2746)
);

HB1xp67_ASAP7_75t_L g2747 ( 
.A(n_2497),
.Y(n_2747)
);

BUFx2_ASAP7_75t_L g2748 ( 
.A(n_2421),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_L g2749 ( 
.A(n_2468),
.B(n_2469),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_L g2750 ( 
.A(n_2469),
.B(n_1800),
.Y(n_2750)
);

CKINVDCx5p33_ASAP7_75t_R g2751 ( 
.A(n_2328),
.Y(n_2751)
);

AO22x2_ASAP7_75t_L g2752 ( 
.A1(n_2614),
.A2(n_2280),
.B1(n_2290),
.B2(n_2273),
.Y(n_2752)
);

BUFx3_ASAP7_75t_L g2753 ( 
.A(n_2320),
.Y(n_2753)
);

OR2x2_ASAP7_75t_SL g2754 ( 
.A(n_2322),
.B(n_2294),
.Y(n_2754)
);

AND2x6_ASAP7_75t_L g2755 ( 
.A(n_2557),
.B(n_1785),
.Y(n_2755)
);

AND2x4_ASAP7_75t_SL g2756 ( 
.A(n_2371),
.B(n_1785),
.Y(n_2756)
);

BUFx6f_ASAP7_75t_L g2757 ( 
.A(n_2454),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_2382),
.Y(n_2758)
);

OAI22xp33_ASAP7_75t_L g2759 ( 
.A1(n_2588),
.A2(n_1795),
.B1(n_1862),
.B2(n_1827),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_2473),
.B(n_1870),
.Y(n_2760)
);

AND2x2_ASAP7_75t_L g2761 ( 
.A(n_2599),
.B(n_2423),
.Y(n_2761)
);

INVxp67_ASAP7_75t_SL g2762 ( 
.A(n_2311),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2382),
.Y(n_2763)
);

AND2x2_ASAP7_75t_L g2764 ( 
.A(n_2599),
.B(n_1779),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2388),
.Y(n_2765)
);

NOR2xp33_ASAP7_75t_L g2766 ( 
.A(n_2409),
.B(n_2430),
.Y(n_2766)
);

INVx2_ASAP7_75t_L g2767 ( 
.A(n_2388),
.Y(n_2767)
);

NOR2xp33_ASAP7_75t_L g2768 ( 
.A(n_2606),
.B(n_1873),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2389),
.Y(n_2769)
);

BUFx6f_ASAP7_75t_L g2770 ( 
.A(n_2454),
.Y(n_2770)
);

AND2x4_ASAP7_75t_L g2771 ( 
.A(n_2436),
.B(n_1700),
.Y(n_2771)
);

INVx2_ASAP7_75t_L g2772 ( 
.A(n_2389),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2391),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2391),
.Y(n_2774)
);

AND3x4_ASAP7_75t_L g2775 ( 
.A(n_2489),
.B(n_71),
.C(n_72),
.Y(n_2775)
);

INVx2_ASAP7_75t_L g2776 ( 
.A(n_2393),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2393),
.Y(n_2777)
);

INVxp67_ASAP7_75t_L g2778 ( 
.A(n_2314),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2403),
.Y(n_2779)
);

HB1xp67_ASAP7_75t_L g2780 ( 
.A(n_2423),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2404),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2355),
.Y(n_2782)
);

INVxp67_ASAP7_75t_L g2783 ( 
.A(n_2346),
.Y(n_2783)
);

CKINVDCx5p33_ASAP7_75t_R g2784 ( 
.A(n_2541),
.Y(n_2784)
);

BUFx6f_ASAP7_75t_L g2785 ( 
.A(n_2454),
.Y(n_2785)
);

AND2x2_ASAP7_75t_SL g2786 ( 
.A(n_2525),
.B(n_1779),
.Y(n_2786)
);

AND2x2_ASAP7_75t_L g2787 ( 
.A(n_2599),
.B(n_1779),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2363),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2417),
.Y(n_2789)
);

INVx2_ASAP7_75t_L g2790 ( 
.A(n_2311),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2446),
.Y(n_2791)
);

HB1xp67_ASAP7_75t_L g2792 ( 
.A(n_2392),
.Y(n_2792)
);

INVx2_ASAP7_75t_SL g2793 ( 
.A(n_2357),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2473),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2478),
.Y(n_2795)
);

NAND2x1p5_ASAP7_75t_L g2796 ( 
.A(n_2323),
.B(n_1774),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2478),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_2510),
.B(n_1882),
.Y(n_2798)
);

NOR2xp33_ASAP7_75t_L g2799 ( 
.A(n_2606),
.B(n_1700),
.Y(n_2799)
);

AND2x2_ASAP7_75t_SL g2800 ( 
.A(n_2545),
.B(n_1774),
.Y(n_2800)
);

NOR2xp33_ASAP7_75t_L g2801 ( 
.A(n_2455),
.B(n_1700),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2510),
.Y(n_2802)
);

INVx4_ASAP7_75t_L g2803 ( 
.A(n_2357),
.Y(n_2803)
);

OAI22xp33_ASAP7_75t_L g2804 ( 
.A1(n_2588),
.A2(n_1768),
.B1(n_1759),
.B2(n_73),
.Y(n_2804)
);

NAND2xp5_ASAP7_75t_L g2805 ( 
.A(n_2514),
.B(n_1735),
.Y(n_2805)
);

AND2x2_ASAP7_75t_L g2806 ( 
.A(n_2392),
.B(n_1735),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2514),
.Y(n_2807)
);

INVx2_ASAP7_75t_L g2808 ( 
.A(n_2312),
.Y(n_2808)
);

INVx2_ASAP7_75t_L g2809 ( 
.A(n_2312),
.Y(n_2809)
);

BUFx2_ASAP7_75t_L g2810 ( 
.A(n_2527),
.Y(n_2810)
);

INVx3_ASAP7_75t_L g2811 ( 
.A(n_2399),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2557),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_L g2813 ( 
.A(n_2512),
.B(n_1757),
.Y(n_2813)
);

NAND3xp33_ASAP7_75t_L g2814 ( 
.A(n_2340),
.B(n_1768),
.C(n_1759),
.Y(n_2814)
);

AND2x6_ASAP7_75t_L g2815 ( 
.A(n_2557),
.B(n_1774),
.Y(n_2815)
);

AND2x4_ASAP7_75t_L g2816 ( 
.A(n_2436),
.B(n_1759),
.Y(n_2816)
);

INVx2_ASAP7_75t_L g2817 ( 
.A(n_2334),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2546),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2546),
.Y(n_2819)
);

AOI22xp5_ASAP7_75t_L g2820 ( 
.A1(n_2609),
.A2(n_1768),
.B1(n_1790),
.B2(n_1774),
.Y(n_2820)
);

AND2x2_ASAP7_75t_L g2821 ( 
.A(n_2411),
.B(n_1757),
.Y(n_2821)
);

AND2x4_ASAP7_75t_L g2822 ( 
.A(n_2372),
.B(n_1775),
.Y(n_2822)
);

BUFx6f_ASAP7_75t_L g2823 ( 
.A(n_2454),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_2512),
.B(n_1761),
.Y(n_2824)
);

BUFx6f_ASAP7_75t_L g2825 ( 
.A(n_2454),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2547),
.Y(n_2826)
);

INVx2_ASAP7_75t_L g2827 ( 
.A(n_2334),
.Y(n_2827)
);

AND2x4_ASAP7_75t_L g2828 ( 
.A(n_2372),
.B(n_1775),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2547),
.Y(n_2829)
);

INVx2_ASAP7_75t_L g2830 ( 
.A(n_2348),
.Y(n_2830)
);

NAND2x1p5_ASAP7_75t_L g2831 ( 
.A(n_2323),
.B(n_1774),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2553),
.Y(n_2832)
);

NAND2x1p5_ASAP7_75t_L g2833 ( 
.A(n_2323),
.B(n_1790),
.Y(n_2833)
);

OAI22xp5_ASAP7_75t_L g2834 ( 
.A1(n_2634),
.A2(n_1781),
.B1(n_1761),
.B2(n_1790),
.Y(n_2834)
);

INVx3_ASAP7_75t_L g2835 ( 
.A(n_2399),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2553),
.Y(n_2836)
);

HB1xp67_ASAP7_75t_L g2837 ( 
.A(n_2411),
.Y(n_2837)
);

AND2x2_ASAP7_75t_L g2838 ( 
.A(n_2535),
.B(n_1781),
.Y(n_2838)
);

OR2x2_ASAP7_75t_SL g2839 ( 
.A(n_2364),
.B(n_2434),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2555),
.Y(n_2840)
);

INVxp67_ASAP7_75t_L g2841 ( 
.A(n_2349),
.Y(n_2841)
);

BUFx6f_ASAP7_75t_L g2842 ( 
.A(n_2463),
.Y(n_2842)
);

NOR2x1p5_ASAP7_75t_L g2843 ( 
.A(n_2405),
.B(n_1717),
.Y(n_2843)
);

AND2x2_ASAP7_75t_L g2844 ( 
.A(n_2535),
.B(n_71),
.Y(n_2844)
);

OAI221xp5_ASAP7_75t_L g2845 ( 
.A1(n_2401),
.A2(n_1790),
.B1(n_1742),
.B2(n_1751),
.C(n_1724),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2555),
.Y(n_2846)
);

INVx2_ASAP7_75t_SL g2847 ( 
.A(n_2405),
.Y(n_2847)
);

NOR2xp33_ASAP7_75t_R g2848 ( 
.A(n_2331),
.B(n_1790),
.Y(n_2848)
);

INVx2_ASAP7_75t_L g2849 ( 
.A(n_2348),
.Y(n_2849)
);

BUFx2_ASAP7_75t_L g2850 ( 
.A(n_2527),
.Y(n_2850)
);

INVx2_ASAP7_75t_L g2851 ( 
.A(n_2350),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2560),
.Y(n_2852)
);

INVx2_ASAP7_75t_L g2853 ( 
.A(n_2350),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_L g2854 ( 
.A(n_2512),
.B(n_1717),
.Y(n_2854)
);

BUFx3_ASAP7_75t_L g2855 ( 
.A(n_2371),
.Y(n_2855)
);

AND2x4_ASAP7_75t_L g2856 ( 
.A(n_2439),
.B(n_1747),
.Y(n_2856)
);

BUFx2_ASAP7_75t_L g2857 ( 
.A(n_2327),
.Y(n_2857)
);

AND2x4_ASAP7_75t_L g2858 ( 
.A(n_2439),
.B(n_2424),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2560),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2562),
.Y(n_2860)
);

AND2x4_ASAP7_75t_L g2861 ( 
.A(n_2424),
.B(n_1747),
.Y(n_2861)
);

NOR2xp33_ASAP7_75t_L g2862 ( 
.A(n_2313),
.B(n_1717),
.Y(n_2862)
);

AND2x6_ASAP7_75t_L g2863 ( 
.A(n_2562),
.B(n_1717),
.Y(n_2863)
);

AND2x4_ASAP7_75t_L g2864 ( 
.A(n_2400),
.B(n_1747),
.Y(n_2864)
);

INVx2_ASAP7_75t_L g2865 ( 
.A(n_2362),
.Y(n_2865)
);

AND2x2_ASAP7_75t_L g2866 ( 
.A(n_2536),
.B(n_72),
.Y(n_2866)
);

AND2x4_ASAP7_75t_L g2867 ( 
.A(n_2400),
.B(n_1747),
.Y(n_2867)
);

INVx4_ASAP7_75t_SL g2868 ( 
.A(n_2387),
.Y(n_2868)
);

BUFx4f_ASAP7_75t_L g2869 ( 
.A(n_2522),
.Y(n_2869)
);

AND2x4_ASAP7_75t_L g2870 ( 
.A(n_2413),
.B(n_1747),
.Y(n_2870)
);

AND2x2_ASAP7_75t_L g2871 ( 
.A(n_2591),
.B(n_2645),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2563),
.Y(n_2872)
);

INVx2_ASAP7_75t_L g2873 ( 
.A(n_2362),
.Y(n_2873)
);

AND2x4_ASAP7_75t_L g2874 ( 
.A(n_2413),
.B(n_1717),
.Y(n_2874)
);

INVx2_ASAP7_75t_L g2875 ( 
.A(n_2365),
.Y(n_2875)
);

INVx1_ASAP7_75t_SL g2876 ( 
.A(n_2513),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2563),
.Y(n_2877)
);

AOI22xp33_ASAP7_75t_L g2878 ( 
.A1(n_2614),
.A2(n_1742),
.B1(n_1751),
.B2(n_1724),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2567),
.Y(n_2879)
);

AOI22xp5_ASAP7_75t_L g2880 ( 
.A1(n_2603),
.A2(n_1742),
.B1(n_1751),
.B2(n_1724),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2567),
.Y(n_2881)
);

INVx2_ASAP7_75t_L g2882 ( 
.A(n_2365),
.Y(n_2882)
);

AOI22xp5_ASAP7_75t_L g2883 ( 
.A1(n_2603),
.A2(n_1742),
.B1(n_1751),
.B2(n_1724),
.Y(n_2883)
);

BUFx3_ASAP7_75t_L g2884 ( 
.A(n_2489),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2571),
.Y(n_2885)
);

BUFx6f_ASAP7_75t_L g2886 ( 
.A(n_2463),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2571),
.Y(n_2887)
);

CKINVDCx8_ASAP7_75t_R g2888 ( 
.A(n_2522),
.Y(n_2888)
);

AND2x4_ASAP7_75t_L g2889 ( 
.A(n_2415),
.B(n_1724),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2487),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2487),
.Y(n_2891)
);

INVx3_ASAP7_75t_L g2892 ( 
.A(n_2399),
.Y(n_2892)
);

NAND2x1p5_ASAP7_75t_L g2893 ( 
.A(n_2337),
.B(n_1742),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2459),
.B(n_1751),
.Y(n_2894)
);

AO21x2_ASAP7_75t_L g2895 ( 
.A1(n_2420),
.A2(n_1765),
.B(n_1756),
.Y(n_2895)
);

INVx4_ASAP7_75t_L g2896 ( 
.A(n_2360),
.Y(n_2896)
);

CKINVDCx5p33_ASAP7_75t_R g2897 ( 
.A(n_2541),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2499),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2499),
.Y(n_2899)
);

INVx1_ASAP7_75t_SL g2900 ( 
.A(n_2513),
.Y(n_2900)
);

NAND2x1p5_ASAP7_75t_L g2901 ( 
.A(n_2337),
.B(n_1756),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_2375),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_L g2903 ( 
.A(n_2625),
.B(n_1756),
.Y(n_2903)
);

INVxp67_ASAP7_75t_L g2904 ( 
.A(n_2643),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2502),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2502),
.Y(n_2906)
);

BUFx6f_ASAP7_75t_L g2907 ( 
.A(n_2463),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_L g2908 ( 
.A(n_2625),
.B(n_1756),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2504),
.Y(n_2909)
);

INVx2_ASAP7_75t_SL g2910 ( 
.A(n_2398),
.Y(n_2910)
);

AND2x4_ASAP7_75t_L g2911 ( 
.A(n_2415),
.B(n_1756),
.Y(n_2911)
);

CKINVDCx20_ASAP7_75t_R g2912 ( 
.A(n_2449),
.Y(n_2912)
);

AND2x2_ASAP7_75t_L g2913 ( 
.A(n_2645),
.B(n_73),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_L g2914 ( 
.A(n_2629),
.B(n_1765),
.Y(n_2914)
);

AND2x4_ASAP7_75t_L g2915 ( 
.A(n_2477),
.B(n_1765),
.Y(n_2915)
);

BUFx6f_ASAP7_75t_L g2916 ( 
.A(n_2463),
.Y(n_2916)
);

AND2x2_ASAP7_75t_L g2917 ( 
.A(n_2648),
.B(n_2659),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2504),
.Y(n_2918)
);

HB1xp67_ASAP7_75t_L g2919 ( 
.A(n_2477),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2506),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2506),
.Y(n_2921)
);

INVx4_ASAP7_75t_L g2922 ( 
.A(n_2449),
.Y(n_2922)
);

INVx2_ASAP7_75t_L g2923 ( 
.A(n_2375),
.Y(n_2923)
);

OAI22xp33_ASAP7_75t_L g2924 ( 
.A1(n_2588),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_2924)
);

INVx4_ASAP7_75t_L g2925 ( 
.A(n_2522),
.Y(n_2925)
);

NOR2xp33_ASAP7_75t_L g2926 ( 
.A(n_2493),
.B(n_1765),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2451),
.Y(n_2927)
);

AND2x4_ASAP7_75t_L g2928 ( 
.A(n_2574),
.B(n_1765),
.Y(n_2928)
);

OR2x2_ASAP7_75t_SL g2929 ( 
.A(n_2434),
.B(n_74),
.Y(n_2929)
);

AOI22xp5_ASAP7_75t_L g2930 ( 
.A1(n_2471),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_2930)
);

INVx2_ASAP7_75t_L g2931 ( 
.A(n_2376),
.Y(n_2931)
);

INVxp67_ASAP7_75t_L g2932 ( 
.A(n_2643),
.Y(n_2932)
);

AND2x4_ASAP7_75t_L g2933 ( 
.A(n_2574),
.B(n_75),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2453),
.Y(n_2934)
);

BUFx6f_ASAP7_75t_L g2935 ( 
.A(n_2463),
.Y(n_2935)
);

OAI22xp33_ASAP7_75t_SL g2936 ( 
.A1(n_2632),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_2629),
.B(n_76),
.Y(n_2937)
);

AND2x4_ASAP7_75t_L g2938 ( 
.A(n_2574),
.B(n_2498),
.Y(n_2938)
);

INVx2_ASAP7_75t_L g2939 ( 
.A(n_2376),
.Y(n_2939)
);

INVx4_ASAP7_75t_L g2940 ( 
.A(n_2522),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2456),
.Y(n_2941)
);

OAI22xp5_ASAP7_75t_L g2942 ( 
.A1(n_2634),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_2942)
);

INVx2_ASAP7_75t_L g2943 ( 
.A(n_2383),
.Y(n_2943)
);

INVx2_ASAP7_75t_L g2944 ( 
.A(n_2383),
.Y(n_2944)
);

INVx2_ASAP7_75t_L g2945 ( 
.A(n_2448),
.Y(n_2945)
);

NAND2x1p5_ASAP7_75t_L g2946 ( 
.A(n_2337),
.B(n_79),
.Y(n_2946)
);

BUFx6f_ASAP7_75t_L g2947 ( 
.A(n_2495),
.Y(n_2947)
);

BUFx2_ASAP7_75t_L g2948 ( 
.A(n_2528),
.Y(n_2948)
);

AND2x4_ASAP7_75t_L g2949 ( 
.A(n_2498),
.B(n_79),
.Y(n_2949)
);

INVx2_ASAP7_75t_SL g2950 ( 
.A(n_2528),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2448),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2452),
.Y(n_2952)
);

AND2x6_ASAP7_75t_L g2953 ( 
.A(n_2642),
.B(n_80),
.Y(n_2953)
);

NAND2x1p5_ASAP7_75t_L g2954 ( 
.A(n_2338),
.B(n_80),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_SL g2955 ( 
.A(n_2550),
.B(n_224),
.Y(n_2955)
);

BUFx2_ASAP7_75t_L g2956 ( 
.A(n_2548),
.Y(n_2956)
);

INVx2_ASAP7_75t_L g2957 ( 
.A(n_2452),
.Y(n_2957)
);

INVx2_ASAP7_75t_L g2958 ( 
.A(n_2465),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2465),
.Y(n_2959)
);

AND2x2_ASAP7_75t_L g2960 ( 
.A(n_2778),
.B(n_2648),
.Y(n_2960)
);

NAND2xp5_ASAP7_75t_SL g2961 ( 
.A(n_2703),
.B(n_2351),
.Y(n_2961)
);

AOI22xp33_ASAP7_75t_L g2962 ( 
.A1(n_2800),
.A2(n_2615),
.B1(n_2646),
.B2(n_2605),
.Y(n_2962)
);

INVx3_ASAP7_75t_L g2963 ( 
.A(n_2815),
.Y(n_2963)
);

NAND2xp5_ASAP7_75t_L g2964 ( 
.A(n_2766),
.B(n_2387),
.Y(n_2964)
);

INVx1_ASAP7_75t_L g2965 ( 
.A(n_2789),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_L g2966 ( 
.A(n_2766),
.B(n_2387),
.Y(n_2966)
);

NOR2xp33_ASAP7_75t_L g2967 ( 
.A(n_2768),
.B(n_2351),
.Y(n_2967)
);

AOI22xp33_ASAP7_75t_L g2968 ( 
.A1(n_2800),
.A2(n_2615),
.B1(n_2646),
.B2(n_2605),
.Y(n_2968)
);

NAND2xp5_ASAP7_75t_L g2969 ( 
.A(n_2749),
.B(n_2387),
.Y(n_2969)
);

INVx2_ASAP7_75t_L g2970 ( 
.A(n_2671),
.Y(n_2970)
);

NOR2xp33_ASAP7_75t_L g2971 ( 
.A(n_2768),
.B(n_2351),
.Y(n_2971)
);

OR2x2_ASAP7_75t_L g2972 ( 
.A(n_2778),
.B(n_2493),
.Y(n_2972)
);

NOR2xp33_ASAP7_75t_L g2973 ( 
.A(n_2799),
.B(n_2329),
.Y(n_2973)
);

AOI22xp5_ASAP7_75t_L g2974 ( 
.A1(n_2685),
.A2(n_2406),
.B1(n_2568),
.B2(n_2329),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_SL g2975 ( 
.A(n_2703),
.B(n_2373),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2791),
.Y(n_2976)
);

AOI22xp33_ASAP7_75t_SL g2977 ( 
.A1(n_2752),
.A2(n_2665),
.B1(n_2651),
.B2(n_2659),
.Y(n_2977)
);

NAND2xp5_ASAP7_75t_L g2978 ( 
.A(n_2749),
.B(n_2387),
.Y(n_2978)
);

INVx2_ASAP7_75t_SL g2979 ( 
.A(n_2687),
.Y(n_2979)
);

INVx8_ASAP7_75t_L g2980 ( 
.A(n_2815),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_2801),
.B(n_2762),
.Y(n_2981)
);

NAND2x1_ASAP7_75t_L g2982 ( 
.A(n_2811),
.B(n_2368),
.Y(n_2982)
);

AOI22xp5_ASAP7_75t_L g2983 ( 
.A1(n_2685),
.A2(n_2542),
.B1(n_2378),
.B2(n_2597),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_L g2984 ( 
.A(n_2801),
.B(n_2762),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_L g2985 ( 
.A(n_2688),
.B(n_2586),
.Y(n_2985)
);

NAND2xp33_ASAP7_75t_SL g2986 ( 
.A(n_2803),
.B(n_2324),
.Y(n_2986)
);

BUFx6f_ASAP7_75t_L g2987 ( 
.A(n_2716),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_L g2988 ( 
.A(n_2681),
.B(n_2474),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_L g2989 ( 
.A(n_2681),
.B(n_2476),
.Y(n_2989)
);

INVx2_ASAP7_75t_L g2990 ( 
.A(n_2683),
.Y(n_2990)
);

AOI22xp5_ASAP7_75t_L g2991 ( 
.A1(n_2799),
.A2(n_2752),
.B1(n_2728),
.B2(n_2694),
.Y(n_2991)
);

INVx2_ASAP7_75t_L g2992 ( 
.A(n_2684),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2668),
.Y(n_2993)
);

AOI22xp5_ASAP7_75t_L g2994 ( 
.A1(n_2752),
.A2(n_2597),
.B1(n_2594),
.B2(n_2583),
.Y(n_2994)
);

AOI22xp33_ASAP7_75t_L g2995 ( 
.A1(n_2871),
.A2(n_2615),
.B1(n_2490),
.B2(n_2651),
.Y(n_2995)
);

NAND2xp5_ASAP7_75t_L g2996 ( 
.A(n_2680),
.B(n_2608),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2680),
.B(n_2572),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2779),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_SL g2999 ( 
.A(n_2728),
.B(n_2428),
.Y(n_2999)
);

BUFx3_ASAP7_75t_L g3000 ( 
.A(n_2730),
.Y(n_3000)
);

NAND2xp5_ASAP7_75t_L g3001 ( 
.A(n_2674),
.B(n_2627),
.Y(n_3001)
);

INVx2_ASAP7_75t_L g3002 ( 
.A(n_2706),
.Y(n_3002)
);

AND2x2_ASAP7_75t_L g3003 ( 
.A(n_2713),
.B(n_2652),
.Y(n_3003)
);

HB1xp67_ASAP7_75t_L g3004 ( 
.A(n_2672),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2781),
.Y(n_3005)
);

NOR2xp33_ASAP7_75t_L g3006 ( 
.A(n_2857),
.B(n_2566),
.Y(n_3006)
);

INVx4_ASAP7_75t_L g3007 ( 
.A(n_2709),
.Y(n_3007)
);

AND2x4_ASAP7_75t_L g3008 ( 
.A(n_2708),
.B(n_2498),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_L g3009 ( 
.A(n_2876),
.B(n_2620),
.Y(n_3009)
);

INVx2_ASAP7_75t_L g3010 ( 
.A(n_2712),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_SL g3011 ( 
.A(n_2729),
.B(n_2353),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2669),
.Y(n_3012)
);

NAND3xp33_ASAP7_75t_SL g3013 ( 
.A(n_2775),
.B(n_2607),
.C(n_2561),
.Y(n_3013)
);

NAND2xp5_ASAP7_75t_L g3014 ( 
.A(n_2876),
.B(n_2620),
.Y(n_3014)
);

OR2x6_ASAP7_75t_L g3015 ( 
.A(n_2904),
.B(n_2511),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2670),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_L g3017 ( 
.A(n_2900),
.B(n_2639),
.Y(n_3017)
);

OR2x2_ASAP7_75t_L g3018 ( 
.A(n_2839),
.B(n_2615),
.Y(n_3018)
);

BUFx4f_ASAP7_75t_L g3019 ( 
.A(n_2677),
.Y(n_3019)
);

NAND2xp5_ASAP7_75t_L g3020 ( 
.A(n_2900),
.B(n_2638),
.Y(n_3020)
);

NAND2xp5_ASAP7_75t_L g3021 ( 
.A(n_2780),
.B(n_2632),
.Y(n_3021)
);

NOR2xp33_ASAP7_75t_L g3022 ( 
.A(n_2754),
.B(n_2580),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_L g3023 ( 
.A(n_2780),
.B(n_2583),
.Y(n_3023)
);

NAND2xp5_ASAP7_75t_L g3024 ( 
.A(n_2792),
.B(n_2583),
.Y(n_3024)
);

INVx2_ASAP7_75t_L g3025 ( 
.A(n_2719),
.Y(n_3025)
);

INVxp67_ASAP7_75t_L g3026 ( 
.A(n_2704),
.Y(n_3026)
);

AOI22xp5_ASAP7_75t_L g3027 ( 
.A1(n_2694),
.A2(n_2597),
.B1(n_2594),
.B2(n_2556),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2792),
.B(n_2594),
.Y(n_3028)
);

AND2x6_ASAP7_75t_SL g3029 ( 
.A(n_2736),
.B(n_2631),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2837),
.B(n_2427),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_L g3031 ( 
.A(n_2837),
.B(n_2612),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_SL g3032 ( 
.A(n_2729),
.B(n_2475),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_2675),
.Y(n_3033)
);

INVxp67_ASAP7_75t_L g3034 ( 
.A(n_2748),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_SL g3035 ( 
.A(n_2677),
.B(n_2460),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_L g3036 ( 
.A(n_2672),
.B(n_2644),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2782),
.B(n_2369),
.Y(n_3037)
);

AND2x2_ASAP7_75t_L g3038 ( 
.A(n_2866),
.B(n_2635),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_2788),
.B(n_2617),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2676),
.Y(n_3040)
);

INVx3_ASAP7_75t_L g3041 ( 
.A(n_2815),
.Y(n_3041)
);

INVx2_ASAP7_75t_SL g3042 ( 
.A(n_2687),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_L g3043 ( 
.A(n_2688),
.B(n_2586),
.Y(n_3043)
);

OR2x2_ASAP7_75t_L g3044 ( 
.A(n_2810),
.B(n_2548),
.Y(n_3044)
);

INVx2_ASAP7_75t_L g3045 ( 
.A(n_2721),
.Y(n_3045)
);

AND2x2_ASAP7_75t_L g3046 ( 
.A(n_2844),
.B(n_2635),
.Y(n_3046)
);

NOR2xp33_ASAP7_75t_L g3047 ( 
.A(n_2850),
.B(n_2607),
.Y(n_3047)
);

AND2x2_ASAP7_75t_L g3048 ( 
.A(n_2949),
.B(n_2635),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_SL g3049 ( 
.A(n_2677),
.B(n_2460),
.Y(n_3049)
);

AOI22xp5_ASAP7_75t_L g3050 ( 
.A1(n_2926),
.A2(n_2556),
.B1(n_2643),
.B2(n_2658),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_L g3051 ( 
.A(n_2689),
.B(n_2586),
.Y(n_3051)
);

INVx2_ASAP7_75t_L g3052 ( 
.A(n_2733),
.Y(n_3052)
);

OR2x2_ASAP7_75t_L g3053 ( 
.A(n_2917),
.B(n_2576),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2686),
.Y(n_3054)
);

INVx2_ASAP7_75t_SL g3055 ( 
.A(n_2687),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2691),
.Y(n_3056)
);

NAND2xp5_ASAP7_75t_SL g3057 ( 
.A(n_2678),
.B(n_2460),
.Y(n_3057)
);

OAI22xp5_ASAP7_75t_L g3058 ( 
.A1(n_2845),
.A2(n_2628),
.B1(n_2595),
.B2(n_2618),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_SL g3059 ( 
.A(n_2678),
.B(n_2658),
.Y(n_3059)
);

AOI22xp33_ASAP7_75t_L g3060 ( 
.A1(n_2746),
.A2(n_2665),
.B1(n_2663),
.B2(n_2655),
.Y(n_3060)
);

NAND2xp5_ASAP7_75t_L g3061 ( 
.A(n_2689),
.B(n_2586),
.Y(n_3061)
);

INVx2_ASAP7_75t_SL g3062 ( 
.A(n_2753),
.Y(n_3062)
);

NOR2xp33_ASAP7_75t_L g3063 ( 
.A(n_2746),
.B(n_2636),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_L g3064 ( 
.A(n_2794),
.B(n_2586),
.Y(n_3064)
);

NAND2xp5_ASAP7_75t_L g3065 ( 
.A(n_2795),
.B(n_2586),
.Y(n_3065)
);

AND2x2_ASAP7_75t_L g3066 ( 
.A(n_2949),
.B(n_2660),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_L g3067 ( 
.A(n_2761),
.B(n_2619),
.Y(n_3067)
);

NOR2x1_ASAP7_75t_L g3068 ( 
.A(n_2843),
.B(n_2576),
.Y(n_3068)
);

O2A1O1Ixp5_ASAP7_75t_L g3069 ( 
.A1(n_2955),
.A2(n_2316),
.B(n_2352),
.C(n_2408),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2737),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2692),
.Y(n_3071)
);

NOR2xp33_ASAP7_75t_L g3072 ( 
.A(n_2667),
.B(n_2636),
.Y(n_3072)
);

NAND2xp33_ASAP7_75t_L g3073 ( 
.A(n_2953),
.B(n_2643),
.Y(n_3073)
);

INVx2_ASAP7_75t_L g3074 ( 
.A(n_2743),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_2695),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2696),
.Y(n_3076)
);

NOR2xp33_ASAP7_75t_L g3077 ( 
.A(n_2667),
.B(n_2636),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2890),
.Y(n_3078)
);

NAND2xp5_ASAP7_75t_L g3079 ( 
.A(n_2797),
.B(n_2802),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_SL g3080 ( 
.A(n_2678),
.B(n_2658),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2838),
.B(n_2660),
.Y(n_3081)
);

NOR2xp33_ASAP7_75t_L g3082 ( 
.A(n_2919),
.B(n_2556),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_SL g3083 ( 
.A(n_2682),
.B(n_2658),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_L g3084 ( 
.A(n_2807),
.B(n_2700),
.Y(n_3084)
);

INVx2_ASAP7_75t_L g3085 ( 
.A(n_2758),
.Y(n_3085)
);

INVx2_ASAP7_75t_SL g3086 ( 
.A(n_2884),
.Y(n_3086)
);

AND2x4_ASAP7_75t_L g3087 ( 
.A(n_2708),
.B(n_2575),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2891),
.Y(n_3088)
);

OAI22xp33_ASAP7_75t_L g3089 ( 
.A1(n_2845),
.A2(n_2658),
.B1(n_2666),
.B2(n_2519),
.Y(n_3089)
);

INVx8_ASAP7_75t_L g3090 ( 
.A(n_2815),
.Y(n_3090)
);

NOR2xp33_ASAP7_75t_L g3091 ( 
.A(n_2919),
.B(n_2416),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_L g3092 ( 
.A(n_2700),
.B(n_2554),
.Y(n_3092)
);

INVx8_ASAP7_75t_L g3093 ( 
.A(n_2815),
.Y(n_3093)
);

AOI22xp5_ASAP7_75t_L g3094 ( 
.A1(n_2926),
.A2(n_2643),
.B1(n_2640),
.B2(n_2649),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_L g3095 ( 
.A(n_2747),
.B(n_2626),
.Y(n_3095)
);

INVx2_ASAP7_75t_L g3096 ( 
.A(n_2765),
.Y(n_3096)
);

NOR2xp33_ASAP7_75t_SL g3097 ( 
.A(n_2953),
.B(n_2643),
.Y(n_3097)
);

AOI22xp5_ASAP7_75t_L g3098 ( 
.A1(n_2953),
.A2(n_2740),
.B1(n_2804),
.B2(n_2775),
.Y(n_3098)
);

NAND2xp5_ASAP7_75t_L g3099 ( 
.A(n_2747),
.B(n_2666),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_L g3100 ( 
.A(n_2937),
.B(n_2600),
.Y(n_3100)
);

NOR2x1p5_ASAP7_75t_L g3101 ( 
.A(n_2702),
.B(n_2664),
.Y(n_3101)
);

NAND2xp33_ASAP7_75t_L g3102 ( 
.A(n_2953),
.B(n_2595),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_2783),
.B(n_2593),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2898),
.Y(n_3104)
);

BUFx6f_ASAP7_75t_L g3105 ( 
.A(n_2716),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_2899),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_2905),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_L g3108 ( 
.A(n_2783),
.B(n_2593),
.Y(n_3108)
);

INVx5_ASAP7_75t_L g3109 ( 
.A(n_2863),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_L g3110 ( 
.A(n_2937),
.B(n_2596),
.Y(n_3110)
);

NOR2xp67_ASAP7_75t_L g3111 ( 
.A(n_2803),
.B(n_2343),
.Y(n_3111)
);

INVxp67_ASAP7_75t_L g3112 ( 
.A(n_2948),
.Y(n_3112)
);

INVx2_ASAP7_75t_L g3113 ( 
.A(n_2767),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_L g3114 ( 
.A(n_2722),
.B(n_2589),
.Y(n_3114)
);

AOI21xp5_ASAP7_75t_L g3115 ( 
.A1(n_2744),
.A2(n_2379),
.B(n_2359),
.Y(n_3115)
);

INVx2_ASAP7_75t_L g3116 ( 
.A(n_2772),
.Y(n_3116)
);

NOR2xp67_ASAP7_75t_L g3117 ( 
.A(n_2690),
.B(n_2343),
.Y(n_3117)
);

INVx2_ASAP7_75t_L g3118 ( 
.A(n_2776),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_L g3119 ( 
.A(n_2673),
.B(n_2598),
.Y(n_3119)
);

BUFx10_ASAP7_75t_L g3120 ( 
.A(n_2702),
.Y(n_3120)
);

OAI22xp33_ASAP7_75t_L g3121 ( 
.A1(n_2930),
.A2(n_2664),
.B1(n_2650),
.B2(n_2540),
.Y(n_3121)
);

NOR2xp33_ASAP7_75t_L g3122 ( 
.A(n_2722),
.B(n_2442),
.Y(n_3122)
);

INVx2_ASAP7_75t_SL g3123 ( 
.A(n_2739),
.Y(n_3123)
);

NOR2xp33_ASAP7_75t_L g3124 ( 
.A(n_2726),
.B(n_2716),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_L g3125 ( 
.A(n_2673),
.B(n_2598),
.Y(n_3125)
);

INVx2_ASAP7_75t_L g3126 ( 
.A(n_2790),
.Y(n_3126)
);

AOI22xp5_ASAP7_75t_L g3127 ( 
.A1(n_2953),
.A2(n_2318),
.B1(n_2517),
.B2(n_2509),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_L g3128 ( 
.A(n_2841),
.B(n_2616),
.Y(n_3128)
);

INVx1_ASAP7_75t_L g3129 ( 
.A(n_2906),
.Y(n_3129)
);

NOR2x1p5_ASAP7_75t_L g3130 ( 
.A(n_2751),
.B(n_2511),
.Y(n_3130)
);

INVx1_ASAP7_75t_L g3131 ( 
.A(n_2909),
.Y(n_3131)
);

NOR2xp33_ASAP7_75t_L g3132 ( 
.A(n_2726),
.B(n_2662),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_2918),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_2920),
.Y(n_3134)
);

NAND2xp5_ASAP7_75t_L g3135 ( 
.A(n_2841),
.B(n_2616),
.Y(n_3135)
);

INVx2_ASAP7_75t_L g3136 ( 
.A(n_2808),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2921),
.Y(n_3137)
);

OR2x2_ASAP7_75t_L g3138 ( 
.A(n_2956),
.B(n_2698),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_L g3139 ( 
.A(n_2723),
.B(n_2578),
.Y(n_3139)
);

INVx2_ASAP7_75t_L g3140 ( 
.A(n_2809),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_2927),
.Y(n_3141)
);

NAND2x1p5_ASAP7_75t_L g3142 ( 
.A(n_2869),
.B(n_2338),
.Y(n_3142)
);

AOI22xp33_ASAP7_75t_L g3143 ( 
.A1(n_2699),
.A2(n_2663),
.B1(n_2655),
.B2(n_2657),
.Y(n_3143)
);

NAND2xp5_ASAP7_75t_L g3144 ( 
.A(n_2938),
.B(n_2590),
.Y(n_3144)
);

BUFx6f_ASAP7_75t_L g3145 ( 
.A(n_2682),
.Y(n_3145)
);

NOR2xp33_ASAP7_75t_SL g3146 ( 
.A(n_2896),
.B(n_2511),
.Y(n_3146)
);

NAND2xp5_ASAP7_75t_L g3147 ( 
.A(n_2938),
.B(n_2584),
.Y(n_3147)
);

OR2x2_ASAP7_75t_L g3148 ( 
.A(n_2715),
.B(n_2657),
.Y(n_3148)
);

NOR2xp33_ASAP7_75t_L g3149 ( 
.A(n_2929),
.B(n_2325),
.Y(n_3149)
);

BUFx2_ASAP7_75t_L g3150 ( 
.A(n_2682),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_L g3151 ( 
.A(n_2818),
.B(n_2565),
.Y(n_3151)
);

NAND2xp5_ASAP7_75t_L g3152 ( 
.A(n_2819),
.B(n_2650),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_2731),
.Y(n_3153)
);

BUFx6f_ASAP7_75t_SL g3154 ( 
.A(n_2896),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_2732),
.Y(n_3155)
);

INVx2_ASAP7_75t_L g3156 ( 
.A(n_2817),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_L g3157 ( 
.A(n_2826),
.B(n_2641),
.Y(n_3157)
);

INVx2_ASAP7_75t_L g3158 ( 
.A(n_2827),
.Y(n_3158)
);

O2A1O1Ixp5_ASAP7_75t_L g3159 ( 
.A1(n_2955),
.A2(n_2450),
.B(n_2529),
.C(n_2531),
.Y(n_3159)
);

INVx2_ASAP7_75t_SL g3160 ( 
.A(n_2739),
.Y(n_3160)
);

INVx3_ASAP7_75t_L g3161 ( 
.A(n_2738),
.Y(n_3161)
);

INVx2_ASAP7_75t_SL g3162 ( 
.A(n_2739),
.Y(n_3162)
);

AOI22xp5_ASAP7_75t_L g3163 ( 
.A1(n_2740),
.A2(n_2319),
.B1(n_2602),
.B2(n_2488),
.Y(n_3163)
);

CKINVDCx5p33_ASAP7_75t_R g3164 ( 
.A(n_2751),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_SL g3165 ( 
.A(n_2697),
.B(n_2533),
.Y(n_3165)
);

INVxp33_ASAP7_75t_L g3166 ( 
.A(n_2745),
.Y(n_3166)
);

NAND2xp5_ASAP7_75t_L g3167 ( 
.A(n_2735),
.B(n_2579),
.Y(n_3167)
);

NOR2xp67_ASAP7_75t_L g3168 ( 
.A(n_2727),
.B(n_2338),
.Y(n_3168)
);

NOR2xp33_ASAP7_75t_L g3169 ( 
.A(n_2710),
.B(n_2637),
.Y(n_3169)
);

INVx3_ASAP7_75t_L g3170 ( 
.A(n_2738),
.Y(n_3170)
);

AND2x2_ASAP7_75t_L g3171 ( 
.A(n_2933),
.B(n_2913),
.Y(n_3171)
);

AOI22xp5_ASAP7_75t_L g3172 ( 
.A1(n_2740),
.A2(n_2319),
.B1(n_2602),
.B2(n_2488),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_L g3173 ( 
.A(n_2741),
.B(n_2602),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_SL g3174 ( 
.A(n_2697),
.B(n_2533),
.Y(n_3174)
);

INVx2_ASAP7_75t_L g3175 ( 
.A(n_2830),
.Y(n_3175)
);

NAND2xp5_ASAP7_75t_SL g3176 ( 
.A(n_2697),
.B(n_2533),
.Y(n_3176)
);

OR2x2_ASAP7_75t_L g3177 ( 
.A(n_2950),
.B(n_2654),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_L g3178 ( 
.A(n_2742),
.B(n_2602),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_2763),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_2769),
.Y(n_3180)
);

NAND2xp33_ASAP7_75t_L g3181 ( 
.A(n_2738),
.B(n_2618),
.Y(n_3181)
);

OR2x2_ASAP7_75t_L g3182 ( 
.A(n_2745),
.B(n_2654),
.Y(n_3182)
);

AOI22xp5_ASAP7_75t_L g3183 ( 
.A1(n_2804),
.A2(n_2319),
.B1(n_2602),
.B2(n_2488),
.Y(n_3183)
);

BUFx3_ASAP7_75t_L g3184 ( 
.A(n_3000),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_3141),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_L g3186 ( 
.A(n_2981),
.B(n_2934),
.Y(n_3186)
);

BUFx12f_ASAP7_75t_L g3187 ( 
.A(n_3164),
.Y(n_3187)
);

AOI22xp33_ASAP7_75t_L g3188 ( 
.A1(n_3098),
.A2(n_2410),
.B1(n_2924),
.B2(n_2942),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_SL g3189 ( 
.A(n_2967),
.B(n_2880),
.Y(n_3189)
);

AOI22xp33_ASAP7_75t_L g3190 ( 
.A1(n_3013),
.A2(n_2410),
.B1(n_2924),
.B2(n_2942),
.Y(n_3190)
);

OR2x2_ASAP7_75t_SL g3191 ( 
.A(n_3018),
.B(n_2745),
.Y(n_3191)
);

CKINVDCx5p33_ASAP7_75t_R g3192 ( 
.A(n_3120),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_2965),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_2976),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_2993),
.Y(n_3195)
);

NAND2xp5_ASAP7_75t_SL g3196 ( 
.A(n_2971),
.B(n_2883),
.Y(n_3196)
);

INVx1_ASAP7_75t_L g3197 ( 
.A(n_2998),
.Y(n_3197)
);

NAND2xp5_ASAP7_75t_L g3198 ( 
.A(n_2981),
.B(n_2984),
.Y(n_3198)
);

NAND2xp5_ASAP7_75t_L g3199 ( 
.A(n_2984),
.B(n_2941),
.Y(n_3199)
);

AND2x2_ASAP7_75t_SL g3200 ( 
.A(n_3097),
.B(n_2869),
.Y(n_3200)
);

OR2x2_ASAP7_75t_L g3201 ( 
.A(n_3001),
.B(n_2812),
.Y(n_3201)
);

BUFx5_ASAP7_75t_L g3202 ( 
.A(n_3008),
.Y(n_3202)
);

AND2x6_ASAP7_75t_L g3203 ( 
.A(n_3183),
.B(n_2708),
.Y(n_3203)
);

NOR2xp33_ASAP7_75t_L g3204 ( 
.A(n_2961),
.B(n_2784),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_3005),
.Y(n_3205)
);

NAND2xp5_ASAP7_75t_SL g3206 ( 
.A(n_2989),
.B(n_2759),
.Y(n_3206)
);

AND2x4_ASAP7_75t_L g3207 ( 
.A(n_3087),
.B(n_2868),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_3012),
.Y(n_3208)
);

BUFx3_ASAP7_75t_L g3209 ( 
.A(n_3086),
.Y(n_3209)
);

BUFx6f_ASAP7_75t_L g3210 ( 
.A(n_3019),
.Y(n_3210)
);

BUFx3_ASAP7_75t_L g3211 ( 
.A(n_3062),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_3016),
.Y(n_3212)
);

INVx5_ASAP7_75t_L g3213 ( 
.A(n_2980),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_3033),
.Y(n_3214)
);

BUFx3_ASAP7_75t_L g3215 ( 
.A(n_3120),
.Y(n_3215)
);

NOR2xp33_ASAP7_75t_L g3216 ( 
.A(n_2973),
.B(n_2784),
.Y(n_3216)
);

NAND2x1p5_ASAP7_75t_L g3217 ( 
.A(n_3109),
.B(n_2925),
.Y(n_3217)
);

AND3x2_ASAP7_75t_SL g3218 ( 
.A(n_3097),
.B(n_2543),
.C(n_2624),
.Y(n_3218)
);

BUFx4f_ASAP7_75t_L g3219 ( 
.A(n_3142),
.Y(n_3219)
);

INVx2_ASAP7_75t_SL g3220 ( 
.A(n_3044),
.Y(n_3220)
);

BUFx2_ASAP7_75t_L g3221 ( 
.A(n_3026),
.Y(n_3221)
);

INVx2_ASAP7_75t_L g3222 ( 
.A(n_2992),
.Y(n_3222)
);

INVx1_ASAP7_75t_L g3223 ( 
.A(n_3040),
.Y(n_3223)
);

INVx2_ASAP7_75t_L g3224 ( 
.A(n_3002),
.Y(n_3224)
);

AND2x6_ASAP7_75t_L g3225 ( 
.A(n_3163),
.B(n_2868),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_3054),
.Y(n_3226)
);

INVx2_ASAP7_75t_L g3227 ( 
.A(n_3010),
.Y(n_3227)
);

NAND2xp5_ASAP7_75t_L g3228 ( 
.A(n_3119),
.B(n_3125),
.Y(n_3228)
);

BUFx3_ASAP7_75t_L g3229 ( 
.A(n_3123),
.Y(n_3229)
);

INVx2_ASAP7_75t_SL g3230 ( 
.A(n_3160),
.Y(n_3230)
);

NOR2x1_ASAP7_75t_L g3231 ( 
.A(n_2997),
.B(n_2855),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_3056),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_3071),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_SL g3234 ( 
.A(n_2988),
.B(n_2759),
.Y(n_3234)
);

BUFx2_ASAP7_75t_L g3235 ( 
.A(n_3034),
.Y(n_3235)
);

CKINVDCx5p33_ASAP7_75t_R g3236 ( 
.A(n_3154),
.Y(n_3236)
);

INVx2_ASAP7_75t_SL g3237 ( 
.A(n_3162),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_3075),
.Y(n_3238)
);

BUFx6f_ASAP7_75t_L g3239 ( 
.A(n_3019),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_3076),
.Y(n_3240)
);

INVx2_ASAP7_75t_SL g3241 ( 
.A(n_2979),
.Y(n_3241)
);

INVxp67_ASAP7_75t_SL g3242 ( 
.A(n_3058),
.Y(n_3242)
);

AOI22xp33_ASAP7_75t_L g3243 ( 
.A1(n_2977),
.A2(n_2488),
.B1(n_2516),
.B2(n_2786),
.Y(n_3243)
);

INVxp67_ASAP7_75t_SL g3244 ( 
.A(n_3058),
.Y(n_3244)
);

INVxp67_ASAP7_75t_L g3245 ( 
.A(n_3082),
.Y(n_3245)
);

INVx1_ASAP7_75t_L g3246 ( 
.A(n_3078),
.Y(n_3246)
);

CKINVDCx5p33_ASAP7_75t_R g3247 ( 
.A(n_3154),
.Y(n_3247)
);

AOI22xp5_ASAP7_75t_SL g3248 ( 
.A1(n_3063),
.A2(n_2936),
.B1(n_2932),
.B2(n_2904),
.Y(n_3248)
);

BUFx3_ASAP7_75t_L g3249 ( 
.A(n_3004),
.Y(n_3249)
);

INVxp67_ASAP7_75t_L g3250 ( 
.A(n_3095),
.Y(n_3250)
);

AOI22xp33_ASAP7_75t_L g3251 ( 
.A1(n_2974),
.A2(n_2488),
.B1(n_2516),
.B2(n_2786),
.Y(n_3251)
);

BUFx3_ASAP7_75t_L g3252 ( 
.A(n_3042),
.Y(n_3252)
);

AOI22xp5_ASAP7_75t_L g3253 ( 
.A1(n_2983),
.A2(n_2991),
.B1(n_3027),
.B2(n_3022),
.Y(n_3253)
);

AO22x1_ASAP7_75t_L g3254 ( 
.A1(n_3149),
.A2(n_2910),
.B1(n_2933),
.B2(n_2897),
.Y(n_3254)
);

INVx3_ASAP7_75t_L g3255 ( 
.A(n_2980),
.Y(n_3255)
);

INVx2_ASAP7_75t_SL g3256 ( 
.A(n_3055),
.Y(n_3256)
);

AOI22xp33_ASAP7_75t_L g3257 ( 
.A1(n_2995),
.A2(n_2488),
.B1(n_2516),
.B2(n_2543),
.Y(n_3257)
);

INVxp67_ASAP7_75t_SL g3258 ( 
.A(n_3102),
.Y(n_3258)
);

CKINVDCx8_ASAP7_75t_R g3259 ( 
.A(n_3029),
.Y(n_3259)
);

INVx2_ASAP7_75t_L g3260 ( 
.A(n_3025),
.Y(n_3260)
);

INVx3_ASAP7_75t_L g3261 ( 
.A(n_2980),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_SL g3262 ( 
.A(n_2996),
.B(n_2925),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_L g3263 ( 
.A(n_3119),
.B(n_2829),
.Y(n_3263)
);

NAND2xp5_ASAP7_75t_L g3264 ( 
.A(n_3125),
.B(n_2832),
.Y(n_3264)
);

AND2x4_ASAP7_75t_L g3265 ( 
.A(n_3087),
.B(n_2868),
.Y(n_3265)
);

INVx2_ASAP7_75t_L g3266 ( 
.A(n_3045),
.Y(n_3266)
);

CKINVDCx6p67_ASAP7_75t_R g3267 ( 
.A(n_3109),
.Y(n_3267)
);

OAI22xp5_ASAP7_75t_L g3268 ( 
.A1(n_3172),
.A2(n_3094),
.B1(n_3050),
.B2(n_2985),
.Y(n_3268)
);

NAND2xp5_ASAP7_75t_L g3269 ( 
.A(n_3103),
.B(n_2836),
.Y(n_3269)
);

INVx3_ASAP7_75t_L g3270 ( 
.A(n_3090),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_3088),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_3104),
.Y(n_3272)
);

AO21x2_ASAP7_75t_L g3273 ( 
.A1(n_3089),
.A2(n_2429),
.B(n_2420),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_3106),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_3107),
.Y(n_3275)
);

INVx1_ASAP7_75t_SL g3276 ( 
.A(n_3150),
.Y(n_3276)
);

INVx1_ASAP7_75t_L g3277 ( 
.A(n_3129),
.Y(n_3277)
);

NOR2xp33_ASAP7_75t_L g3278 ( 
.A(n_3112),
.B(n_2897),
.Y(n_3278)
);

HB1xp67_ASAP7_75t_L g3279 ( 
.A(n_3173),
.Y(n_3279)
);

INVx2_ASAP7_75t_L g3280 ( 
.A(n_3052),
.Y(n_3280)
);

INVx2_ASAP7_75t_L g3281 ( 
.A(n_3070),
.Y(n_3281)
);

CKINVDCx5p33_ASAP7_75t_R g3282 ( 
.A(n_3047),
.Y(n_3282)
);

AOI22xp5_ASAP7_75t_L g3283 ( 
.A1(n_2994),
.A2(n_2932),
.B1(n_2755),
.B2(n_2940),
.Y(n_3283)
);

INVx2_ASAP7_75t_L g3284 ( 
.A(n_3074),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_3131),
.Y(n_3285)
);

AOI22xp5_ASAP7_75t_L g3286 ( 
.A1(n_3073),
.A2(n_2755),
.B1(n_2940),
.B2(n_2734),
.Y(n_3286)
);

NOR2xp33_ASAP7_75t_L g3287 ( 
.A(n_3006),
.B(n_2922),
.Y(n_3287)
);

BUFx2_ASAP7_75t_L g3288 ( 
.A(n_3145),
.Y(n_3288)
);

OR2x2_ASAP7_75t_L g3289 ( 
.A(n_3138),
.B(n_2840),
.Y(n_3289)
);

BUFx4f_ASAP7_75t_L g3290 ( 
.A(n_3142),
.Y(n_3290)
);

INVxp67_ASAP7_75t_L g3291 ( 
.A(n_3099),
.Y(n_3291)
);

INVx2_ASAP7_75t_L g3292 ( 
.A(n_3085),
.Y(n_3292)
);

INVx5_ASAP7_75t_L g3293 ( 
.A(n_3090),
.Y(n_3293)
);

OR2x6_ASAP7_75t_L g3294 ( 
.A(n_3090),
.B(n_2946),
.Y(n_3294)
);

OR2x2_ASAP7_75t_SL g3295 ( 
.A(n_2972),
.B(n_2564),
.Y(n_3295)
);

HB1xp67_ASAP7_75t_L g3296 ( 
.A(n_2960),
.Y(n_3296)
);

AND2x2_ASAP7_75t_L g3297 ( 
.A(n_3171),
.B(n_2858),
.Y(n_3297)
);

INVx5_ASAP7_75t_L g3298 ( 
.A(n_3093),
.Y(n_3298)
);

INVx1_ASAP7_75t_L g3299 ( 
.A(n_3133),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_L g3300 ( 
.A(n_3103),
.B(n_2846),
.Y(n_3300)
);

INVx4_ASAP7_75t_L g3301 ( 
.A(n_3093),
.Y(n_3301)
);

NAND2xp5_ASAP7_75t_L g3302 ( 
.A(n_3108),
.B(n_2852),
.Y(n_3302)
);

INVx1_ASAP7_75t_L g3303 ( 
.A(n_3134),
.Y(n_3303)
);

INVxp67_ASAP7_75t_L g3304 ( 
.A(n_3108),
.Y(n_3304)
);

BUFx2_ASAP7_75t_L g3305 ( 
.A(n_3145),
.Y(n_3305)
);

BUFx2_ASAP7_75t_L g3306 ( 
.A(n_3145),
.Y(n_3306)
);

AOI22xp33_ASAP7_75t_L g3307 ( 
.A1(n_3003),
.A2(n_2602),
.B1(n_2532),
.B2(n_2539),
.Y(n_3307)
);

AOI22x1_ASAP7_75t_L g3308 ( 
.A1(n_3115),
.A2(n_2811),
.B1(n_2892),
.B2(n_2835),
.Y(n_3308)
);

INVx2_ASAP7_75t_SL g3309 ( 
.A(n_3182),
.Y(n_3309)
);

INVx2_ASAP7_75t_SL g3310 ( 
.A(n_3101),
.Y(n_3310)
);

NOR2xp33_ASAP7_75t_L g3311 ( 
.A(n_3072),
.B(n_3077),
.Y(n_3311)
);

INVx1_ASAP7_75t_L g3312 ( 
.A(n_3137),
.Y(n_3312)
);

INVx3_ASAP7_75t_L g3313 ( 
.A(n_3093),
.Y(n_3313)
);

HB1xp67_ASAP7_75t_L g3314 ( 
.A(n_3173),
.Y(n_3314)
);

NOR2xp33_ASAP7_75t_L g3315 ( 
.A(n_3009),
.B(n_2922),
.Y(n_3315)
);

INVx4_ASAP7_75t_L g3316 ( 
.A(n_3109),
.Y(n_3316)
);

INVxp67_ASAP7_75t_L g3317 ( 
.A(n_3128),
.Y(n_3317)
);

AND2x4_ASAP7_75t_L g3318 ( 
.A(n_3008),
.B(n_2771),
.Y(n_3318)
);

BUFx6f_ASAP7_75t_L g3319 ( 
.A(n_2987),
.Y(n_3319)
);

AND2x4_ASAP7_75t_L g3320 ( 
.A(n_3130),
.B(n_2771),
.Y(n_3320)
);

NAND2xp5_ASAP7_75t_L g3321 ( 
.A(n_3128),
.B(n_2859),
.Y(n_3321)
);

AND2x4_ASAP7_75t_L g3322 ( 
.A(n_3015),
.B(n_2816),
.Y(n_3322)
);

NAND2x1p5_ASAP7_75t_L g3323 ( 
.A(n_3109),
.B(n_2963),
.Y(n_3323)
);

INVx2_ASAP7_75t_L g3324 ( 
.A(n_3096),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_3153),
.Y(n_3325)
);

INVx2_ASAP7_75t_L g3326 ( 
.A(n_3113),
.Y(n_3326)
);

AND2x4_ASAP7_75t_L g3327 ( 
.A(n_3015),
.B(n_2816),
.Y(n_3327)
);

INVx1_ASAP7_75t_L g3328 ( 
.A(n_3155),
.Y(n_3328)
);

AND2x4_ASAP7_75t_L g3329 ( 
.A(n_3015),
.B(n_2709),
.Y(n_3329)
);

O2A1O1Ixp5_ASAP7_75t_L g3330 ( 
.A1(n_2975),
.A2(n_2374),
.B(n_2422),
.C(n_2862),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_L g3331 ( 
.A(n_3135),
.B(n_2860),
.Y(n_3331)
);

INVx2_ASAP7_75t_L g3332 ( 
.A(n_3116),
.Y(n_3332)
);

INVx2_ASAP7_75t_L g3333 ( 
.A(n_3118),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3179),
.Y(n_3334)
);

INVx2_ASAP7_75t_L g3335 ( 
.A(n_2970),
.Y(n_3335)
);

BUFx6f_ASAP7_75t_L g3336 ( 
.A(n_2987),
.Y(n_3336)
);

INVx2_ASAP7_75t_SL g3337 ( 
.A(n_3177),
.Y(n_3337)
);

INVx1_ASAP7_75t_L g3338 ( 
.A(n_3180),
.Y(n_3338)
);

INVx1_ASAP7_75t_L g3339 ( 
.A(n_3084),
.Y(n_3339)
);

NAND2xp5_ASAP7_75t_L g3340 ( 
.A(n_3135),
.B(n_2872),
.Y(n_3340)
);

AND2x6_ASAP7_75t_L g3341 ( 
.A(n_2963),
.B(n_2764),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_3079),
.Y(n_3342)
);

BUFx3_ASAP7_75t_L g3343 ( 
.A(n_2987),
.Y(n_3343)
);

NAND2xp5_ASAP7_75t_L g3344 ( 
.A(n_3100),
.B(n_2877),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_3079),
.Y(n_3345)
);

BUFx6f_ASAP7_75t_L g3346 ( 
.A(n_3105),
.Y(n_3346)
);

INVx4_ASAP7_75t_L g3347 ( 
.A(n_3007),
.Y(n_3347)
);

INVx6_ASAP7_75t_L g3348 ( 
.A(n_3105),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_3110),
.B(n_2879),
.Y(n_3349)
);

NOR2x1p5_ASAP7_75t_L g3350 ( 
.A(n_3067),
.B(n_2711),
.Y(n_3350)
);

HB1xp67_ASAP7_75t_L g3351 ( 
.A(n_3092),
.Y(n_3351)
);

NAND2x1p5_ASAP7_75t_L g3352 ( 
.A(n_3041),
.B(n_2757),
.Y(n_3352)
);

INVxp67_ASAP7_75t_L g3353 ( 
.A(n_3091),
.Y(n_3353)
);

BUFx6f_ASAP7_75t_L g3354 ( 
.A(n_3105),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_SL g3355 ( 
.A(n_3039),
.B(n_2757),
.Y(n_3355)
);

HB1xp67_ASAP7_75t_L g3356 ( 
.A(n_3178),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_2990),
.Y(n_3357)
);

INVx5_ASAP7_75t_L g3358 ( 
.A(n_3041),
.Y(n_3358)
);

INVx2_ASAP7_75t_L g3359 ( 
.A(n_3126),
.Y(n_3359)
);

AND2x2_ASAP7_75t_L g3360 ( 
.A(n_3066),
.B(n_2858),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_L g3361 ( 
.A(n_2985),
.B(n_2881),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3136),
.Y(n_3362)
);

INVx1_ASAP7_75t_L g3363 ( 
.A(n_3140),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_L g3364 ( 
.A(n_3043),
.B(n_2885),
.Y(n_3364)
);

NAND2xp5_ASAP7_75t_SL g3365 ( 
.A(n_3030),
.B(n_2757),
.Y(n_3365)
);

AOI22xp5_ASAP7_75t_L g3366 ( 
.A1(n_3122),
.A2(n_3132),
.B1(n_3032),
.B2(n_3146),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_3156),
.Y(n_3367)
);

BUFx3_ASAP7_75t_L g3368 ( 
.A(n_3124),
.Y(n_3368)
);

BUFx3_ASAP7_75t_L g3369 ( 
.A(n_3161),
.Y(n_3369)
);

OAI21x1_ASAP7_75t_L g3370 ( 
.A1(n_3069),
.A2(n_2431),
.B(n_2429),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_L g3371 ( 
.A(n_3043),
.B(n_2887),
.Y(n_3371)
);

NOR2x1p5_ASAP7_75t_L g3372 ( 
.A(n_3014),
.B(n_2711),
.Y(n_3372)
);

OR2x2_ASAP7_75t_L g3373 ( 
.A(n_3053),
.B(n_2773),
.Y(n_3373)
);

INVx2_ASAP7_75t_L g3374 ( 
.A(n_3158),
.Y(n_3374)
);

BUFx3_ASAP7_75t_L g3375 ( 
.A(n_3161),
.Y(n_3375)
);

INVx3_ASAP7_75t_L g3376 ( 
.A(n_3007),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_3175),
.Y(n_3377)
);

BUFx12f_ASAP7_75t_L g3378 ( 
.A(n_3038),
.Y(n_3378)
);

INVx2_ASAP7_75t_SL g3379 ( 
.A(n_3170),
.Y(n_3379)
);

INVx2_ASAP7_75t_SL g3380 ( 
.A(n_3170),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_3021),
.Y(n_3381)
);

NAND2xp5_ASAP7_75t_L g3382 ( 
.A(n_3051),
.B(n_2774),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_L g3383 ( 
.A(n_3051),
.B(n_2777),
.Y(n_3383)
);

AOI22xp5_ASAP7_75t_L g3384 ( 
.A1(n_3146),
.A2(n_2755),
.B1(n_2734),
.B2(n_2863),
.Y(n_3384)
);

INVx2_ASAP7_75t_SL g3385 ( 
.A(n_3068),
.Y(n_3385)
);

HB1xp67_ASAP7_75t_L g3386 ( 
.A(n_3178),
.Y(n_3386)
);

AND2x2_ASAP7_75t_L g3387 ( 
.A(n_3048),
.B(n_3046),
.Y(n_3387)
);

INVx2_ASAP7_75t_L g3388 ( 
.A(n_3151),
.Y(n_3388)
);

CKINVDCx11_ASAP7_75t_R g3389 ( 
.A(n_3166),
.Y(n_3389)
);

INVx1_ASAP7_75t_L g3390 ( 
.A(n_3139),
.Y(n_3390)
);

AND3x2_ASAP7_75t_SL g3391 ( 
.A(n_2962),
.B(n_2936),
.C(n_2888),
.Y(n_3391)
);

CKINVDCx5p33_ASAP7_75t_R g3392 ( 
.A(n_3169),
.Y(n_3392)
);

NOR2xp67_ASAP7_75t_L g3393 ( 
.A(n_3111),
.B(n_2793),
.Y(n_3393)
);

INVx2_ASAP7_75t_L g3394 ( 
.A(n_3139),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_3167),
.Y(n_3395)
);

INVx3_ASAP7_75t_L g3396 ( 
.A(n_2982),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_L g3397 ( 
.A(n_3061),
.B(n_2849),
.Y(n_3397)
);

AOI21xp5_ASAP7_75t_L g3398 ( 
.A1(n_3258),
.A2(n_3181),
.B(n_2330),
.Y(n_3398)
);

NAND3xp33_ASAP7_75t_L g3399 ( 
.A(n_3190),
.B(n_3159),
.C(n_2537),
.Y(n_3399)
);

OA22x2_ASAP7_75t_L g3400 ( 
.A1(n_3253),
.A2(n_2999),
.B1(n_3127),
.B2(n_3036),
.Y(n_3400)
);

OAI22xp5_ASAP7_75t_L g3401 ( 
.A1(n_3188),
.A2(n_3061),
.B1(n_2966),
.B2(n_2964),
.Y(n_3401)
);

AOI21xp5_ASAP7_75t_L g3402 ( 
.A1(n_3258),
.A2(n_2330),
.B(n_2986),
.Y(n_3402)
);

O2A1O1Ixp33_ASAP7_75t_SL g3403 ( 
.A1(n_3234),
.A2(n_2912),
.B(n_3049),
.C(n_3035),
.Y(n_3403)
);

OAI21xp33_ASAP7_75t_L g3404 ( 
.A1(n_3242),
.A2(n_3244),
.B(n_3206),
.Y(n_3404)
);

BUFx6f_ASAP7_75t_L g3405 ( 
.A(n_3210),
.Y(n_3405)
);

INVx2_ASAP7_75t_L g3406 ( 
.A(n_3222),
.Y(n_3406)
);

AOI21xp5_ASAP7_75t_L g3407 ( 
.A1(n_3242),
.A2(n_2978),
.B(n_2969),
.Y(n_3407)
);

AOI21xp5_ASAP7_75t_L g3408 ( 
.A1(n_3244),
.A2(n_2978),
.B(n_2969),
.Y(n_3408)
);

OAI22xp5_ASAP7_75t_L g3409 ( 
.A1(n_3245),
.A2(n_2966),
.B1(n_2964),
.B2(n_3023),
.Y(n_3409)
);

AOI21xp5_ASAP7_75t_L g3410 ( 
.A1(n_3198),
.A2(n_2862),
.B(n_2359),
.Y(n_3410)
);

NAND2xp5_ASAP7_75t_L g3411 ( 
.A(n_3351),
.B(n_3167),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_3246),
.Y(n_3412)
);

AND2x2_ASAP7_75t_L g3413 ( 
.A(n_3387),
.B(n_3024),
.Y(n_3413)
);

NAND2x1p5_ASAP7_75t_L g3414 ( 
.A(n_3210),
.B(n_3239),
.Y(n_3414)
);

AOI21xp5_ASAP7_75t_L g3415 ( 
.A1(n_3198),
.A2(n_2814),
.B(n_2379),
.Y(n_3415)
);

NOR2xp33_ASAP7_75t_L g3416 ( 
.A(n_3282),
.B(n_2912),
.Y(n_3416)
);

AOI21x1_ASAP7_75t_L g3417 ( 
.A1(n_3189),
.A2(n_3080),
.B(n_3059),
.Y(n_3417)
);

BUFx6f_ASAP7_75t_L g3418 ( 
.A(n_3210),
.Y(n_3418)
);

BUFx6f_ASAP7_75t_L g3419 ( 
.A(n_3239),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_L g3420 ( 
.A(n_3250),
.B(n_3304),
.Y(n_3420)
);

CKINVDCx5p33_ASAP7_75t_R g3421 ( 
.A(n_3187),
.Y(n_3421)
);

BUFx6f_ASAP7_75t_L g3422 ( 
.A(n_3239),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_3271),
.Y(n_3423)
);

O2A1O1Ixp33_ASAP7_75t_L g3424 ( 
.A1(n_3196),
.A2(n_3121),
.B(n_3028),
.C(n_2523),
.Y(n_3424)
);

AOI22xp5_ASAP7_75t_L g3425 ( 
.A1(n_3251),
.A2(n_3114),
.B1(n_3031),
.B2(n_2661),
.Y(n_3425)
);

NAND2xp5_ASAP7_75t_L g3426 ( 
.A(n_3250),
.B(n_3020),
.Y(n_3426)
);

OAI21x1_ASAP7_75t_L g3427 ( 
.A1(n_3308),
.A2(n_2432),
.B(n_2431),
.Y(n_3427)
);

NAND2xp5_ASAP7_75t_L g3428 ( 
.A(n_3304),
.B(n_3017),
.Y(n_3428)
);

INVx3_ASAP7_75t_L g3429 ( 
.A(n_3316),
.Y(n_3429)
);

NAND2xp5_ASAP7_75t_L g3430 ( 
.A(n_3317),
.B(n_3081),
.Y(n_3430)
);

NAND2xp5_ASAP7_75t_L g3431 ( 
.A(n_3317),
.B(n_3147),
.Y(n_3431)
);

AOI21xp5_ASAP7_75t_L g3432 ( 
.A1(n_3200),
.A2(n_2814),
.B(n_3064),
.Y(n_3432)
);

INVx3_ASAP7_75t_L g3433 ( 
.A(n_3316),
.Y(n_3433)
);

BUFx2_ASAP7_75t_L g3434 ( 
.A(n_3249),
.Y(n_3434)
);

NAND2x1_ASAP7_75t_L g3435 ( 
.A(n_3396),
.B(n_3064),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_SL g3436 ( 
.A(n_3392),
.B(n_3144),
.Y(n_3436)
);

INVx1_ASAP7_75t_L g3437 ( 
.A(n_3272),
.Y(n_3437)
);

AOI21xp5_ASAP7_75t_L g3438 ( 
.A1(n_3384),
.A2(n_3065),
.B(n_3165),
.Y(n_3438)
);

AOI221xp5_ASAP7_75t_L g3439 ( 
.A1(n_3339),
.A2(n_2534),
.B1(n_3185),
.B2(n_3194),
.C(n_3193),
.Y(n_3439)
);

HB1xp67_ASAP7_75t_L g3440 ( 
.A(n_3245),
.Y(n_3440)
);

NAND2xp5_ASAP7_75t_L g3441 ( 
.A(n_3228),
.B(n_3037),
.Y(n_3441)
);

AOI21xp5_ASAP7_75t_L g3442 ( 
.A1(n_3273),
.A2(n_3065),
.B(n_3174),
.Y(n_3442)
);

AOI22xp33_ASAP7_75t_L g3443 ( 
.A1(n_3243),
.A2(n_2968),
.B1(n_3060),
.B2(n_3148),
.Y(n_3443)
);

OAI22xp5_ASAP7_75t_L g3444 ( 
.A1(n_3353),
.A2(n_2946),
.B1(n_2954),
.B2(n_2533),
.Y(n_3444)
);

NAND2xp5_ASAP7_75t_L g3445 ( 
.A(n_3228),
.B(n_3157),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_SL g3446 ( 
.A(n_3366),
.B(n_3168),
.Y(n_3446)
);

NAND2xp5_ASAP7_75t_SL g3447 ( 
.A(n_3231),
.B(n_2770),
.Y(n_3447)
);

NAND2xp5_ASAP7_75t_L g3448 ( 
.A(n_3353),
.B(n_2701),
.Y(n_3448)
);

AOI21xp5_ASAP7_75t_L g3449 ( 
.A1(n_3273),
.A2(n_3176),
.B(n_2854),
.Y(n_3449)
);

AOI21xp5_ASAP7_75t_L g3450 ( 
.A1(n_3330),
.A2(n_2854),
.B(n_2395),
.Y(n_3450)
);

A2O1A1Ixp33_ASAP7_75t_L g3451 ( 
.A1(n_3248),
.A2(n_2581),
.B(n_2552),
.C(n_2610),
.Y(n_3451)
);

AOI21xp5_ASAP7_75t_L g3452 ( 
.A1(n_3330),
.A2(n_2395),
.B(n_2394),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_L g3453 ( 
.A(n_3390),
.B(n_2707),
.Y(n_3453)
);

INVx2_ASAP7_75t_L g3454 ( 
.A(n_3224),
.Y(n_3454)
);

OAI21x1_ASAP7_75t_L g3455 ( 
.A1(n_3370),
.A2(n_2435),
.B(n_2432),
.Y(n_3455)
);

NAND2xp5_ASAP7_75t_L g3456 ( 
.A(n_3395),
.B(n_2714),
.Y(n_3456)
);

A2O1A1Ixp33_ASAP7_75t_SL g3457 ( 
.A1(n_3287),
.A2(n_2526),
.B(n_2538),
.C(n_2633),
.Y(n_3457)
);

BUFx6f_ASAP7_75t_L g3458 ( 
.A(n_3389),
.Y(n_3458)
);

NAND2xp5_ASAP7_75t_L g3459 ( 
.A(n_3201),
.B(n_2717),
.Y(n_3459)
);

NOR2xp33_ASAP7_75t_L g3460 ( 
.A(n_3216),
.B(n_2847),
.Y(n_3460)
);

AOI21xp5_ASAP7_75t_L g3461 ( 
.A1(n_3294),
.A2(n_2402),
.B(n_2394),
.Y(n_3461)
);

AOI21x1_ASAP7_75t_L g3462 ( 
.A1(n_3254),
.A2(n_3083),
.B(n_3152),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_SL g3463 ( 
.A(n_3311),
.B(n_3315),
.Y(n_3463)
);

OA22x2_ASAP7_75t_L g3464 ( 
.A1(n_3310),
.A2(n_3011),
.B1(n_2720),
.B2(n_2718),
.Y(n_3464)
);

NAND2xp5_ASAP7_75t_SL g3465 ( 
.A(n_3358),
.B(n_2770),
.Y(n_3465)
);

NAND2xp5_ASAP7_75t_SL g3466 ( 
.A(n_3358),
.B(n_2770),
.Y(n_3466)
);

O2A1O1Ixp33_ASAP7_75t_SL g3467 ( 
.A1(n_3204),
.A2(n_3057),
.B(n_2633),
.C(n_2538),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_SL g3468 ( 
.A(n_3358),
.B(n_2785),
.Y(n_3468)
);

O2A1O1Ixp5_ASAP7_75t_L g3469 ( 
.A1(n_3355),
.A2(n_2613),
.B(n_2526),
.C(n_2585),
.Y(n_3469)
);

NAND2x1p5_ASAP7_75t_L g3470 ( 
.A(n_3213),
.B(n_2785),
.Y(n_3470)
);

INVx2_ASAP7_75t_SL g3471 ( 
.A(n_3184),
.Y(n_3471)
);

NAND2xp5_ASAP7_75t_L g3472 ( 
.A(n_3291),
.B(n_2851),
.Y(n_3472)
);

NOR2xp33_ASAP7_75t_L g3473 ( 
.A(n_3278),
.B(n_3209),
.Y(n_3473)
);

AO32x1_ASAP7_75t_L g3474 ( 
.A1(n_3337),
.A2(n_2834),
.A3(n_2438),
.B1(n_2440),
.B2(n_2437),
.Y(n_3474)
);

OAI22xp5_ASAP7_75t_L g3475 ( 
.A1(n_3295),
.A2(n_2954),
.B1(n_2533),
.B2(n_2878),
.Y(n_3475)
);

INVx2_ASAP7_75t_L g3476 ( 
.A(n_3227),
.Y(n_3476)
);

OR2x6_ASAP7_75t_SL g3477 ( 
.A(n_3236),
.B(n_2903),
.Y(n_3477)
);

AOI21xp5_ASAP7_75t_L g3478 ( 
.A1(n_3294),
.A2(n_2402),
.B(n_2744),
.Y(n_3478)
);

AOI21xp5_ASAP7_75t_L g3479 ( 
.A1(n_3294),
.A2(n_2760),
.B(n_2750),
.Y(n_3479)
);

INVx2_ASAP7_75t_L g3480 ( 
.A(n_3260),
.Y(n_3480)
);

AOI21xp5_ASAP7_75t_L g3481 ( 
.A1(n_3358),
.A2(n_2760),
.B(n_2750),
.Y(n_3481)
);

OAI22xp5_ASAP7_75t_L g3482 ( 
.A1(n_3307),
.A2(n_2878),
.B1(n_2526),
.B2(n_2550),
.Y(n_3482)
);

AOI21x1_ASAP7_75t_L g3483 ( 
.A1(n_3365),
.A2(n_2908),
.B(n_2903),
.Y(n_3483)
);

A2O1A1Ixp33_ASAP7_75t_L g3484 ( 
.A1(n_3248),
.A2(n_2621),
.B(n_2622),
.C(n_3117),
.Y(n_3484)
);

OAI22xp5_ASAP7_75t_L g3485 ( 
.A1(n_3259),
.A2(n_2544),
.B1(n_2549),
.B2(n_2820),
.Y(n_3485)
);

NAND2xp5_ASAP7_75t_L g3486 ( 
.A(n_3291),
.B(n_2853),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_L g3487 ( 
.A(n_3394),
.B(n_2865),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_3274),
.Y(n_3488)
);

INVx2_ASAP7_75t_L g3489 ( 
.A(n_3266),
.Y(n_3489)
);

INVx2_ASAP7_75t_L g3490 ( 
.A(n_3280),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_L g3491 ( 
.A(n_3342),
.B(n_2873),
.Y(n_3491)
);

OAI22xp5_ASAP7_75t_SL g3492 ( 
.A1(n_3378),
.A2(n_3143),
.B1(n_2426),
.B2(n_2710),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_SL g3493 ( 
.A(n_3329),
.B(n_2785),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_3275),
.Y(n_3494)
);

INVx2_ASAP7_75t_L g3495 ( 
.A(n_3281),
.Y(n_3495)
);

BUFx3_ASAP7_75t_L g3496 ( 
.A(n_3211),
.Y(n_3496)
);

INVx1_ASAP7_75t_SL g3497 ( 
.A(n_3368),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_L g3498 ( 
.A(n_3345),
.B(n_2875),
.Y(n_3498)
);

BUFx3_ASAP7_75t_L g3499 ( 
.A(n_3215),
.Y(n_3499)
);

INVx4_ASAP7_75t_L g3500 ( 
.A(n_3347),
.Y(n_3500)
);

NOR2xp33_ASAP7_75t_L g3501 ( 
.A(n_3252),
.B(n_225),
.Y(n_3501)
);

AOI21xp5_ASAP7_75t_L g3502 ( 
.A1(n_3382),
.A2(n_2798),
.B(n_2437),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_SL g3503 ( 
.A(n_3329),
.B(n_2823),
.Y(n_3503)
);

CKINVDCx20_ASAP7_75t_R g3504 ( 
.A(n_3247),
.Y(n_3504)
);

AND2x4_ASAP7_75t_L g3505 ( 
.A(n_3322),
.B(n_2928),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_L g3506 ( 
.A(n_3296),
.B(n_2882),
.Y(n_3506)
);

NOR2xp33_ASAP7_75t_L g3507 ( 
.A(n_3221),
.B(n_226),
.Y(n_3507)
);

AOI22xp5_ASAP7_75t_L g3508 ( 
.A1(n_3268),
.A2(n_2755),
.B1(n_2863),
.B2(n_2319),
.Y(n_3508)
);

OAI22xp5_ASAP7_75t_L g3509 ( 
.A1(n_3257),
.A2(n_3350),
.B1(n_3235),
.B2(n_3283),
.Y(n_3509)
);

AOI22xp5_ASAP7_75t_L g3510 ( 
.A1(n_3268),
.A2(n_2755),
.B1(n_2863),
.B2(n_2319),
.Y(n_3510)
);

OAI22xp5_ASAP7_75t_L g3511 ( 
.A1(n_3286),
.A2(n_3372),
.B1(n_3290),
.B2(n_3219),
.Y(n_3511)
);

NAND2xp5_ASAP7_75t_L g3512 ( 
.A(n_3373),
.B(n_3388),
.Y(n_3512)
);

NOR2xp33_ASAP7_75t_L g3513 ( 
.A(n_3241),
.B(n_227),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_3277),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_L g3515 ( 
.A(n_3220),
.B(n_2902),
.Y(n_3515)
);

AOI21xp5_ASAP7_75t_L g3516 ( 
.A1(n_3382),
.A2(n_2798),
.B(n_2438),
.Y(n_3516)
);

AOI21xp5_ASAP7_75t_L g3517 ( 
.A1(n_3383),
.A2(n_2440),
.B(n_2435),
.Y(n_3517)
);

OA22x2_ASAP7_75t_L g3518 ( 
.A1(n_3262),
.A2(n_2630),
.B1(n_2623),
.B2(n_2822),
.Y(n_3518)
);

INVx2_ASAP7_75t_SL g3519 ( 
.A(n_3229),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_SL g3520 ( 
.A(n_3219),
.B(n_2823),
.Y(n_3520)
);

O2A1O1Ixp33_ASAP7_75t_L g3521 ( 
.A1(n_3256),
.A2(n_2505),
.B(n_2915),
.C(n_2894),
.Y(n_3521)
);

NOR2x1_ASAP7_75t_L g3522 ( 
.A(n_3369),
.B(n_2908),
.Y(n_3522)
);

INVx2_ASAP7_75t_L g3523 ( 
.A(n_3284),
.Y(n_3523)
);

NAND2xp5_ASAP7_75t_L g3524 ( 
.A(n_3381),
.B(n_2923),
.Y(n_3524)
);

AOI21xp5_ASAP7_75t_L g3525 ( 
.A1(n_3383),
.A2(n_2914),
.B(n_2834),
.Y(n_3525)
);

AOI22xp33_ASAP7_75t_L g3526 ( 
.A1(n_3225),
.A2(n_2319),
.B1(n_2630),
.B2(n_2931),
.Y(n_3526)
);

OAI21x1_ASAP7_75t_L g3527 ( 
.A1(n_3323),
.A2(n_2370),
.B(n_2914),
.Y(n_3527)
);

AOI21xp5_ASAP7_75t_L g3528 ( 
.A1(n_3213),
.A2(n_2520),
.B(n_2813),
.Y(n_3528)
);

OAI22xp5_ASAP7_75t_L g3529 ( 
.A1(n_3290),
.A2(n_2621),
.B1(n_2622),
.B2(n_2835),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_SL g3530 ( 
.A(n_3376),
.B(n_2823),
.Y(n_3530)
);

AND2x2_ASAP7_75t_L g3531 ( 
.A(n_3297),
.B(n_2928),
.Y(n_3531)
);

NAND2xp5_ASAP7_75t_L g3532 ( 
.A(n_3276),
.B(n_2939),
.Y(n_3532)
);

NAND2xp5_ASAP7_75t_L g3533 ( 
.A(n_3276),
.B(n_2943),
.Y(n_3533)
);

O2A1O1Ixp33_ASAP7_75t_SL g3534 ( 
.A1(n_3376),
.A2(n_2894),
.B(n_2892),
.C(n_2705),
.Y(n_3534)
);

AOI21xp5_ASAP7_75t_L g3535 ( 
.A1(n_3213),
.A2(n_2824),
.B(n_2813),
.Y(n_3535)
);

CKINVDCx5p33_ASAP7_75t_R g3536 ( 
.A(n_3192),
.Y(n_3536)
);

AND2x2_ASAP7_75t_L g3537 ( 
.A(n_3360),
.B(n_2787),
.Y(n_3537)
);

BUFx4f_ASAP7_75t_L g3538 ( 
.A(n_3267),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_L g3539 ( 
.A(n_3186),
.B(n_2944),
.Y(n_3539)
);

OAI22xp5_ASAP7_75t_L g3540 ( 
.A1(n_3347),
.A2(n_2915),
.B1(n_2642),
.B2(n_2656),
.Y(n_3540)
);

AOI21xp5_ASAP7_75t_L g3541 ( 
.A1(n_3213),
.A2(n_2824),
.B(n_2656),
.Y(n_3541)
);

O2A1O1Ixp33_ASAP7_75t_L g3542 ( 
.A1(n_3195),
.A2(n_2821),
.B(n_2806),
.C(n_2461),
.Y(n_3542)
);

NOR2xp33_ASAP7_75t_L g3543 ( 
.A(n_3375),
.B(n_227),
.Y(n_3543)
);

AOI22x1_ASAP7_75t_L g3544 ( 
.A1(n_3396),
.A2(n_2679),
.B1(n_2705),
.B2(n_2893),
.Y(n_3544)
);

O2A1O1Ixp33_ASAP7_75t_SL g3545 ( 
.A1(n_3379),
.A2(n_2679),
.B(n_2480),
.C(n_2481),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_3285),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_SL g3547 ( 
.A(n_3319),
.B(n_2825),
.Y(n_3547)
);

BUFx6f_ASAP7_75t_L g3548 ( 
.A(n_3319),
.Y(n_3548)
);

INVx2_ASAP7_75t_L g3549 ( 
.A(n_3292),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3299),
.Y(n_3550)
);

OR2x2_ASAP7_75t_L g3551 ( 
.A(n_3289),
.B(n_2951),
.Y(n_3551)
);

O2A1O1Ixp33_ASAP7_75t_L g3552 ( 
.A1(n_3197),
.A2(n_2822),
.B(n_2828),
.C(n_2577),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_L g3553 ( 
.A(n_3186),
.B(n_2863),
.Y(n_3553)
);

O2A1O1Ixp33_ASAP7_75t_L g3554 ( 
.A1(n_3205),
.A2(n_2828),
.B(n_2889),
.C(n_2874),
.Y(n_3554)
);

INVx2_ASAP7_75t_L g3555 ( 
.A(n_3324),
.Y(n_3555)
);

NAND2xp5_ASAP7_75t_L g3556 ( 
.A(n_3199),
.B(n_2377),
.Y(n_3556)
);

OR2x6_ASAP7_75t_SL g3557 ( 
.A(n_3199),
.B(n_2623),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_L g3558 ( 
.A(n_3208),
.B(n_2377),
.Y(n_3558)
);

AND2x2_ASAP7_75t_L g3559 ( 
.A(n_3212),
.B(n_2907),
.Y(n_3559)
);

NOR2xp67_ASAP7_75t_L g3560 ( 
.A(n_3230),
.B(n_2825),
.Y(n_3560)
);

AOI22xp5_ASAP7_75t_L g3561 ( 
.A1(n_3203),
.A2(n_2470),
.B1(n_2472),
.B2(n_2462),
.Y(n_3561)
);

NOR2xp33_ASAP7_75t_L g3562 ( 
.A(n_3237),
.B(n_228),
.Y(n_3562)
);

BUFx6f_ASAP7_75t_L g3563 ( 
.A(n_3319),
.Y(n_3563)
);

INVx2_ASAP7_75t_L g3564 ( 
.A(n_3326),
.Y(n_3564)
);

INVx2_ASAP7_75t_SL g3565 ( 
.A(n_3348),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_SL g3566 ( 
.A(n_3336),
.B(n_2825),
.Y(n_3566)
);

AND2x2_ASAP7_75t_L g3567 ( 
.A(n_3214),
.B(n_2907),
.Y(n_3567)
);

CKINVDCx5p33_ASAP7_75t_R g3568 ( 
.A(n_3343),
.Y(n_3568)
);

AOI21xp5_ASAP7_75t_L g3569 ( 
.A1(n_3293),
.A2(n_2656),
.B(n_2642),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_L g3570 ( 
.A(n_3223),
.B(n_2377),
.Y(n_3570)
);

OAI321xp33_ASAP7_75t_L g3571 ( 
.A1(n_3397),
.A2(n_2693),
.A3(n_2642),
.B1(n_2656),
.B2(n_2959),
.C(n_2952),
.Y(n_3571)
);

CKINVDCx5p33_ASAP7_75t_R g3572 ( 
.A(n_3288),
.Y(n_3572)
);

NOR2xp33_ASAP7_75t_L g3573 ( 
.A(n_3320),
.B(n_228),
.Y(n_3573)
);

AND2x2_ASAP7_75t_L g3574 ( 
.A(n_3226),
.B(n_2907),
.Y(n_3574)
);

INVx3_ASAP7_75t_L g3575 ( 
.A(n_3336),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_L g3576 ( 
.A(n_3232),
.B(n_2377),
.Y(n_3576)
);

INVx5_ASAP7_75t_L g3577 ( 
.A(n_3203),
.Y(n_3577)
);

OAI22xp5_ASAP7_75t_L g3578 ( 
.A1(n_3320),
.A2(n_2642),
.B1(n_2656),
.B2(n_2396),
.Y(n_3578)
);

AOI21xp5_ASAP7_75t_L g3579 ( 
.A1(n_3293),
.A2(n_2604),
.B(n_2805),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_3233),
.B(n_2377),
.Y(n_3580)
);

NOR2xp33_ASAP7_75t_L g3581 ( 
.A(n_3348),
.B(n_229),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_L g3582 ( 
.A(n_3238),
.B(n_3240),
.Y(n_3582)
);

OR2x2_ASAP7_75t_L g3583 ( 
.A(n_3303),
.B(n_2693),
.Y(n_3583)
);

INVx4_ASAP7_75t_L g3584 ( 
.A(n_3336),
.Y(n_3584)
);

AOI21xp5_ASAP7_75t_L g3585 ( 
.A1(n_3293),
.A2(n_2604),
.B(n_2805),
.Y(n_3585)
);

INVx2_ASAP7_75t_L g3586 ( 
.A(n_3332),
.Y(n_3586)
);

CKINVDCx10_ASAP7_75t_R g3587 ( 
.A(n_3393),
.Y(n_3587)
);

AOI22xp5_ASAP7_75t_L g3588 ( 
.A1(n_3203),
.A2(n_2470),
.B1(n_2472),
.B2(n_2462),
.Y(n_3588)
);

NAND2xp5_ASAP7_75t_L g3589 ( 
.A(n_3312),
.B(n_2377),
.Y(n_3589)
);

AOI21xp5_ASAP7_75t_L g3590 ( 
.A1(n_3293),
.A2(n_2604),
.B(n_2895),
.Y(n_3590)
);

NAND2xp5_ASAP7_75t_L g3591 ( 
.A(n_3325),
.B(n_3328),
.Y(n_3591)
);

BUFx2_ASAP7_75t_L g3592 ( 
.A(n_3305),
.Y(n_3592)
);

AOI21xp5_ASAP7_75t_L g3593 ( 
.A1(n_3298),
.A2(n_3349),
.B(n_3344),
.Y(n_3593)
);

AO21x1_ASAP7_75t_L g3594 ( 
.A1(n_3269),
.A2(n_2889),
.B(n_2874),
.Y(n_3594)
);

NOR2xp33_ASAP7_75t_L g3595 ( 
.A(n_3380),
.B(n_3334),
.Y(n_3595)
);

INVxp67_ASAP7_75t_SL g3596 ( 
.A(n_3269),
.Y(n_3596)
);

OAI22xp5_ASAP7_75t_L g3597 ( 
.A1(n_3298),
.A2(n_2396),
.B1(n_2508),
.B2(n_2358),
.Y(n_3597)
);

AOI21x1_ASAP7_75t_L g3598 ( 
.A1(n_3306),
.A2(n_2370),
.B(n_2443),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_L g3599 ( 
.A(n_3338),
.B(n_2842),
.Y(n_3599)
);

NAND2xp5_ASAP7_75t_L g3600 ( 
.A(n_3300),
.B(n_2842),
.Y(n_3600)
);

NOR2xp33_ASAP7_75t_L g3601 ( 
.A(n_3346),
.B(n_229),
.Y(n_3601)
);

INVx2_ASAP7_75t_L g3602 ( 
.A(n_3333),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_L g3603 ( 
.A(n_3300),
.B(n_2842),
.Y(n_3603)
);

OAI22xp5_ASAP7_75t_L g3604 ( 
.A1(n_3298),
.A2(n_2396),
.B1(n_2508),
.B2(n_2358),
.Y(n_3604)
);

AOI22xp5_ASAP7_75t_L g3605 ( 
.A1(n_3203),
.A2(n_2470),
.B1(n_2472),
.B2(n_2462),
.Y(n_3605)
);

INVxp67_ASAP7_75t_SL g3606 ( 
.A(n_3302),
.Y(n_3606)
);

INVx4_ASAP7_75t_L g3607 ( 
.A(n_3346),
.Y(n_3607)
);

HB1xp67_ASAP7_75t_L g3608 ( 
.A(n_3279),
.Y(n_3608)
);

AOI22xp5_ASAP7_75t_L g3609 ( 
.A1(n_3322),
.A2(n_2470),
.B1(n_2472),
.B2(n_2462),
.Y(n_3609)
);

AOI22xp5_ASAP7_75t_L g3610 ( 
.A1(n_3327),
.A2(n_2470),
.B1(n_2472),
.B2(n_2462),
.Y(n_3610)
);

AND2x2_ASAP7_75t_L g3611 ( 
.A(n_3309),
.B(n_2886),
.Y(n_3611)
);

NOR2x1_ASAP7_75t_L g3612 ( 
.A(n_3255),
.B(n_2895),
.Y(n_3612)
);

OAI22xp5_ASAP7_75t_L g3613 ( 
.A1(n_3298),
.A2(n_2508),
.B1(n_2358),
.B2(n_2339),
.Y(n_3613)
);

AO21x1_ASAP7_75t_L g3614 ( 
.A1(n_3302),
.A2(n_2911),
.B(n_2585),
.Y(n_3614)
);

AOI22xp33_ASAP7_75t_L g3615 ( 
.A1(n_3225),
.A2(n_2447),
.B1(n_2585),
.B2(n_2945),
.Y(n_3615)
);

OAI22xp5_ASAP7_75t_L g3616 ( 
.A1(n_3255),
.A2(n_2339),
.B1(n_2447),
.B2(n_2911),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_3412),
.Y(n_3617)
);

AOI21xp5_ASAP7_75t_L g3618 ( 
.A1(n_3402),
.A2(n_3331),
.B(n_3321),
.Y(n_3618)
);

BUFx6f_ASAP7_75t_L g3619 ( 
.A(n_3538),
.Y(n_3619)
);

AND2x2_ASAP7_75t_L g3620 ( 
.A(n_3434),
.B(n_3279),
.Y(n_3620)
);

OAI21x1_ASAP7_75t_L g3621 ( 
.A1(n_3590),
.A2(n_3323),
.B(n_3217),
.Y(n_3621)
);

AOI21x1_ASAP7_75t_L g3622 ( 
.A1(n_3462),
.A2(n_3349),
.B(n_3344),
.Y(n_3622)
);

AND2x2_ASAP7_75t_L g3623 ( 
.A(n_3413),
.B(n_3314),
.Y(n_3623)
);

INVx1_ASAP7_75t_L g3624 ( 
.A(n_3423),
.Y(n_3624)
);

INVx2_ASAP7_75t_L g3625 ( 
.A(n_3406),
.Y(n_3625)
);

NOR2xp33_ASAP7_75t_SL g3626 ( 
.A(n_3497),
.B(n_3301),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_L g3627 ( 
.A(n_3440),
.B(n_3386),
.Y(n_3627)
);

OAI21x1_ASAP7_75t_L g3628 ( 
.A1(n_3579),
.A2(n_3217),
.B(n_3352),
.Y(n_3628)
);

INVx2_ASAP7_75t_SL g3629 ( 
.A(n_3496),
.Y(n_3629)
);

OR2x2_ASAP7_75t_L g3630 ( 
.A(n_3420),
.B(n_3314),
.Y(n_3630)
);

AOI21x1_ASAP7_75t_L g3631 ( 
.A1(n_3447),
.A2(n_3331),
.B(n_3321),
.Y(n_3631)
);

OAI21x1_ASAP7_75t_L g3632 ( 
.A1(n_3585),
.A2(n_3352),
.B(n_3340),
.Y(n_3632)
);

OAI21xp5_ASAP7_75t_L g3633 ( 
.A1(n_3399),
.A2(n_3340),
.B(n_3264),
.Y(n_3633)
);

NAND2xp5_ASAP7_75t_L g3634 ( 
.A(n_3411),
.B(n_3445),
.Y(n_3634)
);

INVx4_ASAP7_75t_L g3635 ( 
.A(n_3500),
.Y(n_3635)
);

OAI21x1_ASAP7_75t_SL g3636 ( 
.A1(n_3500),
.A2(n_3264),
.B(n_3263),
.Y(n_3636)
);

INVx4_ASAP7_75t_L g3637 ( 
.A(n_3538),
.Y(n_3637)
);

OAI21xp5_ASAP7_75t_L g3638 ( 
.A1(n_3399),
.A2(n_3263),
.B(n_3356),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3437),
.Y(n_3639)
);

OAI21x1_ASAP7_75t_L g3640 ( 
.A1(n_3398),
.A2(n_3397),
.B(n_3270),
.Y(n_3640)
);

AOI21xp5_ASAP7_75t_L g3641 ( 
.A1(n_3404),
.A2(n_3327),
.B(n_3356),
.Y(n_3641)
);

OAI21x1_ASAP7_75t_L g3642 ( 
.A1(n_3483),
.A2(n_3270),
.B(n_3261),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_3488),
.Y(n_3643)
);

AOI31xp67_ASAP7_75t_L g3644 ( 
.A1(n_3400),
.A2(n_3364),
.A3(n_3371),
.B(n_3361),
.Y(n_3644)
);

OAI21xp5_ASAP7_75t_L g3645 ( 
.A1(n_3404),
.A2(n_3451),
.B(n_3484),
.Y(n_3645)
);

AOI21x1_ASAP7_75t_L g3646 ( 
.A1(n_3446),
.A2(n_3385),
.B(n_3364),
.Y(n_3646)
);

AND2x4_ASAP7_75t_L g3647 ( 
.A(n_3577),
.B(n_3386),
.Y(n_3647)
);

AOI22xp33_ASAP7_75t_L g3648 ( 
.A1(n_3492),
.A2(n_3225),
.B1(n_3391),
.B2(n_3362),
.Y(n_3648)
);

NAND2x1p5_ASAP7_75t_L g3649 ( 
.A(n_3577),
.B(n_3301),
.Y(n_3649)
);

OAI22xp5_ASAP7_75t_L g3650 ( 
.A1(n_3508),
.A2(n_3261),
.B1(n_3313),
.B2(n_3191),
.Y(n_3650)
);

OAI21x1_ASAP7_75t_L g3651 ( 
.A1(n_3449),
.A2(n_3598),
.B(n_3450),
.Y(n_3651)
);

AND2x2_ASAP7_75t_L g3652 ( 
.A(n_3592),
.B(n_3346),
.Y(n_3652)
);

AOI22xp5_ASAP7_75t_L g3653 ( 
.A1(n_3509),
.A2(n_3225),
.B1(n_3341),
.B2(n_3265),
.Y(n_3653)
);

OAI21x1_ASAP7_75t_L g3654 ( 
.A1(n_3452),
.A2(n_3313),
.B(n_3361),
.Y(n_3654)
);

BUFx8_ASAP7_75t_L g3655 ( 
.A(n_3458),
.Y(n_3655)
);

NAND2xp5_ASAP7_75t_L g3656 ( 
.A(n_3441),
.B(n_3371),
.Y(n_3656)
);

AO31x2_ASAP7_75t_L g3657 ( 
.A1(n_3614),
.A2(n_3363),
.A3(n_3367),
.B(n_3357),
.Y(n_3657)
);

INVxp67_ASAP7_75t_L g3658 ( 
.A(n_3463),
.Y(n_3658)
);

INVx2_ASAP7_75t_L g3659 ( 
.A(n_3454),
.Y(n_3659)
);

INVx5_ASAP7_75t_L g3660 ( 
.A(n_3577),
.Y(n_3660)
);

A2O1A1Ixp33_ASAP7_75t_L g3661 ( 
.A1(n_3424),
.A2(n_3391),
.B(n_3265),
.C(n_3207),
.Y(n_3661)
);

INVx2_ASAP7_75t_L g3662 ( 
.A(n_3476),
.Y(n_3662)
);

AND2x2_ASAP7_75t_L g3663 ( 
.A(n_3572),
.B(n_3537),
.Y(n_3663)
);

NAND2xp5_ASAP7_75t_L g3664 ( 
.A(n_3430),
.B(n_3341),
.Y(n_3664)
);

AOI21xp5_ASAP7_75t_L g3665 ( 
.A1(n_3481),
.A2(n_2500),
.B(n_3207),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_L g3666 ( 
.A(n_3426),
.B(n_3341),
.Y(n_3666)
);

INVx1_ASAP7_75t_L g3667 ( 
.A(n_3494),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3608),
.B(n_3341),
.Y(n_3668)
);

INVx2_ASAP7_75t_L g3669 ( 
.A(n_3480),
.Y(n_3669)
);

AOI21x1_ASAP7_75t_L g3670 ( 
.A1(n_3417),
.A2(n_3377),
.B(n_3359),
.Y(n_3670)
);

AOI22xp5_ASAP7_75t_L g3671 ( 
.A1(n_3508),
.A2(n_2470),
.B1(n_2472),
.B2(n_2462),
.Y(n_3671)
);

AOI21xp5_ASAP7_75t_L g3672 ( 
.A1(n_3479),
.A2(n_2725),
.B(n_2724),
.Y(n_3672)
);

AO31x2_ASAP7_75t_L g3673 ( 
.A1(n_3594),
.A2(n_3335),
.A3(n_3374),
.B(n_3218),
.Y(n_3673)
);

NAND2xp5_ASAP7_75t_L g3674 ( 
.A(n_3431),
.B(n_3354),
.Y(n_3674)
);

OAI21xp5_ASAP7_75t_L g3675 ( 
.A1(n_3522),
.A2(n_2867),
.B(n_2864),
.Y(n_3675)
);

OAI21x1_ASAP7_75t_L g3676 ( 
.A1(n_3427),
.A2(n_2725),
.B(n_2724),
.Y(n_3676)
);

OAI21xp5_ASAP7_75t_L g3677 ( 
.A1(n_3475),
.A2(n_2867),
.B(n_2864),
.Y(n_3677)
);

AOI21xp5_ASAP7_75t_SL g3678 ( 
.A1(n_3511),
.A2(n_3354),
.B(n_3318),
.Y(n_3678)
);

AOI21xp5_ASAP7_75t_L g3679 ( 
.A1(n_3569),
.A2(n_3218),
.B(n_3354),
.Y(n_3679)
);

INVx3_ASAP7_75t_L g3680 ( 
.A(n_3548),
.Y(n_3680)
);

NAND2xp5_ASAP7_75t_L g3681 ( 
.A(n_3448),
.B(n_3202),
.Y(n_3681)
);

OAI21x1_ASAP7_75t_L g3682 ( 
.A1(n_3528),
.A2(n_2486),
.B(n_2443),
.Y(n_3682)
);

NAND2xp5_ASAP7_75t_L g3683 ( 
.A(n_3596),
.B(n_3202),
.Y(n_3683)
);

INVx1_ASAP7_75t_SL g3684 ( 
.A(n_3568),
.Y(n_3684)
);

AO22x2_ASAP7_75t_L g3685 ( 
.A1(n_3606),
.A2(n_2958),
.B1(n_2957),
.B2(n_3318),
.Y(n_3685)
);

AO31x2_ASAP7_75t_L g3686 ( 
.A1(n_3442),
.A2(n_3401),
.A3(n_3432),
.B(n_3444),
.Y(n_3686)
);

NAND2xp5_ASAP7_75t_L g3687 ( 
.A(n_3428),
.B(n_3202),
.Y(n_3687)
);

O2A1O1Ixp33_ASAP7_75t_SL g3688 ( 
.A1(n_3504),
.A2(n_231),
.B(n_232),
.C(n_230),
.Y(n_3688)
);

NAND2xp5_ASAP7_75t_SL g3689 ( 
.A(n_3593),
.B(n_3202),
.Y(n_3689)
);

OAI21xp5_ASAP7_75t_L g3690 ( 
.A1(n_3410),
.A2(n_2870),
.B(n_2592),
.Y(n_3690)
);

NOR2xp67_ASAP7_75t_L g3691 ( 
.A(n_3429),
.B(n_2886),
.Y(n_3691)
);

AOI21xp5_ASAP7_75t_L g3692 ( 
.A1(n_3534),
.A2(n_2916),
.B(n_2886),
.Y(n_3692)
);

HB1xp67_ASAP7_75t_L g3693 ( 
.A(n_3595),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3514),
.Y(n_3694)
);

AND2x2_ASAP7_75t_L g3695 ( 
.A(n_3519),
.B(n_3202),
.Y(n_3695)
);

INVx1_ASAP7_75t_L g3696 ( 
.A(n_3546),
.Y(n_3696)
);

OAI21xp5_ASAP7_75t_L g3697 ( 
.A1(n_3457),
.A2(n_2870),
.B(n_2592),
.Y(n_3697)
);

OAI21xp5_ASAP7_75t_L g3698 ( 
.A1(n_3467),
.A2(n_2856),
.B(n_2893),
.Y(n_3698)
);

AOI21xp5_ASAP7_75t_L g3699 ( 
.A1(n_3415),
.A2(n_2935),
.B(n_2916),
.Y(n_3699)
);

OAI21x1_ASAP7_75t_L g3700 ( 
.A1(n_3455),
.A2(n_2486),
.B(n_2901),
.Y(n_3700)
);

AO21x1_ASAP7_75t_L g3701 ( 
.A1(n_3436),
.A2(n_2756),
.B(n_2861),
.Y(n_3701)
);

OAI21x1_ASAP7_75t_L g3702 ( 
.A1(n_3527),
.A2(n_3541),
.B(n_3535),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_L g3703 ( 
.A(n_3506),
.B(n_80),
.Y(n_3703)
);

AND2x2_ASAP7_75t_L g3704 ( 
.A(n_3471),
.B(n_2916),
.Y(n_3704)
);

NOR2xp67_ASAP7_75t_L g3705 ( 
.A(n_3429),
.B(n_2935),
.Y(n_3705)
);

OR2x2_ASAP7_75t_L g3706 ( 
.A(n_3550),
.B(n_81),
.Y(n_3706)
);

OAI21x1_ASAP7_75t_L g3707 ( 
.A1(n_3612),
.A2(n_2486),
.B(n_2901),
.Y(n_3707)
);

AOI21xp5_ASAP7_75t_L g3708 ( 
.A1(n_3525),
.A2(n_2947),
.B(n_2935),
.Y(n_3708)
);

NAND3x1_ASAP7_75t_L g3709 ( 
.A(n_3473),
.B(n_81),
.C(n_82),
.Y(n_3709)
);

INVxp67_ASAP7_75t_SL g3710 ( 
.A(n_3553),
.Y(n_3710)
);

NAND3x1_ASAP7_75t_L g3711 ( 
.A(n_3507),
.B(n_3416),
.C(n_3501),
.Y(n_3711)
);

INVx1_ASAP7_75t_L g3712 ( 
.A(n_3582),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_L g3713 ( 
.A(n_3557),
.B(n_81),
.Y(n_3713)
);

INVx1_ASAP7_75t_L g3714 ( 
.A(n_3591),
.Y(n_3714)
);

AOI22xp5_ASAP7_75t_L g3715 ( 
.A1(n_3510),
.A2(n_2861),
.B1(n_2551),
.B2(n_2653),
.Y(n_3715)
);

OAI21x1_ASAP7_75t_L g3716 ( 
.A1(n_3478),
.A2(n_2831),
.B(n_2796),
.Y(n_3716)
);

INVx1_ASAP7_75t_SL g3717 ( 
.A(n_3499),
.Y(n_3717)
);

OAI21x1_ASAP7_75t_SL g3718 ( 
.A1(n_3542),
.A2(n_2483),
.B(n_2457),
.Y(n_3718)
);

INVx2_ASAP7_75t_SL g3719 ( 
.A(n_3458),
.Y(n_3719)
);

O2A1O1Ixp5_ASAP7_75t_L g3720 ( 
.A1(n_3601),
.A2(n_2856),
.B(n_2339),
.C(n_2483),
.Y(n_3720)
);

OAI21x1_ASAP7_75t_L g3721 ( 
.A1(n_3461),
.A2(n_3469),
.B(n_3521),
.Y(n_3721)
);

NAND2xp5_ASAP7_75t_L g3722 ( 
.A(n_3409),
.B(n_82),
.Y(n_3722)
);

AND2x2_ASAP7_75t_L g3723 ( 
.A(n_3477),
.B(n_2947),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_3600),
.Y(n_3724)
);

AOI21x1_ASAP7_75t_L g3725 ( 
.A1(n_3530),
.A2(n_2484),
.B(n_2466),
.Y(n_3725)
);

OAI22xp5_ASAP7_75t_L g3726 ( 
.A1(n_3510),
.A2(n_2831),
.B1(n_2833),
.B2(n_2796),
.Y(n_3726)
);

OAI21x1_ASAP7_75t_L g3727 ( 
.A1(n_3502),
.A2(n_2833),
.B(n_2441),
.Y(n_3727)
);

NAND2xp5_ASAP7_75t_SL g3728 ( 
.A(n_3548),
.B(n_2947),
.Y(n_3728)
);

NAND2xp5_ASAP7_75t_L g3729 ( 
.A(n_3512),
.B(n_83),
.Y(n_3729)
);

OAI21x1_ASAP7_75t_L g3730 ( 
.A1(n_3516),
.A2(n_2441),
.B(n_2433),
.Y(n_3730)
);

AOI21x1_ASAP7_75t_L g3731 ( 
.A1(n_3560),
.A2(n_2484),
.B(n_2466),
.Y(n_3731)
);

OAI21xp5_ASAP7_75t_L g3732 ( 
.A1(n_3485),
.A2(n_2570),
.B(n_2569),
.Y(n_3732)
);

AO21x1_ASAP7_75t_L g3733 ( 
.A1(n_3543),
.A2(n_2483),
.B(n_2457),
.Y(n_3733)
);

AND2x6_ASAP7_75t_L g3734 ( 
.A(n_3561),
.B(n_3588),
.Y(n_3734)
);

AOI21x1_ASAP7_75t_L g3735 ( 
.A1(n_3532),
.A2(n_2492),
.B(n_2485),
.Y(n_3735)
);

NOR2x1_ASAP7_75t_SL g3736 ( 
.A(n_3540),
.B(n_2495),
.Y(n_3736)
);

AO31x2_ASAP7_75t_L g3737 ( 
.A1(n_3482),
.A2(n_3517),
.A3(n_3438),
.B(n_3408),
.Y(n_3737)
);

O2A1O1Ixp5_ASAP7_75t_L g3738 ( 
.A1(n_3581),
.A2(n_2491),
.B(n_2457),
.C(n_2433),
.Y(n_3738)
);

NAND2xp5_ASAP7_75t_L g3739 ( 
.A(n_3439),
.B(n_83),
.Y(n_3739)
);

INVx4_ASAP7_75t_L g3740 ( 
.A(n_3548),
.Y(n_3740)
);

AOI21xp5_ASAP7_75t_L g3741 ( 
.A1(n_3561),
.A2(n_2390),
.B(n_2368),
.Y(n_3741)
);

INVx1_ASAP7_75t_SL g3742 ( 
.A(n_3460),
.Y(n_3742)
);

BUFx5_ASAP7_75t_L g3743 ( 
.A(n_3559),
.Y(n_3743)
);

AND2x2_ASAP7_75t_L g3744 ( 
.A(n_3567),
.B(n_83),
.Y(n_3744)
);

NAND3xp33_ASAP7_75t_L g3745 ( 
.A(n_3599),
.B(n_2496),
.C(n_2495),
.Y(n_3745)
);

OAI21x1_ASAP7_75t_L g3746 ( 
.A1(n_3544),
.A2(n_2441),
.B(n_2433),
.Y(n_3746)
);

INVx5_ASAP7_75t_L g3747 ( 
.A(n_3563),
.Y(n_3747)
);

NAND3xp33_ASAP7_75t_L g3748 ( 
.A(n_3552),
.B(n_2496),
.C(n_2495),
.Y(n_3748)
);

AOI21xp5_ASAP7_75t_L g3749 ( 
.A1(n_3588),
.A2(n_2390),
.B(n_2368),
.Y(n_3749)
);

OAI21x1_ASAP7_75t_L g3750 ( 
.A1(n_3518),
.A2(n_2458),
.B(n_2445),
.Y(n_3750)
);

NAND2xp5_ASAP7_75t_L g3751 ( 
.A(n_3459),
.B(n_84),
.Y(n_3751)
);

HB1xp67_ASAP7_75t_L g3752 ( 
.A(n_3574),
.Y(n_3752)
);

OAI21x1_ASAP7_75t_L g3753 ( 
.A1(n_3433),
.A2(n_2458),
.B(n_2445),
.Y(n_3753)
);

AOI21xp5_ASAP7_75t_L g3754 ( 
.A1(n_3605),
.A2(n_2390),
.B(n_2397),
.Y(n_3754)
);

BUFx6f_ASAP7_75t_L g3755 ( 
.A(n_3563),
.Y(n_3755)
);

NAND2xp5_ASAP7_75t_L g3756 ( 
.A(n_3603),
.B(n_84),
.Y(n_3756)
);

A2O1A1Ixp33_ASAP7_75t_L g3757 ( 
.A1(n_3605),
.A2(n_2445),
.B(n_2482),
.C(n_2458),
.Y(n_3757)
);

INVx2_ASAP7_75t_L g3758 ( 
.A(n_3489),
.Y(n_3758)
);

OAI21x1_ASAP7_75t_L g3759 ( 
.A1(n_3433),
.A2(n_3407),
.B(n_3435),
.Y(n_3759)
);

AOI21xp5_ASAP7_75t_L g3760 ( 
.A1(n_3545),
.A2(n_3403),
.B(n_3571),
.Y(n_3760)
);

NAND2xp5_ASAP7_75t_L g3761 ( 
.A(n_3533),
.B(n_84),
.Y(n_3761)
);

AO31x2_ASAP7_75t_L g3762 ( 
.A1(n_3490),
.A2(n_2491),
.A3(n_2492),
.B(n_2485),
.Y(n_3762)
);

INVx1_ASAP7_75t_SL g3763 ( 
.A(n_3587),
.Y(n_3763)
);

OAI21x1_ASAP7_75t_L g3764 ( 
.A1(n_3464),
.A2(n_2494),
.B(n_2482),
.Y(n_3764)
);

OAI21x1_ASAP7_75t_L g3765 ( 
.A1(n_3554),
.A2(n_2494),
.B(n_2482),
.Y(n_3765)
);

BUFx2_ASAP7_75t_L g3766 ( 
.A(n_3458),
.Y(n_3766)
);

NAND2xp5_ASAP7_75t_L g3767 ( 
.A(n_3551),
.B(n_85),
.Y(n_3767)
);

AO21x1_ASAP7_75t_L g3768 ( 
.A1(n_3562),
.A2(n_2491),
.B(n_85),
.Y(n_3768)
);

HB1xp67_ASAP7_75t_L g3769 ( 
.A(n_3583),
.Y(n_3769)
);

NAND2xp5_ASAP7_75t_L g3770 ( 
.A(n_3472),
.B(n_85),
.Y(n_3770)
);

AOI21x1_ASAP7_75t_L g3771 ( 
.A1(n_3547),
.A2(n_2503),
.B(n_2501),
.Y(n_3771)
);

OAI21x1_ASAP7_75t_L g3772 ( 
.A1(n_3578),
.A2(n_2507),
.B(n_2494),
.Y(n_3772)
);

NOR4xp25_ASAP7_75t_L g3773 ( 
.A(n_3513),
.B(n_88),
.C(n_86),
.D(n_87),
.Y(n_3773)
);

BUFx10_ASAP7_75t_L g3774 ( 
.A(n_3536),
.Y(n_3774)
);

AO31x2_ASAP7_75t_L g3775 ( 
.A1(n_3495),
.A2(n_2501),
.A3(n_2503),
.B(n_2647),
.Y(n_3775)
);

AO31x2_ASAP7_75t_L g3776 ( 
.A1(n_3523),
.A2(n_2647),
.A3(n_2653),
.B(n_2397),
.Y(n_3776)
);

AOI21x1_ASAP7_75t_SL g3777 ( 
.A1(n_3587),
.A2(n_87),
.B(n_89),
.Y(n_3777)
);

AO31x2_ASAP7_75t_L g3778 ( 
.A1(n_3549),
.A2(n_2582),
.A3(n_2587),
.B(n_2573),
.Y(n_3778)
);

OAI21xp5_ASAP7_75t_L g3779 ( 
.A1(n_3573),
.A2(n_2507),
.B(n_2558),
.Y(n_3779)
);

NAND2x1p5_ASAP7_75t_L g3780 ( 
.A(n_3405),
.B(n_2496),
.Y(n_3780)
);

NAND2xp5_ASAP7_75t_L g3781 ( 
.A(n_3486),
.B(n_87),
.Y(n_3781)
);

OAI21xp5_ASAP7_75t_L g3782 ( 
.A1(n_3529),
.A2(n_3425),
.B(n_3609),
.Y(n_3782)
);

AOI221x1_ASAP7_75t_L g3783 ( 
.A1(n_3515),
.A2(n_2495),
.B1(n_2496),
.B2(n_2559),
.C(n_2507),
.Y(n_3783)
);

INVx3_ASAP7_75t_L g3784 ( 
.A(n_3563),
.Y(n_3784)
);

AND2x2_ASAP7_75t_L g3785 ( 
.A(n_3531),
.B(n_89),
.Y(n_3785)
);

NAND2xp5_ASAP7_75t_L g3786 ( 
.A(n_3539),
.B(n_89),
.Y(n_3786)
);

OAI21xp5_ASAP7_75t_L g3787 ( 
.A1(n_3425),
.A2(n_2582),
.B(n_2573),
.Y(n_3787)
);

BUFx6f_ASAP7_75t_L g3788 ( 
.A(n_3405),
.Y(n_3788)
);

A2O1A1Ixp33_ASAP7_75t_L g3789 ( 
.A1(n_3609),
.A2(n_2496),
.B(n_2587),
.C(n_2848),
.Y(n_3789)
);

INVx2_ASAP7_75t_SL g3790 ( 
.A(n_3565),
.Y(n_3790)
);

OAI21x1_ASAP7_75t_L g3791 ( 
.A1(n_3465),
.A2(n_3468),
.B(n_3466),
.Y(n_3791)
);

NAND2xp5_ASAP7_75t_L g3792 ( 
.A(n_3556),
.B(n_90),
.Y(n_3792)
);

OAI21x1_ASAP7_75t_L g3793 ( 
.A1(n_3597),
.A2(n_2848),
.B(n_90),
.Y(n_3793)
);

AOI21xp5_ASAP7_75t_L g3794 ( 
.A1(n_3474),
.A2(n_91),
.B(n_92),
.Y(n_3794)
);

OAI21x1_ASAP7_75t_SL g3795 ( 
.A1(n_3558),
.A2(n_241),
.B(n_233),
.Y(n_3795)
);

AOI22xp5_ASAP7_75t_L g3796 ( 
.A1(n_3492),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_3796)
);

AOI21x1_ASAP7_75t_L g3797 ( 
.A1(n_3566),
.A2(n_91),
.B(n_92),
.Y(n_3797)
);

OAI21x1_ASAP7_75t_L g3798 ( 
.A1(n_3604),
.A2(n_93),
.B(n_94),
.Y(n_3798)
);

AOI31xp67_ASAP7_75t_L g3799 ( 
.A1(n_3493),
.A2(n_96),
.A3(n_93),
.B(n_95),
.Y(n_3799)
);

OAI21x1_ASAP7_75t_SL g3800 ( 
.A1(n_3570),
.A2(n_247),
.B(n_238),
.Y(n_3800)
);

INVx2_ASAP7_75t_L g3801 ( 
.A(n_3555),
.Y(n_3801)
);

OAI21x1_ASAP7_75t_L g3802 ( 
.A1(n_3613),
.A2(n_3470),
.B(n_3610),
.Y(n_3802)
);

OAI21x1_ASAP7_75t_SL g3803 ( 
.A1(n_3576),
.A2(n_247),
.B(n_238),
.Y(n_3803)
);

OAI21x1_ASAP7_75t_L g3804 ( 
.A1(n_3470),
.A2(n_95),
.B(n_96),
.Y(n_3804)
);

OAI21x1_ASAP7_75t_L g3805 ( 
.A1(n_3610),
.A2(n_3616),
.B(n_3526),
.Y(n_3805)
);

NAND2xp5_ASAP7_75t_L g3806 ( 
.A(n_3453),
.B(n_96),
.Y(n_3806)
);

OAI21xp5_ASAP7_75t_L g3807 ( 
.A1(n_3503),
.A2(n_97),
.B(n_98),
.Y(n_3807)
);

AOI21xp5_ASAP7_75t_L g3808 ( 
.A1(n_3474),
.A2(n_99),
.B(n_100),
.Y(n_3808)
);

INVx1_ASAP7_75t_L g3809 ( 
.A(n_3456),
.Y(n_3809)
);

AOI21x1_ASAP7_75t_SL g3810 ( 
.A1(n_3580),
.A2(n_99),
.B(n_100),
.Y(n_3810)
);

AND2x4_ASAP7_75t_L g3811 ( 
.A(n_3611),
.B(n_99),
.Y(n_3811)
);

AO31x2_ASAP7_75t_L g3812 ( 
.A1(n_3564),
.A2(n_3602),
.A3(n_3586),
.B(n_3491),
.Y(n_3812)
);

NAND2xp5_ASAP7_75t_SL g3813 ( 
.A(n_3584),
.B(n_230),
.Y(n_3813)
);

AO31x2_ASAP7_75t_L g3814 ( 
.A1(n_3498),
.A2(n_3589),
.A3(n_3524),
.B(n_3487),
.Y(n_3814)
);

AO31x2_ASAP7_75t_L g3815 ( 
.A1(n_3474),
.A2(n_102),
.A3(n_100),
.B(n_101),
.Y(n_3815)
);

AOI21xp5_ASAP7_75t_L g3816 ( 
.A1(n_3520),
.A2(n_101),
.B(n_102),
.Y(n_3816)
);

INVx1_ASAP7_75t_L g3817 ( 
.A(n_3575),
.Y(n_3817)
);

OAI21xp5_ASAP7_75t_L g3818 ( 
.A1(n_3414),
.A2(n_102),
.B(n_103),
.Y(n_3818)
);

OAI21xp33_ASAP7_75t_L g3819 ( 
.A1(n_3575),
.A2(n_103),
.B(n_104),
.Y(n_3819)
);

OAI21x1_ASAP7_75t_L g3820 ( 
.A1(n_3615),
.A2(n_103),
.B(n_104),
.Y(n_3820)
);

OAI21xp5_ASAP7_75t_L g3821 ( 
.A1(n_3607),
.A2(n_104),
.B(n_105),
.Y(n_3821)
);

AND2x4_ASAP7_75t_L g3822 ( 
.A(n_3584),
.B(n_105),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_3607),
.Y(n_3823)
);

OAI21x1_ASAP7_75t_L g3824 ( 
.A1(n_3443),
.A2(n_105),
.B(n_106),
.Y(n_3824)
);

AND2x2_ASAP7_75t_L g3825 ( 
.A(n_3505),
.B(n_106),
.Y(n_3825)
);

AOI21xp5_ASAP7_75t_L g3826 ( 
.A1(n_3505),
.A2(n_106),
.B(n_107),
.Y(n_3826)
);

BUFx2_ASAP7_75t_L g3827 ( 
.A(n_3405),
.Y(n_3827)
);

BUFx6f_ASAP7_75t_L g3828 ( 
.A(n_3418),
.Y(n_3828)
);

INVx3_ASAP7_75t_L g3829 ( 
.A(n_3418),
.Y(n_3829)
);

OAI21x1_ASAP7_75t_L g3830 ( 
.A1(n_3418),
.A2(n_107),
.B(n_108),
.Y(n_3830)
);

OAI21x1_ASAP7_75t_L g3831 ( 
.A1(n_3419),
.A2(n_107),
.B(n_108),
.Y(n_3831)
);

NOR2xp67_ASAP7_75t_L g3832 ( 
.A(n_3422),
.B(n_231),
.Y(n_3832)
);

INVx4_ASAP7_75t_L g3833 ( 
.A(n_3422),
.Y(n_3833)
);

INVx2_ASAP7_75t_SL g3834 ( 
.A(n_3419),
.Y(n_3834)
);

A2O1A1Ixp33_ASAP7_75t_L g3835 ( 
.A1(n_3419),
.A2(n_110),
.B(n_108),
.C(n_109),
.Y(n_3835)
);

NAND2xp5_ASAP7_75t_L g3836 ( 
.A(n_3422),
.B(n_111),
.Y(n_3836)
);

INVx2_ASAP7_75t_L g3837 ( 
.A(n_3421),
.Y(n_3837)
);

AO22x2_ASAP7_75t_L g3838 ( 
.A1(n_3596),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_3838)
);

INVx2_ASAP7_75t_L g3839 ( 
.A(n_3406),
.Y(n_3839)
);

OAI21x1_ASAP7_75t_L g3840 ( 
.A1(n_3590),
.A2(n_111),
.B(n_112),
.Y(n_3840)
);

O2A1O1Ixp5_ASAP7_75t_L g3841 ( 
.A1(n_3463),
.A2(n_115),
.B(n_113),
.C(n_114),
.Y(n_3841)
);

NAND2xp5_ASAP7_75t_L g3842 ( 
.A(n_3440),
.B(n_113),
.Y(n_3842)
);

NAND2xp5_ASAP7_75t_SL g3843 ( 
.A(n_3577),
.B(n_234),
.Y(n_3843)
);

NOR2xp33_ASAP7_75t_SL g3844 ( 
.A(n_3497),
.B(n_114),
.Y(n_3844)
);

NAND2xp5_ASAP7_75t_L g3845 ( 
.A(n_3440),
.B(n_114),
.Y(n_3845)
);

NAND2xp5_ASAP7_75t_L g3846 ( 
.A(n_3724),
.B(n_234),
.Y(n_3846)
);

CKINVDCx5p33_ASAP7_75t_R g3847 ( 
.A(n_3655),
.Y(n_3847)
);

OAI21x1_ASAP7_75t_SL g3848 ( 
.A1(n_3713),
.A2(n_115),
.B(n_116),
.Y(n_3848)
);

AOI21xp5_ASAP7_75t_L g3849 ( 
.A1(n_3645),
.A2(n_123),
.B(n_115),
.Y(n_3849)
);

OAI21xp5_ASAP7_75t_L g3850 ( 
.A1(n_3796),
.A2(n_116),
.B(n_117),
.Y(n_3850)
);

AND2x2_ASAP7_75t_L g3851 ( 
.A(n_3620),
.B(n_116),
.Y(n_3851)
);

OR2x6_ASAP7_75t_L g3852 ( 
.A(n_3678),
.B(n_117),
.Y(n_3852)
);

NAND3xp33_ASAP7_75t_L g3853 ( 
.A(n_3796),
.B(n_117),
.C(n_118),
.Y(n_3853)
);

NOR2xp67_ASAP7_75t_L g3854 ( 
.A(n_3658),
.B(n_118),
.Y(n_3854)
);

CKINVDCx11_ASAP7_75t_R g3855 ( 
.A(n_3774),
.Y(n_3855)
);

NAND2xp5_ASAP7_75t_L g3856 ( 
.A(n_3724),
.B(n_235),
.Y(n_3856)
);

INVxp67_ASAP7_75t_SL g3857 ( 
.A(n_3683),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_L g3858 ( 
.A(n_3627),
.B(n_235),
.Y(n_3858)
);

NOR2xp33_ASAP7_75t_L g3859 ( 
.A(n_3742),
.B(n_236),
.Y(n_3859)
);

NAND3xp33_ASAP7_75t_SL g3860 ( 
.A(n_3844),
.B(n_119),
.C(n_120),
.Y(n_3860)
);

NOR4xp25_ASAP7_75t_L g3861 ( 
.A(n_3711),
.B(n_122),
.C(n_119),
.D(n_121),
.Y(n_3861)
);

INVx1_ASAP7_75t_L g3862 ( 
.A(n_3617),
.Y(n_3862)
);

AOI21xp5_ASAP7_75t_L g3863 ( 
.A1(n_3760),
.A2(n_129),
.B(n_121),
.Y(n_3863)
);

AOI21xp5_ASAP7_75t_L g3864 ( 
.A1(n_3689),
.A2(n_129),
.B(n_121),
.Y(n_3864)
);

NAND2xp5_ASAP7_75t_L g3865 ( 
.A(n_3630),
.B(n_236),
.Y(n_3865)
);

NAND2xp5_ASAP7_75t_L g3866 ( 
.A(n_3623),
.B(n_237),
.Y(n_3866)
);

A2O1A1Ixp33_ASAP7_75t_L g3867 ( 
.A1(n_3739),
.A2(n_124),
.B(n_122),
.C(n_123),
.Y(n_3867)
);

AOI21xp5_ASAP7_75t_L g3868 ( 
.A1(n_3618),
.A2(n_132),
.B(n_124),
.Y(n_3868)
);

OR2x6_ASAP7_75t_L g3869 ( 
.A(n_3766),
.B(n_124),
.Y(n_3869)
);

AND2x4_ASAP7_75t_L g3870 ( 
.A(n_3710),
.B(n_125),
.Y(n_3870)
);

OAI22x1_ASAP7_75t_L g3871 ( 
.A1(n_3693),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.Y(n_3871)
);

BUFx3_ASAP7_75t_L g3872 ( 
.A(n_3655),
.Y(n_3872)
);

O2A1O1Ixp33_ASAP7_75t_SL g3873 ( 
.A1(n_3763),
.A2(n_128),
.B(n_126),
.C(n_127),
.Y(n_3873)
);

AOI21xp5_ASAP7_75t_L g3874 ( 
.A1(n_3782),
.A2(n_137),
.B(n_126),
.Y(n_3874)
);

NOR2xp67_ASAP7_75t_SL g3875 ( 
.A(n_3619),
.B(n_237),
.Y(n_3875)
);

AOI21xp5_ASAP7_75t_L g3876 ( 
.A1(n_3722),
.A2(n_138),
.B(n_129),
.Y(n_3876)
);

OAI21xp5_ASAP7_75t_L g3877 ( 
.A1(n_3709),
.A2(n_130),
.B(n_131),
.Y(n_3877)
);

OAI21xp5_ASAP7_75t_L g3878 ( 
.A1(n_3773),
.A2(n_130),
.B(n_131),
.Y(n_3878)
);

INVx2_ASAP7_75t_L g3879 ( 
.A(n_3812),
.Y(n_3879)
);

INVx2_ASAP7_75t_L g3880 ( 
.A(n_3812),
.Y(n_3880)
);

OR2x2_ASAP7_75t_L g3881 ( 
.A(n_3769),
.B(n_130),
.Y(n_3881)
);

INVx1_ASAP7_75t_L g3882 ( 
.A(n_3617),
.Y(n_3882)
);

AOI21xp5_ASAP7_75t_L g3883 ( 
.A1(n_3641),
.A2(n_141),
.B(n_131),
.Y(n_3883)
);

INVx2_ASAP7_75t_L g3884 ( 
.A(n_3812),
.Y(n_3884)
);

A2O1A1Ixp33_ASAP7_75t_L g3885 ( 
.A1(n_3819),
.A2(n_135),
.B(n_133),
.C(n_134),
.Y(n_3885)
);

AO31x2_ASAP7_75t_L g3886 ( 
.A1(n_3733),
.A2(n_137),
.A3(n_134),
.B(n_136),
.Y(n_3886)
);

CKINVDCx20_ASAP7_75t_R g3887 ( 
.A(n_3774),
.Y(n_3887)
);

BUFx2_ASAP7_75t_L g3888 ( 
.A(n_3652),
.Y(n_3888)
);

OAI22xp5_ASAP7_75t_L g3889 ( 
.A1(n_3648),
.A2(n_137),
.B1(n_134),
.B2(n_136),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3624),
.Y(n_3890)
);

CKINVDCx11_ASAP7_75t_R g3891 ( 
.A(n_3684),
.Y(n_3891)
);

INVx2_ASAP7_75t_L g3892 ( 
.A(n_3625),
.Y(n_3892)
);

OAI21x1_ASAP7_75t_L g3893 ( 
.A1(n_3622),
.A2(n_139),
.B(n_140),
.Y(n_3893)
);

AND2x2_ASAP7_75t_L g3894 ( 
.A(n_3752),
.B(n_139),
.Y(n_3894)
);

AND2x2_ASAP7_75t_L g3895 ( 
.A(n_3663),
.B(n_139),
.Y(n_3895)
);

OAI21xp5_ASAP7_75t_L g3896 ( 
.A1(n_3841),
.A2(n_140),
.B(n_141),
.Y(n_3896)
);

OAI21x1_ASAP7_75t_L g3897 ( 
.A1(n_3670),
.A2(n_140),
.B(n_141),
.Y(n_3897)
);

NAND2xp5_ASAP7_75t_L g3898 ( 
.A(n_3634),
.B(n_3712),
.Y(n_3898)
);

OAI21x1_ASAP7_75t_L g3899 ( 
.A1(n_3651),
.A2(n_142),
.B(n_143),
.Y(n_3899)
);

CKINVDCx6p67_ASAP7_75t_R g3900 ( 
.A(n_3717),
.Y(n_3900)
);

INVxp67_ASAP7_75t_SL g3901 ( 
.A(n_3681),
.Y(n_3901)
);

AOI21xp5_ASAP7_75t_L g3902 ( 
.A1(n_3672),
.A2(n_150),
.B(n_142),
.Y(n_3902)
);

OAI21x1_ASAP7_75t_L g3903 ( 
.A1(n_3721),
.A2(n_142),
.B(n_143),
.Y(n_3903)
);

AOI21xp5_ASAP7_75t_L g3904 ( 
.A1(n_3741),
.A2(n_143),
.B(n_144),
.Y(n_3904)
);

NAND2x1p5_ASAP7_75t_L g3905 ( 
.A(n_3637),
.B(n_239),
.Y(n_3905)
);

AOI21xp5_ASAP7_75t_L g3906 ( 
.A1(n_3749),
.A2(n_144),
.B(n_145),
.Y(n_3906)
);

INVx1_ASAP7_75t_L g3907 ( 
.A(n_3624),
.Y(n_3907)
);

OAI21xp5_ASAP7_75t_L g3908 ( 
.A1(n_3794),
.A2(n_144),
.B(n_145),
.Y(n_3908)
);

AO21x2_ASAP7_75t_L g3909 ( 
.A1(n_3808),
.A2(n_145),
.B(n_146),
.Y(n_3909)
);

INVx2_ASAP7_75t_L g3910 ( 
.A(n_3659),
.Y(n_3910)
);

NAND2xp5_ASAP7_75t_L g3911 ( 
.A(n_3712),
.B(n_239),
.Y(n_3911)
);

AO31x2_ASAP7_75t_L g3912 ( 
.A1(n_3783),
.A2(n_148),
.A3(n_146),
.B(n_147),
.Y(n_3912)
);

BUFx2_ASAP7_75t_R g3913 ( 
.A(n_3674),
.Y(n_3913)
);

INVx2_ASAP7_75t_L g3914 ( 
.A(n_3662),
.Y(n_3914)
);

OAI21x1_ASAP7_75t_L g3915 ( 
.A1(n_3702),
.A2(n_146),
.B(n_147),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3639),
.Y(n_3916)
);

INVx3_ASAP7_75t_L g3917 ( 
.A(n_3635),
.Y(n_3917)
);

AND2x2_ASAP7_75t_L g3918 ( 
.A(n_3743),
.B(n_148),
.Y(n_3918)
);

INVx2_ASAP7_75t_L g3919 ( 
.A(n_3669),
.Y(n_3919)
);

INVx1_ASAP7_75t_L g3920 ( 
.A(n_3639),
.Y(n_3920)
);

OAI22x1_ASAP7_75t_L g3921 ( 
.A1(n_3811),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_3921)
);

OAI22xp33_ASAP7_75t_L g3922 ( 
.A1(n_3653),
.A2(n_151),
.B1(n_149),
.B2(n_150),
.Y(n_3922)
);

AO31x2_ASAP7_75t_L g3923 ( 
.A1(n_3736),
.A2(n_152),
.A3(n_149),
.B(n_151),
.Y(n_3923)
);

NAND2xp5_ASAP7_75t_L g3924 ( 
.A(n_3714),
.B(n_240),
.Y(n_3924)
);

INVx2_ASAP7_75t_L g3925 ( 
.A(n_3758),
.Y(n_3925)
);

OAI22x1_ASAP7_75t_L g3926 ( 
.A1(n_3811),
.A2(n_3714),
.B1(n_3719),
.B2(n_3822),
.Y(n_3926)
);

OA21x2_ASAP7_75t_L g3927 ( 
.A1(n_3759),
.A2(n_151),
.B(n_152),
.Y(n_3927)
);

AO21x2_ASAP7_75t_L g3928 ( 
.A1(n_3770),
.A2(n_152),
.B(n_153),
.Y(n_3928)
);

OAI21x1_ASAP7_75t_L g3929 ( 
.A1(n_3646),
.A2(n_153),
.B(n_154),
.Y(n_3929)
);

O2A1O1Ixp33_ASAP7_75t_L g3930 ( 
.A1(n_3688),
.A2(n_155),
.B(n_153),
.C(n_154),
.Y(n_3930)
);

AND2x4_ASAP7_75t_L g3931 ( 
.A(n_3647),
.B(n_155),
.Y(n_3931)
);

BUFx3_ASAP7_75t_L g3932 ( 
.A(n_3629),
.Y(n_3932)
);

O2A1O1Ixp33_ASAP7_75t_SL g3933 ( 
.A1(n_3813),
.A2(n_157),
.B(n_155),
.C(n_156),
.Y(n_3933)
);

A2O1A1Ixp33_ASAP7_75t_L g3934 ( 
.A1(n_3826),
.A2(n_158),
.B(n_156),
.C(n_157),
.Y(n_3934)
);

BUFx6f_ASAP7_75t_L g3935 ( 
.A(n_3619),
.Y(n_3935)
);

O2A1O1Ixp5_ASAP7_75t_L g3936 ( 
.A1(n_3768),
.A2(n_158),
.B(n_156),
.C(n_157),
.Y(n_3936)
);

AOI21xp5_ASAP7_75t_L g3937 ( 
.A1(n_3754),
.A2(n_158),
.B(n_159),
.Y(n_3937)
);

AOI21xp5_ASAP7_75t_L g3938 ( 
.A1(n_3708),
.A2(n_159),
.B(n_160),
.Y(n_3938)
);

INVx2_ASAP7_75t_L g3939 ( 
.A(n_3801),
.Y(n_3939)
);

INVx2_ASAP7_75t_L g3940 ( 
.A(n_3839),
.Y(n_3940)
);

A2O1A1Ixp33_ASAP7_75t_L g3941 ( 
.A1(n_3821),
.A2(n_161),
.B(n_159),
.C(n_160),
.Y(n_3941)
);

AOI21x1_ASAP7_75t_L g3942 ( 
.A1(n_3838),
.A2(n_160),
.B(n_161),
.Y(n_3942)
);

INVx3_ASAP7_75t_L g3943 ( 
.A(n_3635),
.Y(n_3943)
);

OAI21xp5_ASAP7_75t_L g3944 ( 
.A1(n_3835),
.A2(n_162),
.B(n_163),
.Y(n_3944)
);

BUFx10_ASAP7_75t_L g3945 ( 
.A(n_3619),
.Y(n_3945)
);

INVx2_ASAP7_75t_SL g3946 ( 
.A(n_3790),
.Y(n_3946)
);

A2O1A1Ixp33_ASAP7_75t_L g3947 ( 
.A1(n_3633),
.A2(n_3818),
.B(n_3832),
.C(n_3638),
.Y(n_3947)
);

A2O1A1Ixp33_ASAP7_75t_L g3948 ( 
.A1(n_3832),
.A2(n_165),
.B(n_163),
.C(n_164),
.Y(n_3948)
);

AOI21xp33_ASAP7_75t_L g3949 ( 
.A1(n_3838),
.A2(n_163),
.B(n_164),
.Y(n_3949)
);

INVx5_ASAP7_75t_L g3950 ( 
.A(n_3637),
.Y(n_3950)
);

NOR2xp33_ASAP7_75t_L g3951 ( 
.A(n_3837),
.B(n_242),
.Y(n_3951)
);

OR2x2_ASAP7_75t_L g3952 ( 
.A(n_3809),
.B(n_165),
.Y(n_3952)
);

O2A1O1Ixp33_ASAP7_75t_L g3953 ( 
.A1(n_3843),
.A2(n_168),
.B(n_166),
.C(n_167),
.Y(n_3953)
);

AND2x2_ASAP7_75t_L g3954 ( 
.A(n_3743),
.B(n_166),
.Y(n_3954)
);

INVx1_ASAP7_75t_L g3955 ( 
.A(n_3643),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_L g3956 ( 
.A(n_3656),
.B(n_242),
.Y(n_3956)
);

AO31x2_ASAP7_75t_L g3957 ( 
.A1(n_3679),
.A2(n_168),
.A3(n_166),
.B(n_167),
.Y(n_3957)
);

NAND2xp5_ASAP7_75t_L g3958 ( 
.A(n_3809),
.B(n_243),
.Y(n_3958)
);

INVx2_ASAP7_75t_L g3959 ( 
.A(n_3643),
.Y(n_3959)
);

AOI22xp5_ASAP7_75t_L g3960 ( 
.A1(n_3734),
.A2(n_169),
.B1(n_167),
.B2(n_168),
.Y(n_3960)
);

AOI21xp5_ASAP7_75t_L g3961 ( 
.A1(n_3665),
.A2(n_169),
.B(n_170),
.Y(n_3961)
);

OAI21x1_ASAP7_75t_L g3962 ( 
.A1(n_3654),
.A2(n_169),
.B(n_170),
.Y(n_3962)
);

INVx1_ASAP7_75t_SL g3963 ( 
.A(n_3695),
.Y(n_3963)
);

INVx1_ASAP7_75t_L g3964 ( 
.A(n_3667),
.Y(n_3964)
);

AOI21xp5_ASAP7_75t_L g3965 ( 
.A1(n_3692),
.A2(n_3699),
.B(n_3748),
.Y(n_3965)
);

AOI21xp5_ASAP7_75t_L g3966 ( 
.A1(n_3720),
.A2(n_170),
.B(n_171),
.Y(n_3966)
);

INVx2_ASAP7_75t_SL g3967 ( 
.A(n_3755),
.Y(n_3967)
);

A2O1A1Ixp33_ASAP7_75t_L g3968 ( 
.A1(n_3661),
.A2(n_173),
.B(n_171),
.C(n_172),
.Y(n_3968)
);

AOI21xp5_ASAP7_75t_L g3969 ( 
.A1(n_3690),
.A2(n_171),
.B(n_172),
.Y(n_3969)
);

OAI22xp5_ASAP7_75t_L g3970 ( 
.A1(n_3671),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_3970)
);

INVx1_ASAP7_75t_L g3971 ( 
.A(n_3667),
.Y(n_3971)
);

NAND2x1p5_ASAP7_75t_L g3972 ( 
.A(n_3747),
.B(n_243),
.Y(n_3972)
);

AND3x4_ASAP7_75t_L g3973 ( 
.A(n_3822),
.B(n_173),
.C(n_175),
.Y(n_3973)
);

AND2x6_ASAP7_75t_L g3974 ( 
.A(n_3647),
.B(n_244),
.Y(n_3974)
);

AO21x1_ASAP7_75t_L g3975 ( 
.A1(n_3842),
.A2(n_176),
.B(n_177),
.Y(n_3975)
);

BUFx6f_ASAP7_75t_L g3976 ( 
.A(n_3788),
.Y(n_3976)
);

INVx1_ASAP7_75t_L g3977 ( 
.A(n_3694),
.Y(n_3977)
);

INVx2_ASAP7_75t_L g3978 ( 
.A(n_3694),
.Y(n_3978)
);

AO21x2_ASAP7_75t_L g3979 ( 
.A1(n_3781),
.A2(n_176),
.B(n_177),
.Y(n_3979)
);

OAI22xp5_ASAP7_75t_L g3980 ( 
.A1(n_3671),
.A2(n_178),
.B1(n_176),
.B2(n_177),
.Y(n_3980)
);

INVx1_ASAP7_75t_SL g3981 ( 
.A(n_3827),
.Y(n_3981)
);

AND2x4_ASAP7_75t_L g3982 ( 
.A(n_3668),
.B(n_178),
.Y(n_3982)
);

INVx1_ASAP7_75t_L g3983 ( 
.A(n_3696),
.Y(n_3983)
);

AND2x2_ASAP7_75t_L g3984 ( 
.A(n_3743),
.B(n_178),
.Y(n_3984)
);

BUFx6f_ASAP7_75t_L g3985 ( 
.A(n_3788),
.Y(n_3985)
);

OAI21x1_ASAP7_75t_L g3986 ( 
.A1(n_3628),
.A2(n_179),
.B(n_180),
.Y(n_3986)
);

AOI22xp5_ASAP7_75t_L g3987 ( 
.A1(n_3734),
.A2(n_182),
.B1(n_180),
.B2(n_181),
.Y(n_3987)
);

O2A1O1Ixp33_ASAP7_75t_SL g3988 ( 
.A1(n_3845),
.A2(n_182),
.B(n_180),
.C(n_181),
.Y(n_3988)
);

A2O1A1Ixp33_ASAP7_75t_L g3989 ( 
.A1(n_3807),
.A2(n_183),
.B(n_181),
.C(n_182),
.Y(n_3989)
);

NAND2xp5_ASAP7_75t_L g3990 ( 
.A(n_3687),
.B(n_244),
.Y(n_3990)
);

INVx1_ASAP7_75t_L g3991 ( 
.A(n_3696),
.Y(n_3991)
);

O2A1O1Ixp33_ASAP7_75t_SL g3992 ( 
.A1(n_3756),
.A2(n_185),
.B(n_183),
.C(n_184),
.Y(n_3992)
);

OAI21x1_ASAP7_75t_L g3993 ( 
.A1(n_3632),
.A2(n_184),
.B(n_185),
.Y(n_3993)
);

A2O1A1Ixp33_ASAP7_75t_L g3994 ( 
.A1(n_3816),
.A2(n_187),
.B(n_184),
.C(n_186),
.Y(n_3994)
);

INVx1_ASAP7_75t_L g3995 ( 
.A(n_3814),
.Y(n_3995)
);

A2O1A1Ixp33_ASAP7_75t_L g3996 ( 
.A1(n_3779),
.A2(n_189),
.B(n_186),
.C(n_188),
.Y(n_3996)
);

AOI21xp5_ASAP7_75t_L g3997 ( 
.A1(n_3738),
.A2(n_188),
.B(n_189),
.Y(n_3997)
);

OAI21x1_ASAP7_75t_SL g3998 ( 
.A1(n_3636),
.A2(n_188),
.B(n_189),
.Y(n_3998)
);

O2A1O1Ixp33_ASAP7_75t_SL g3999 ( 
.A1(n_3806),
.A2(n_193),
.B(n_191),
.C(n_192),
.Y(n_3999)
);

O2A1O1Ixp33_ASAP7_75t_SL g4000 ( 
.A1(n_3751),
.A2(n_3706),
.B(n_3767),
.C(n_3703),
.Y(n_4000)
);

AOI21xp5_ASAP7_75t_L g4001 ( 
.A1(n_3757),
.A2(n_191),
.B(n_193),
.Y(n_4001)
);

NOR2xp33_ASAP7_75t_L g4002 ( 
.A(n_3626),
.B(n_245),
.Y(n_4002)
);

AOI21xp5_ASAP7_75t_L g4003 ( 
.A1(n_3789),
.A2(n_193),
.B(n_194),
.Y(n_4003)
);

AOI21xp5_ASAP7_75t_L g4004 ( 
.A1(n_3698),
.A2(n_194),
.B(n_195),
.Y(n_4004)
);

AND2x4_ASAP7_75t_L g4005 ( 
.A(n_3817),
.B(n_3723),
.Y(n_4005)
);

AOI21xp5_ASAP7_75t_L g4006 ( 
.A1(n_3697),
.A2(n_195),
.B(n_196),
.Y(n_4006)
);

OAI21xp5_ASAP7_75t_L g4007 ( 
.A1(n_3644),
.A2(n_195),
.B(n_196),
.Y(n_4007)
);

INVx1_ASAP7_75t_L g4008 ( 
.A(n_3631),
.Y(n_4008)
);

OR2x2_ASAP7_75t_L g4009 ( 
.A(n_3666),
.B(n_197),
.Y(n_4009)
);

NAND2xp33_ASAP7_75t_SL g4010 ( 
.A(n_3740),
.B(n_198),
.Y(n_4010)
);

OAI21xp5_ASAP7_75t_L g4011 ( 
.A1(n_3840),
.A2(n_199),
.B(n_200),
.Y(n_4011)
);

INVx1_ASAP7_75t_L g4012 ( 
.A(n_3814),
.Y(n_4012)
);

AOI21xp5_ASAP7_75t_L g4013 ( 
.A1(n_3726),
.A2(n_199),
.B(n_200),
.Y(n_4013)
);

OAI21x1_ASAP7_75t_L g4014 ( 
.A1(n_3642),
.A2(n_199),
.B(n_200),
.Y(n_4014)
);

OAI21x1_ASAP7_75t_L g4015 ( 
.A1(n_3640),
.A2(n_3621),
.B(n_3735),
.Y(n_4015)
);

OR2x2_ASAP7_75t_L g4016 ( 
.A(n_3664),
.B(n_201),
.Y(n_4016)
);

OAI21x1_ASAP7_75t_L g4017 ( 
.A1(n_3802),
.A2(n_201),
.B(n_202),
.Y(n_4017)
);

O2A1O1Ixp33_ASAP7_75t_L g4018 ( 
.A1(n_3761),
.A2(n_3786),
.B(n_3729),
.C(n_3795),
.Y(n_4018)
);

OAI22x1_ASAP7_75t_L g4019 ( 
.A1(n_3660),
.A2(n_203),
.B1(n_201),
.B2(n_202),
.Y(n_4019)
);

O2A1O1Ixp33_ASAP7_75t_SL g4020 ( 
.A1(n_3836),
.A2(n_204),
.B(n_202),
.C(n_203),
.Y(n_4020)
);

NAND2xp5_ASAP7_75t_L g4021 ( 
.A(n_3814),
.B(n_3743),
.Y(n_4021)
);

O2A1O1Ixp33_ASAP7_75t_L g4022 ( 
.A1(n_3800),
.A2(n_205),
.B(n_203),
.C(n_204),
.Y(n_4022)
);

AOI22xp5_ASAP7_75t_L g4023 ( 
.A1(n_3734),
.A2(n_206),
.B1(n_204),
.B2(n_205),
.Y(n_4023)
);

NAND2x1p5_ASAP7_75t_L g4024 ( 
.A(n_3747),
.B(n_245),
.Y(n_4024)
);

CKINVDCx5p33_ASAP7_75t_R g4025 ( 
.A(n_3755),
.Y(n_4025)
);

INVx2_ASAP7_75t_SL g4026 ( 
.A(n_3755),
.Y(n_4026)
);

AND2x2_ASAP7_75t_L g4027 ( 
.A(n_3743),
.B(n_205),
.Y(n_4027)
);

INVx2_ASAP7_75t_L g4028 ( 
.A(n_3959),
.Y(n_4028)
);

AOI22xp33_ASAP7_75t_L g4029 ( 
.A1(n_3853),
.A2(n_3734),
.B1(n_3824),
.B2(n_3732),
.Y(n_4029)
);

OAI21x1_ASAP7_75t_L g4030 ( 
.A1(n_3965),
.A2(n_4015),
.B(n_4008),
.Y(n_4030)
);

NAND2x1p5_ASAP7_75t_L g4031 ( 
.A(n_3950),
.B(n_3660),
.Y(n_4031)
);

CKINVDCx6p67_ASAP7_75t_R g4032 ( 
.A(n_3872),
.Y(n_4032)
);

INVx1_ASAP7_75t_L g4033 ( 
.A(n_3890),
.Y(n_4033)
);

INVxp67_ASAP7_75t_L g4034 ( 
.A(n_4008),
.Y(n_4034)
);

AOI22xp33_ASAP7_75t_SL g4035 ( 
.A1(n_3850),
.A2(n_3685),
.B1(n_3785),
.B2(n_3803),
.Y(n_4035)
);

AOI22xp33_ASAP7_75t_L g4036 ( 
.A1(n_3877),
.A2(n_3744),
.B1(n_3715),
.B2(n_3820),
.Y(n_4036)
);

AO31x2_ASAP7_75t_L g4037 ( 
.A1(n_3995),
.A2(n_3650),
.A3(n_3701),
.B(n_3817),
.Y(n_4037)
);

AND2x4_ASAP7_75t_L g4038 ( 
.A(n_4005),
.B(n_3823),
.Y(n_4038)
);

NAND2xp5_ASAP7_75t_L g4039 ( 
.A(n_3901),
.B(n_3737),
.Y(n_4039)
);

OR2x2_ASAP7_75t_L g4040 ( 
.A(n_3898),
.B(n_3737),
.Y(n_4040)
);

OAI22xp5_ASAP7_75t_L g4041 ( 
.A1(n_3960),
.A2(n_3715),
.B1(n_3792),
.B2(n_3685),
.Y(n_4041)
);

CKINVDCx5p33_ASAP7_75t_R g4042 ( 
.A(n_3891),
.Y(n_4042)
);

INVx1_ASAP7_75t_L g4043 ( 
.A(n_3890),
.Y(n_4043)
);

INVx1_ASAP7_75t_L g4044 ( 
.A(n_3907),
.Y(n_4044)
);

AOI21xp5_ASAP7_75t_L g4045 ( 
.A1(n_4021),
.A2(n_3660),
.B(n_3718),
.Y(n_4045)
);

OR2x2_ASAP7_75t_L g4046 ( 
.A(n_3963),
.B(n_3737),
.Y(n_4046)
);

OAI21x1_ASAP7_75t_L g4047 ( 
.A1(n_4012),
.A2(n_3791),
.B(n_3823),
.Y(n_4047)
);

OA21x2_ASAP7_75t_L g4048 ( 
.A1(n_4012),
.A2(n_3805),
.B(n_3682),
.Y(n_4048)
);

OAI21x1_ASAP7_75t_L g4049 ( 
.A1(n_3917),
.A2(n_3725),
.B(n_3810),
.Y(n_4049)
);

OR2x2_ASAP7_75t_L g4050 ( 
.A(n_3857),
.B(n_3686),
.Y(n_4050)
);

INVx1_ASAP7_75t_L g4051 ( 
.A(n_3907),
.Y(n_4051)
);

AND2x2_ASAP7_75t_L g4052 ( 
.A(n_3888),
.B(n_3704),
.Y(n_4052)
);

INVx1_ASAP7_75t_L g4053 ( 
.A(n_3964),
.Y(n_4053)
);

AND2x2_ASAP7_75t_L g4054 ( 
.A(n_3981),
.B(n_3680),
.Y(n_4054)
);

O2A1O1Ixp33_ASAP7_75t_SL g4055 ( 
.A1(n_3887),
.A2(n_3777),
.B(n_3834),
.C(n_3784),
.Y(n_4055)
);

OR2x2_ASAP7_75t_L g4056 ( 
.A(n_3978),
.B(n_3964),
.Y(n_4056)
);

BUFx2_ASAP7_75t_L g4057 ( 
.A(n_4005),
.Y(n_4057)
);

INVx3_ASAP7_75t_L g4058 ( 
.A(n_3917),
.Y(n_4058)
);

INVx6_ASAP7_75t_L g4059 ( 
.A(n_3950),
.Y(n_4059)
);

INVx1_ASAP7_75t_SL g4060 ( 
.A(n_3900),
.Y(n_4060)
);

OAI21x1_ASAP7_75t_L g4061 ( 
.A1(n_3943),
.A2(n_3731),
.B(n_3707),
.Y(n_4061)
);

BUFx2_ASAP7_75t_R g4062 ( 
.A(n_3847),
.Y(n_4062)
);

OR2x2_ASAP7_75t_L g4063 ( 
.A(n_3971),
.B(n_3686),
.Y(n_4063)
);

AOI22xp33_ASAP7_75t_L g4064 ( 
.A1(n_3975),
.A2(n_3825),
.B1(n_3677),
.B2(n_3787),
.Y(n_4064)
);

AND2x2_ASAP7_75t_L g4065 ( 
.A(n_3932),
.B(n_3680),
.Y(n_4065)
);

OAI21x1_ASAP7_75t_L g4066 ( 
.A1(n_3943),
.A2(n_3771),
.B(n_3784),
.Y(n_4066)
);

AOI22xp33_ASAP7_75t_L g4067 ( 
.A1(n_3874),
.A2(n_3798),
.B1(n_3793),
.B2(n_3675),
.Y(n_4067)
);

INVx1_ASAP7_75t_L g4068 ( 
.A(n_3971),
.Y(n_4068)
);

INVx2_ASAP7_75t_SL g4069 ( 
.A(n_3946),
.Y(n_4069)
);

INVx3_ASAP7_75t_L g4070 ( 
.A(n_3931),
.Y(n_4070)
);

AND2x4_ASAP7_75t_L g4071 ( 
.A(n_3870),
.B(n_3686),
.Y(n_4071)
);

A2O1A1Ixp33_ASAP7_75t_L g4072 ( 
.A1(n_3849),
.A2(n_3863),
.B(n_3930),
.C(n_3936),
.Y(n_4072)
);

NAND2xp5_ASAP7_75t_L g4073 ( 
.A(n_3977),
.B(n_3815),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_3977),
.Y(n_4074)
);

NAND2x1_ASAP7_75t_L g4075 ( 
.A(n_3927),
.B(n_3740),
.Y(n_4075)
);

OAI21xp5_ASAP7_75t_L g4076 ( 
.A1(n_3861),
.A2(n_3799),
.B(n_3830),
.Y(n_4076)
);

OAI22xp5_ASAP7_75t_L g4077 ( 
.A1(n_3987),
.A2(n_3797),
.B1(n_3691),
.B2(n_3705),
.Y(n_4077)
);

INVx2_ASAP7_75t_L g4078 ( 
.A(n_3879),
.Y(n_4078)
);

OAI21xp5_ASAP7_75t_L g4079 ( 
.A1(n_3947),
.A2(n_3831),
.B(n_3804),
.Y(n_4079)
);

HB1xp67_ASAP7_75t_L g4080 ( 
.A(n_3927),
.Y(n_4080)
);

BUFx2_ASAP7_75t_SL g4081 ( 
.A(n_3931),
.Y(n_4081)
);

OAI21x1_ASAP7_75t_L g4082 ( 
.A1(n_3880),
.A2(n_3772),
.B(n_3676),
.Y(n_4082)
);

BUFx8_ASAP7_75t_SL g4083 ( 
.A(n_4025),
.Y(n_4083)
);

INVx1_ASAP7_75t_L g4084 ( 
.A(n_3862),
.Y(n_4084)
);

INVx2_ASAP7_75t_L g4085 ( 
.A(n_3884),
.Y(n_4085)
);

BUFx3_ASAP7_75t_L g4086 ( 
.A(n_3855),
.Y(n_4086)
);

O2A1O1Ixp33_ASAP7_75t_SL g4087 ( 
.A1(n_4002),
.A2(n_3941),
.B(n_3951),
.C(n_3866),
.Y(n_4087)
);

INVx2_ASAP7_75t_L g4088 ( 
.A(n_3892),
.Y(n_4088)
);

INVx1_ASAP7_75t_L g4089 ( 
.A(n_3882),
.Y(n_4089)
);

OR2x2_ASAP7_75t_L g4090 ( 
.A(n_3916),
.B(n_3920),
.Y(n_4090)
);

OA21x2_ASAP7_75t_L g4091 ( 
.A1(n_3846),
.A2(n_3750),
.B(n_3730),
.Y(n_4091)
);

AOI22xp33_ASAP7_75t_L g4092 ( 
.A1(n_3944),
.A2(n_3764),
.B1(n_3745),
.B2(n_3765),
.Y(n_4092)
);

AOI22xp5_ASAP7_75t_L g4093 ( 
.A1(n_3973),
.A2(n_3691),
.B1(n_3705),
.B2(n_3829),
.Y(n_4093)
);

BUFx2_ASAP7_75t_L g4094 ( 
.A(n_3982),
.Y(n_4094)
);

BUFx2_ASAP7_75t_R g4095 ( 
.A(n_3928),
.Y(n_4095)
);

AOI22xp33_ASAP7_75t_L g4096 ( 
.A1(n_3860),
.A2(n_3649),
.B1(n_3828),
.B2(n_3788),
.Y(n_4096)
);

OAI21x1_ASAP7_75t_L g4097 ( 
.A1(n_3903),
.A2(n_3829),
.B(n_3753),
.Y(n_4097)
);

HB1xp67_ASAP7_75t_L g4098 ( 
.A(n_3955),
.Y(n_4098)
);

BUFx2_ASAP7_75t_L g4099 ( 
.A(n_3982),
.Y(n_4099)
);

OAI21x1_ASAP7_75t_L g4100 ( 
.A1(n_3962),
.A2(n_3727),
.B(n_3700),
.Y(n_4100)
);

AOI22x1_ASAP7_75t_L g4101 ( 
.A1(n_3868),
.A2(n_3833),
.B1(n_3828),
.B2(n_3780),
.Y(n_4101)
);

OR2x2_ASAP7_75t_L g4102 ( 
.A(n_3983),
.B(n_3657),
.Y(n_4102)
);

HB1xp67_ASAP7_75t_L g4103 ( 
.A(n_3991),
.Y(n_4103)
);

AND2x4_ASAP7_75t_L g4104 ( 
.A(n_3870),
.B(n_3833),
.Y(n_4104)
);

OAI21x1_ASAP7_75t_L g4105 ( 
.A1(n_3899),
.A2(n_3716),
.B(n_3746),
.Y(n_4105)
);

AND2x2_ASAP7_75t_L g4106 ( 
.A(n_3851),
.B(n_3747),
.Y(n_4106)
);

AO21x2_ASAP7_75t_L g4107 ( 
.A1(n_4007),
.A2(n_3728),
.B(n_3815),
.Y(n_4107)
);

AND2x2_ASAP7_75t_L g4108 ( 
.A(n_3967),
.B(n_3828),
.Y(n_4108)
);

OA21x2_ASAP7_75t_L g4109 ( 
.A1(n_3856),
.A2(n_3815),
.B(n_3657),
.Y(n_4109)
);

INVxp67_ASAP7_75t_SL g4110 ( 
.A(n_3990),
.Y(n_4110)
);

NOR2xp67_ASAP7_75t_L g4111 ( 
.A(n_3950),
.B(n_206),
.Y(n_4111)
);

OAI21x1_ASAP7_75t_L g4112 ( 
.A1(n_3893),
.A2(n_3657),
.B(n_3673),
.Y(n_4112)
);

OAI22xp5_ASAP7_75t_L g4113 ( 
.A1(n_4023),
.A2(n_3673),
.B1(n_248),
.B2(n_249),
.Y(n_4113)
);

INVx2_ASAP7_75t_L g4114 ( 
.A(n_3910),
.Y(n_4114)
);

NOR2xp67_ASAP7_75t_L g4115 ( 
.A(n_3926),
.B(n_206),
.Y(n_4115)
);

INVx2_ASAP7_75t_L g4116 ( 
.A(n_3914),
.Y(n_4116)
);

AO21x2_ASAP7_75t_L g4117 ( 
.A1(n_3942),
.A2(n_3673),
.B(n_3762),
.Y(n_4117)
);

INVx2_ASAP7_75t_SL g4118 ( 
.A(n_3945),
.Y(n_4118)
);

BUFx2_ASAP7_75t_L g4119 ( 
.A(n_3974),
.Y(n_4119)
);

INVx1_ASAP7_75t_L g4120 ( 
.A(n_3952),
.Y(n_4120)
);

INVx1_ASAP7_75t_L g4121 ( 
.A(n_3919),
.Y(n_4121)
);

INVx1_ASAP7_75t_L g4122 ( 
.A(n_3925),
.Y(n_4122)
);

A2O1A1Ixp33_ASAP7_75t_L g4123 ( 
.A1(n_3883),
.A2(n_209),
.B(n_207),
.C(n_208),
.Y(n_4123)
);

AND2x2_ASAP7_75t_L g4124 ( 
.A(n_4026),
.B(n_3776),
.Y(n_4124)
);

A2O1A1Ixp33_ASAP7_75t_L g4125 ( 
.A1(n_3969),
.A2(n_210),
.B(n_207),
.C(n_209),
.Y(n_4125)
);

OAI21x1_ASAP7_75t_L g4126 ( 
.A1(n_3929),
.A2(n_3776),
.B(n_3762),
.Y(n_4126)
);

OAI21x1_ASAP7_75t_L g4127 ( 
.A1(n_3915),
.A2(n_3776),
.B(n_3762),
.Y(n_4127)
);

INVx1_ASAP7_75t_L g4128 ( 
.A(n_3939),
.Y(n_4128)
);

HB1xp67_ASAP7_75t_L g4129 ( 
.A(n_3886),
.Y(n_4129)
);

OAI21xp5_ASAP7_75t_L g4130 ( 
.A1(n_3961),
.A2(n_207),
.B(n_209),
.Y(n_4130)
);

OAI21x1_ASAP7_75t_L g4131 ( 
.A1(n_4014),
.A2(n_3775),
.B(n_3778),
.Y(n_4131)
);

INVx1_ASAP7_75t_L g4132 ( 
.A(n_3940),
.Y(n_4132)
);

AND2x2_ASAP7_75t_L g4133 ( 
.A(n_3894),
.B(n_3775),
.Y(n_4133)
);

INVx3_ASAP7_75t_SL g4134 ( 
.A(n_3869),
.Y(n_4134)
);

INVx2_ASAP7_75t_L g4135 ( 
.A(n_4009),
.Y(n_4135)
);

INVx1_ASAP7_75t_L g4136 ( 
.A(n_3911),
.Y(n_4136)
);

INVx1_ASAP7_75t_L g4137 ( 
.A(n_3924),
.Y(n_4137)
);

A2O1A1Ixp33_ASAP7_75t_L g4138 ( 
.A1(n_3968),
.A2(n_212),
.B(n_210),
.C(n_211),
.Y(n_4138)
);

NAND2xp5_ASAP7_75t_L g4139 ( 
.A(n_3958),
.B(n_3775),
.Y(n_4139)
);

INVx2_ASAP7_75t_L g4140 ( 
.A(n_4016),
.Y(n_4140)
);

OAI21x1_ASAP7_75t_L g4141 ( 
.A1(n_4017),
.A2(n_3778),
.B(n_210),
.Y(n_4141)
);

HB1xp67_ASAP7_75t_L g4142 ( 
.A(n_3886),
.Y(n_4142)
);

OAI21x1_ASAP7_75t_L g4143 ( 
.A1(n_3993),
.A2(n_3778),
.B(n_211),
.Y(n_4143)
);

OAI21xp5_ASAP7_75t_L g4144 ( 
.A1(n_4003),
.A2(n_212),
.B(n_213),
.Y(n_4144)
);

AOI22xp33_ASAP7_75t_L g4145 ( 
.A1(n_3949),
.A2(n_214),
.B1(n_212),
.B2(n_213),
.Y(n_4145)
);

OAI22xp5_ASAP7_75t_L g4146 ( 
.A1(n_3996),
.A2(n_249),
.B1(n_250),
.B2(n_246),
.Y(n_4146)
);

OA21x2_ASAP7_75t_L g4147 ( 
.A1(n_3858),
.A2(n_3865),
.B(n_3956),
.Y(n_4147)
);

NAND2xp5_ASAP7_75t_L g4148 ( 
.A(n_3886),
.B(n_213),
.Y(n_4148)
);

AND2x2_ASAP7_75t_L g4149 ( 
.A(n_3895),
.B(n_215),
.Y(n_4149)
);

AOI22xp33_ASAP7_75t_L g4150 ( 
.A1(n_3878),
.A2(n_217),
.B1(n_215),
.B2(n_216),
.Y(n_4150)
);

INVx1_ASAP7_75t_L g4151 ( 
.A(n_3881),
.Y(n_4151)
);

OAI21x1_ASAP7_75t_L g4152 ( 
.A1(n_3897),
.A2(n_215),
.B(n_216),
.Y(n_4152)
);

OAI21x1_ASAP7_75t_L g4153 ( 
.A1(n_3998),
.A2(n_4018),
.B(n_3997),
.Y(n_4153)
);

AND2x6_ASAP7_75t_L g4154 ( 
.A(n_3918),
.B(n_250),
.Y(n_4154)
);

AND2x2_ASAP7_75t_L g4155 ( 
.A(n_3954),
.B(n_216),
.Y(n_4155)
);

AND2x4_ASAP7_75t_L g4156 ( 
.A(n_3984),
.B(n_217),
.Y(n_4156)
);

INVx3_ASAP7_75t_L g4157 ( 
.A(n_3976),
.Y(n_4157)
);

NAND2xp5_ASAP7_75t_SL g4158 ( 
.A(n_3935),
.B(n_251),
.Y(n_4158)
);

NAND2xp5_ASAP7_75t_L g4159 ( 
.A(n_4027),
.B(n_217),
.Y(n_4159)
);

NAND2x1p5_ASAP7_75t_L g4160 ( 
.A(n_3976),
.B(n_252),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_3957),
.Y(n_4161)
);

AND2x2_ASAP7_75t_L g4162 ( 
.A(n_3976),
.B(n_252),
.Y(n_4162)
);

BUFx12f_ASAP7_75t_L g4163 ( 
.A(n_3869),
.Y(n_4163)
);

AND2x4_ASAP7_75t_L g4164 ( 
.A(n_3974),
.B(n_253),
.Y(n_4164)
);

AOI22xp33_ASAP7_75t_L g4165 ( 
.A1(n_3896),
.A2(n_256),
.B1(n_254),
.B2(n_255),
.Y(n_4165)
);

AOI222xp33_ASAP7_75t_L g4166 ( 
.A1(n_3871),
.A2(n_256),
.B1(n_258),
.B2(n_254),
.C1(n_255),
.C2(n_257),
.Y(n_4166)
);

AOI22xp33_ASAP7_75t_L g4167 ( 
.A1(n_3979),
.A2(n_259),
.B1(n_257),
.B2(n_258),
.Y(n_4167)
);

OA21x2_ASAP7_75t_L g4168 ( 
.A1(n_3986),
.A2(n_3966),
.B(n_4004),
.Y(n_4168)
);

A2O1A1Ixp33_ASAP7_75t_L g4169 ( 
.A1(n_3876),
.A2(n_261),
.B(n_259),
.C(n_260),
.Y(n_4169)
);

NAND2xp5_ASAP7_75t_SL g4170 ( 
.A(n_3935),
.B(n_260),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_3957),
.Y(n_4171)
);

OAI21x1_ASAP7_75t_L g4172 ( 
.A1(n_3864),
.A2(n_261),
.B(n_262),
.Y(n_4172)
);

OAI21x1_ASAP7_75t_L g4173 ( 
.A1(n_4013),
.A2(n_263),
.B(n_264),
.Y(n_4173)
);

INVx6_ASAP7_75t_L g4174 ( 
.A(n_3945),
.Y(n_4174)
);

OAI21xp33_ASAP7_75t_L g4175 ( 
.A1(n_3867),
.A2(n_263),
.B(n_264),
.Y(n_4175)
);

OAI22xp5_ASAP7_75t_L g4176 ( 
.A1(n_3885),
.A2(n_267),
.B1(n_265),
.B2(n_266),
.Y(n_4176)
);

OAI21x1_ASAP7_75t_L g4177 ( 
.A1(n_4006),
.A2(n_265),
.B(n_266),
.Y(n_4177)
);

INVx2_ASAP7_75t_L g4178 ( 
.A(n_3923),
.Y(n_4178)
);

INVx3_ASAP7_75t_L g4179 ( 
.A(n_3985),
.Y(n_4179)
);

INVx1_ASAP7_75t_L g4180 ( 
.A(n_3957),
.Y(n_4180)
);

AOI221xp5_ASAP7_75t_L g4181 ( 
.A1(n_3873),
.A2(n_269),
.B1(n_267),
.B2(n_268),
.C(n_270),
.Y(n_4181)
);

INVx3_ASAP7_75t_L g4182 ( 
.A(n_4174),
.Y(n_4182)
);

OAI21x1_ASAP7_75t_L g4183 ( 
.A1(n_4030),
.A2(n_3848),
.B(n_3902),
.Y(n_4183)
);

OA21x2_ASAP7_75t_L g4184 ( 
.A1(n_4039),
.A2(n_3908),
.B(n_3854),
.Y(n_4184)
);

NAND2xp5_ASAP7_75t_L g4185 ( 
.A(n_4080),
.B(n_4000),
.Y(n_4185)
);

OAI21x1_ASAP7_75t_L g4186 ( 
.A1(n_4047),
.A2(n_3938),
.B(n_3937),
.Y(n_4186)
);

AND2x2_ASAP7_75t_L g4187 ( 
.A(n_4057),
.B(n_3985),
.Y(n_4187)
);

NAND2x1p5_ASAP7_75t_L g4188 ( 
.A(n_4164),
.B(n_3985),
.Y(n_4188)
);

OAI21xp5_ASAP7_75t_L g4189 ( 
.A1(n_4113),
.A2(n_3948),
.B(n_4022),
.Y(n_4189)
);

AND2x2_ASAP7_75t_L g4190 ( 
.A(n_4054),
.B(n_3935),
.Y(n_4190)
);

NAND2xp5_ASAP7_75t_L g4191 ( 
.A(n_4080),
.B(n_3923),
.Y(n_4191)
);

OAI21x1_ASAP7_75t_L g4192 ( 
.A1(n_4039),
.A2(n_3906),
.B(n_3904),
.Y(n_4192)
);

NAND2xp5_ASAP7_75t_L g4193 ( 
.A(n_4098),
.B(n_3923),
.Y(n_4193)
);

AO21x2_ASAP7_75t_L g4194 ( 
.A1(n_4148),
.A2(n_3859),
.B(n_3922),
.Y(n_4194)
);

OR2x2_ASAP7_75t_L g4195 ( 
.A(n_4151),
.B(n_3909),
.Y(n_4195)
);

INVx1_ASAP7_75t_L g4196 ( 
.A(n_4098),
.Y(n_4196)
);

NAND2xp5_ASAP7_75t_L g4197 ( 
.A(n_4103),
.B(n_3974),
.Y(n_4197)
);

INVx4_ASAP7_75t_L g4198 ( 
.A(n_4042),
.Y(n_4198)
);

HB1xp67_ASAP7_75t_L g4199 ( 
.A(n_4103),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_4090),
.Y(n_4200)
);

HB1xp67_ASAP7_75t_L g4201 ( 
.A(n_4063),
.Y(n_4201)
);

OAI21x1_ASAP7_75t_L g4202 ( 
.A1(n_4073),
.A2(n_4112),
.B(n_4050),
.Y(n_4202)
);

NAND2xp5_ASAP7_75t_L g4203 ( 
.A(n_4034),
.B(n_3974),
.Y(n_4203)
);

OR2x2_ASAP7_75t_L g4204 ( 
.A(n_4120),
.B(n_3912),
.Y(n_4204)
);

OA21x2_ASAP7_75t_L g4205 ( 
.A1(n_4034),
.A2(n_4011),
.B(n_4001),
.Y(n_4205)
);

AO21x2_ASAP7_75t_L g4206 ( 
.A1(n_4148),
.A2(n_3988),
.B(n_3999),
.Y(n_4206)
);

NAND2xp5_ASAP7_75t_L g4207 ( 
.A(n_4110),
.B(n_3912),
.Y(n_4207)
);

OR2x2_ASAP7_75t_L g4208 ( 
.A(n_4040),
.B(n_3912),
.Y(n_4208)
);

NAND2xp5_ASAP7_75t_L g4209 ( 
.A(n_4110),
.B(n_3992),
.Y(n_4209)
);

CKINVDCx11_ASAP7_75t_R g4210 ( 
.A(n_4032),
.Y(n_4210)
);

OAI21x1_ASAP7_75t_SL g4211 ( 
.A1(n_4069),
.A2(n_3953),
.B(n_3889),
.Y(n_4211)
);

AOI21xp5_ASAP7_75t_L g4212 ( 
.A1(n_4113),
.A2(n_3980),
.B(n_3970),
.Y(n_4212)
);

OAI21x1_ASAP7_75t_L g4213 ( 
.A1(n_4073),
.A2(n_4045),
.B(n_4139),
.Y(n_4213)
);

AOI21xp5_ASAP7_75t_L g4214 ( 
.A1(n_4087),
.A2(n_3852),
.B(n_4010),
.Y(n_4214)
);

INVx1_ASAP7_75t_L g4215 ( 
.A(n_4033),
.Y(n_4215)
);

OA21x2_ASAP7_75t_L g4216 ( 
.A1(n_4078),
.A2(n_3989),
.B(n_3934),
.Y(n_4216)
);

HB1xp67_ASAP7_75t_L g4217 ( 
.A(n_4056),
.Y(n_4217)
);

INVx1_ASAP7_75t_L g4218 ( 
.A(n_4043),
.Y(n_4218)
);

INVx2_ASAP7_75t_L g4219 ( 
.A(n_4124),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_4044),
.Y(n_4220)
);

BUFx12f_ASAP7_75t_L g4221 ( 
.A(n_4163),
.Y(n_4221)
);

AO31x2_ASAP7_75t_L g4222 ( 
.A1(n_4161),
.A2(n_4171),
.A3(n_4180),
.B(n_4178),
.Y(n_4222)
);

AO21x2_ASAP7_75t_L g4223 ( 
.A1(n_4129),
.A2(n_4020),
.B(n_3994),
.Y(n_4223)
);

INVx1_ASAP7_75t_L g4224 ( 
.A(n_4051),
.Y(n_4224)
);

NOR2xp33_ASAP7_75t_L g4225 ( 
.A(n_4062),
.B(n_3905),
.Y(n_4225)
);

INVx2_ASAP7_75t_L g4226 ( 
.A(n_4102),
.Y(n_4226)
);

AO31x2_ASAP7_75t_L g4227 ( 
.A1(n_4041),
.A2(n_4019),
.A3(n_3921),
.B(n_3913),
.Y(n_4227)
);

CKINVDCx5p33_ASAP7_75t_R g4228 ( 
.A(n_4083),
.Y(n_4228)
);

INVx2_ASAP7_75t_L g4229 ( 
.A(n_4094),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_4053),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_4068),
.Y(n_4231)
);

BUFx2_ASAP7_75t_L g4232 ( 
.A(n_4086),
.Y(n_4232)
);

INVx4_ASAP7_75t_SL g4233 ( 
.A(n_4134),
.Y(n_4233)
);

NAND2x1p5_ASAP7_75t_L g4234 ( 
.A(n_4164),
.B(n_3875),
.Y(n_4234)
);

INVx3_ASAP7_75t_L g4235 ( 
.A(n_4174),
.Y(n_4235)
);

CKINVDCx20_ASAP7_75t_R g4236 ( 
.A(n_4060),
.Y(n_4236)
);

INVx1_ASAP7_75t_L g4237 ( 
.A(n_4074),
.Y(n_4237)
);

NAND2xp5_ASAP7_75t_L g4238 ( 
.A(n_4071),
.B(n_3972),
.Y(n_4238)
);

AOI22xp5_ASAP7_75t_L g4239 ( 
.A1(n_4175),
.A2(n_3852),
.B1(n_3933),
.B2(n_4024),
.Y(n_4239)
);

AOI21xp5_ASAP7_75t_L g4240 ( 
.A1(n_4075),
.A2(n_268),
.B(n_269),
.Y(n_4240)
);

AND2x2_ASAP7_75t_L g4241 ( 
.A(n_4052),
.B(n_270),
.Y(n_4241)
);

OAI21x1_ASAP7_75t_L g4242 ( 
.A1(n_4045),
.A2(n_271),
.B(n_272),
.Y(n_4242)
);

OAI22xp5_ASAP7_75t_L g4243 ( 
.A1(n_4064),
.A2(n_274),
.B1(n_272),
.B2(n_273),
.Y(n_4243)
);

NAND2xp5_ASAP7_75t_L g4244 ( 
.A(n_4071),
.B(n_275),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_4084),
.Y(n_4245)
);

OAI21x1_ASAP7_75t_L g4246 ( 
.A1(n_4139),
.A2(n_275),
.B(n_277),
.Y(n_4246)
);

INVx1_ASAP7_75t_L g4247 ( 
.A(n_4089),
.Y(n_4247)
);

NAND2xp5_ASAP7_75t_L g4248 ( 
.A(n_4129),
.B(n_277),
.Y(n_4248)
);

BUFx10_ASAP7_75t_L g4249 ( 
.A(n_4059),
.Y(n_4249)
);

AO21x2_ASAP7_75t_L g4250 ( 
.A1(n_4142),
.A2(n_278),
.B(n_279),
.Y(n_4250)
);

NOR2xp33_ASAP7_75t_L g4251 ( 
.A(n_4062),
.B(n_278),
.Y(n_4251)
);

NAND2xp5_ASAP7_75t_SL g4252 ( 
.A(n_4119),
.B(n_4060),
.Y(n_4252)
);

INVx1_ASAP7_75t_L g4253 ( 
.A(n_4142),
.Y(n_4253)
);

AND2x4_ASAP7_75t_L g4254 ( 
.A(n_4070),
.B(n_4099),
.Y(n_4254)
);

HB1xp67_ASAP7_75t_L g4255 ( 
.A(n_4109),
.Y(n_4255)
);

NAND2xp5_ASAP7_75t_L g4256 ( 
.A(n_4147),
.B(n_279),
.Y(n_4256)
);

INVx1_ASAP7_75t_L g4257 ( 
.A(n_4028),
.Y(n_4257)
);

HB1xp67_ASAP7_75t_L g4258 ( 
.A(n_4109),
.Y(n_4258)
);

OA21x2_ASAP7_75t_L g4259 ( 
.A1(n_4085),
.A2(n_280),
.B(n_282),
.Y(n_4259)
);

AO21x2_ASAP7_75t_L g4260 ( 
.A1(n_4159),
.A2(n_280),
.B(n_282),
.Y(n_4260)
);

INVx2_ASAP7_75t_L g4261 ( 
.A(n_4088),
.Y(n_4261)
);

OR2x2_ASAP7_75t_L g4262 ( 
.A(n_4136),
.B(n_283),
.Y(n_4262)
);

NAND2xp5_ASAP7_75t_L g4263 ( 
.A(n_4147),
.B(n_283),
.Y(n_4263)
);

OAI21x1_ASAP7_75t_SL g4264 ( 
.A1(n_4159),
.A2(n_284),
.B(n_285),
.Y(n_4264)
);

NAND2xp5_ASAP7_75t_L g4265 ( 
.A(n_4137),
.B(n_284),
.Y(n_4265)
);

OR2x2_ASAP7_75t_L g4266 ( 
.A(n_4135),
.B(n_285),
.Y(n_4266)
);

OA21x2_ASAP7_75t_L g4267 ( 
.A1(n_4046),
.A2(n_286),
.B(n_287),
.Y(n_4267)
);

CKINVDCx5p33_ASAP7_75t_R g4268 ( 
.A(n_4134),
.Y(n_4268)
);

NAND2xp5_ASAP7_75t_L g4269 ( 
.A(n_4133),
.B(n_286),
.Y(n_4269)
);

INVx1_ASAP7_75t_L g4270 ( 
.A(n_4140),
.Y(n_4270)
);

AOI21xp5_ASAP7_75t_L g4271 ( 
.A1(n_4041),
.A2(n_288),
.B(n_289),
.Y(n_4271)
);

INVx2_ASAP7_75t_L g4272 ( 
.A(n_4114),
.Y(n_4272)
);

AND2x2_ASAP7_75t_L g4273 ( 
.A(n_4065),
.B(n_288),
.Y(n_4273)
);

AO21x2_ASAP7_75t_L g4274 ( 
.A1(n_4117),
.A2(n_289),
.B(n_290),
.Y(n_4274)
);

INVx2_ASAP7_75t_L g4275 ( 
.A(n_4116),
.Y(n_4275)
);

AOI21xp5_ASAP7_75t_L g4276 ( 
.A1(n_4146),
.A2(n_291),
.B(n_292),
.Y(n_4276)
);

NOR2xp33_ASAP7_75t_L g4277 ( 
.A(n_4070),
.B(n_291),
.Y(n_4277)
);

NAND2xp5_ASAP7_75t_L g4278 ( 
.A(n_4037),
.B(n_292),
.Y(n_4278)
);

HB1xp67_ASAP7_75t_L g4279 ( 
.A(n_4107),
.Y(n_4279)
);

AO31x2_ASAP7_75t_L g4280 ( 
.A1(n_4077),
.A2(n_295),
.A3(n_293),
.B(n_294),
.Y(n_4280)
);

OAI21x1_ASAP7_75t_L g4281 ( 
.A1(n_4058),
.A2(n_293),
.B(n_294),
.Y(n_4281)
);

INVx3_ASAP7_75t_L g4282 ( 
.A(n_4174),
.Y(n_4282)
);

AND2x2_ASAP7_75t_L g4283 ( 
.A(n_4108),
.B(n_295),
.Y(n_4283)
);

BUFx6f_ASAP7_75t_L g4284 ( 
.A(n_4160),
.Y(n_4284)
);

OAI22xp5_ASAP7_75t_L g4285 ( 
.A1(n_4064),
.A2(n_298),
.B1(n_296),
.B2(n_297),
.Y(n_4285)
);

OA21x2_ASAP7_75t_L g4286 ( 
.A1(n_4066),
.A2(n_4082),
.B(n_4061),
.Y(n_4286)
);

INVx1_ASAP7_75t_SL g4287 ( 
.A(n_4081),
.Y(n_4287)
);

OAI21x1_ASAP7_75t_L g4288 ( 
.A1(n_4058),
.A2(n_297),
.B(n_299),
.Y(n_4288)
);

OAI21x1_ASAP7_75t_SL g4289 ( 
.A1(n_4118),
.A2(n_4079),
.B(n_4076),
.Y(n_4289)
);

INVx1_ASAP7_75t_L g4290 ( 
.A(n_4121),
.Y(n_4290)
);

AOI21xp5_ASAP7_75t_L g4291 ( 
.A1(n_4146),
.A2(n_299),
.B(n_300),
.Y(n_4291)
);

OAI21x1_ASAP7_75t_L g4292 ( 
.A1(n_4126),
.A2(n_300),
.B(n_301),
.Y(n_4292)
);

AOI21xp5_ASAP7_75t_L g4293 ( 
.A1(n_4176),
.A2(n_303),
.B(n_304),
.Y(n_4293)
);

AND2x4_ASAP7_75t_L g4294 ( 
.A(n_4104),
.B(n_303),
.Y(n_4294)
);

OAI21x1_ASAP7_75t_L g4295 ( 
.A1(n_4127),
.A2(n_304),
.B(n_305),
.Y(n_4295)
);

AOI21x1_ASAP7_75t_L g4296 ( 
.A1(n_4115),
.A2(n_307),
.B(n_308),
.Y(n_4296)
);

AND2x2_ASAP7_75t_L g4297 ( 
.A(n_4106),
.B(n_307),
.Y(n_4297)
);

INVx1_ASAP7_75t_L g4298 ( 
.A(n_4122),
.Y(n_4298)
);

INVx4_ASAP7_75t_SL g4299 ( 
.A(n_4154),
.Y(n_4299)
);

AOI21xp5_ASAP7_75t_L g4300 ( 
.A1(n_4176),
.A2(n_308),
.B(n_309),
.Y(n_4300)
);

OAI21x1_ASAP7_75t_L g4301 ( 
.A1(n_4131),
.A2(n_309),
.B(n_310),
.Y(n_4301)
);

OAI21x1_ASAP7_75t_SL g4302 ( 
.A1(n_4079),
.A2(n_312),
.B(n_313),
.Y(n_4302)
);

OR2x6_ASAP7_75t_L g4303 ( 
.A(n_4111),
.B(n_312),
.Y(n_4303)
);

OAI21x1_ASAP7_75t_L g4304 ( 
.A1(n_4100),
.A2(n_314),
.B(n_315),
.Y(n_4304)
);

INVx1_ASAP7_75t_L g4305 ( 
.A(n_4128),
.Y(n_4305)
);

OAI21x1_ASAP7_75t_L g4306 ( 
.A1(n_4031),
.A2(n_314),
.B(n_316),
.Y(n_4306)
);

NAND2xp5_ASAP7_75t_L g4307 ( 
.A(n_4037),
.B(n_317),
.Y(n_4307)
);

NAND2xp5_ASAP7_75t_L g4308 ( 
.A(n_4037),
.B(n_317),
.Y(n_4308)
);

OA21x2_ASAP7_75t_L g4309 ( 
.A1(n_4132),
.A2(n_319),
.B(n_320),
.Y(n_4309)
);

INVx2_ASAP7_75t_L g4310 ( 
.A(n_4048),
.Y(n_4310)
);

BUFx3_ASAP7_75t_L g4311 ( 
.A(n_4149),
.Y(n_4311)
);

AO31x2_ASAP7_75t_L g4312 ( 
.A1(n_4077),
.A2(n_322),
.A3(n_320),
.B(n_321),
.Y(n_4312)
);

OAI21x1_ASAP7_75t_L g4313 ( 
.A1(n_4031),
.A2(n_321),
.B(n_322),
.Y(n_4313)
);

HB1xp67_ASAP7_75t_L g4314 ( 
.A(n_4107),
.Y(n_4314)
);

NOR2xp33_ASAP7_75t_L g4315 ( 
.A(n_4156),
.B(n_323),
.Y(n_4315)
);

AND2x2_ASAP7_75t_L g4316 ( 
.A(n_4038),
.B(n_323),
.Y(n_4316)
);

INVx2_ASAP7_75t_L g4317 ( 
.A(n_4048),
.Y(n_4317)
);

AO222x2_ASAP7_75t_L g4318 ( 
.A1(n_4155),
.A2(n_326),
.B1(n_329),
.B2(n_324),
.C1(n_325),
.C2(n_328),
.Y(n_4318)
);

INVx1_ASAP7_75t_L g4319 ( 
.A(n_4095),
.Y(n_4319)
);

OA21x2_ASAP7_75t_L g4320 ( 
.A1(n_4153),
.A2(n_324),
.B(n_326),
.Y(n_4320)
);

OA21x2_ASAP7_75t_L g4321 ( 
.A1(n_4105),
.A2(n_328),
.B(n_329),
.Y(n_4321)
);

AO21x2_ASAP7_75t_L g4322 ( 
.A1(n_4117),
.A2(n_330),
.B(n_331),
.Y(n_4322)
);

INVx3_ASAP7_75t_L g4323 ( 
.A(n_4038),
.Y(n_4323)
);

BUFx4f_ASAP7_75t_L g4324 ( 
.A(n_4160),
.Y(n_4324)
);

NAND2xp5_ASAP7_75t_L g4325 ( 
.A(n_4091),
.B(n_330),
.Y(n_4325)
);

OAI21x1_ASAP7_75t_L g4326 ( 
.A1(n_4157),
.A2(n_331),
.B(n_332),
.Y(n_4326)
);

AOI21xp5_ASAP7_75t_L g4327 ( 
.A1(n_4072),
.A2(n_332),
.B(n_333),
.Y(n_4327)
);

OR2x2_ASAP7_75t_L g4328 ( 
.A(n_4157),
.B(n_4179),
.Y(n_4328)
);

INVx1_ASAP7_75t_L g4329 ( 
.A(n_4095),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_4091),
.Y(n_4330)
);

BUFx3_ASAP7_75t_L g4331 ( 
.A(n_4156),
.Y(n_4331)
);

INVx1_ASAP7_75t_L g4332 ( 
.A(n_4104),
.Y(n_4332)
);

BUFx8_ASAP7_75t_L g4333 ( 
.A(n_4162),
.Y(n_4333)
);

INVx2_ASAP7_75t_L g4334 ( 
.A(n_4049),
.Y(n_4334)
);

AND2x4_ASAP7_75t_L g4335 ( 
.A(n_4179),
.B(n_333),
.Y(n_4335)
);

INVx2_ASAP7_75t_L g4336 ( 
.A(n_4097),
.Y(n_4336)
);

AOI21xp5_ASAP7_75t_L g4337 ( 
.A1(n_4055),
.A2(n_334),
.B(n_335),
.Y(n_4337)
);

BUFx2_ASAP7_75t_L g4338 ( 
.A(n_4154),
.Y(n_4338)
);

AND2x4_ASAP7_75t_L g4339 ( 
.A(n_4093),
.B(n_334),
.Y(n_4339)
);

BUFx8_ASAP7_75t_L g4340 ( 
.A(n_4154),
.Y(n_4340)
);

OAI21x1_ASAP7_75t_L g4341 ( 
.A1(n_4092),
.A2(n_335),
.B(n_336),
.Y(n_4341)
);

OA21x2_ASAP7_75t_L g4342 ( 
.A1(n_4092),
.A2(n_337),
.B(n_338),
.Y(n_4342)
);

BUFx6f_ASAP7_75t_L g4343 ( 
.A(n_4172),
.Y(n_4343)
);

INVx2_ASAP7_75t_L g4344 ( 
.A(n_4143),
.Y(n_4344)
);

HB1xp67_ASAP7_75t_L g4345 ( 
.A(n_4168),
.Y(n_4345)
);

AND2x2_ASAP7_75t_L g4346 ( 
.A(n_4059),
.B(n_337),
.Y(n_4346)
);

INVx1_ASAP7_75t_L g4347 ( 
.A(n_4256),
.Y(n_4347)
);

OAI22xp5_ASAP7_75t_L g4348 ( 
.A1(n_4287),
.A2(n_4338),
.B1(n_4307),
.B2(n_4308),
.Y(n_4348)
);

AOI22xp33_ASAP7_75t_L g4349 ( 
.A1(n_4205),
.A2(n_4168),
.B1(n_4035),
.B2(n_4154),
.Y(n_4349)
);

NOR2x1p5_ASAP7_75t_L g4350 ( 
.A(n_4268),
.B(n_4154),
.Y(n_4350)
);

CKINVDCx5p33_ASAP7_75t_R g4351 ( 
.A(n_4228),
.Y(n_4351)
);

OAI22xp5_ASAP7_75t_L g4352 ( 
.A1(n_4287),
.A2(n_4035),
.B1(n_4150),
.B2(n_4096),
.Y(n_4352)
);

INVx1_ASAP7_75t_L g4353 ( 
.A(n_4256),
.Y(n_4353)
);

INVx1_ASAP7_75t_L g4354 ( 
.A(n_4263),
.Y(n_4354)
);

INVx4_ASAP7_75t_L g4355 ( 
.A(n_4233),
.Y(n_4355)
);

HB1xp67_ASAP7_75t_L g4356 ( 
.A(n_4325),
.Y(n_4356)
);

AOI22xp33_ASAP7_75t_SL g4357 ( 
.A1(n_4319),
.A2(n_4144),
.B1(n_4130),
.B2(n_4076),
.Y(n_4357)
);

NOR2xp33_ASAP7_75t_L g4358 ( 
.A(n_4198),
.B(n_4158),
.Y(n_4358)
);

OAI22xp5_ASAP7_75t_L g4359 ( 
.A1(n_4278),
.A2(n_4150),
.B1(n_4096),
.B2(n_4029),
.Y(n_4359)
);

INVx3_ASAP7_75t_L g4360 ( 
.A(n_4254),
.Y(n_4360)
);

AOI22xp33_ASAP7_75t_L g4361 ( 
.A1(n_4205),
.A2(n_4144),
.B1(n_4181),
.B2(n_4130),
.Y(n_4361)
);

INVx5_ASAP7_75t_L g4362 ( 
.A(n_4221),
.Y(n_4362)
);

AOI22xp33_ASAP7_75t_L g4363 ( 
.A1(n_4189),
.A2(n_4181),
.B1(n_4165),
.B2(n_4036),
.Y(n_4363)
);

CKINVDCx5p33_ASAP7_75t_R g4364 ( 
.A(n_4210),
.Y(n_4364)
);

NOR2x1p5_ASAP7_75t_L g4365 ( 
.A(n_4198),
.B(n_4059),
.Y(n_4365)
);

BUFx3_ASAP7_75t_L g4366 ( 
.A(n_4333),
.Y(n_4366)
);

OAI22xp5_ASAP7_75t_L g4367 ( 
.A1(n_4278),
.A2(n_4029),
.B1(n_4036),
.B2(n_4165),
.Y(n_4367)
);

BUFx6f_ASAP7_75t_L g4368 ( 
.A(n_4232),
.Y(n_4368)
);

INVx2_ASAP7_75t_L g4369 ( 
.A(n_4343),
.Y(n_4369)
);

NOR2xp33_ASAP7_75t_L g4370 ( 
.A(n_4236),
.B(n_4170),
.Y(n_4370)
);

AOI222xp33_ASAP7_75t_L g4371 ( 
.A1(n_4318),
.A2(n_4167),
.B1(n_4138),
.B2(n_4145),
.C1(n_4169),
.C2(n_4125),
.Y(n_4371)
);

AOI22xp5_ASAP7_75t_L g4372 ( 
.A1(n_4243),
.A2(n_4166),
.B1(n_4167),
.B2(n_4067),
.Y(n_4372)
);

AOI22xp33_ASAP7_75t_L g4373 ( 
.A1(n_4189),
.A2(n_4166),
.B1(n_4177),
.B2(n_4067),
.Y(n_4373)
);

AOI22xp33_ASAP7_75t_L g4374 ( 
.A1(n_4216),
.A2(n_4101),
.B1(n_4145),
.B2(n_4141),
.Y(n_4374)
);

AOI22xp33_ASAP7_75t_L g4375 ( 
.A1(n_4216),
.A2(n_4173),
.B1(n_4152),
.B2(n_4123),
.Y(n_4375)
);

OAI22xp5_ASAP7_75t_L g4376 ( 
.A1(n_4307),
.A2(n_341),
.B1(n_339),
.B2(n_340),
.Y(n_4376)
);

OAI22xp33_ASAP7_75t_L g4377 ( 
.A1(n_4308),
.A2(n_342),
.B1(n_339),
.B2(n_340),
.Y(n_4377)
);

NOR2xp33_ASAP7_75t_L g4378 ( 
.A(n_4225),
.B(n_342),
.Y(n_4378)
);

AOI22xp33_ASAP7_75t_L g4379 ( 
.A1(n_4184),
.A2(n_345),
.B1(n_343),
.B2(n_344),
.Y(n_4379)
);

AOI22xp5_ASAP7_75t_L g4380 ( 
.A1(n_4243),
.A2(n_346),
.B1(n_343),
.B2(n_345),
.Y(n_4380)
);

NAND2xp5_ASAP7_75t_L g4381 ( 
.A(n_4263),
.B(n_346),
.Y(n_4381)
);

AOI22xp33_ASAP7_75t_L g4382 ( 
.A1(n_4184),
.A2(n_349),
.B1(n_347),
.B2(n_348),
.Y(n_4382)
);

AOI22xp33_ASAP7_75t_L g4383 ( 
.A1(n_4194),
.A2(n_4342),
.B1(n_4223),
.B2(n_4329),
.Y(n_4383)
);

AOI22xp33_ASAP7_75t_L g4384 ( 
.A1(n_4194),
.A2(n_350),
.B1(n_347),
.B2(n_348),
.Y(n_4384)
);

AOI22xp33_ASAP7_75t_SL g4385 ( 
.A1(n_4345),
.A2(n_352),
.B1(n_350),
.B2(n_351),
.Y(n_4385)
);

OAI21xp33_ASAP7_75t_L g4386 ( 
.A1(n_4327),
.A2(n_351),
.B(n_352),
.Y(n_4386)
);

CKINVDCx16_ASAP7_75t_R g4387 ( 
.A(n_4311),
.Y(n_4387)
);

AOI22xp33_ASAP7_75t_L g4388 ( 
.A1(n_4342),
.A2(n_4223),
.B1(n_4206),
.B2(n_4274),
.Y(n_4388)
);

INVx2_ASAP7_75t_L g4389 ( 
.A(n_4343),
.Y(n_4389)
);

INVx2_ASAP7_75t_L g4390 ( 
.A(n_4343),
.Y(n_4390)
);

AOI22xp33_ASAP7_75t_SL g4391 ( 
.A1(n_4289),
.A2(n_355),
.B1(n_353),
.B2(n_354),
.Y(n_4391)
);

INVx1_ASAP7_75t_L g4392 ( 
.A(n_4195),
.Y(n_4392)
);

AOI22xp33_ASAP7_75t_L g4393 ( 
.A1(n_4206),
.A2(n_357),
.B1(n_353),
.B2(n_356),
.Y(n_4393)
);

AOI22xp33_ASAP7_75t_L g4394 ( 
.A1(n_4274),
.A2(n_361),
.B1(n_358),
.B2(n_359),
.Y(n_4394)
);

AOI22xp33_ASAP7_75t_SL g4395 ( 
.A1(n_4185),
.A2(n_361),
.B1(n_358),
.B2(n_359),
.Y(n_4395)
);

AOI221xp5_ASAP7_75t_SL g4396 ( 
.A1(n_4327),
.A2(n_365),
.B1(n_362),
.B2(n_364),
.C(n_366),
.Y(n_4396)
);

AOI22xp33_ASAP7_75t_SL g4397 ( 
.A1(n_4185),
.A2(n_368),
.B1(n_362),
.B2(n_367),
.Y(n_4397)
);

BUFx2_ASAP7_75t_L g4398 ( 
.A(n_4233),
.Y(n_4398)
);

AOI22xp33_ASAP7_75t_L g4399 ( 
.A1(n_4322),
.A2(n_369),
.B1(n_367),
.B2(n_368),
.Y(n_4399)
);

CKINVDCx5p33_ASAP7_75t_R g4400 ( 
.A(n_4333),
.Y(n_4400)
);

INVx3_ASAP7_75t_L g4401 ( 
.A(n_4254),
.Y(n_4401)
);

INVx1_ASAP7_75t_L g4402 ( 
.A(n_4248),
.Y(n_4402)
);

NAND2xp5_ASAP7_75t_L g4403 ( 
.A(n_4209),
.B(n_369),
.Y(n_4403)
);

AND2x4_ASAP7_75t_L g4404 ( 
.A(n_4229),
.B(n_4332),
.Y(n_4404)
);

AOI22xp5_ASAP7_75t_L g4405 ( 
.A1(n_4285),
.A2(n_4271),
.B1(n_4250),
.B2(n_4322),
.Y(n_4405)
);

CKINVDCx5p33_ASAP7_75t_R g4406 ( 
.A(n_4251),
.Y(n_4406)
);

INVx1_ASAP7_75t_L g4407 ( 
.A(n_4248),
.Y(n_4407)
);

OAI22xp5_ASAP7_75t_L g4408 ( 
.A1(n_4337),
.A2(n_4234),
.B1(n_4325),
.B2(n_4212),
.Y(n_4408)
);

AOI22xp33_ASAP7_75t_L g4409 ( 
.A1(n_4285),
.A2(n_372),
.B1(n_370),
.B2(n_371),
.Y(n_4409)
);

INVx3_ASAP7_75t_L g4410 ( 
.A(n_4249),
.Y(n_4410)
);

AOI22xp5_ASAP7_75t_SL g4411 ( 
.A1(n_4214),
.A2(n_373),
.B1(n_370),
.B2(n_372),
.Y(n_4411)
);

AOI22xp33_ASAP7_75t_L g4412 ( 
.A1(n_4267),
.A2(n_375),
.B1(n_373),
.B2(n_374),
.Y(n_4412)
);

INVx4_ASAP7_75t_SL g4413 ( 
.A(n_4280),
.Y(n_4413)
);

AND2x2_ASAP7_75t_L g4414 ( 
.A(n_4182),
.B(n_375),
.Y(n_4414)
);

NAND2xp5_ASAP7_75t_L g4415 ( 
.A(n_4209),
.B(n_376),
.Y(n_4415)
);

INVx4_ASAP7_75t_L g4416 ( 
.A(n_4320),
.Y(n_4416)
);

BUFx6f_ASAP7_75t_L g4417 ( 
.A(n_4304),
.Y(n_4417)
);

AND2x2_ASAP7_75t_L g4418 ( 
.A(n_4182),
.B(n_4235),
.Y(n_4418)
);

AOI22xp33_ASAP7_75t_SL g4419 ( 
.A1(n_4340),
.A2(n_378),
.B1(n_376),
.B2(n_377),
.Y(n_4419)
);

INVx1_ASAP7_75t_L g4420 ( 
.A(n_4245),
.Y(n_4420)
);

OAI22xp5_ASAP7_75t_L g4421 ( 
.A1(n_4234),
.A2(n_379),
.B1(n_377),
.B2(n_378),
.Y(n_4421)
);

NAND2xp5_ASAP7_75t_SL g4422 ( 
.A(n_4235),
.B(n_379),
.Y(n_4422)
);

INVx3_ASAP7_75t_L g4423 ( 
.A(n_4249),
.Y(n_4423)
);

OAI22xp5_ASAP7_75t_L g4424 ( 
.A1(n_4212),
.A2(n_4203),
.B1(n_4197),
.B2(n_4324),
.Y(n_4424)
);

BUFx3_ASAP7_75t_L g4425 ( 
.A(n_4331),
.Y(n_4425)
);

NAND2xp5_ASAP7_75t_L g4426 ( 
.A(n_4260),
.B(n_380),
.Y(n_4426)
);

INVx2_ASAP7_75t_L g4427 ( 
.A(n_4242),
.Y(n_4427)
);

AND2x6_ASAP7_75t_L g4428 ( 
.A(n_4294),
.B(n_380),
.Y(n_4428)
);

INVx1_ASAP7_75t_L g4429 ( 
.A(n_4247),
.Y(n_4429)
);

OAI22xp5_ASAP7_75t_L g4430 ( 
.A1(n_4203),
.A2(n_383),
.B1(n_381),
.B2(n_382),
.Y(n_4430)
);

OAI22xp5_ASAP7_75t_L g4431 ( 
.A1(n_4197),
.A2(n_384),
.B1(n_382),
.B2(n_383),
.Y(n_4431)
);

INVx1_ASAP7_75t_L g4432 ( 
.A(n_4253),
.Y(n_4432)
);

OAI22xp5_ASAP7_75t_L g4433 ( 
.A1(n_4324),
.A2(n_386),
.B1(n_384),
.B2(n_385),
.Y(n_4433)
);

INVx1_ASAP7_75t_L g4434 ( 
.A(n_4200),
.Y(n_4434)
);

BUFx4f_ASAP7_75t_SL g4435 ( 
.A(n_4273),
.Y(n_4435)
);

INVx1_ASAP7_75t_L g4436 ( 
.A(n_4204),
.Y(n_4436)
);

INVx1_ASAP7_75t_L g4437 ( 
.A(n_4215),
.Y(n_4437)
);

BUFx8_ASAP7_75t_SL g4438 ( 
.A(n_4297),
.Y(n_4438)
);

HB1xp67_ASAP7_75t_L g4439 ( 
.A(n_4279),
.Y(n_4439)
);

INVx2_ASAP7_75t_L g4440 ( 
.A(n_4334),
.Y(n_4440)
);

INVx1_ASAP7_75t_L g4441 ( 
.A(n_4218),
.Y(n_4441)
);

OAI22xp5_ASAP7_75t_L g4442 ( 
.A1(n_4214),
.A2(n_388),
.B1(n_386),
.B2(n_387),
.Y(n_4442)
);

AOI22xp33_ASAP7_75t_L g4443 ( 
.A1(n_4267),
.A2(n_389),
.B1(n_387),
.B2(n_388),
.Y(n_4443)
);

AOI22xp33_ASAP7_75t_L g4444 ( 
.A1(n_4344),
.A2(n_392),
.B1(n_390),
.B2(n_391),
.Y(n_4444)
);

AND2x2_ASAP7_75t_L g4445 ( 
.A(n_4282),
.B(n_390),
.Y(n_4445)
);

AOI22xp33_ASAP7_75t_SL g4446 ( 
.A1(n_4340),
.A2(n_395),
.B1(n_393),
.B2(n_394),
.Y(n_4446)
);

INVx1_ASAP7_75t_L g4447 ( 
.A(n_4220),
.Y(n_4447)
);

OAI222xp33_ASAP7_75t_L g4448 ( 
.A1(n_4208),
.A2(n_393),
.B1(n_394),
.B2(n_396),
.C1(n_397),
.C2(n_398),
.Y(n_4448)
);

NOR2x1_ASAP7_75t_L g4449 ( 
.A(n_4294),
.B(n_4244),
.Y(n_4449)
);

INVx3_ASAP7_75t_L g4450 ( 
.A(n_4282),
.Y(n_4450)
);

INVx8_ASAP7_75t_L g4451 ( 
.A(n_4335),
.Y(n_4451)
);

INVx1_ASAP7_75t_L g4452 ( 
.A(n_4224),
.Y(n_4452)
);

OAI22xp5_ASAP7_75t_L g4453 ( 
.A1(n_4238),
.A2(n_4244),
.B1(n_4240),
.B2(n_4269),
.Y(n_4453)
);

AOI21xp33_ASAP7_75t_SL g4454 ( 
.A1(n_4252),
.A2(n_398),
.B(n_400),
.Y(n_4454)
);

INVx1_ASAP7_75t_L g4455 ( 
.A(n_4230),
.Y(n_4455)
);

HB1xp67_ASAP7_75t_L g4456 ( 
.A(n_4314),
.Y(n_4456)
);

INVx1_ASAP7_75t_L g4457 ( 
.A(n_4231),
.Y(n_4457)
);

OAI21xp5_ASAP7_75t_SL g4458 ( 
.A1(n_4239),
.A2(n_400),
.B(n_401),
.Y(n_4458)
);

INVx1_ASAP7_75t_L g4459 ( 
.A(n_4237),
.Y(n_4459)
);

OAI21xp33_ASAP7_75t_L g4460 ( 
.A1(n_4191),
.A2(n_402),
.B(n_403),
.Y(n_4460)
);

INVxp67_ASAP7_75t_L g4461 ( 
.A(n_4238),
.Y(n_4461)
);

AOI22xp33_ASAP7_75t_L g4462 ( 
.A1(n_4320),
.A2(n_4250),
.B1(n_4299),
.B2(n_4211),
.Y(n_4462)
);

INVx1_ASAP7_75t_L g4463 ( 
.A(n_4270),
.Y(n_4463)
);

AND2x2_ASAP7_75t_L g4464 ( 
.A(n_4323),
.B(n_403),
.Y(n_4464)
);

OAI22xp5_ASAP7_75t_L g4465 ( 
.A1(n_4240),
.A2(n_407),
.B1(n_405),
.B2(n_406),
.Y(n_4465)
);

AOI22xp33_ASAP7_75t_SL g4466 ( 
.A1(n_4255),
.A2(n_408),
.B1(n_405),
.B2(n_406),
.Y(n_4466)
);

OAI22xp33_ASAP7_75t_L g4467 ( 
.A1(n_4269),
.A2(n_411),
.B1(n_409),
.B2(n_410),
.Y(n_4467)
);

OAI22xp5_ASAP7_75t_L g4468 ( 
.A1(n_4188),
.A2(n_411),
.B1(n_409),
.B2(n_410),
.Y(n_4468)
);

BUFx4f_ASAP7_75t_SL g4469 ( 
.A(n_4283),
.Y(n_4469)
);

AOI22xp33_ASAP7_75t_SL g4470 ( 
.A1(n_4258),
.A2(n_414),
.B1(n_412),
.B2(n_413),
.Y(n_4470)
);

AOI22xp33_ASAP7_75t_L g4471 ( 
.A1(n_4299),
.A2(n_415),
.B1(n_412),
.B2(n_414),
.Y(n_4471)
);

AOI22xp33_ASAP7_75t_L g4472 ( 
.A1(n_4293),
.A2(n_418),
.B1(n_416),
.B2(n_417),
.Y(n_4472)
);

AOI22xp33_ASAP7_75t_L g4473 ( 
.A1(n_4293),
.A2(n_419),
.B1(n_417),
.B2(n_418),
.Y(n_4473)
);

HB1xp67_ASAP7_75t_SL g4474 ( 
.A(n_4339),
.Y(n_4474)
);

NAND2xp5_ASAP7_75t_L g4475 ( 
.A(n_4260),
.B(n_419),
.Y(n_4475)
);

INVx1_ASAP7_75t_L g4476 ( 
.A(n_4217),
.Y(n_4476)
);

AOI22xp33_ASAP7_75t_L g4477 ( 
.A1(n_4300),
.A2(n_4291),
.B1(n_4276),
.B2(n_4309),
.Y(n_4477)
);

INVx5_ASAP7_75t_SL g4478 ( 
.A(n_4303),
.Y(n_4478)
);

AND2x2_ASAP7_75t_L g4479 ( 
.A(n_4323),
.B(n_420),
.Y(n_4479)
);

OAI22xp5_ASAP7_75t_L g4480 ( 
.A1(n_4239),
.A2(n_422),
.B1(n_420),
.B2(n_421),
.Y(n_4480)
);

OAI22xp33_ASAP7_75t_SL g4481 ( 
.A1(n_4207),
.A2(n_424),
.B1(n_421),
.B2(n_423),
.Y(n_4481)
);

HB1xp67_ASAP7_75t_L g4482 ( 
.A(n_4191),
.Y(n_4482)
);

INVx1_ASAP7_75t_L g4483 ( 
.A(n_4290),
.Y(n_4483)
);

AOI22xp33_ASAP7_75t_L g4484 ( 
.A1(n_4300),
.A2(n_425),
.B1(n_423),
.B2(n_424),
.Y(n_4484)
);

BUFx4f_ASAP7_75t_SL g4485 ( 
.A(n_4241),
.Y(n_4485)
);

AOI22xp33_ASAP7_75t_L g4486 ( 
.A1(n_4276),
.A2(n_427),
.B1(n_425),
.B2(n_426),
.Y(n_4486)
);

INVx1_ASAP7_75t_L g4487 ( 
.A(n_4298),
.Y(n_4487)
);

OAI22xp5_ASAP7_75t_L g4488 ( 
.A1(n_4291),
.A2(n_430),
.B1(n_428),
.B2(n_429),
.Y(n_4488)
);

AND2x2_ASAP7_75t_L g4489 ( 
.A(n_4187),
.B(n_430),
.Y(n_4489)
);

INVx2_ASAP7_75t_L g4490 ( 
.A(n_4309),
.Y(n_4490)
);

OAI21xp5_ASAP7_75t_SL g4491 ( 
.A1(n_4339),
.A2(n_432),
.B(n_433),
.Y(n_4491)
);

INVx1_ASAP7_75t_L g4492 ( 
.A(n_4305),
.Y(n_4492)
);

AOI22xp33_ASAP7_75t_SL g4493 ( 
.A1(n_4302),
.A2(n_436),
.B1(n_434),
.B2(n_435),
.Y(n_4493)
);

INVx2_ASAP7_75t_L g4494 ( 
.A(n_4259),
.Y(n_4494)
);

OAI22xp5_ASAP7_75t_L g4495 ( 
.A1(n_4188),
.A2(n_437),
.B1(n_434),
.B2(n_436),
.Y(n_4495)
);

OAI222xp33_ASAP7_75t_L g4496 ( 
.A1(n_4207),
.A2(n_437),
.B1(n_438),
.B2(n_439),
.C1(n_440),
.C2(n_441),
.Y(n_4496)
);

AND2x2_ASAP7_75t_L g4497 ( 
.A(n_4190),
.B(n_438),
.Y(n_4497)
);

AOI22xp33_ASAP7_75t_L g4498 ( 
.A1(n_4321),
.A2(n_443),
.B1(n_440),
.B2(n_442),
.Y(n_4498)
);

BUFx2_ASAP7_75t_L g4499 ( 
.A(n_4335),
.Y(n_4499)
);

BUFx4f_ASAP7_75t_SL g4500 ( 
.A(n_4316),
.Y(n_4500)
);

OAI21xp5_ASAP7_75t_SL g4501 ( 
.A1(n_4315),
.A2(n_442),
.B(n_443),
.Y(n_4501)
);

AOI22xp33_ASAP7_75t_L g4502 ( 
.A1(n_4321),
.A2(n_446),
.B1(n_444),
.B2(n_445),
.Y(n_4502)
);

AND2x2_ASAP7_75t_L g4503 ( 
.A(n_4328),
.B(n_4199),
.Y(n_4503)
);

OAI22xp5_ASAP7_75t_L g4504 ( 
.A1(n_4277),
.A2(n_448),
.B1(n_445),
.B2(n_447),
.Y(n_4504)
);

INVx1_ASAP7_75t_L g4505 ( 
.A(n_4356),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_4437),
.Y(n_4506)
);

OAI21xp5_ASAP7_75t_L g4507 ( 
.A1(n_4349),
.A2(n_4192),
.B(n_4183),
.Y(n_4507)
);

INVx2_ASAP7_75t_L g4508 ( 
.A(n_4413),
.Y(n_4508)
);

AND2x2_ASAP7_75t_L g4509 ( 
.A(n_4387),
.B(n_4196),
.Y(n_4509)
);

AOI21xp5_ASAP7_75t_L g4510 ( 
.A1(n_4388),
.A2(n_4193),
.B(n_4265),
.Y(n_4510)
);

AND2x2_ASAP7_75t_L g4511 ( 
.A(n_4418),
.B(n_4336),
.Y(n_4511)
);

INVx1_ASAP7_75t_L g4512 ( 
.A(n_4441),
.Y(n_4512)
);

OR2x2_ASAP7_75t_L g4513 ( 
.A(n_4402),
.B(n_4265),
.Y(n_4513)
);

INVx1_ASAP7_75t_L g4514 ( 
.A(n_4447),
.Y(n_4514)
);

OAI21xp5_ASAP7_75t_L g4515 ( 
.A1(n_4458),
.A2(n_4213),
.B(n_4341),
.Y(n_4515)
);

INVx2_ASAP7_75t_L g4516 ( 
.A(n_4413),
.Y(n_4516)
);

NOR2xp33_ASAP7_75t_SL g4517 ( 
.A(n_4364),
.B(n_4400),
.Y(n_4517)
);

HB1xp67_ASAP7_75t_L g4518 ( 
.A(n_4416),
.Y(n_4518)
);

INVx2_ASAP7_75t_L g4519 ( 
.A(n_4413),
.Y(n_4519)
);

NAND2xp5_ASAP7_75t_L g4520 ( 
.A(n_4361),
.B(n_4357),
.Y(n_4520)
);

AOI21x1_ASAP7_75t_L g4521 ( 
.A1(n_4398),
.A2(n_4330),
.B(n_4193),
.Y(n_4521)
);

OA21x2_ASAP7_75t_L g4522 ( 
.A1(n_4383),
.A2(n_4202),
.B(n_4310),
.Y(n_4522)
);

NOR2xp33_ASAP7_75t_L g4523 ( 
.A(n_4355),
.B(n_4262),
.Y(n_4523)
);

INVx1_ASAP7_75t_L g4524 ( 
.A(n_4452),
.Y(n_4524)
);

BUFx3_ASAP7_75t_L g4525 ( 
.A(n_4366),
.Y(n_4525)
);

INVx2_ASAP7_75t_L g4526 ( 
.A(n_4416),
.Y(n_4526)
);

AND2x2_ASAP7_75t_L g4527 ( 
.A(n_4360),
.B(n_4286),
.Y(n_4527)
);

AOI21xp5_ASAP7_75t_SL g4528 ( 
.A1(n_4442),
.A2(n_4303),
.B(n_4259),
.Y(n_4528)
);

AND2x2_ASAP7_75t_L g4529 ( 
.A(n_4360),
.B(n_4286),
.Y(n_4529)
);

NAND2xp5_ASAP7_75t_L g4530 ( 
.A(n_4481),
.B(n_4246),
.Y(n_4530)
);

HB1xp67_ASAP7_75t_L g4531 ( 
.A(n_4439),
.Y(n_4531)
);

AO21x2_ASAP7_75t_L g4532 ( 
.A1(n_4403),
.A2(n_4317),
.B(n_4264),
.Y(n_4532)
);

BUFx2_ASAP7_75t_L g4533 ( 
.A(n_4438),
.Y(n_4533)
);

NAND2xp5_ASAP7_75t_L g4534 ( 
.A(n_4407),
.B(n_4201),
.Y(n_4534)
);

INVx4_ASAP7_75t_L g4535 ( 
.A(n_4362),
.Y(n_4535)
);

INVx2_ASAP7_75t_L g4536 ( 
.A(n_4490),
.Y(n_4536)
);

INVx1_ASAP7_75t_L g4537 ( 
.A(n_4455),
.Y(n_4537)
);

INVx1_ASAP7_75t_L g4538 ( 
.A(n_4457),
.Y(n_4538)
);

INVx2_ASAP7_75t_L g4539 ( 
.A(n_4494),
.Y(n_4539)
);

INVx1_ASAP7_75t_L g4540 ( 
.A(n_4459),
.Y(n_4540)
);

AND2x2_ASAP7_75t_L g4541 ( 
.A(n_4499),
.B(n_4346),
.Y(n_4541)
);

OR2x2_ASAP7_75t_L g4542 ( 
.A(n_4476),
.B(n_4219),
.Y(n_4542)
);

AND2x2_ASAP7_75t_L g4543 ( 
.A(n_4368),
.B(n_4227),
.Y(n_4543)
);

INVx1_ASAP7_75t_L g4544 ( 
.A(n_4420),
.Y(n_4544)
);

INVx1_ASAP7_75t_L g4545 ( 
.A(n_4429),
.Y(n_4545)
);

BUFx2_ASAP7_75t_R g4546 ( 
.A(n_4351),
.Y(n_4546)
);

INVx2_ASAP7_75t_L g4547 ( 
.A(n_4417),
.Y(n_4547)
);

INVx3_ASAP7_75t_L g4548 ( 
.A(n_4355),
.Y(n_4548)
);

OR2x6_ASAP7_75t_L g4549 ( 
.A(n_4458),
.B(n_4303),
.Y(n_4549)
);

BUFx2_ASAP7_75t_L g4550 ( 
.A(n_4368),
.Y(n_4550)
);

INVx2_ASAP7_75t_L g4551 ( 
.A(n_4417),
.Y(n_4551)
);

HB1xp67_ASAP7_75t_L g4552 ( 
.A(n_4456),
.Y(n_4552)
);

INVx3_ASAP7_75t_L g4553 ( 
.A(n_4368),
.Y(n_4553)
);

HB1xp67_ASAP7_75t_L g4554 ( 
.A(n_4482),
.Y(n_4554)
);

BUFx3_ASAP7_75t_L g4555 ( 
.A(n_4362),
.Y(n_4555)
);

AND2x2_ASAP7_75t_L g4556 ( 
.A(n_4401),
.B(n_4227),
.Y(n_4556)
);

INVx3_ASAP7_75t_L g4557 ( 
.A(n_4401),
.Y(n_4557)
);

AND2x2_ASAP7_75t_L g4558 ( 
.A(n_4410),
.B(n_4423),
.Y(n_4558)
);

AND2x2_ASAP7_75t_L g4559 ( 
.A(n_4410),
.B(n_4227),
.Y(n_4559)
);

OAI21x1_ASAP7_75t_L g4560 ( 
.A1(n_4450),
.A2(n_4226),
.B(n_4257),
.Y(n_4560)
);

OA21x2_ASAP7_75t_L g4561 ( 
.A1(n_4462),
.A2(n_4186),
.B(n_4292),
.Y(n_4561)
);

OA21x2_ASAP7_75t_L g4562 ( 
.A1(n_4369),
.A2(n_4295),
.B(n_4301),
.Y(n_4562)
);

INVxp67_ASAP7_75t_SL g4563 ( 
.A(n_4474),
.Y(n_4563)
);

INVx1_ASAP7_75t_L g4564 ( 
.A(n_4483),
.Y(n_4564)
);

INVx1_ASAP7_75t_L g4565 ( 
.A(n_4487),
.Y(n_4565)
);

NAND2xp5_ASAP7_75t_L g4566 ( 
.A(n_4347),
.B(n_4353),
.Y(n_4566)
);

AOI22xp5_ASAP7_75t_L g4567 ( 
.A1(n_4372),
.A2(n_4266),
.B1(n_4284),
.B2(n_4272),
.Y(n_4567)
);

INVx3_ASAP7_75t_L g4568 ( 
.A(n_4362),
.Y(n_4568)
);

INVx3_ASAP7_75t_L g4569 ( 
.A(n_4362),
.Y(n_4569)
);

AND2x2_ASAP7_75t_L g4570 ( 
.A(n_4365),
.B(n_4284),
.Y(n_4570)
);

NOR2x1_ASAP7_75t_L g4571 ( 
.A(n_4415),
.B(n_4284),
.Y(n_4571)
);

NOR2xp33_ASAP7_75t_L g4572 ( 
.A(n_4485),
.B(n_4296),
.Y(n_4572)
);

NAND2xp5_ASAP7_75t_L g4573 ( 
.A(n_4354),
.B(n_4280),
.Y(n_4573)
);

AND2x2_ASAP7_75t_L g4574 ( 
.A(n_4425),
.B(n_4280),
.Y(n_4574)
);

AND2x4_ASAP7_75t_L g4575 ( 
.A(n_4350),
.B(n_4312),
.Y(n_4575)
);

NAND4xp25_ASAP7_75t_L g4576 ( 
.A(n_4363),
.B(n_4312),
.C(n_4288),
.D(n_4281),
.Y(n_4576)
);

AND2x2_ASAP7_75t_L g4577 ( 
.A(n_4423),
.B(n_4312),
.Y(n_4577)
);

INVx1_ASAP7_75t_L g4578 ( 
.A(n_4492),
.Y(n_4578)
);

AO31x2_ASAP7_75t_L g4579 ( 
.A1(n_4348),
.A2(n_4261),
.A3(n_4275),
.B(n_4222),
.Y(n_4579)
);

INVx3_ASAP7_75t_L g4580 ( 
.A(n_4417),
.Y(n_4580)
);

NOR2xp33_ASAP7_75t_L g4581 ( 
.A(n_4435),
.B(n_4306),
.Y(n_4581)
);

INVx2_ASAP7_75t_L g4582 ( 
.A(n_4427),
.Y(n_4582)
);

AND2x4_ASAP7_75t_L g4583 ( 
.A(n_4450),
.B(n_4222),
.Y(n_4583)
);

INVx1_ASAP7_75t_L g4584 ( 
.A(n_4463),
.Y(n_4584)
);

INVx2_ASAP7_75t_L g4585 ( 
.A(n_4449),
.Y(n_4585)
);

AND2x2_ASAP7_75t_L g4586 ( 
.A(n_4503),
.B(n_4313),
.Y(n_4586)
);

INVxp67_ASAP7_75t_L g4587 ( 
.A(n_4358),
.Y(n_4587)
);

NAND2xp5_ASAP7_75t_L g4588 ( 
.A(n_4379),
.B(n_4222),
.Y(n_4588)
);

INVx1_ASAP7_75t_L g4589 ( 
.A(n_4434),
.Y(n_4589)
);

NOR2x1_ASAP7_75t_L g4590 ( 
.A(n_4501),
.B(n_4408),
.Y(n_4590)
);

INVx2_ASAP7_75t_L g4591 ( 
.A(n_4440),
.Y(n_4591)
);

BUFx2_ASAP7_75t_L g4592 ( 
.A(n_4469),
.Y(n_4592)
);

INVx2_ASAP7_75t_SL g4593 ( 
.A(n_4451),
.Y(n_4593)
);

AND2x2_ASAP7_75t_L g4594 ( 
.A(n_4404),
.B(n_4326),
.Y(n_4594)
);

INVx1_ASAP7_75t_L g4595 ( 
.A(n_4432),
.Y(n_4595)
);

OA21x2_ASAP7_75t_L g4596 ( 
.A1(n_4389),
.A2(n_449),
.B(n_450),
.Y(n_4596)
);

AND2x2_ASAP7_75t_L g4597 ( 
.A(n_4404),
.B(n_450),
.Y(n_4597)
);

OA21x2_ASAP7_75t_L g4598 ( 
.A1(n_4390),
.A2(n_451),
.B(n_452),
.Y(n_4598)
);

INVx1_ASAP7_75t_L g4599 ( 
.A(n_4426),
.Y(n_4599)
);

INVx1_ASAP7_75t_L g4600 ( 
.A(n_4475),
.Y(n_4600)
);

BUFx3_ASAP7_75t_L g4601 ( 
.A(n_4428),
.Y(n_4601)
);

AND2x4_ASAP7_75t_L g4602 ( 
.A(n_4461),
.B(n_451),
.Y(n_4602)
);

INVx3_ASAP7_75t_L g4603 ( 
.A(n_4451),
.Y(n_4603)
);

AO21x2_ASAP7_75t_L g4604 ( 
.A1(n_4381),
.A2(n_452),
.B(n_454),
.Y(n_4604)
);

INVx2_ASAP7_75t_L g4605 ( 
.A(n_4464),
.Y(n_4605)
);

OR2x6_ASAP7_75t_L g4606 ( 
.A(n_4491),
.B(n_454),
.Y(n_4606)
);

HB1xp67_ASAP7_75t_L g4607 ( 
.A(n_4453),
.Y(n_4607)
);

OAI211xp5_ASAP7_75t_L g4608 ( 
.A1(n_4391),
.A2(n_457),
.B(n_455),
.C(n_456),
.Y(n_4608)
);

INVx2_ASAP7_75t_SL g4609 ( 
.A(n_4451),
.Y(n_4609)
);

INVx2_ASAP7_75t_L g4610 ( 
.A(n_4479),
.Y(n_4610)
);

INVx2_ASAP7_75t_L g4611 ( 
.A(n_4478),
.Y(n_4611)
);

INVx1_ASAP7_75t_L g4612 ( 
.A(n_4436),
.Y(n_4612)
);

INVx1_ASAP7_75t_L g4613 ( 
.A(n_4392),
.Y(n_4613)
);

AND2x4_ASAP7_75t_L g4614 ( 
.A(n_4489),
.B(n_457),
.Y(n_4614)
);

AO21x2_ASAP7_75t_L g4615 ( 
.A1(n_4405),
.A2(n_458),
.B(n_460),
.Y(n_4615)
);

OR2x6_ASAP7_75t_L g4616 ( 
.A(n_4491),
.B(n_458),
.Y(n_4616)
);

OA21x2_ASAP7_75t_L g4617 ( 
.A1(n_4373),
.A2(n_460),
.B(n_461),
.Y(n_4617)
);

INVx2_ASAP7_75t_L g4618 ( 
.A(n_4478),
.Y(n_4618)
);

INVx3_ASAP7_75t_L g4619 ( 
.A(n_4428),
.Y(n_4619)
);

INVx1_ASAP7_75t_L g4620 ( 
.A(n_4376),
.Y(n_4620)
);

BUFx6f_ASAP7_75t_L g4621 ( 
.A(n_4414),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_4367),
.Y(n_4622)
);

INVx1_ASAP7_75t_L g4623 ( 
.A(n_4445),
.Y(n_4623)
);

INVx2_ASAP7_75t_L g4624 ( 
.A(n_4478),
.Y(n_4624)
);

INVx1_ASAP7_75t_L g4625 ( 
.A(n_4359),
.Y(n_4625)
);

NAND2xp5_ASAP7_75t_L g4626 ( 
.A(n_4382),
.B(n_461),
.Y(n_4626)
);

OR2x2_ASAP7_75t_L g4627 ( 
.A(n_4424),
.B(n_462),
.Y(n_4627)
);

AND2x2_ASAP7_75t_L g4628 ( 
.A(n_4497),
.B(n_462),
.Y(n_4628)
);

AOI21x1_ASAP7_75t_L g4629 ( 
.A1(n_4352),
.A2(n_463),
.B(n_464),
.Y(n_4629)
);

OAI21xp5_ASAP7_75t_L g4630 ( 
.A1(n_4477),
.A2(n_464),
.B(n_465),
.Y(n_4630)
);

INVx1_ASAP7_75t_L g4631 ( 
.A(n_4377),
.Y(n_4631)
);

BUFx2_ASAP7_75t_L g4632 ( 
.A(n_4500),
.Y(n_4632)
);

INVx1_ASAP7_75t_L g4633 ( 
.A(n_4460),
.Y(n_4633)
);

INVx1_ASAP7_75t_L g4634 ( 
.A(n_4480),
.Y(n_4634)
);

AO21x1_ASAP7_75t_SL g4635 ( 
.A1(n_4374),
.A2(n_466),
.B(n_468),
.Y(n_4635)
);

AO21x2_ASAP7_75t_L g4636 ( 
.A1(n_4378),
.A2(n_4480),
.B(n_4467),
.Y(n_4636)
);

AND2x2_ASAP7_75t_L g4637 ( 
.A(n_4370),
.B(n_469),
.Y(n_4637)
);

INVx1_ASAP7_75t_L g4638 ( 
.A(n_4431),
.Y(n_4638)
);

AO21x2_ASAP7_75t_L g4639 ( 
.A1(n_4496),
.A2(n_4448),
.B(n_4430),
.Y(n_4639)
);

INVx1_ASAP7_75t_L g4640 ( 
.A(n_4488),
.Y(n_4640)
);

INVx2_ASAP7_75t_L g4641 ( 
.A(n_4428),
.Y(n_4641)
);

BUFx2_ASAP7_75t_SL g4642 ( 
.A(n_4428),
.Y(n_4642)
);

AOI21x1_ASAP7_75t_L g4643 ( 
.A1(n_4421),
.A2(n_469),
.B(n_470),
.Y(n_4643)
);

INVx2_ASAP7_75t_L g4644 ( 
.A(n_4422),
.Y(n_4644)
);

OA21x2_ASAP7_75t_L g4645 ( 
.A1(n_4396),
.A2(n_4384),
.B(n_4375),
.Y(n_4645)
);

INVx1_ASAP7_75t_L g4646 ( 
.A(n_4488),
.Y(n_4646)
);

BUFx4f_ASAP7_75t_SL g4647 ( 
.A(n_4419),
.Y(n_4647)
);

INVx2_ASAP7_75t_L g4648 ( 
.A(n_4406),
.Y(n_4648)
);

HB1xp67_ASAP7_75t_L g4649 ( 
.A(n_4518),
.Y(n_4649)
);

INVx1_ASAP7_75t_L g4650 ( 
.A(n_4531),
.Y(n_4650)
);

OR2x2_ASAP7_75t_L g4651 ( 
.A(n_4607),
.B(n_4501),
.Y(n_4651)
);

INVx3_ASAP7_75t_L g4652 ( 
.A(n_4525),
.Y(n_4652)
);

BUFx2_ASAP7_75t_L g4653 ( 
.A(n_4590),
.Y(n_4653)
);

NAND2xp5_ASAP7_75t_L g4654 ( 
.A(n_4602),
.B(n_4411),
.Y(n_4654)
);

AND2x2_ASAP7_75t_L g4655 ( 
.A(n_4563),
.B(n_4396),
.Y(n_4655)
);

OAI21xp5_ASAP7_75t_L g4656 ( 
.A1(n_4528),
.A2(n_4386),
.B(n_4395),
.Y(n_4656)
);

INVx1_ASAP7_75t_SL g4657 ( 
.A(n_4546),
.Y(n_4657)
);

AND2x2_ASAP7_75t_L g4658 ( 
.A(n_4509),
.B(n_4397),
.Y(n_4658)
);

AND2x4_ASAP7_75t_L g4659 ( 
.A(n_4553),
.B(n_4393),
.Y(n_4659)
);

BUFx2_ASAP7_75t_L g4660 ( 
.A(n_4592),
.Y(n_4660)
);

INVx2_ASAP7_75t_L g4661 ( 
.A(n_4606),
.Y(n_4661)
);

INVx1_ASAP7_75t_L g4662 ( 
.A(n_4536),
.Y(n_4662)
);

INVx1_ASAP7_75t_L g4663 ( 
.A(n_4536),
.Y(n_4663)
);

HB1xp67_ASAP7_75t_L g4664 ( 
.A(n_4518),
.Y(n_4664)
);

OAI21xp33_ASAP7_75t_L g4665 ( 
.A1(n_4520),
.A2(n_4385),
.B(n_4446),
.Y(n_4665)
);

NAND2xp5_ASAP7_75t_L g4666 ( 
.A(n_4602),
.B(n_4371),
.Y(n_4666)
);

AOI22xp33_ASAP7_75t_L g4667 ( 
.A1(n_4645),
.A2(n_4371),
.B1(n_4443),
.B2(n_4412),
.Y(n_4667)
);

AND2x2_ASAP7_75t_L g4668 ( 
.A(n_4509),
.B(n_4454),
.Y(n_4668)
);

AND2x2_ASAP7_75t_L g4669 ( 
.A(n_4603),
.B(n_4468),
.Y(n_4669)
);

AND2x2_ASAP7_75t_L g4670 ( 
.A(n_4603),
.B(n_4495),
.Y(n_4670)
);

OAI22xp5_ASAP7_75t_SL g4671 ( 
.A1(n_4647),
.A2(n_4493),
.B1(n_4470),
.B2(n_4466),
.Y(n_4671)
);

BUFx2_ASAP7_75t_L g4672 ( 
.A(n_4533),
.Y(n_4672)
);

NAND2xp5_ASAP7_75t_L g4673 ( 
.A(n_4602),
.B(n_4498),
.Y(n_4673)
);

INVx1_ASAP7_75t_L g4674 ( 
.A(n_4539),
.Y(n_4674)
);

INVxp67_ASAP7_75t_SL g4675 ( 
.A(n_4607),
.Y(n_4675)
);

INVx1_ASAP7_75t_L g4676 ( 
.A(n_4531),
.Y(n_4676)
);

AND2x2_ASAP7_75t_L g4677 ( 
.A(n_4603),
.B(n_4550),
.Y(n_4677)
);

OR2x2_ASAP7_75t_L g4678 ( 
.A(n_4513),
.B(n_4465),
.Y(n_4678)
);

AND2x2_ASAP7_75t_L g4679 ( 
.A(n_4553),
.B(n_4502),
.Y(n_4679)
);

INVx1_ASAP7_75t_L g4680 ( 
.A(n_4552),
.Y(n_4680)
);

AND2x2_ASAP7_75t_L g4681 ( 
.A(n_4553),
.B(n_4444),
.Y(n_4681)
);

BUFx2_ASAP7_75t_L g4682 ( 
.A(n_4632),
.Y(n_4682)
);

INVxp67_ASAP7_75t_L g4683 ( 
.A(n_4635),
.Y(n_4683)
);

INVx1_ASAP7_75t_L g4684 ( 
.A(n_4552),
.Y(n_4684)
);

INVx1_ASAP7_75t_L g4685 ( 
.A(n_4539),
.Y(n_4685)
);

BUFx2_ASAP7_75t_L g4686 ( 
.A(n_4525),
.Y(n_4686)
);

INVx2_ASAP7_75t_L g4687 ( 
.A(n_4606),
.Y(n_4687)
);

NAND2xp5_ASAP7_75t_L g4688 ( 
.A(n_4639),
.B(n_4504),
.Y(n_4688)
);

INVx1_ASAP7_75t_L g4689 ( 
.A(n_4554),
.Y(n_4689)
);

HB1xp67_ASAP7_75t_L g4690 ( 
.A(n_4526),
.Y(n_4690)
);

INVx2_ASAP7_75t_L g4691 ( 
.A(n_4606),
.Y(n_4691)
);

INVx1_ASAP7_75t_L g4692 ( 
.A(n_4554),
.Y(n_4692)
);

INVxp67_ASAP7_75t_L g4693 ( 
.A(n_4517),
.Y(n_4693)
);

AOI21xp5_ASAP7_75t_SL g4694 ( 
.A1(n_4616),
.A2(n_4433),
.B(n_4380),
.Y(n_4694)
);

AND2x2_ASAP7_75t_L g4695 ( 
.A(n_4558),
.B(n_4471),
.Y(n_4695)
);

AND2x2_ASAP7_75t_L g4696 ( 
.A(n_4558),
.B(n_4394),
.Y(n_4696)
);

BUFx3_ASAP7_75t_L g4697 ( 
.A(n_4555),
.Y(n_4697)
);

AND2x2_ASAP7_75t_L g4698 ( 
.A(n_4570),
.B(n_4399),
.Y(n_4698)
);

BUFx3_ASAP7_75t_L g4699 ( 
.A(n_4555),
.Y(n_4699)
);

BUFx2_ASAP7_75t_L g4700 ( 
.A(n_4568),
.Y(n_4700)
);

INVx2_ASAP7_75t_L g4701 ( 
.A(n_4616),
.Y(n_4701)
);

NAND2xp5_ASAP7_75t_L g4702 ( 
.A(n_4639),
.B(n_4472),
.Y(n_4702)
);

INVx2_ASAP7_75t_L g4703 ( 
.A(n_4616),
.Y(n_4703)
);

HB1xp67_ASAP7_75t_L g4704 ( 
.A(n_4526),
.Y(n_4704)
);

INVx2_ASAP7_75t_L g4705 ( 
.A(n_4596),
.Y(n_4705)
);

INVx2_ASAP7_75t_L g4706 ( 
.A(n_4596),
.Y(n_4706)
);

AND2x2_ASAP7_75t_L g4707 ( 
.A(n_4586),
.B(n_4486),
.Y(n_4707)
);

HB1xp67_ASAP7_75t_L g4708 ( 
.A(n_4532),
.Y(n_4708)
);

AND2x2_ASAP7_75t_L g4709 ( 
.A(n_4593),
.B(n_4473),
.Y(n_4709)
);

INVx1_ASAP7_75t_L g4710 ( 
.A(n_4506),
.Y(n_4710)
);

OR2x2_ASAP7_75t_L g4711 ( 
.A(n_4566),
.B(n_4484),
.Y(n_4711)
);

AND2x2_ASAP7_75t_L g4712 ( 
.A(n_4593),
.B(n_4409),
.Y(n_4712)
);

INVx1_ASAP7_75t_L g4713 ( 
.A(n_4512),
.Y(n_4713)
);

INVx1_ASAP7_75t_L g4714 ( 
.A(n_4514),
.Y(n_4714)
);

INVx1_ASAP7_75t_L g4715 ( 
.A(n_4524),
.Y(n_4715)
);

AO31x2_ASAP7_75t_L g4716 ( 
.A1(n_4508),
.A2(n_691),
.A3(n_473),
.B(n_470),
.Y(n_4716)
);

NAND2xp5_ASAP7_75t_L g4717 ( 
.A(n_4645),
.B(n_472),
.Y(n_4717)
);

OR2x2_ASAP7_75t_L g4718 ( 
.A(n_4505),
.B(n_474),
.Y(n_4718)
);

AND2x2_ASAP7_75t_L g4719 ( 
.A(n_4609),
.B(n_691),
.Y(n_4719)
);

INVx5_ASAP7_75t_L g4720 ( 
.A(n_4535),
.Y(n_4720)
);

INVx1_ASAP7_75t_L g4721 ( 
.A(n_4537),
.Y(n_4721)
);

AND2x2_ASAP7_75t_L g4722 ( 
.A(n_4609),
.B(n_476),
.Y(n_4722)
);

AND2x2_ASAP7_75t_L g4723 ( 
.A(n_4557),
.B(n_690),
.Y(n_4723)
);

AND2x2_ASAP7_75t_L g4724 ( 
.A(n_4557),
.B(n_690),
.Y(n_4724)
);

AND2x2_ASAP7_75t_L g4725 ( 
.A(n_4557),
.B(n_477),
.Y(n_4725)
);

BUFx4f_ASAP7_75t_SL g4726 ( 
.A(n_4535),
.Y(n_4726)
);

INVx2_ASAP7_75t_L g4727 ( 
.A(n_4596),
.Y(n_4727)
);

HB1xp67_ASAP7_75t_L g4728 ( 
.A(n_4532),
.Y(n_4728)
);

INVx1_ASAP7_75t_L g4729 ( 
.A(n_4538),
.Y(n_4729)
);

INVx2_ASAP7_75t_L g4730 ( 
.A(n_4598),
.Y(n_4730)
);

INVx2_ASAP7_75t_L g4731 ( 
.A(n_4598),
.Y(n_4731)
);

NOR2xp33_ASAP7_75t_L g4732 ( 
.A(n_4535),
.B(n_478),
.Y(n_4732)
);

INVx1_ASAP7_75t_L g4733 ( 
.A(n_4540),
.Y(n_4733)
);

AND2x2_ASAP7_75t_L g4734 ( 
.A(n_4523),
.B(n_689),
.Y(n_4734)
);

BUFx2_ASAP7_75t_L g4735 ( 
.A(n_4568),
.Y(n_4735)
);

INVx1_ASAP7_75t_L g4736 ( 
.A(n_4544),
.Y(n_4736)
);

AOI22xp33_ASAP7_75t_L g4737 ( 
.A1(n_4645),
.A2(n_480),
.B1(n_478),
.B2(n_479),
.Y(n_4737)
);

INVx1_ASAP7_75t_L g4738 ( 
.A(n_4545),
.Y(n_4738)
);

HB1xp67_ASAP7_75t_L g4739 ( 
.A(n_4541),
.Y(n_4739)
);

INVx1_ASAP7_75t_SL g4740 ( 
.A(n_4647),
.Y(n_4740)
);

INVx2_ASAP7_75t_L g4741 ( 
.A(n_4598),
.Y(n_4741)
);

INVxp67_ASAP7_75t_L g4742 ( 
.A(n_4642),
.Y(n_4742)
);

INVx2_ASAP7_75t_L g4743 ( 
.A(n_4549),
.Y(n_4743)
);

BUFx4f_ASAP7_75t_SL g4744 ( 
.A(n_4648),
.Y(n_4744)
);

OR2x2_ASAP7_75t_L g4745 ( 
.A(n_4640),
.B(n_479),
.Y(n_4745)
);

INVx2_ASAP7_75t_L g4746 ( 
.A(n_4549),
.Y(n_4746)
);

NAND2xp5_ASAP7_75t_L g4747 ( 
.A(n_4636),
.B(n_480),
.Y(n_4747)
);

HB1xp67_ASAP7_75t_L g4748 ( 
.A(n_4562),
.Y(n_4748)
);

INVx1_ASAP7_75t_L g4749 ( 
.A(n_4564),
.Y(n_4749)
);

INVx3_ASAP7_75t_L g4750 ( 
.A(n_4621),
.Y(n_4750)
);

INVx2_ASAP7_75t_L g4751 ( 
.A(n_4549),
.Y(n_4751)
);

INVx3_ASAP7_75t_L g4752 ( 
.A(n_4621),
.Y(n_4752)
);

INVx2_ASAP7_75t_L g4753 ( 
.A(n_4615),
.Y(n_4753)
);

INVx1_ASAP7_75t_L g4754 ( 
.A(n_4565),
.Y(n_4754)
);

AND2x2_ASAP7_75t_L g4755 ( 
.A(n_4523),
.B(n_4511),
.Y(n_4755)
);

BUFx3_ASAP7_75t_L g4756 ( 
.A(n_4568),
.Y(n_4756)
);

OR2x2_ASAP7_75t_L g4757 ( 
.A(n_4646),
.B(n_481),
.Y(n_4757)
);

INVx1_ASAP7_75t_L g4758 ( 
.A(n_4578),
.Y(n_4758)
);

NOR2xp33_ASAP7_75t_L g4759 ( 
.A(n_4569),
.B(n_481),
.Y(n_4759)
);

INVx2_ASAP7_75t_L g4760 ( 
.A(n_4615),
.Y(n_4760)
);

HB1xp67_ASAP7_75t_L g4761 ( 
.A(n_4562),
.Y(n_4761)
);

NOR2x1_ASAP7_75t_R g4762 ( 
.A(n_4653),
.B(n_4569),
.Y(n_4762)
);

INVx2_ASAP7_75t_L g4763 ( 
.A(n_4653),
.Y(n_4763)
);

INVx3_ASAP7_75t_L g4764 ( 
.A(n_4651),
.Y(n_4764)
);

AND2x2_ASAP7_75t_L g4765 ( 
.A(n_4686),
.B(n_4569),
.Y(n_4765)
);

INVx1_ASAP7_75t_L g4766 ( 
.A(n_4747),
.Y(n_4766)
);

BUFx6f_ASAP7_75t_L g4767 ( 
.A(n_4717),
.Y(n_4767)
);

INVx2_ASAP7_75t_L g4768 ( 
.A(n_4753),
.Y(n_4768)
);

AND2x2_ASAP7_75t_L g4769 ( 
.A(n_4686),
.B(n_4548),
.Y(n_4769)
);

AND2x4_ASAP7_75t_L g4770 ( 
.A(n_4652),
.B(n_4543),
.Y(n_4770)
);

INVx2_ASAP7_75t_L g4771 ( 
.A(n_4753),
.Y(n_4771)
);

NOR2xp33_ASAP7_75t_L g4772 ( 
.A(n_4657),
.B(n_4652),
.Y(n_4772)
);

AND2x4_ASAP7_75t_L g4773 ( 
.A(n_4652),
.B(n_4548),
.Y(n_4773)
);

NAND2xp5_ASAP7_75t_L g4774 ( 
.A(n_4675),
.B(n_4636),
.Y(n_4774)
);

HB1xp67_ASAP7_75t_L g4775 ( 
.A(n_4660),
.Y(n_4775)
);

INVxp67_ASAP7_75t_L g4776 ( 
.A(n_4672),
.Y(n_4776)
);

HB1xp67_ASAP7_75t_L g4777 ( 
.A(n_4660),
.Y(n_4777)
);

BUFx2_ASAP7_75t_L g4778 ( 
.A(n_4651),
.Y(n_4778)
);

AND2x2_ASAP7_75t_L g4779 ( 
.A(n_4672),
.B(n_4682),
.Y(n_4779)
);

AND2x2_ASAP7_75t_L g4780 ( 
.A(n_4682),
.B(n_4548),
.Y(n_4780)
);

AND2x2_ASAP7_75t_L g4781 ( 
.A(n_4755),
.B(n_4648),
.Y(n_4781)
);

INVx3_ASAP7_75t_L g4782 ( 
.A(n_4659),
.Y(n_4782)
);

AND2x2_ASAP7_75t_L g4783 ( 
.A(n_4755),
.B(n_4587),
.Y(n_4783)
);

INVx1_ASAP7_75t_L g4784 ( 
.A(n_4708),
.Y(n_4784)
);

HB1xp67_ASAP7_75t_L g4785 ( 
.A(n_4739),
.Y(n_4785)
);

AND2x2_ASAP7_75t_L g4786 ( 
.A(n_4668),
.B(n_4577),
.Y(n_4786)
);

BUFx2_ASAP7_75t_L g4787 ( 
.A(n_4728),
.Y(n_4787)
);

INVx1_ASAP7_75t_L g4788 ( 
.A(n_4761),
.Y(n_4788)
);

OR2x2_ASAP7_75t_L g4789 ( 
.A(n_4666),
.B(n_4534),
.Y(n_4789)
);

BUFx3_ASAP7_75t_L g4790 ( 
.A(n_4734),
.Y(n_4790)
);

AO21x2_ASAP7_75t_L g4791 ( 
.A1(n_4688),
.A2(n_4516),
.B(n_4508),
.Y(n_4791)
);

OR2x2_ASAP7_75t_L g4792 ( 
.A(n_4650),
.B(n_4589),
.Y(n_4792)
);

AND2x2_ASAP7_75t_L g4793 ( 
.A(n_4668),
.B(n_4581),
.Y(n_4793)
);

INVx2_ASAP7_75t_L g4794 ( 
.A(n_4760),
.Y(n_4794)
);

NAND2xp5_ASAP7_75t_L g4795 ( 
.A(n_4723),
.B(n_4605),
.Y(n_4795)
);

AND2x2_ASAP7_75t_L g4796 ( 
.A(n_4693),
.B(n_4581),
.Y(n_4796)
);

NAND2xp5_ASAP7_75t_L g4797 ( 
.A(n_4737),
.B(n_4634),
.Y(n_4797)
);

HB1xp67_ASAP7_75t_L g4798 ( 
.A(n_4649),
.Y(n_4798)
);

AO21x2_ASAP7_75t_L g4799 ( 
.A1(n_4702),
.A2(n_4519),
.B(n_4516),
.Y(n_4799)
);

INVx1_ASAP7_75t_L g4800 ( 
.A(n_4748),
.Y(n_4800)
);

OR2x2_ASAP7_75t_L g4801 ( 
.A(n_4650),
.B(n_4595),
.Y(n_4801)
);

INVx1_ASAP7_75t_L g4802 ( 
.A(n_4664),
.Y(n_4802)
);

NAND2xp5_ASAP7_75t_L g4803 ( 
.A(n_4723),
.B(n_4605),
.Y(n_4803)
);

INVx2_ASAP7_75t_L g4804 ( 
.A(n_4760),
.Y(n_4804)
);

NAND2xp5_ASAP7_75t_L g4805 ( 
.A(n_4724),
.B(n_4610),
.Y(n_4805)
);

INVx2_ASAP7_75t_L g4806 ( 
.A(n_4705),
.Y(n_4806)
);

NAND2xp5_ASAP7_75t_L g4807 ( 
.A(n_4724),
.B(n_4610),
.Y(n_4807)
);

AND2x2_ASAP7_75t_L g4808 ( 
.A(n_4750),
.B(n_4594),
.Y(n_4808)
);

NAND2xp5_ASAP7_75t_L g4809 ( 
.A(n_4725),
.B(n_4510),
.Y(n_4809)
);

BUFx3_ASAP7_75t_L g4810 ( 
.A(n_4734),
.Y(n_4810)
);

INVx2_ASAP7_75t_L g4811 ( 
.A(n_4705),
.Y(n_4811)
);

AOI22xp33_ASAP7_75t_L g4812 ( 
.A1(n_4667),
.A2(n_4617),
.B1(n_4625),
.B2(n_4622),
.Y(n_4812)
);

OR2x2_ASAP7_75t_L g4813 ( 
.A(n_4676),
.B(n_4612),
.Y(n_4813)
);

INVx3_ASAP7_75t_L g4814 ( 
.A(n_4659),
.Y(n_4814)
);

AND2x2_ASAP7_75t_L g4815 ( 
.A(n_4750),
.B(n_4511),
.Y(n_4815)
);

INVx4_ASAP7_75t_L g4816 ( 
.A(n_4720),
.Y(n_4816)
);

INVx2_ASAP7_75t_L g4817 ( 
.A(n_4706),
.Y(n_4817)
);

INVx1_ASAP7_75t_L g4818 ( 
.A(n_4676),
.Y(n_4818)
);

INVx1_ASAP7_75t_L g4819 ( 
.A(n_4680),
.Y(n_4819)
);

AND2x4_ASAP7_75t_L g4820 ( 
.A(n_4750),
.B(n_4611),
.Y(n_4820)
);

INVx2_ASAP7_75t_L g4821 ( 
.A(n_4706),
.Y(n_4821)
);

HB1xp67_ASAP7_75t_L g4822 ( 
.A(n_4740),
.Y(n_4822)
);

NAND2xp5_ASAP7_75t_L g4823 ( 
.A(n_4725),
.B(n_4638),
.Y(n_4823)
);

INVx1_ASAP7_75t_L g4824 ( 
.A(n_4680),
.Y(n_4824)
);

INVx2_ASAP7_75t_L g4825 ( 
.A(n_4727),
.Y(n_4825)
);

BUFx2_ASAP7_75t_L g4826 ( 
.A(n_4752),
.Y(n_4826)
);

INVx2_ASAP7_75t_L g4827 ( 
.A(n_4727),
.Y(n_4827)
);

OR2x2_ASAP7_75t_L g4828 ( 
.A(n_4684),
.B(n_4584),
.Y(n_4828)
);

OR2x2_ASAP7_75t_L g4829 ( 
.A(n_4684),
.B(n_4613),
.Y(n_4829)
);

NAND2xp5_ASAP7_75t_L g4830 ( 
.A(n_4655),
.B(n_4665),
.Y(n_4830)
);

INVx1_ASAP7_75t_L g4831 ( 
.A(n_4689),
.Y(n_4831)
);

INVx1_ASAP7_75t_L g4832 ( 
.A(n_4689),
.Y(n_4832)
);

INVx2_ASAP7_75t_L g4833 ( 
.A(n_4730),
.Y(n_4833)
);

HB1xp67_ASAP7_75t_L g4834 ( 
.A(n_4690),
.Y(n_4834)
);

INVx2_ASAP7_75t_L g4835 ( 
.A(n_4782),
.Y(n_4835)
);

NAND2xp5_ASAP7_75t_L g4836 ( 
.A(n_4790),
.B(n_4655),
.Y(n_4836)
);

AND2x2_ASAP7_75t_L g4837 ( 
.A(n_4779),
.B(n_4677),
.Y(n_4837)
);

AND2x2_ASAP7_75t_L g4838 ( 
.A(n_4779),
.B(n_4677),
.Y(n_4838)
);

NAND2xp5_ASAP7_75t_L g4839 ( 
.A(n_4790),
.B(n_4658),
.Y(n_4839)
);

INVxp67_ASAP7_75t_SL g4840 ( 
.A(n_4774),
.Y(n_4840)
);

AND2x2_ASAP7_75t_L g4841 ( 
.A(n_4822),
.B(n_4752),
.Y(n_4841)
);

AOI21xp5_ASAP7_75t_SL g4842 ( 
.A1(n_4762),
.A2(n_4732),
.B(n_4656),
.Y(n_4842)
);

INVx1_ASAP7_75t_L g4843 ( 
.A(n_4775),
.Y(n_4843)
);

INVxp67_ASAP7_75t_SL g4844 ( 
.A(n_4790),
.Y(n_4844)
);

INVx1_ASAP7_75t_L g4845 ( 
.A(n_4777),
.Y(n_4845)
);

OAI221xp5_ASAP7_75t_L g4846 ( 
.A1(n_4812),
.A2(n_4507),
.B1(n_4528),
.B2(n_4576),
.C(n_4515),
.Y(n_4846)
);

HB1xp67_ASAP7_75t_L g4847 ( 
.A(n_4810),
.Y(n_4847)
);

AND2x2_ASAP7_75t_L g4848 ( 
.A(n_4778),
.B(n_4752),
.Y(n_4848)
);

INVx1_ASAP7_75t_L g4849 ( 
.A(n_4782),
.Y(n_4849)
);

NAND2xp5_ASAP7_75t_L g4850 ( 
.A(n_4810),
.B(n_4658),
.Y(n_4850)
);

AOI221xp5_ASAP7_75t_L g4851 ( 
.A1(n_4778),
.A2(n_4707),
.B1(n_4694),
.B2(n_4556),
.C(n_4600),
.Y(n_4851)
);

INVx2_ASAP7_75t_L g4852 ( 
.A(n_4782),
.Y(n_4852)
);

AND2x2_ASAP7_75t_L g4853 ( 
.A(n_4783),
.B(n_4669),
.Y(n_4853)
);

AND2x2_ASAP7_75t_L g4854 ( 
.A(n_4783),
.B(n_4669),
.Y(n_4854)
);

AND2x2_ASAP7_75t_L g4855 ( 
.A(n_4781),
.B(n_4670),
.Y(n_4855)
);

INVx2_ASAP7_75t_L g4856 ( 
.A(n_4782),
.Y(n_4856)
);

INVx1_ASAP7_75t_L g4857 ( 
.A(n_4814),
.Y(n_4857)
);

AND2x2_ASAP7_75t_L g4858 ( 
.A(n_4781),
.B(n_4670),
.Y(n_4858)
);

INVx1_ASAP7_75t_L g4859 ( 
.A(n_4814),
.Y(n_4859)
);

INVx2_ASAP7_75t_L g4860 ( 
.A(n_4814),
.Y(n_4860)
);

NAND4xp25_ASAP7_75t_L g4861 ( 
.A(n_4772),
.B(n_4697),
.C(n_4699),
.D(n_4742),
.Y(n_4861)
);

OR2x2_ASAP7_75t_L g4862 ( 
.A(n_4764),
.B(n_4692),
.Y(n_4862)
);

NAND2x1_ASAP7_75t_SL g4863 ( 
.A(n_4770),
.B(n_4704),
.Y(n_4863)
);

AND2x2_ASAP7_75t_L g4864 ( 
.A(n_4780),
.B(n_4695),
.Y(n_4864)
);

AND2x4_ASAP7_75t_L g4865 ( 
.A(n_4770),
.B(n_4697),
.Y(n_4865)
);

INVx1_ASAP7_75t_L g4866 ( 
.A(n_4814),
.Y(n_4866)
);

NAND2xp5_ASAP7_75t_L g4867 ( 
.A(n_4810),
.B(n_4696),
.Y(n_4867)
);

NAND2xp5_ASAP7_75t_L g4868 ( 
.A(n_4776),
.B(n_4696),
.Y(n_4868)
);

NAND2xp5_ASAP7_75t_L g4869 ( 
.A(n_4780),
.B(n_4745),
.Y(n_4869)
);

AND2x4_ASAP7_75t_L g4870 ( 
.A(n_4770),
.B(n_4699),
.Y(n_4870)
);

AND2x2_ASAP7_75t_L g4871 ( 
.A(n_4786),
.B(n_4695),
.Y(n_4871)
);

INVx1_ASAP7_75t_SL g4872 ( 
.A(n_4786),
.Y(n_4872)
);

NAND3xp33_ASAP7_75t_L g4873 ( 
.A(n_4830),
.B(n_4764),
.C(n_4767),
.Y(n_4873)
);

NAND2xp5_ASAP7_75t_SL g4874 ( 
.A(n_4770),
.B(n_4621),
.Y(n_4874)
);

AND2x2_ASAP7_75t_L g4875 ( 
.A(n_4764),
.B(n_4712),
.Y(n_4875)
);

NAND2xp5_ASAP7_75t_SL g4876 ( 
.A(n_4769),
.B(n_4621),
.Y(n_4876)
);

AND2x2_ASAP7_75t_L g4877 ( 
.A(n_4764),
.B(n_4712),
.Y(n_4877)
);

AND2x2_ASAP7_75t_L g4878 ( 
.A(n_4815),
.B(n_4709),
.Y(n_4878)
);

INVx1_ASAP7_75t_L g4879 ( 
.A(n_4785),
.Y(n_4879)
);

NAND2xp5_ASAP7_75t_L g4880 ( 
.A(n_4769),
.B(n_4745),
.Y(n_4880)
);

INVx1_ASAP7_75t_L g4881 ( 
.A(n_4834),
.Y(n_4881)
);

INVx2_ASAP7_75t_SL g4882 ( 
.A(n_4765),
.Y(n_4882)
);

INVx1_ASAP7_75t_L g4883 ( 
.A(n_4787),
.Y(n_4883)
);

INVx1_ASAP7_75t_SL g4884 ( 
.A(n_4793),
.Y(n_4884)
);

INVx1_ASAP7_75t_L g4885 ( 
.A(n_4787),
.Y(n_4885)
);

INVx1_ASAP7_75t_L g4886 ( 
.A(n_4806),
.Y(n_4886)
);

OR2x2_ASAP7_75t_L g4887 ( 
.A(n_4763),
.B(n_4692),
.Y(n_4887)
);

INVx2_ASAP7_75t_L g4888 ( 
.A(n_4768),
.Y(n_4888)
);

INVx2_ASAP7_75t_L g4889 ( 
.A(n_4768),
.Y(n_4889)
);

AND2x2_ASAP7_75t_L g4890 ( 
.A(n_4815),
.B(n_4709),
.Y(n_4890)
);

NAND2xp5_ASAP7_75t_L g4891 ( 
.A(n_4763),
.B(n_4757),
.Y(n_4891)
);

AND2x2_ASAP7_75t_L g4892 ( 
.A(n_4765),
.B(n_4756),
.Y(n_4892)
);

AND2x2_ASAP7_75t_L g4893 ( 
.A(n_4808),
.B(n_4756),
.Y(n_4893)
);

OR2x2_ASAP7_75t_L g4894 ( 
.A(n_4763),
.B(n_4711),
.Y(n_4894)
);

BUFx2_ASAP7_75t_L g4895 ( 
.A(n_4863),
.Y(n_4895)
);

AND2x4_ASAP7_75t_L g4896 ( 
.A(n_4835),
.B(n_4773),
.Y(n_4896)
);

INVx1_ASAP7_75t_L g4897 ( 
.A(n_4847),
.Y(n_4897)
);

NOR2xp67_ASAP7_75t_L g4898 ( 
.A(n_4882),
.B(n_4683),
.Y(n_4898)
);

INVx2_ASAP7_75t_SL g4899 ( 
.A(n_4863),
.Y(n_4899)
);

OR2x2_ASAP7_75t_L g4900 ( 
.A(n_4894),
.B(n_4789),
.Y(n_4900)
);

NAND2xp5_ASAP7_75t_L g4901 ( 
.A(n_4855),
.B(n_4793),
.Y(n_4901)
);

INVx1_ASAP7_75t_L g4902 ( 
.A(n_4844),
.Y(n_4902)
);

INVx2_ASAP7_75t_L g4903 ( 
.A(n_4888),
.Y(n_4903)
);

INVx1_ASAP7_75t_L g4904 ( 
.A(n_4835),
.Y(n_4904)
);

INVx1_ASAP7_75t_L g4905 ( 
.A(n_4852),
.Y(n_4905)
);

AND2x2_ASAP7_75t_L g4906 ( 
.A(n_4855),
.B(n_4808),
.Y(n_4906)
);

INVx2_ASAP7_75t_L g4907 ( 
.A(n_4888),
.Y(n_4907)
);

AND2x2_ASAP7_75t_L g4908 ( 
.A(n_4858),
.B(n_4773),
.Y(n_4908)
);

AND2x4_ASAP7_75t_SL g4909 ( 
.A(n_4865),
.B(n_4773),
.Y(n_4909)
);

AND2x2_ASAP7_75t_L g4910 ( 
.A(n_4858),
.B(n_4773),
.Y(n_4910)
);

INVx1_ASAP7_75t_L g4911 ( 
.A(n_4886),
.Y(n_4911)
);

INVx1_ASAP7_75t_L g4912 ( 
.A(n_4886),
.Y(n_4912)
);

NOR2xp33_ASAP7_75t_L g4913 ( 
.A(n_4861),
.B(n_4744),
.Y(n_4913)
);

INVxp67_ASAP7_75t_L g4914 ( 
.A(n_4853),
.Y(n_4914)
);

INVx1_ASAP7_75t_L g4915 ( 
.A(n_4852),
.Y(n_4915)
);

INVx1_ASAP7_75t_L g4916 ( 
.A(n_4856),
.Y(n_4916)
);

INVx1_ASAP7_75t_L g4917 ( 
.A(n_4856),
.Y(n_4917)
);

NAND2xp5_ASAP7_75t_L g4918 ( 
.A(n_4853),
.B(n_4661),
.Y(n_4918)
);

INVx2_ASAP7_75t_L g4919 ( 
.A(n_4889),
.Y(n_4919)
);

INVx1_ASAP7_75t_L g4920 ( 
.A(n_4860),
.Y(n_4920)
);

INVx1_ASAP7_75t_SL g4921 ( 
.A(n_4854),
.Y(n_4921)
);

HB1xp67_ASAP7_75t_L g4922 ( 
.A(n_4854),
.Y(n_4922)
);

AND2x2_ASAP7_75t_L g4923 ( 
.A(n_4864),
.B(n_4796),
.Y(n_4923)
);

AND2x4_ASAP7_75t_SL g4924 ( 
.A(n_4865),
.B(n_4796),
.Y(n_4924)
);

INVx1_ASAP7_75t_L g4925 ( 
.A(n_4860),
.Y(n_4925)
);

INVx2_ASAP7_75t_L g4926 ( 
.A(n_4889),
.Y(n_4926)
);

INVx2_ASAP7_75t_L g4927 ( 
.A(n_4862),
.Y(n_4927)
);

AND2x2_ASAP7_75t_L g4928 ( 
.A(n_4864),
.B(n_4820),
.Y(n_4928)
);

INVx1_ASAP7_75t_L g4929 ( 
.A(n_4857),
.Y(n_4929)
);

INVx1_ASAP7_75t_L g4930 ( 
.A(n_4857),
.Y(n_4930)
);

AND2x2_ASAP7_75t_L g4931 ( 
.A(n_4837),
.B(n_4820),
.Y(n_4931)
);

INVx1_ASAP7_75t_L g4932 ( 
.A(n_4859),
.Y(n_4932)
);

INVx2_ASAP7_75t_L g4933 ( 
.A(n_4862),
.Y(n_4933)
);

INVx1_ASAP7_75t_L g4934 ( 
.A(n_4859),
.Y(n_4934)
);

AND2x4_ASAP7_75t_L g4935 ( 
.A(n_4865),
.B(n_4611),
.Y(n_4935)
);

INVx1_ASAP7_75t_L g4936 ( 
.A(n_4848),
.Y(n_4936)
);

NAND2xp5_ASAP7_75t_L g4937 ( 
.A(n_4837),
.B(n_4661),
.Y(n_4937)
);

OR2x2_ASAP7_75t_L g4938 ( 
.A(n_4894),
.B(n_4789),
.Y(n_4938)
);

AND2x4_ASAP7_75t_L g4939 ( 
.A(n_4870),
.B(n_4618),
.Y(n_4939)
);

NAND2xp5_ASAP7_75t_L g4940 ( 
.A(n_4838),
.B(n_4687),
.Y(n_4940)
);

AND2x2_ASAP7_75t_L g4941 ( 
.A(n_4838),
.B(n_4820),
.Y(n_4941)
);

AND2x2_ASAP7_75t_L g4942 ( 
.A(n_4878),
.B(n_4820),
.Y(n_4942)
);

AND2x2_ASAP7_75t_L g4943 ( 
.A(n_4878),
.B(n_4826),
.Y(n_4943)
);

AND2x2_ASAP7_75t_L g4944 ( 
.A(n_4890),
.B(n_4826),
.Y(n_4944)
);

INVx2_ASAP7_75t_L g4945 ( 
.A(n_4848),
.Y(n_4945)
);

BUFx2_ASAP7_75t_L g4946 ( 
.A(n_4875),
.Y(n_4946)
);

AND2x2_ASAP7_75t_L g4947 ( 
.A(n_4890),
.B(n_4798),
.Y(n_4947)
);

INVx1_ASAP7_75t_L g4948 ( 
.A(n_4875),
.Y(n_4948)
);

INVx1_ASAP7_75t_L g4949 ( 
.A(n_4877),
.Y(n_4949)
);

INVx1_ASAP7_75t_L g4950 ( 
.A(n_4849),
.Y(n_4950)
);

INVx1_ASAP7_75t_L g4951 ( 
.A(n_4946),
.Y(n_4951)
);

INVx1_ASAP7_75t_L g4952 ( 
.A(n_4946),
.Y(n_4952)
);

AND2x2_ASAP7_75t_L g4953 ( 
.A(n_4928),
.B(n_4871),
.Y(n_4953)
);

AND2x2_ASAP7_75t_L g4954 ( 
.A(n_4928),
.B(n_4871),
.Y(n_4954)
);

AND2x4_ASAP7_75t_SL g4955 ( 
.A(n_4908),
.B(n_4870),
.Y(n_4955)
);

INVx1_ASAP7_75t_L g4956 ( 
.A(n_4922),
.Y(n_4956)
);

INVx2_ASAP7_75t_L g4957 ( 
.A(n_4895),
.Y(n_4957)
);

NOR2xp33_ASAP7_75t_SL g4958 ( 
.A(n_4923),
.B(n_4884),
.Y(n_4958)
);

INVx1_ASAP7_75t_L g4959 ( 
.A(n_4895),
.Y(n_4959)
);

AND2x2_ASAP7_75t_L g4960 ( 
.A(n_4923),
.B(n_4892),
.Y(n_4960)
);

HB1xp67_ASAP7_75t_L g4961 ( 
.A(n_4943),
.Y(n_4961)
);

AND2x2_ASAP7_75t_L g4962 ( 
.A(n_4943),
.B(n_4892),
.Y(n_4962)
);

AND2x2_ASAP7_75t_L g4963 ( 
.A(n_4944),
.B(n_4942),
.Y(n_4963)
);

INVx1_ASAP7_75t_L g4964 ( 
.A(n_4944),
.Y(n_4964)
);

INVx1_ASAP7_75t_L g4965 ( 
.A(n_4947),
.Y(n_4965)
);

AND2x2_ASAP7_75t_L g4966 ( 
.A(n_4942),
.B(n_4893),
.Y(n_4966)
);

AND2x2_ASAP7_75t_L g4967 ( 
.A(n_4931),
.B(n_4893),
.Y(n_4967)
);

INVx2_ASAP7_75t_L g4968 ( 
.A(n_4899),
.Y(n_4968)
);

INVx2_ASAP7_75t_L g4969 ( 
.A(n_4899),
.Y(n_4969)
);

INVx2_ASAP7_75t_L g4970 ( 
.A(n_4900),
.Y(n_4970)
);

OR2x2_ASAP7_75t_L g4971 ( 
.A(n_4921),
.B(n_4839),
.Y(n_4971)
);

AND2x2_ASAP7_75t_L g4972 ( 
.A(n_4931),
.B(n_4841),
.Y(n_4972)
);

INVx2_ASAP7_75t_L g4973 ( 
.A(n_4900),
.Y(n_4973)
);

NOR2x1_ASAP7_75t_L g4974 ( 
.A(n_4948),
.B(n_4873),
.Y(n_4974)
);

INVx1_ASAP7_75t_L g4975 ( 
.A(n_4938),
.Y(n_4975)
);

INVx1_ASAP7_75t_L g4976 ( 
.A(n_4938),
.Y(n_4976)
);

AND2x2_ASAP7_75t_L g4977 ( 
.A(n_4941),
.B(n_4841),
.Y(n_4977)
);

NAND2xp5_ASAP7_75t_L g4978 ( 
.A(n_4941),
.B(n_4882),
.Y(n_4978)
);

OR2x2_ASAP7_75t_L g4979 ( 
.A(n_4948),
.B(n_4850),
.Y(n_4979)
);

AND2x2_ASAP7_75t_L g4980 ( 
.A(n_4906),
.B(n_4877),
.Y(n_4980)
);

AND2x4_ASAP7_75t_SL g4981 ( 
.A(n_4908),
.B(n_4870),
.Y(n_4981)
);

INVx1_ASAP7_75t_L g4982 ( 
.A(n_4947),
.Y(n_4982)
);

AO21x1_ASAP7_75t_L g4983 ( 
.A1(n_4911),
.A2(n_4885),
.B(n_4883),
.Y(n_4983)
);

AND2x2_ASAP7_75t_L g4984 ( 
.A(n_4906),
.B(n_4910),
.Y(n_4984)
);

AND2x4_ASAP7_75t_L g4985 ( 
.A(n_4910),
.B(n_4866),
.Y(n_4985)
);

INVx1_ASAP7_75t_L g4986 ( 
.A(n_4903),
.Y(n_4986)
);

AND2x2_ASAP7_75t_L g4987 ( 
.A(n_4924),
.B(n_4872),
.Y(n_4987)
);

NAND2xp5_ASAP7_75t_L g4988 ( 
.A(n_4924),
.B(n_4880),
.Y(n_4988)
);

AND2x4_ASAP7_75t_L g4989 ( 
.A(n_4909),
.B(n_4876),
.Y(n_4989)
);

OR2x2_ASAP7_75t_L g4990 ( 
.A(n_4949),
.B(n_4867),
.Y(n_4990)
);

AND2x2_ASAP7_75t_L g4991 ( 
.A(n_4909),
.B(n_4869),
.Y(n_4991)
);

AND2x4_ASAP7_75t_L g4992 ( 
.A(n_4896),
.B(n_4935),
.Y(n_4992)
);

OR2x2_ASAP7_75t_L g4993 ( 
.A(n_4949),
.B(n_4836),
.Y(n_4993)
);

AND2x2_ASAP7_75t_L g4994 ( 
.A(n_4914),
.B(n_4879),
.Y(n_4994)
);

INVx2_ASAP7_75t_L g4995 ( 
.A(n_4903),
.Y(n_4995)
);

OR2x2_ASAP7_75t_L g4996 ( 
.A(n_4901),
.B(n_4945),
.Y(n_4996)
);

AND2x2_ASAP7_75t_L g4997 ( 
.A(n_4945),
.B(n_4874),
.Y(n_4997)
);

AND2x2_ASAP7_75t_L g4998 ( 
.A(n_4936),
.B(n_4881),
.Y(n_4998)
);

INVxp67_ASAP7_75t_L g4999 ( 
.A(n_4918),
.Y(n_4999)
);

INVxp67_ASAP7_75t_L g5000 ( 
.A(n_4898),
.Y(n_5000)
);

AOI22xp5_ASAP7_75t_L g5001 ( 
.A1(n_4970),
.A2(n_4846),
.B1(n_4973),
.B2(n_4767),
.Y(n_5001)
);

NAND2xp5_ASAP7_75t_L g5002 ( 
.A(n_4962),
.B(n_4896),
.Y(n_5002)
);

AND2x2_ASAP7_75t_L g5003 ( 
.A(n_4953),
.B(n_4935),
.Y(n_5003)
);

INVx1_ASAP7_75t_L g5004 ( 
.A(n_4953),
.Y(n_5004)
);

INVx1_ASAP7_75t_L g5005 ( 
.A(n_4954),
.Y(n_5005)
);

AND2x2_ASAP7_75t_L g5006 ( 
.A(n_4954),
.B(n_4935),
.Y(n_5006)
);

NAND2xp5_ASAP7_75t_L g5007 ( 
.A(n_4962),
.B(n_4960),
.Y(n_5007)
);

INVx1_ASAP7_75t_L g5008 ( 
.A(n_4980),
.Y(n_5008)
);

OR2x2_ASAP7_75t_L g5009 ( 
.A(n_4961),
.B(n_4868),
.Y(n_5009)
);

OR2x2_ASAP7_75t_L g5010 ( 
.A(n_4970),
.B(n_4937),
.Y(n_5010)
);

AND2x2_ASAP7_75t_L g5011 ( 
.A(n_4960),
.B(n_4980),
.Y(n_5011)
);

OR2x2_ASAP7_75t_L g5012 ( 
.A(n_4973),
.B(n_4940),
.Y(n_5012)
);

INVx1_ASAP7_75t_L g5013 ( 
.A(n_4984),
.Y(n_5013)
);

HB1xp67_ASAP7_75t_L g5014 ( 
.A(n_4984),
.Y(n_5014)
);

INVx2_ASAP7_75t_L g5015 ( 
.A(n_4992),
.Y(n_5015)
);

NOR2xp33_ASAP7_75t_L g5016 ( 
.A(n_4958),
.B(n_4896),
.Y(n_5016)
);

NAND2xp5_ASAP7_75t_L g5017 ( 
.A(n_4966),
.B(n_4939),
.Y(n_5017)
);

HB1xp67_ASAP7_75t_L g5018 ( 
.A(n_4963),
.Y(n_5018)
);

INVx1_ASAP7_75t_L g5019 ( 
.A(n_4963),
.Y(n_5019)
);

INVx3_ASAP7_75t_L g5020 ( 
.A(n_4992),
.Y(n_5020)
);

AND2x2_ASAP7_75t_L g5021 ( 
.A(n_4966),
.B(n_4939),
.Y(n_5021)
);

AND2x2_ASAP7_75t_L g5022 ( 
.A(n_4967),
.B(n_4939),
.Y(n_5022)
);

INVx1_ASAP7_75t_L g5023 ( 
.A(n_4983),
.Y(n_5023)
);

AND2x2_ASAP7_75t_L g5024 ( 
.A(n_4967),
.B(n_4902),
.Y(n_5024)
);

AND2x2_ASAP7_75t_L g5025 ( 
.A(n_4972),
.B(n_4897),
.Y(n_5025)
);

HB1xp67_ASAP7_75t_L g5026 ( 
.A(n_4972),
.Y(n_5026)
);

INVx1_ASAP7_75t_L g5027 ( 
.A(n_4983),
.Y(n_5027)
);

NAND2xp5_ASAP7_75t_L g5028 ( 
.A(n_4977),
.B(n_4851),
.Y(n_5028)
);

INVx1_ASAP7_75t_L g5029 ( 
.A(n_4975),
.Y(n_5029)
);

AND2x2_ASAP7_75t_L g5030 ( 
.A(n_4977),
.B(n_4955),
.Y(n_5030)
);

INVx1_ASAP7_75t_L g5031 ( 
.A(n_4975),
.Y(n_5031)
);

INVx1_ASAP7_75t_L g5032 ( 
.A(n_4976),
.Y(n_5032)
);

NAND2xp5_ASAP7_75t_L g5033 ( 
.A(n_4992),
.B(n_4891),
.Y(n_5033)
);

INVx1_ASAP7_75t_L g5034 ( 
.A(n_4976),
.Y(n_5034)
);

INVx1_ASAP7_75t_L g5035 ( 
.A(n_4971),
.Y(n_5035)
);

AND2x4_ASAP7_75t_L g5036 ( 
.A(n_4955),
.B(n_4915),
.Y(n_5036)
);

AND2x2_ASAP7_75t_L g5037 ( 
.A(n_4981),
.B(n_4843),
.Y(n_5037)
);

NAND2xp5_ASAP7_75t_L g5038 ( 
.A(n_4987),
.B(n_4654),
.Y(n_5038)
);

AND2x2_ASAP7_75t_L g5039 ( 
.A(n_4981),
.B(n_4845),
.Y(n_5039)
);

OR2x2_ASAP7_75t_L g5040 ( 
.A(n_4971),
.B(n_4927),
.Y(n_5040)
);

NAND2xp5_ASAP7_75t_L g5041 ( 
.A(n_4987),
.B(n_4687),
.Y(n_5041)
);

NOR2xp33_ASAP7_75t_L g5042 ( 
.A(n_4964),
.B(n_4927),
.Y(n_5042)
);

AND2x2_ASAP7_75t_L g5043 ( 
.A(n_4991),
.B(n_4933),
.Y(n_5043)
);

INVx1_ASAP7_75t_L g5044 ( 
.A(n_4996),
.Y(n_5044)
);

AND2x2_ASAP7_75t_L g5045 ( 
.A(n_4991),
.B(n_4933),
.Y(n_5045)
);

AND2x2_ASAP7_75t_L g5046 ( 
.A(n_4965),
.B(n_4913),
.Y(n_5046)
);

AND2x2_ASAP7_75t_L g5047 ( 
.A(n_4982),
.B(n_4904),
.Y(n_5047)
);

BUFx2_ASAP7_75t_L g5048 ( 
.A(n_4985),
.Y(n_5048)
);

INVx1_ASAP7_75t_L g5049 ( 
.A(n_4996),
.Y(n_5049)
);

HB1xp67_ASAP7_75t_L g5050 ( 
.A(n_4951),
.Y(n_5050)
);

INVx1_ASAP7_75t_L g5051 ( 
.A(n_4951),
.Y(n_5051)
);

AND2x2_ASAP7_75t_L g5052 ( 
.A(n_4985),
.B(n_4905),
.Y(n_5052)
);

INVx1_ASAP7_75t_L g5053 ( 
.A(n_4990),
.Y(n_5053)
);

OR2x2_ASAP7_75t_L g5054 ( 
.A(n_5007),
.B(n_4990),
.Y(n_5054)
);

AOI22xp5_ASAP7_75t_L g5055 ( 
.A1(n_5023),
.A2(n_5027),
.B1(n_4840),
.B2(n_4767),
.Y(n_5055)
);

BUFx2_ASAP7_75t_L g5056 ( 
.A(n_5011),
.Y(n_5056)
);

AND2x2_ASAP7_75t_L g5057 ( 
.A(n_5011),
.B(n_4989),
.Y(n_5057)
);

INVx1_ASAP7_75t_L g5058 ( 
.A(n_5014),
.Y(n_5058)
);

NAND3xp33_ASAP7_75t_L g5059 ( 
.A(n_5040),
.B(n_4986),
.C(n_4959),
.Y(n_5059)
);

AND2x2_ASAP7_75t_L g5060 ( 
.A(n_5030),
.B(n_4989),
.Y(n_5060)
);

AND2x4_ASAP7_75t_L g5061 ( 
.A(n_5021),
.B(n_4985),
.Y(n_5061)
);

INVx2_ASAP7_75t_L g5062 ( 
.A(n_5021),
.Y(n_5062)
);

NAND2xp5_ASAP7_75t_SL g5063 ( 
.A(n_5022),
.B(n_5003),
.Y(n_5063)
);

NAND4xp25_ASAP7_75t_SL g5064 ( 
.A(n_5017),
.B(n_4842),
.C(n_4978),
.D(n_4988),
.Y(n_5064)
);

NAND2xp5_ASAP7_75t_L g5065 ( 
.A(n_5022),
.B(n_4997),
.Y(n_5065)
);

BUFx2_ASAP7_75t_L g5066 ( 
.A(n_5003),
.Y(n_5066)
);

AND2x4_ASAP7_75t_L g5067 ( 
.A(n_5006),
.B(n_4989),
.Y(n_5067)
);

INVx1_ASAP7_75t_L g5068 ( 
.A(n_5018),
.Y(n_5068)
);

AND2x2_ASAP7_75t_L g5069 ( 
.A(n_5030),
.B(n_4997),
.Y(n_5069)
);

INVx1_ASAP7_75t_L g5070 ( 
.A(n_5026),
.Y(n_5070)
);

INVx1_ASAP7_75t_L g5071 ( 
.A(n_5048),
.Y(n_5071)
);

AND2x2_ASAP7_75t_L g5072 ( 
.A(n_5006),
.B(n_4998),
.Y(n_5072)
);

INVx1_ASAP7_75t_SL g5073 ( 
.A(n_5040),
.Y(n_5073)
);

OR2x2_ASAP7_75t_L g5074 ( 
.A(n_5002),
.B(n_4979),
.Y(n_5074)
);

AND2x2_ASAP7_75t_L g5075 ( 
.A(n_5043),
.B(n_4998),
.Y(n_5075)
);

INVx1_ASAP7_75t_L g5076 ( 
.A(n_5043),
.Y(n_5076)
);

OR2x2_ASAP7_75t_L g5077 ( 
.A(n_5019),
.B(n_4979),
.Y(n_5077)
);

INVx1_ASAP7_75t_L g5078 ( 
.A(n_5045),
.Y(n_5078)
);

OAI22xp33_ASAP7_75t_SL g5079 ( 
.A1(n_5020),
.A2(n_4766),
.B1(n_4811),
.B2(n_4806),
.Y(n_5079)
);

INVx1_ASAP7_75t_L g5080 ( 
.A(n_5045),
.Y(n_5080)
);

INVx1_ASAP7_75t_L g5081 ( 
.A(n_5020),
.Y(n_5081)
);

INVx1_ASAP7_75t_L g5082 ( 
.A(n_5020),
.Y(n_5082)
);

INVx1_ASAP7_75t_L g5083 ( 
.A(n_5024),
.Y(n_5083)
);

INVx1_ASAP7_75t_L g5084 ( 
.A(n_5024),
.Y(n_5084)
);

OR2x2_ASAP7_75t_L g5085 ( 
.A(n_5013),
.B(n_4993),
.Y(n_5085)
);

OR2x2_ASAP7_75t_L g5086 ( 
.A(n_5004),
.B(n_4993),
.Y(n_5086)
);

AND2x2_ASAP7_75t_L g5087 ( 
.A(n_5025),
.B(n_4994),
.Y(n_5087)
);

NAND2xp5_ASAP7_75t_L g5088 ( 
.A(n_5036),
.B(n_4952),
.Y(n_5088)
);

INVx1_ASAP7_75t_L g5089 ( 
.A(n_5052),
.Y(n_5089)
);

INVx1_ASAP7_75t_L g5090 ( 
.A(n_5052),
.Y(n_5090)
);

OR2x2_ASAP7_75t_L g5091 ( 
.A(n_5005),
.B(n_4956),
.Y(n_5091)
);

OR2x2_ASAP7_75t_L g5092 ( 
.A(n_5008),
.B(n_4956),
.Y(n_5092)
);

NAND2xp5_ASAP7_75t_L g5093 ( 
.A(n_5036),
.B(n_4968),
.Y(n_5093)
);

AND2x2_ASAP7_75t_L g5094 ( 
.A(n_5025),
.B(n_4994),
.Y(n_5094)
);

INVx1_ASAP7_75t_SL g5095 ( 
.A(n_5010),
.Y(n_5095)
);

INVx1_ASAP7_75t_L g5096 ( 
.A(n_5012),
.Y(n_5096)
);

OR2x2_ASAP7_75t_L g5097 ( 
.A(n_5009),
.B(n_4823),
.Y(n_5097)
);

INVxp67_ASAP7_75t_SL g5098 ( 
.A(n_5016),
.Y(n_5098)
);

INVx1_ASAP7_75t_L g5099 ( 
.A(n_5036),
.Y(n_5099)
);

OR2x2_ASAP7_75t_L g5100 ( 
.A(n_5033),
.B(n_4957),
.Y(n_5100)
);

NAND2xp5_ASAP7_75t_L g5101 ( 
.A(n_5075),
.B(n_5057),
.Y(n_5101)
);

NAND2xp5_ASAP7_75t_L g5102 ( 
.A(n_5067),
.B(n_5016),
.Y(n_5102)
);

INVx1_ASAP7_75t_SL g5103 ( 
.A(n_5056),
.Y(n_5103)
);

INVxp67_ASAP7_75t_L g5104 ( 
.A(n_5066),
.Y(n_5104)
);

AND2x2_ASAP7_75t_L g5105 ( 
.A(n_5069),
.B(n_5037),
.Y(n_5105)
);

NOR2xp33_ASAP7_75t_L g5106 ( 
.A(n_5073),
.B(n_5044),
.Y(n_5106)
);

INVx1_ASAP7_75t_L g5107 ( 
.A(n_5087),
.Y(n_5107)
);

INVx1_ASAP7_75t_L g5108 ( 
.A(n_5094),
.Y(n_5108)
);

AND2x2_ASAP7_75t_L g5109 ( 
.A(n_5072),
.B(n_5037),
.Y(n_5109)
);

NAND2xp5_ASAP7_75t_L g5110 ( 
.A(n_5067),
.B(n_5061),
.Y(n_5110)
);

INVx1_ASAP7_75t_L g5111 ( 
.A(n_5065),
.Y(n_5111)
);

INVx1_ASAP7_75t_L g5112 ( 
.A(n_5054),
.Y(n_5112)
);

INVx2_ASAP7_75t_L g5113 ( 
.A(n_5061),
.Y(n_5113)
);

NAND2xp5_ASAP7_75t_L g5114 ( 
.A(n_5073),
.B(n_5060),
.Y(n_5114)
);

OR2x2_ASAP7_75t_L g5115 ( 
.A(n_5095),
.B(n_5049),
.Y(n_5115)
);

NAND2xp5_ASAP7_75t_L g5116 ( 
.A(n_5095),
.B(n_5015),
.Y(n_5116)
);

AND2x2_ASAP7_75t_L g5117 ( 
.A(n_5062),
.B(n_5039),
.Y(n_5117)
);

INVx1_ASAP7_75t_L g5118 ( 
.A(n_5076),
.Y(n_5118)
);

INVx1_ASAP7_75t_L g5119 ( 
.A(n_5078),
.Y(n_5119)
);

NAND2xp5_ASAP7_75t_L g5120 ( 
.A(n_5080),
.B(n_5015),
.Y(n_5120)
);

HB1xp67_ASAP7_75t_L g5121 ( 
.A(n_5059),
.Y(n_5121)
);

INVx1_ASAP7_75t_L g5122 ( 
.A(n_5093),
.Y(n_5122)
);

INVx3_ASAP7_75t_L g5123 ( 
.A(n_5077),
.Y(n_5123)
);

INVx1_ASAP7_75t_L g5124 ( 
.A(n_5085),
.Y(n_5124)
);

OR2x2_ASAP7_75t_L g5125 ( 
.A(n_5063),
.B(n_5035),
.Y(n_5125)
);

INVx1_ASAP7_75t_L g5126 ( 
.A(n_5086),
.Y(n_5126)
);

INVx1_ASAP7_75t_L g5127 ( 
.A(n_5074),
.Y(n_5127)
);

O2A1O1Ixp5_ASAP7_75t_L g5128 ( 
.A1(n_5059),
.A2(n_4885),
.B(n_4883),
.C(n_4957),
.Y(n_5128)
);

INVx2_ASAP7_75t_L g5129 ( 
.A(n_5100),
.Y(n_5129)
);

OAI22xp5_ASAP7_75t_L g5130 ( 
.A1(n_5083),
.A2(n_5000),
.B1(n_5038),
.B2(n_5028),
.Y(n_5130)
);

INVx1_ASAP7_75t_L g5131 ( 
.A(n_5084),
.Y(n_5131)
);

OR2x2_ASAP7_75t_L g5132 ( 
.A(n_5089),
.B(n_5053),
.Y(n_5132)
);

AND2x2_ASAP7_75t_L g5133 ( 
.A(n_5090),
.B(n_5039),
.Y(n_5133)
);

NAND2xp5_ASAP7_75t_L g5134 ( 
.A(n_5098),
.B(n_5042),
.Y(n_5134)
);

INVx2_ASAP7_75t_L g5135 ( 
.A(n_5097),
.Y(n_5135)
);

AND2x2_ASAP7_75t_L g5136 ( 
.A(n_5058),
.B(n_5047),
.Y(n_5136)
);

INVx2_ASAP7_75t_L g5137 ( 
.A(n_5099),
.Y(n_5137)
);

NAND2xp5_ASAP7_75t_L g5138 ( 
.A(n_5096),
.B(n_5042),
.Y(n_5138)
);

INVx1_ASAP7_75t_SL g5139 ( 
.A(n_5091),
.Y(n_5139)
);

NAND2xp5_ASAP7_75t_L g5140 ( 
.A(n_5105),
.B(n_5050),
.Y(n_5140)
);

AOI32xp33_ASAP7_75t_L g5141 ( 
.A1(n_5121),
.A2(n_4974),
.A3(n_4959),
.B1(n_5071),
.B2(n_4800),
.Y(n_5141)
);

OAI21xp33_ASAP7_75t_L g5142 ( 
.A1(n_5114),
.A2(n_4842),
.B(n_5001),
.Y(n_5142)
);

NAND2xp5_ASAP7_75t_L g5143 ( 
.A(n_5123),
.B(n_5047),
.Y(n_5143)
);

INVx1_ASAP7_75t_SL g5144 ( 
.A(n_5109),
.Y(n_5144)
);

AND2x2_ASAP7_75t_L g5145 ( 
.A(n_5117),
.B(n_5068),
.Y(n_5145)
);

INVxp33_ASAP7_75t_L g5146 ( 
.A(n_5106),
.Y(n_5146)
);

AOI21xp5_ASAP7_75t_L g5147 ( 
.A1(n_5121),
.A2(n_5088),
.B(n_5079),
.Y(n_5147)
);

INVxp67_ASAP7_75t_L g5148 ( 
.A(n_5106),
.Y(n_5148)
);

OR2x2_ASAP7_75t_L g5149 ( 
.A(n_5123),
.B(n_5092),
.Y(n_5149)
);

O2A1O1Ixp33_ASAP7_75t_L g5150 ( 
.A1(n_5128),
.A2(n_5079),
.B(n_4969),
.C(n_4968),
.Y(n_5150)
);

INVx1_ASAP7_75t_L g5151 ( 
.A(n_5123),
.Y(n_5151)
);

INVx1_ASAP7_75t_L g5152 ( 
.A(n_5101),
.Y(n_5152)
);

OR2x2_ASAP7_75t_L g5153 ( 
.A(n_5110),
.B(n_5041),
.Y(n_5153)
);

INVx1_ASAP7_75t_L g5154 ( 
.A(n_5134),
.Y(n_5154)
);

NAND2xp33_ASAP7_75t_L g5155 ( 
.A(n_5103),
.B(n_5070),
.Y(n_5155)
);

AOI322xp5_ASAP7_75t_L g5156 ( 
.A1(n_5116),
.A2(n_4766),
.A3(n_4986),
.B1(n_4995),
.B2(n_4919),
.C1(n_4926),
.C2(n_4907),
.Y(n_5156)
);

NAND2xp5_ASAP7_75t_L g5157 ( 
.A(n_5104),
.B(n_4969),
.Y(n_5157)
);

INVx1_ASAP7_75t_L g5158 ( 
.A(n_5133),
.Y(n_5158)
);

INVx1_ASAP7_75t_L g5159 ( 
.A(n_5129),
.Y(n_5159)
);

INVx1_ASAP7_75t_L g5160 ( 
.A(n_5129),
.Y(n_5160)
);

INVx2_ASAP7_75t_L g5161 ( 
.A(n_5113),
.Y(n_5161)
);

O2A1O1Ixp5_ASAP7_75t_L g5162 ( 
.A1(n_5128),
.A2(n_4816),
.B(n_4916),
.C(n_4915),
.Y(n_5162)
);

NAND2xp5_ASAP7_75t_L g5163 ( 
.A(n_5104),
.B(n_5029),
.Y(n_5163)
);

AND2x2_ASAP7_75t_L g5164 ( 
.A(n_5136),
.B(n_4999),
.Y(n_5164)
);

INVx1_ASAP7_75t_L g5165 ( 
.A(n_5125),
.Y(n_5165)
);

OAI21xp33_ASAP7_75t_L g5166 ( 
.A1(n_5102),
.A2(n_5064),
.B(n_5046),
.Y(n_5166)
);

OAI21xp33_ASAP7_75t_SL g5167 ( 
.A1(n_5139),
.A2(n_4800),
.B(n_4788),
.Y(n_5167)
);

OR2x2_ASAP7_75t_L g5168 ( 
.A(n_5113),
.B(n_4795),
.Y(n_5168)
);

OAI21xp5_ASAP7_75t_L g5169 ( 
.A1(n_5127),
.A2(n_5138),
.B(n_5112),
.Y(n_5169)
);

AND2x4_ASAP7_75t_L g5170 ( 
.A(n_5137),
.B(n_5081),
.Y(n_5170)
);

NAND2xp5_ASAP7_75t_L g5171 ( 
.A(n_5135),
.B(n_5031),
.Y(n_5171)
);

O2A1O1Ixp33_ASAP7_75t_L g5172 ( 
.A1(n_5115),
.A2(n_5082),
.B(n_5032),
.C(n_5034),
.Y(n_5172)
);

OAI21xp5_ASAP7_75t_L g5173 ( 
.A1(n_5124),
.A2(n_5055),
.B(n_5051),
.Y(n_5173)
);

O2A1O1Ixp33_ASAP7_75t_L g5174 ( 
.A1(n_5150),
.A2(n_5130),
.B(n_5135),
.C(n_5120),
.Y(n_5174)
);

INVx1_ASAP7_75t_L g5175 ( 
.A(n_5143),
.Y(n_5175)
);

OAI21xp5_ASAP7_75t_L g5176 ( 
.A1(n_5147),
.A2(n_5126),
.B(n_5137),
.Y(n_5176)
);

INVx1_ASAP7_75t_SL g5177 ( 
.A(n_5149),
.Y(n_5177)
);

INVx1_ASAP7_75t_SL g5178 ( 
.A(n_5144),
.Y(n_5178)
);

INVx1_ASAP7_75t_L g5179 ( 
.A(n_5140),
.Y(n_5179)
);

INVx1_ASAP7_75t_L g5180 ( 
.A(n_5170),
.Y(n_5180)
);

INVx2_ASAP7_75t_L g5181 ( 
.A(n_5170),
.Y(n_5181)
);

INVx1_ASAP7_75t_L g5182 ( 
.A(n_5153),
.Y(n_5182)
);

AOI21xp5_ASAP7_75t_L g5183 ( 
.A1(n_5155),
.A2(n_5108),
.B(n_5107),
.Y(n_5183)
);

O2A1O1Ixp33_ASAP7_75t_L g5184 ( 
.A1(n_5167),
.A2(n_5111),
.B(n_5122),
.C(n_5132),
.Y(n_5184)
);

INVx1_ASAP7_75t_L g5185 ( 
.A(n_5161),
.Y(n_5185)
);

OR2x2_ASAP7_75t_L g5186 ( 
.A(n_5159),
.B(n_4803),
.Y(n_5186)
);

OAI22xp33_ASAP7_75t_L g5187 ( 
.A1(n_5146),
.A2(n_5055),
.B1(n_4767),
.B2(n_4788),
.Y(n_5187)
);

OR2x2_ASAP7_75t_L g5188 ( 
.A(n_5160),
.B(n_4805),
.Y(n_5188)
);

AOI32xp33_ASAP7_75t_L g5189 ( 
.A1(n_5145),
.A2(n_5119),
.A3(n_5118),
.B1(n_5131),
.B2(n_4920),
.Y(n_5189)
);

OAI222xp33_ASAP7_75t_L g5190 ( 
.A1(n_5141),
.A2(n_4887),
.B1(n_4925),
.B2(n_4917),
.C1(n_4811),
.C2(n_4806),
.Y(n_5190)
);

AND2x2_ASAP7_75t_L g5191 ( 
.A(n_5164),
.B(n_5046),
.Y(n_5191)
);

NAND2xp5_ASAP7_75t_L g5192 ( 
.A(n_5156),
.B(n_4995),
.Y(n_5192)
);

INVx1_ASAP7_75t_L g5193 ( 
.A(n_5168),
.Y(n_5193)
);

AOI221xp5_ASAP7_75t_L g5194 ( 
.A1(n_5151),
.A2(n_4912),
.B1(n_4911),
.B2(n_4916),
.C(n_4811),
.Y(n_5194)
);

O2A1O1Ixp5_ASAP7_75t_L g5195 ( 
.A1(n_5162),
.A2(n_4816),
.B(n_4912),
.C(n_4929),
.Y(n_5195)
);

AOI21xp5_ASAP7_75t_L g5196 ( 
.A1(n_5171),
.A2(n_4932),
.B(n_4930),
.Y(n_5196)
);

OAI222xp33_ASAP7_75t_L g5197 ( 
.A1(n_5148),
.A2(n_4887),
.B1(n_4821),
.B2(n_4817),
.C1(n_4833),
.C2(n_4827),
.Y(n_5197)
);

AND2x2_ASAP7_75t_L g5198 ( 
.A(n_5158),
.B(n_4802),
.Y(n_5198)
);

NAND2xp5_ASAP7_75t_L g5199 ( 
.A(n_5165),
.B(n_4767),
.Y(n_5199)
);

NAND2xp5_ASAP7_75t_L g5200 ( 
.A(n_5152),
.B(n_4767),
.Y(n_5200)
);

NOR2xp33_ASAP7_75t_L g5201 ( 
.A(n_5157),
.B(n_4907),
.Y(n_5201)
);

INVx2_ASAP7_75t_L g5202 ( 
.A(n_5154),
.Y(n_5202)
);

INVx1_ASAP7_75t_L g5203 ( 
.A(n_5163),
.Y(n_5203)
);

OAI221xp5_ASAP7_75t_L g5204 ( 
.A1(n_5167),
.A2(n_4934),
.B1(n_4784),
.B2(n_4950),
.C(n_4809),
.Y(n_5204)
);

AOI211xp5_ASAP7_75t_L g5205 ( 
.A1(n_5172),
.A2(n_4784),
.B(n_4926),
.C(n_4919),
.Y(n_5205)
);

OAI21xp33_ASAP7_75t_L g5206 ( 
.A1(n_5166),
.A2(n_4802),
.B(n_4818),
.Y(n_5206)
);

AOI33xp33_ASAP7_75t_L g5207 ( 
.A1(n_5142),
.A2(n_4831),
.A3(n_4818),
.B1(n_4832),
.B2(n_4824),
.B3(n_4819),
.Y(n_5207)
);

AOI221xp5_ASAP7_75t_L g5208 ( 
.A1(n_5173),
.A2(n_4825),
.B1(n_4827),
.B2(n_4821),
.C(n_4817),
.Y(n_5208)
);

INVx1_ASAP7_75t_L g5209 ( 
.A(n_5169),
.Y(n_5209)
);

NAND2xp5_ASAP7_75t_L g5210 ( 
.A(n_5144),
.B(n_4691),
.Y(n_5210)
);

AOI22xp5_ASAP7_75t_L g5211 ( 
.A1(n_5159),
.A2(n_4821),
.B1(n_4825),
.B2(n_4817),
.Y(n_5211)
);

NOR3xp33_ASAP7_75t_L g5212 ( 
.A(n_5174),
.B(n_4771),
.C(n_4768),
.Y(n_5212)
);

INVx2_ASAP7_75t_L g5213 ( 
.A(n_5191),
.Y(n_5213)
);

INVx1_ASAP7_75t_L g5214 ( 
.A(n_5211),
.Y(n_5214)
);

NOR2xp33_ASAP7_75t_L g5215 ( 
.A(n_5177),
.B(n_5181),
.Y(n_5215)
);

NAND2xp5_ASAP7_75t_L g5216 ( 
.A(n_5178),
.B(n_4825),
.Y(n_5216)
);

INVx1_ASAP7_75t_L g5217 ( 
.A(n_5186),
.Y(n_5217)
);

NAND3xp33_ASAP7_75t_L g5218 ( 
.A(n_5176),
.B(n_4833),
.C(n_4827),
.Y(n_5218)
);

AOI211xp5_ASAP7_75t_L g5219 ( 
.A1(n_5187),
.A2(n_4762),
.B(n_4824),
.C(n_4819),
.Y(n_5219)
);

NOR2xp33_ASAP7_75t_L g5220 ( 
.A(n_5197),
.B(n_4833),
.Y(n_5220)
);

INVx1_ASAP7_75t_L g5221 ( 
.A(n_5188),
.Y(n_5221)
);

AOI21xp5_ASAP7_75t_L g5222 ( 
.A1(n_5184),
.A2(n_5183),
.B(n_5190),
.Y(n_5222)
);

INVx3_ASAP7_75t_L g5223 ( 
.A(n_5178),
.Y(n_5223)
);

O2A1O1Ixp5_ASAP7_75t_L g5224 ( 
.A1(n_5201),
.A2(n_4816),
.B(n_4832),
.C(n_4831),
.Y(n_5224)
);

OAI21xp33_ASAP7_75t_L g5225 ( 
.A1(n_5209),
.A2(n_4807),
.B(n_4746),
.Y(n_5225)
);

AOI21xp5_ASAP7_75t_L g5226 ( 
.A1(n_5199),
.A2(n_4816),
.B(n_4813),
.Y(n_5226)
);

OR2x2_ASAP7_75t_L g5227 ( 
.A(n_5180),
.B(n_4791),
.Y(n_5227)
);

AOI22xp33_ASAP7_75t_L g5228 ( 
.A1(n_5208),
.A2(n_4771),
.B1(n_4804),
.B2(n_4794),
.Y(n_5228)
);

OAI211xp5_ASAP7_75t_L g5229 ( 
.A1(n_5189),
.A2(n_5205),
.B(n_5206),
.C(n_5194),
.Y(n_5229)
);

AND2x4_ASAP7_75t_L g5230 ( 
.A(n_5182),
.B(n_4618),
.Y(n_5230)
);

A2O1A1Ixp33_ASAP7_75t_L g5231 ( 
.A1(n_5205),
.A2(n_4794),
.B(n_4804),
.C(n_4771),
.Y(n_5231)
);

OAI22xp5_ASAP7_75t_L g5232 ( 
.A1(n_5200),
.A2(n_4829),
.B1(n_4813),
.B2(n_4801),
.Y(n_5232)
);

INVx1_ASAP7_75t_L g5233 ( 
.A(n_5185),
.Y(n_5233)
);

NOR2xp67_ASAP7_75t_L g5234 ( 
.A(n_5196),
.B(n_4720),
.Y(n_5234)
);

NAND2xp5_ASAP7_75t_L g5235 ( 
.A(n_5193),
.B(n_4791),
.Y(n_5235)
);

O2A1O1Ixp33_ASAP7_75t_L g5236 ( 
.A1(n_5192),
.A2(n_4804),
.B(n_4794),
.C(n_4829),
.Y(n_5236)
);

AOI211xp5_ASAP7_75t_L g5237 ( 
.A1(n_5204),
.A2(n_4792),
.B(n_4828),
.C(n_4801),
.Y(n_5237)
);

XNOR2x2_ASAP7_75t_L g5238 ( 
.A(n_5179),
.B(n_4792),
.Y(n_5238)
);

OAI32xp33_ASAP7_75t_L g5239 ( 
.A1(n_5210),
.A2(n_5202),
.A3(n_5203),
.B1(n_5175),
.B2(n_5198),
.Y(n_5239)
);

AOI22xp33_ASAP7_75t_L g5240 ( 
.A1(n_5207),
.A2(n_4799),
.B1(n_4791),
.B2(n_4685),
.Y(n_5240)
);

OAI22xp33_ASAP7_75t_L g5241 ( 
.A1(n_5195),
.A2(n_4726),
.B1(n_4718),
.B2(n_4720),
.Y(n_5241)
);

AND2x2_ASAP7_75t_L g5242 ( 
.A(n_5191),
.B(n_4791),
.Y(n_5242)
);

INVx1_ASAP7_75t_L g5243 ( 
.A(n_5191),
.Y(n_5243)
);

NOR2xp33_ASAP7_75t_SL g5244 ( 
.A(n_5191),
.B(n_4759),
.Y(n_5244)
);

INVx1_ASAP7_75t_L g5245 ( 
.A(n_5191),
.Y(n_5245)
);

OAI22xp5_ASAP7_75t_L g5246 ( 
.A1(n_5177),
.A2(n_4828),
.B1(n_4700),
.B2(n_4735),
.Y(n_5246)
);

INVx2_ASAP7_75t_SL g5247 ( 
.A(n_5191),
.Y(n_5247)
);

OAI21xp5_ASAP7_75t_L g5248 ( 
.A1(n_5176),
.A2(n_4519),
.B(n_4685),
.Y(n_5248)
);

AOI22xp5_ASAP7_75t_L g5249 ( 
.A1(n_5208),
.A2(n_4799),
.B1(n_4662),
.B2(n_4674),
.Y(n_5249)
);

AOI21xp33_ASAP7_75t_L g5250 ( 
.A1(n_5201),
.A2(n_4799),
.B(n_4663),
.Y(n_5250)
);

NAND2xp5_ASAP7_75t_L g5251 ( 
.A(n_5191),
.B(n_4799),
.Y(n_5251)
);

INVx1_ASAP7_75t_L g5252 ( 
.A(n_5191),
.Y(n_5252)
);

INVx2_ASAP7_75t_L g5253 ( 
.A(n_5191),
.Y(n_5253)
);

NAND2x1p5_ASAP7_75t_L g5254 ( 
.A(n_5191),
.B(n_4720),
.Y(n_5254)
);

OAI22xp33_ASAP7_75t_L g5255 ( 
.A1(n_5177),
.A2(n_4718),
.B1(n_4720),
.B2(n_4580),
.Y(n_5255)
);

NAND2xp5_ASAP7_75t_L g5256 ( 
.A(n_5191),
.B(n_4691),
.Y(n_5256)
);

NAND2xp5_ASAP7_75t_L g5257 ( 
.A(n_5191),
.B(n_4701),
.Y(n_5257)
);

INVx1_ASAP7_75t_L g5258 ( 
.A(n_5191),
.Y(n_5258)
);

INVx1_ASAP7_75t_L g5259 ( 
.A(n_5238),
.Y(n_5259)
);

O2A1O1Ixp33_ASAP7_75t_L g5260 ( 
.A1(n_5223),
.A2(n_5216),
.B(n_5239),
.C(n_5251),
.Y(n_5260)
);

INVx1_ASAP7_75t_L g5261 ( 
.A(n_5242),
.Y(n_5261)
);

OAI221xp5_ASAP7_75t_L g5262 ( 
.A1(n_5223),
.A2(n_4700),
.B1(n_4735),
.B2(n_4746),
.C(n_4743),
.Y(n_5262)
);

AND2x2_ASAP7_75t_L g5263 ( 
.A(n_5247),
.B(n_4743),
.Y(n_5263)
);

OAI22xp33_ASAP7_75t_L g5264 ( 
.A1(n_5218),
.A2(n_5244),
.B1(n_5233),
.B2(n_5243),
.Y(n_5264)
);

OR2x2_ASAP7_75t_L g5265 ( 
.A(n_5256),
.B(n_4751),
.Y(n_5265)
);

AOI321xp33_ASAP7_75t_L g5266 ( 
.A1(n_5222),
.A2(n_5212),
.A3(n_5215),
.B1(n_5246),
.B2(n_5219),
.C(n_5236),
.Y(n_5266)
);

NAND2xp5_ASAP7_75t_SL g5267 ( 
.A(n_5213),
.B(n_4585),
.Y(n_5267)
);

AOI221xp5_ASAP7_75t_L g5268 ( 
.A1(n_5220),
.A2(n_4797),
.B1(n_4751),
.B2(n_4580),
.C(n_4714),
.Y(n_5268)
);

AOI22xp33_ASAP7_75t_L g5269 ( 
.A1(n_5214),
.A2(n_4730),
.B1(n_4741),
.B2(n_4731),
.Y(n_5269)
);

OAI211xp5_ASAP7_75t_L g5270 ( 
.A1(n_5229),
.A2(n_4713),
.B(n_4714),
.C(n_4710),
.Y(n_5270)
);

AND2x2_ASAP7_75t_L g5271 ( 
.A(n_5253),
.B(n_4624),
.Y(n_5271)
);

NOR2xp33_ASAP7_75t_SL g5272 ( 
.A(n_5245),
.B(n_4719),
.Y(n_5272)
);

AOI221xp5_ASAP7_75t_L g5273 ( 
.A1(n_5250),
.A2(n_4797),
.B1(n_4580),
.B2(n_4715),
.C(n_4713),
.Y(n_5273)
);

AOI211xp5_ASAP7_75t_L g5274 ( 
.A1(n_5252),
.A2(n_4694),
.B(n_4572),
.C(n_4757),
.Y(n_5274)
);

NAND2xp5_ASAP7_75t_L g5275 ( 
.A(n_5230),
.B(n_4701),
.Y(n_5275)
);

INVx1_ASAP7_75t_L g5276 ( 
.A(n_5227),
.Y(n_5276)
);

INVx1_ASAP7_75t_L g5277 ( 
.A(n_5258),
.Y(n_5277)
);

AND2x2_ASAP7_75t_L g5278 ( 
.A(n_5230),
.B(n_4624),
.Y(n_5278)
);

AOI221xp5_ASAP7_75t_L g5279 ( 
.A1(n_5235),
.A2(n_4721),
.B1(n_4729),
.B2(n_4715),
.C(n_4710),
.Y(n_5279)
);

NOR3xp33_ASAP7_75t_L g5280 ( 
.A(n_5217),
.B(n_4703),
.C(n_4731),
.Y(n_5280)
);

O2A1O1Ixp33_ASAP7_75t_L g5281 ( 
.A1(n_5221),
.A2(n_4703),
.B(n_4627),
.C(n_4559),
.Y(n_5281)
);

OAI21xp33_ASAP7_75t_SL g5282 ( 
.A1(n_5234),
.A2(n_5240),
.B(n_5232),
.Y(n_5282)
);

AOI22xp5_ASAP7_75t_L g5283 ( 
.A1(n_5225),
.A2(n_4572),
.B1(n_4659),
.B2(n_4551),
.Y(n_5283)
);

OAI211xp5_ASAP7_75t_L g5284 ( 
.A1(n_5226),
.A2(n_4729),
.B(n_4733),
.C(n_4721),
.Y(n_5284)
);

NAND2xp5_ASAP7_75t_L g5285 ( 
.A(n_5255),
.B(n_4547),
.Y(n_5285)
);

AOI221x1_ASAP7_75t_L g5286 ( 
.A1(n_5248),
.A2(n_4733),
.B1(n_4749),
.B2(n_4738),
.C(n_4736),
.Y(n_5286)
);

INVx1_ASAP7_75t_L g5287 ( 
.A(n_5257),
.Y(n_5287)
);

INVx2_ASAP7_75t_L g5288 ( 
.A(n_5254),
.Y(n_5288)
);

AOI21xp5_ASAP7_75t_L g5289 ( 
.A1(n_5231),
.A2(n_4758),
.B(n_4754),
.Y(n_5289)
);

NOR2x1_ASAP7_75t_L g5290 ( 
.A(n_5241),
.B(n_4719),
.Y(n_5290)
);

OAI32xp33_ASAP7_75t_L g5291 ( 
.A1(n_5228),
.A2(n_5237),
.A3(n_4585),
.B1(n_5224),
.B2(n_4722),
.Y(n_5291)
);

AOI221xp5_ASAP7_75t_L g5292 ( 
.A1(n_5249),
.A2(n_4599),
.B1(n_4551),
.B2(n_4547),
.C(n_4741),
.Y(n_5292)
);

AOI22xp5_ASAP7_75t_L g5293 ( 
.A1(n_5216),
.A2(n_4722),
.B1(n_4679),
.B2(n_4637),
.Y(n_5293)
);

OAI32xp33_ASAP7_75t_L g5294 ( 
.A1(n_5223),
.A2(n_4711),
.A3(n_4619),
.B1(n_4559),
.B2(n_4678),
.Y(n_5294)
);

INVx1_ASAP7_75t_SL g5295 ( 
.A(n_5238),
.Y(n_5295)
);

OAI22xp33_ASAP7_75t_L g5296 ( 
.A1(n_5216),
.A2(n_4573),
.B1(n_4582),
.B2(n_4678),
.Y(n_5296)
);

AOI22xp5_ASAP7_75t_L g5297 ( 
.A1(n_5216),
.A2(n_4679),
.B1(n_4637),
.B2(n_4681),
.Y(n_5297)
);

INVx1_ASAP7_75t_L g5298 ( 
.A(n_5238),
.Y(n_5298)
);

NAND2xp5_ASAP7_75t_L g5299 ( 
.A(n_5223),
.B(n_4681),
.Y(n_5299)
);

AOI221xp5_ASAP7_75t_L g5300 ( 
.A1(n_5239),
.A2(n_4529),
.B1(n_4527),
.B2(n_4707),
.C(n_4582),
.Y(n_5300)
);

AOI21xp5_ASAP7_75t_L g5301 ( 
.A1(n_5216),
.A2(n_4529),
.B(n_4527),
.Y(n_5301)
);

NAND2xp5_ASAP7_75t_L g5302 ( 
.A(n_5223),
.B(n_4619),
.Y(n_5302)
);

AOI21xp5_ASAP7_75t_L g5303 ( 
.A1(n_5216),
.A2(n_4673),
.B(n_4522),
.Y(n_5303)
);

OAI22xp33_ASAP7_75t_L g5304 ( 
.A1(n_5216),
.A2(n_4522),
.B1(n_4619),
.B2(n_4601),
.Y(n_5304)
);

NAND2xp5_ASAP7_75t_SL g5305 ( 
.A(n_5223),
.B(n_4556),
.Y(n_5305)
);

NAND2xp5_ASAP7_75t_L g5306 ( 
.A(n_5223),
.B(n_4574),
.Y(n_5306)
);

NAND2xp5_ASAP7_75t_L g5307 ( 
.A(n_5223),
.B(n_4698),
.Y(n_5307)
);

AOI221xp5_ASAP7_75t_L g5308 ( 
.A1(n_5239),
.A2(n_4630),
.B1(n_4671),
.B2(n_4698),
.C(n_4583),
.Y(n_5308)
);

INVx2_ASAP7_75t_SL g5309 ( 
.A(n_5223),
.Y(n_5309)
);

NAND2xp5_ASAP7_75t_L g5310 ( 
.A(n_5223),
.B(n_4641),
.Y(n_5310)
);

OAI21xp5_ASAP7_75t_L g5311 ( 
.A1(n_5307),
.A2(n_4522),
.B(n_4575),
.Y(n_5311)
);

NAND3xp33_ASAP7_75t_L g5312 ( 
.A(n_5259),
.B(n_4601),
.C(n_4641),
.Y(n_5312)
);

NAND2xp5_ASAP7_75t_L g5313 ( 
.A(n_5297),
.B(n_4604),
.Y(n_5313)
);

OAI211xp5_ASAP7_75t_L g5314 ( 
.A1(n_5298),
.A2(n_4521),
.B(n_4620),
.C(n_4561),
.Y(n_5314)
);

NAND2xp5_ASAP7_75t_L g5315 ( 
.A(n_5293),
.B(n_4604),
.Y(n_5315)
);

O2A1O1Ixp33_ASAP7_75t_SL g5316 ( 
.A1(n_5309),
.A2(n_4623),
.B(n_4644),
.C(n_4631),
.Y(n_5316)
);

OAI31xp33_ASAP7_75t_L g5317 ( 
.A1(n_5295),
.A2(n_4575),
.A3(n_4628),
.B(n_4583),
.Y(n_5317)
);

NOR4xp25_ASAP7_75t_L g5318 ( 
.A(n_5260),
.B(n_4628),
.C(n_4597),
.D(n_4588),
.Y(n_5318)
);

AOI221xp5_ASAP7_75t_L g5319 ( 
.A1(n_5264),
.A2(n_4575),
.B1(n_4583),
.B2(n_4633),
.C(n_4530),
.Y(n_5319)
);

NOR3xp33_ASAP7_75t_L g5320 ( 
.A(n_5261),
.B(n_4629),
.C(n_4571),
.Y(n_5320)
);

NOR2x1_ASAP7_75t_L g5321 ( 
.A(n_5277),
.B(n_4561),
.Y(n_5321)
);

OR2x2_ASAP7_75t_L g5322 ( 
.A(n_5299),
.B(n_4579),
.Y(n_5322)
);

OAI221xp5_ASAP7_75t_L g5323 ( 
.A1(n_5266),
.A2(n_4561),
.B1(n_4644),
.B2(n_4617),
.C(n_4608),
.Y(n_5323)
);

AOI21xp5_ASAP7_75t_L g5324 ( 
.A1(n_5302),
.A2(n_4614),
.B(n_4617),
.Y(n_5324)
);

NOR4xp25_ASAP7_75t_SL g5325 ( 
.A(n_5305),
.B(n_4579),
.C(n_4614),
.D(n_4716),
.Y(n_5325)
);

AOI22xp5_ASAP7_75t_L g5326 ( 
.A1(n_5272),
.A2(n_4614),
.B1(n_4591),
.B2(n_4567),
.Y(n_5326)
);

AOI211xp5_ASAP7_75t_L g5327 ( 
.A1(n_5291),
.A2(n_4626),
.B(n_4591),
.C(n_4560),
.Y(n_5327)
);

NAND3xp33_ASAP7_75t_SL g5328 ( 
.A(n_5287),
.B(n_4542),
.C(n_4716),
.Y(n_5328)
);

AOI221xp5_ASAP7_75t_L g5329 ( 
.A1(n_5282),
.A2(n_4579),
.B1(n_4716),
.B2(n_4562),
.C(n_4643),
.Y(n_5329)
);

NOR2xp33_ASAP7_75t_L g5330 ( 
.A(n_5306),
.B(n_4560),
.Y(n_5330)
);

INVx1_ASAP7_75t_L g5331 ( 
.A(n_5278),
.Y(n_5331)
);

INVx1_ASAP7_75t_L g5332 ( 
.A(n_5263),
.Y(n_5332)
);

AOI211xp5_ASAP7_75t_SL g5333 ( 
.A1(n_5288),
.A2(n_484),
.B(n_482),
.C(n_483),
.Y(n_5333)
);

NOR2x1_ASAP7_75t_SL g5334 ( 
.A(n_5310),
.B(n_4579),
.Y(n_5334)
);

AOI22xp33_ASAP7_75t_L g5335 ( 
.A1(n_5280),
.A2(n_5303),
.B1(n_5300),
.B2(n_5269),
.Y(n_5335)
);

OAI211xp5_ASAP7_75t_SL g5336 ( 
.A1(n_5276),
.A2(n_485),
.B(n_483),
.C(n_484),
.Y(n_5336)
);

OAI221xp5_ASAP7_75t_SL g5337 ( 
.A1(n_5262),
.A2(n_4716),
.B1(n_486),
.B2(n_487),
.C(n_488),
.Y(n_5337)
);

AOI21xp5_ASAP7_75t_L g5338 ( 
.A1(n_5267),
.A2(n_4716),
.B(n_485),
.Y(n_5338)
);

AOI21xp5_ASAP7_75t_L g5339 ( 
.A1(n_5285),
.A2(n_487),
.B(n_488),
.Y(n_5339)
);

NAND2xp5_ASAP7_75t_L g5340 ( 
.A(n_5274),
.B(n_688),
.Y(n_5340)
);

NAND2xp5_ASAP7_75t_L g5341 ( 
.A(n_5274),
.B(n_688),
.Y(n_5341)
);

AOI21xp5_ASAP7_75t_L g5342 ( 
.A1(n_5271),
.A2(n_489),
.B(n_490),
.Y(n_5342)
);

NOR3xp33_ASAP7_75t_SL g5343 ( 
.A(n_5275),
.B(n_687),
.C(n_489),
.Y(n_5343)
);

AOI221xp5_ASAP7_75t_L g5344 ( 
.A1(n_5294),
.A2(n_491),
.B1(n_492),
.B2(n_493),
.C(n_494),
.Y(n_5344)
);

AOI21xp33_ASAP7_75t_L g5345 ( 
.A1(n_5265),
.A2(n_491),
.B(n_492),
.Y(n_5345)
);

AOI21xp33_ASAP7_75t_L g5346 ( 
.A1(n_5292),
.A2(n_493),
.B(n_494),
.Y(n_5346)
);

NOR2xp33_ASAP7_75t_L g5347 ( 
.A(n_5283),
.B(n_496),
.Y(n_5347)
);

AOI221xp5_ASAP7_75t_SL g5348 ( 
.A1(n_5289),
.A2(n_497),
.B1(n_498),
.B2(n_499),
.C(n_500),
.Y(n_5348)
);

NOR2xp33_ASAP7_75t_L g5349 ( 
.A(n_5296),
.B(n_497),
.Y(n_5349)
);

AOI221xp5_ASAP7_75t_SL g5350 ( 
.A1(n_5335),
.A2(n_5301),
.B1(n_5279),
.B2(n_5273),
.C(n_5268),
.Y(n_5350)
);

AND2x2_ASAP7_75t_L g5351 ( 
.A(n_5318),
.B(n_5290),
.Y(n_5351)
);

AOI21xp5_ASAP7_75t_L g5352 ( 
.A1(n_5340),
.A2(n_5270),
.B(n_5304),
.Y(n_5352)
);

AOI221xp5_ASAP7_75t_L g5353 ( 
.A1(n_5312),
.A2(n_5281),
.B1(n_5308),
.B2(n_5284),
.C(n_5286),
.Y(n_5353)
);

INVx1_ASAP7_75t_L g5354 ( 
.A(n_5322),
.Y(n_5354)
);

INVx1_ASAP7_75t_L g5355 ( 
.A(n_5332),
.Y(n_5355)
);

INVx1_ASAP7_75t_L g5356 ( 
.A(n_5343),
.Y(n_5356)
);

NAND3xp33_ASAP7_75t_L g5357 ( 
.A(n_5331),
.B(n_500),
.C(n_501),
.Y(n_5357)
);

NOR3x1_ASAP7_75t_L g5358 ( 
.A(n_5341),
.B(n_502),
.C(n_503),
.Y(n_5358)
);

OAI221xp5_ASAP7_75t_L g5359 ( 
.A1(n_5317),
.A2(n_503),
.B1(n_504),
.B2(n_505),
.C(n_506),
.Y(n_5359)
);

NAND2xp5_ASAP7_75t_L g5360 ( 
.A(n_5321),
.B(n_504),
.Y(n_5360)
);

OAI21xp33_ASAP7_75t_L g5361 ( 
.A1(n_5336),
.A2(n_507),
.B(n_508),
.Y(n_5361)
);

OAI21xp33_ASAP7_75t_L g5362 ( 
.A1(n_5313),
.A2(n_509),
.B(n_510),
.Y(n_5362)
);

AOI21xp5_ASAP7_75t_L g5363 ( 
.A1(n_5346),
.A2(n_509),
.B(n_511),
.Y(n_5363)
);

INVx1_ASAP7_75t_L g5364 ( 
.A(n_5334),
.Y(n_5364)
);

OAI22xp5_ASAP7_75t_L g5365 ( 
.A1(n_5314),
.A2(n_687),
.B1(n_512),
.B2(n_513),
.Y(n_5365)
);

OAI322xp33_ASAP7_75t_L g5366 ( 
.A1(n_5347),
.A2(n_511),
.A3(n_512),
.B1(n_514),
.B2(n_515),
.C1(n_517),
.C2(n_518),
.Y(n_5366)
);

NAND4xp25_ASAP7_75t_L g5367 ( 
.A(n_5348),
.B(n_514),
.C(n_515),
.D(n_518),
.Y(n_5367)
);

AOI22xp5_ASAP7_75t_L g5368 ( 
.A1(n_5330),
.A2(n_519),
.B1(n_520),
.B2(n_521),
.Y(n_5368)
);

NAND3xp33_ASAP7_75t_L g5369 ( 
.A(n_5333),
.B(n_521),
.C(n_522),
.Y(n_5369)
);

AOI21xp5_ASAP7_75t_L g5370 ( 
.A1(n_5339),
.A2(n_523),
.B(n_524),
.Y(n_5370)
);

OAI21xp33_ASAP7_75t_L g5371 ( 
.A1(n_5319),
.A2(n_523),
.B(n_524),
.Y(n_5371)
);

XOR2x2_ASAP7_75t_L g5372 ( 
.A(n_5337),
.B(n_525),
.Y(n_5372)
);

NOR3xp33_ASAP7_75t_L g5373 ( 
.A(n_5345),
.B(n_525),
.C(n_526),
.Y(n_5373)
);

AOI211xp5_ASAP7_75t_L g5374 ( 
.A1(n_5344),
.A2(n_527),
.B(n_528),
.C(n_529),
.Y(n_5374)
);

NAND2xp5_ASAP7_75t_L g5375 ( 
.A(n_5325),
.B(n_528),
.Y(n_5375)
);

NAND2xp5_ASAP7_75t_L g5376 ( 
.A(n_5311),
.B(n_529),
.Y(n_5376)
);

AOI211xp5_ASAP7_75t_L g5377 ( 
.A1(n_5349),
.A2(n_530),
.B(n_531),
.C(n_532),
.Y(n_5377)
);

AOI211xp5_ASAP7_75t_SL g5378 ( 
.A1(n_5342),
.A2(n_685),
.B(n_531),
.C(n_533),
.Y(n_5378)
);

INVx1_ASAP7_75t_L g5379 ( 
.A(n_5315),
.Y(n_5379)
);

OAI211xp5_ASAP7_75t_SL g5380 ( 
.A1(n_5327),
.A2(n_530),
.B(n_533),
.C(n_534),
.Y(n_5380)
);

OAI211xp5_ASAP7_75t_SL g5381 ( 
.A1(n_5338),
.A2(n_534),
.B(n_536),
.C(n_537),
.Y(n_5381)
);

INVx1_ASAP7_75t_L g5382 ( 
.A(n_5328),
.Y(n_5382)
);

OAI211xp5_ASAP7_75t_SL g5383 ( 
.A1(n_5382),
.A2(n_5329),
.B(n_5316),
.C(n_5323),
.Y(n_5383)
);

NOR5xp2_ASAP7_75t_L g5384 ( 
.A(n_5359),
.B(n_5324),
.C(n_5326),
.D(n_5320),
.E(n_539),
.Y(n_5384)
);

AOI222xp33_ASAP7_75t_L g5385 ( 
.A1(n_5364),
.A2(n_536),
.B1(n_537),
.B2(n_538),
.C1(n_540),
.C2(n_541),
.Y(n_5385)
);

INVx1_ASAP7_75t_L g5386 ( 
.A(n_5360),
.Y(n_5386)
);

NOR2xp33_ASAP7_75t_L g5387 ( 
.A(n_5375),
.B(n_541),
.Y(n_5387)
);

NAND2xp5_ASAP7_75t_L g5388 ( 
.A(n_5356),
.B(n_542),
.Y(n_5388)
);

AO21x1_ASAP7_75t_L g5389 ( 
.A1(n_5351),
.A2(n_543),
.B(n_544),
.Y(n_5389)
);

AND2x2_ASAP7_75t_L g5390 ( 
.A(n_5358),
.B(n_543),
.Y(n_5390)
);

INVx1_ASAP7_75t_L g5391 ( 
.A(n_5372),
.Y(n_5391)
);

NOR2xp67_ASAP7_75t_L g5392 ( 
.A(n_5367),
.B(n_544),
.Y(n_5392)
);

INVxp67_ASAP7_75t_SL g5393 ( 
.A(n_5355),
.Y(n_5393)
);

NOR3xp33_ASAP7_75t_L g5394 ( 
.A(n_5354),
.B(n_545),
.C(n_546),
.Y(n_5394)
);

NAND2xp5_ASAP7_75t_SL g5395 ( 
.A(n_5353),
.B(n_545),
.Y(n_5395)
);

OR2x2_ASAP7_75t_L g5396 ( 
.A(n_5369),
.B(n_546),
.Y(n_5396)
);

NAND4xp25_ASAP7_75t_SL g5397 ( 
.A(n_5350),
.B(n_547),
.C(n_548),
.D(n_549),
.Y(n_5397)
);

OAI21xp33_ASAP7_75t_L g5398 ( 
.A1(n_5361),
.A2(n_548),
.B(n_550),
.Y(n_5398)
);

NAND2xp5_ASAP7_75t_SL g5399 ( 
.A(n_5352),
.B(n_5365),
.Y(n_5399)
);

NAND4xp25_ASAP7_75t_L g5400 ( 
.A(n_5378),
.B(n_550),
.C(n_551),
.D(n_552),
.Y(n_5400)
);

OAI211xp5_ASAP7_75t_L g5401 ( 
.A1(n_5379),
.A2(n_551),
.B(n_552),
.C(n_554),
.Y(n_5401)
);

AOI221x1_ASAP7_75t_L g5402 ( 
.A1(n_5371),
.A2(n_555),
.B1(n_556),
.B2(n_558),
.C(n_559),
.Y(n_5402)
);

NOR4xp25_ASAP7_75t_L g5403 ( 
.A(n_5380),
.B(n_559),
.C(n_560),
.D(n_561),
.Y(n_5403)
);

INVx1_ASAP7_75t_L g5404 ( 
.A(n_5376),
.Y(n_5404)
);

NOR2xp33_ASAP7_75t_L g5405 ( 
.A(n_5381),
.B(n_560),
.Y(n_5405)
);

NAND2xp5_ASAP7_75t_SL g5406 ( 
.A(n_5368),
.B(n_5377),
.Y(n_5406)
);

OAI211xp5_ASAP7_75t_L g5407 ( 
.A1(n_5362),
.A2(n_561),
.B(n_562),
.C(n_563),
.Y(n_5407)
);

AOI211xp5_ASAP7_75t_L g5408 ( 
.A1(n_5366),
.A2(n_562),
.B(n_563),
.C(n_564),
.Y(n_5408)
);

NAND4xp25_ASAP7_75t_L g5409 ( 
.A(n_5373),
.B(n_564),
.C(n_565),
.D(n_566),
.Y(n_5409)
);

NOR2x1_ASAP7_75t_L g5410 ( 
.A(n_5397),
.B(n_5357),
.Y(n_5410)
);

OAI221xp5_ASAP7_75t_L g5411 ( 
.A1(n_5393),
.A2(n_5374),
.B1(n_5370),
.B2(n_5363),
.C(n_569),
.Y(n_5411)
);

O2A1O1Ixp33_ASAP7_75t_L g5412 ( 
.A1(n_5399),
.A2(n_566),
.B(n_567),
.C(n_568),
.Y(n_5412)
);

NAND3xp33_ASAP7_75t_SL g5413 ( 
.A(n_5389),
.B(n_567),
.C(n_569),
.Y(n_5413)
);

NOR4xp25_ASAP7_75t_L g5414 ( 
.A(n_5383),
.B(n_570),
.C(n_571),
.D(n_572),
.Y(n_5414)
);

NAND3xp33_ASAP7_75t_L g5415 ( 
.A(n_5387),
.B(n_571),
.C(n_573),
.Y(n_5415)
);

NOR4xp75_ASAP7_75t_L g5416 ( 
.A(n_5395),
.B(n_573),
.C(n_574),
.D(n_575),
.Y(n_5416)
);

NAND3xp33_ASAP7_75t_L g5417 ( 
.A(n_5386),
.B(n_574),
.C(n_575),
.Y(n_5417)
);

NAND2xp5_ASAP7_75t_SL g5418 ( 
.A(n_5392),
.B(n_577),
.Y(n_5418)
);

NAND4xp75_ASAP7_75t_L g5419 ( 
.A(n_5391),
.B(n_578),
.C(n_579),
.D(n_580),
.Y(n_5419)
);

NAND2xp5_ASAP7_75t_L g5420 ( 
.A(n_5390),
.B(n_578),
.Y(n_5420)
);

NOR5xp2_ASAP7_75t_L g5421 ( 
.A(n_5401),
.B(n_579),
.C(n_580),
.D(n_581),
.E(n_582),
.Y(n_5421)
);

NAND4xp75_ASAP7_75t_L g5422 ( 
.A(n_5404),
.B(n_581),
.C(n_582),
.D(n_583),
.Y(n_5422)
);

INVx1_ASAP7_75t_L g5423 ( 
.A(n_5388),
.Y(n_5423)
);

NOR3xp33_ASAP7_75t_SL g5424 ( 
.A(n_5400),
.B(n_583),
.C(n_584),
.Y(n_5424)
);

O2A1O1Ixp5_ASAP7_75t_SL g5425 ( 
.A1(n_5406),
.A2(n_584),
.B(n_585),
.C(n_586),
.Y(n_5425)
);

OAI21xp33_ASAP7_75t_SL g5426 ( 
.A1(n_5405),
.A2(n_587),
.B(n_588),
.Y(n_5426)
);

NAND4xp25_ASAP7_75t_L g5427 ( 
.A(n_5384),
.B(n_588),
.C(n_589),
.D(n_591),
.Y(n_5427)
);

AOI21xp5_ASAP7_75t_L g5428 ( 
.A1(n_5385),
.A2(n_589),
.B(n_592),
.Y(n_5428)
);

NOR2x1_ASAP7_75t_L g5429 ( 
.A(n_5409),
.B(n_592),
.Y(n_5429)
);

NAND5xp2_ASAP7_75t_L g5430 ( 
.A(n_5408),
.B(n_593),
.C(n_594),
.D(n_595),
.E(n_596),
.Y(n_5430)
);

INVx1_ASAP7_75t_L g5431 ( 
.A(n_5396),
.Y(n_5431)
);

AOI221xp5_ASAP7_75t_L g5432 ( 
.A1(n_5403),
.A2(n_593),
.B1(n_595),
.B2(n_597),
.C(n_598),
.Y(n_5432)
);

NOR3xp33_ASAP7_75t_L g5433 ( 
.A(n_5394),
.B(n_597),
.C(n_599),
.Y(n_5433)
);

NAND4xp25_ASAP7_75t_SL g5434 ( 
.A(n_5402),
.B(n_599),
.C(n_600),
.D(n_601),
.Y(n_5434)
);

NOR5xp2_ASAP7_75t_L g5435 ( 
.A(n_5407),
.B(n_603),
.C(n_604),
.D(n_605),
.E(n_606),
.Y(n_5435)
);

INVx1_ASAP7_75t_L g5436 ( 
.A(n_5398),
.Y(n_5436)
);

NOR2xp33_ASAP7_75t_SL g5437 ( 
.A(n_5393),
.B(n_603),
.Y(n_5437)
);

NAND3xp33_ASAP7_75t_L g5438 ( 
.A(n_5393),
.B(n_604),
.C(n_605),
.Y(n_5438)
);

AOI211x1_ASAP7_75t_L g5439 ( 
.A1(n_5389),
.A2(n_606),
.B(n_607),
.C(n_608),
.Y(n_5439)
);

INVx3_ASAP7_75t_L g5440 ( 
.A(n_5390),
.Y(n_5440)
);

INVx2_ASAP7_75t_L g5441 ( 
.A(n_5439),
.Y(n_5441)
);

AOI22xp5_ASAP7_75t_L g5442 ( 
.A1(n_5440),
.A2(n_607),
.B1(n_608),
.B2(n_609),
.Y(n_5442)
);

AND2x4_ASAP7_75t_L g5443 ( 
.A(n_5440),
.B(n_609),
.Y(n_5443)
);

INVx1_ASAP7_75t_L g5444 ( 
.A(n_5420),
.Y(n_5444)
);

AOI22xp5_ASAP7_75t_L g5445 ( 
.A1(n_5427),
.A2(n_611),
.B1(n_613),
.B2(n_614),
.Y(n_5445)
);

NAND2xp5_ASAP7_75t_L g5446 ( 
.A(n_5431),
.B(n_613),
.Y(n_5446)
);

AOI22xp5_ASAP7_75t_L g5447 ( 
.A1(n_5410),
.A2(n_615),
.B1(n_616),
.B2(n_617),
.Y(n_5447)
);

NAND2xp5_ASAP7_75t_L g5448 ( 
.A(n_5423),
.B(n_615),
.Y(n_5448)
);

INVx3_ASAP7_75t_L g5449 ( 
.A(n_5419),
.Y(n_5449)
);

AND2x4_ASAP7_75t_L g5450 ( 
.A(n_5416),
.B(n_616),
.Y(n_5450)
);

INVx2_ASAP7_75t_L g5451 ( 
.A(n_5422),
.Y(n_5451)
);

NOR2x1_ASAP7_75t_L g5452 ( 
.A(n_5413),
.B(n_618),
.Y(n_5452)
);

NOR2x1_ASAP7_75t_L g5453 ( 
.A(n_5415),
.B(n_619),
.Y(n_5453)
);

NOR4xp25_ASAP7_75t_L g5454 ( 
.A(n_5418),
.B(n_5426),
.C(n_5411),
.D(n_5436),
.Y(n_5454)
);

INVxp33_ASAP7_75t_SL g5455 ( 
.A(n_5414),
.Y(n_5455)
);

AOI221xp5_ASAP7_75t_L g5456 ( 
.A1(n_5434),
.A2(n_619),
.B1(n_620),
.B2(n_621),
.C(n_622),
.Y(n_5456)
);

NOR2x1_ASAP7_75t_L g5457 ( 
.A(n_5438),
.B(n_620),
.Y(n_5457)
);

NOR2x1_ASAP7_75t_L g5458 ( 
.A(n_5417),
.B(n_621),
.Y(n_5458)
);

NOR2x1_ASAP7_75t_L g5459 ( 
.A(n_5430),
.B(n_622),
.Y(n_5459)
);

INVx1_ASAP7_75t_L g5460 ( 
.A(n_5429),
.Y(n_5460)
);

INVx1_ASAP7_75t_L g5461 ( 
.A(n_5437),
.Y(n_5461)
);

NOR2x1_ASAP7_75t_L g5462 ( 
.A(n_5412),
.B(n_623),
.Y(n_5462)
);

INVx1_ASAP7_75t_L g5463 ( 
.A(n_5424),
.Y(n_5463)
);

INVx1_ASAP7_75t_L g5464 ( 
.A(n_5433),
.Y(n_5464)
);

INVx1_ASAP7_75t_L g5465 ( 
.A(n_5428),
.Y(n_5465)
);

NAND4xp25_ASAP7_75t_L g5466 ( 
.A(n_5432),
.B(n_624),
.C(n_625),
.D(n_626),
.Y(n_5466)
);

AOI22xp5_ASAP7_75t_L g5467 ( 
.A1(n_5421),
.A2(n_624),
.B1(n_625),
.B2(n_627),
.Y(n_5467)
);

AND2x4_ASAP7_75t_L g5468 ( 
.A(n_5435),
.B(n_628),
.Y(n_5468)
);

AND2x2_ASAP7_75t_L g5469 ( 
.A(n_5425),
.B(n_628),
.Y(n_5469)
);

HB1xp67_ASAP7_75t_L g5470 ( 
.A(n_5443),
.Y(n_5470)
);

NOR3xp33_ASAP7_75t_L g5471 ( 
.A(n_5444),
.B(n_629),
.C(n_630),
.Y(n_5471)
);

NAND4xp75_ASAP7_75t_L g5472 ( 
.A(n_5460),
.B(n_630),
.C(n_631),
.D(n_633),
.Y(n_5472)
);

XNOR2x1_ASAP7_75t_L g5473 ( 
.A(n_5459),
.B(n_633),
.Y(n_5473)
);

OR2x2_ASAP7_75t_L g5474 ( 
.A(n_5441),
.B(n_634),
.Y(n_5474)
);

NOR2x1_ASAP7_75t_L g5475 ( 
.A(n_5461),
.B(n_634),
.Y(n_5475)
);

NAND4xp25_ASAP7_75t_SL g5476 ( 
.A(n_5456),
.B(n_636),
.C(n_637),
.D(n_638),
.Y(n_5476)
);

NOR2xp67_ASAP7_75t_L g5477 ( 
.A(n_5450),
.B(n_5468),
.Y(n_5477)
);

AND4x1_ASAP7_75t_L g5478 ( 
.A(n_5454),
.B(n_636),
.C(n_638),
.D(n_639),
.Y(n_5478)
);

AOI211x1_ASAP7_75t_SL g5479 ( 
.A1(n_5451),
.A2(n_639),
.B(n_640),
.C(n_641),
.Y(n_5479)
);

AND2x2_ASAP7_75t_L g5480 ( 
.A(n_5452),
.B(n_640),
.Y(n_5480)
);

NAND3x1_ASAP7_75t_L g5481 ( 
.A(n_5449),
.B(n_641),
.C(n_642),
.Y(n_5481)
);

NOR2x1_ASAP7_75t_L g5482 ( 
.A(n_5465),
.B(n_5463),
.Y(n_5482)
);

INVx1_ASAP7_75t_L g5483 ( 
.A(n_5446),
.Y(n_5483)
);

AND2x4_ASAP7_75t_L g5484 ( 
.A(n_5464),
.B(n_642),
.Y(n_5484)
);

NAND3xp33_ASAP7_75t_SL g5485 ( 
.A(n_5445),
.B(n_643),
.C(n_644),
.Y(n_5485)
);

INVx1_ASAP7_75t_L g5486 ( 
.A(n_5448),
.Y(n_5486)
);

AND2x4_ASAP7_75t_L g5487 ( 
.A(n_5453),
.B(n_644),
.Y(n_5487)
);

INVx2_ASAP7_75t_SL g5488 ( 
.A(n_5457),
.Y(n_5488)
);

NAND2xp5_ASAP7_75t_L g5489 ( 
.A(n_5455),
.B(n_685),
.Y(n_5489)
);

AND2x4_ASAP7_75t_L g5490 ( 
.A(n_5458),
.B(n_645),
.Y(n_5490)
);

NOR2xp33_ASAP7_75t_L g5491 ( 
.A(n_5470),
.B(n_5469),
.Y(n_5491)
);

AOI211xp5_ASAP7_75t_L g5492 ( 
.A1(n_5477),
.A2(n_5466),
.B(n_5467),
.C(n_5447),
.Y(n_5492)
);

NAND5xp2_ASAP7_75t_L g5493 ( 
.A(n_5480),
.B(n_5442),
.C(n_5462),
.D(n_647),
.E(n_648),
.Y(n_5493)
);

AND2x4_ASAP7_75t_L g5494 ( 
.A(n_5482),
.B(n_645),
.Y(n_5494)
);

OAI22xp5_ASAP7_75t_L g5495 ( 
.A1(n_5474),
.A2(n_646),
.B1(n_648),
.B2(n_649),
.Y(n_5495)
);

INVx1_ASAP7_75t_L g5496 ( 
.A(n_5473),
.Y(n_5496)
);

AND2x2_ASAP7_75t_L g5497 ( 
.A(n_5488),
.B(n_646),
.Y(n_5497)
);

OAI21xp5_ASAP7_75t_SL g5498 ( 
.A1(n_5479),
.A2(n_650),
.B(n_651),
.Y(n_5498)
);

NOR3xp33_ASAP7_75t_L g5499 ( 
.A(n_5483),
.B(n_650),
.C(n_652),
.Y(n_5499)
);

INVx1_ASAP7_75t_L g5500 ( 
.A(n_5475),
.Y(n_5500)
);

INVx1_ASAP7_75t_L g5501 ( 
.A(n_5490),
.Y(n_5501)
);

NOR3x1_ASAP7_75t_L g5502 ( 
.A(n_5472),
.B(n_652),
.C(n_653),
.Y(n_5502)
);

OAI22xp33_ASAP7_75t_L g5503 ( 
.A1(n_5486),
.A2(n_653),
.B1(n_655),
.B2(n_656),
.Y(n_5503)
);

AND3x4_ASAP7_75t_L g5504 ( 
.A(n_5494),
.B(n_5478),
.C(n_5487),
.Y(n_5504)
);

NAND4xp25_ASAP7_75t_L g5505 ( 
.A(n_5491),
.B(n_5471),
.C(n_5485),
.D(n_5489),
.Y(n_5505)
);

NAND2x1p5_ASAP7_75t_L g5506 ( 
.A(n_5501),
.B(n_5484),
.Y(n_5506)
);

NOR3xp33_ASAP7_75t_SL g5507 ( 
.A(n_5496),
.B(n_5500),
.C(n_5493),
.Y(n_5507)
);

NAND3xp33_ASAP7_75t_SL g5508 ( 
.A(n_5492),
.B(n_5481),
.C(n_5476),
.Y(n_5508)
);

INVx3_ASAP7_75t_L g5509 ( 
.A(n_5497),
.Y(n_5509)
);

AND2x2_ASAP7_75t_L g5510 ( 
.A(n_5502),
.B(n_655),
.Y(n_5510)
);

INVx1_ASAP7_75t_L g5511 ( 
.A(n_5506),
.Y(n_5511)
);

INVx1_ASAP7_75t_L g5512 ( 
.A(n_5504),
.Y(n_5512)
);

INVx1_ASAP7_75t_L g5513 ( 
.A(n_5509),
.Y(n_5513)
);

OAI22xp5_ASAP7_75t_L g5514 ( 
.A1(n_5507),
.A2(n_5498),
.B1(n_5495),
.B2(n_5499),
.Y(n_5514)
);

OR2x6_ASAP7_75t_L g5515 ( 
.A(n_5511),
.B(n_5513),
.Y(n_5515)
);

INVx2_ASAP7_75t_L g5516 ( 
.A(n_5512),
.Y(n_5516)
);

CKINVDCx20_ASAP7_75t_R g5517 ( 
.A(n_5515),
.Y(n_5517)
);

NAND2xp5_ASAP7_75t_L g5518 ( 
.A(n_5516),
.B(n_5505),
.Y(n_5518)
);

OAI22xp5_ASAP7_75t_SL g5519 ( 
.A1(n_5517),
.A2(n_5514),
.B1(n_5508),
.B2(n_5510),
.Y(n_5519)
);

INVx1_ASAP7_75t_L g5520 ( 
.A(n_5518),
.Y(n_5520)
);

AOI221xp5_ASAP7_75t_L g5521 ( 
.A1(n_5520),
.A2(n_5503),
.B1(n_658),
.B2(n_659),
.C(n_660),
.Y(n_5521)
);

AOI21x1_ASAP7_75t_L g5522 ( 
.A1(n_5521),
.A2(n_5519),
.B(n_658),
.Y(n_5522)
);

INVx1_ASAP7_75t_L g5523 ( 
.A(n_5522),
.Y(n_5523)
);

OAI331xp33_ASAP7_75t_L g5524 ( 
.A1(n_5523),
.A2(n_657),
.A3(n_659),
.B1(n_660),
.B2(n_661),
.B3(n_662),
.C1(n_663),
.Y(n_5524)
);

INVx1_ASAP7_75t_L g5525 ( 
.A(n_5524),
.Y(n_5525)
);

OA21x2_ASAP7_75t_L g5526 ( 
.A1(n_5525),
.A2(n_657),
.B(n_661),
.Y(n_5526)
);

BUFx2_ASAP7_75t_L g5527 ( 
.A(n_5526),
.Y(n_5527)
);

BUFx2_ASAP7_75t_L g5528 ( 
.A(n_5526),
.Y(n_5528)
);

OR2x6_ASAP7_75t_L g5529 ( 
.A(n_5527),
.B(n_662),
.Y(n_5529)
);

OAI21x1_ASAP7_75t_L g5530 ( 
.A1(n_5528),
.A2(n_663),
.B(n_664),
.Y(n_5530)
);

OAI221xp5_ASAP7_75t_R g5531 ( 
.A1(n_5529),
.A2(n_5530),
.B1(n_667),
.B2(n_668),
.C(n_669),
.Y(n_5531)
);

AOI221xp5_ASAP7_75t_L g5532 ( 
.A1(n_5529),
.A2(n_665),
.B1(n_667),
.B2(n_668),
.C(n_669),
.Y(n_5532)
);

AOI22xp33_ASAP7_75t_L g5533 ( 
.A1(n_5532),
.A2(n_665),
.B1(n_670),
.B2(n_671),
.Y(n_5533)
);

AOI211xp5_ASAP7_75t_L g5534 ( 
.A1(n_5533),
.A2(n_5531),
.B(n_671),
.C(n_672),
.Y(n_5534)
);


endmodule