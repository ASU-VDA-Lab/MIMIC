module fake_jpeg_17378_n_39 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_39);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_39;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_13),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_14),
.B(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_18),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_18),
.A2(n_4),
.B1(n_11),
.B2(n_8),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_22),
.A2(n_20),
.B1(n_17),
.B2(n_19),
.Y(n_26)
);

INVx3_ASAP7_75t_SL g23 ( 
.A(n_16),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_24),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_0),
.Y(n_24)
);

NOR2x1_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_0),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_25),
.A2(n_26),
.B(n_27),
.C(n_3),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_21),
.A2(n_15),
.B(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_24),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_1),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_30),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_29),
.B(n_2),
.Y(n_31)
);

NOR2x1_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_32),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_2),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_25),
.B1(n_33),
.B2(n_34),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_36),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_34),
.Y(n_38)
);

BUFx24_ASAP7_75t_SL g39 ( 
.A(n_38),
.Y(n_39)
);


endmodule