module fake_jpeg_6275_n_273 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_273);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_273;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx2_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx11_ASAP7_75t_SL g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_9),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_36),
.Y(n_43)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_12),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_21),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_40),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_24),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_44),
.B(n_49),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_25),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_50),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_25),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_56),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_32),
.A2(n_24),
.B1(n_15),
.B2(n_16),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_53),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_21),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_35),
.A2(n_24),
.B1(n_15),
.B2(n_16),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_SL g74 ( 
.A(n_57),
.B(n_58),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_32),
.B(n_30),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_23),
.Y(n_59)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_62),
.B(n_64),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_23),
.Y(n_65)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_33),
.B(n_26),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_30),
.Y(n_80)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_70),
.Y(n_88)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_76),
.B(n_80),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_78),
.A2(n_28),
.B1(n_55),
.B2(n_45),
.Y(n_89)
);

OA21x2_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_31),
.B(n_33),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_50),
.B(n_72),
.C(n_58),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_63),
.A2(n_17),
.B1(n_28),
.B2(n_27),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_52),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_87),
.Y(n_96)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_18),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g121 ( 
.A1(n_89),
.A2(n_82),
.B1(n_18),
.B2(n_19),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_74),
.A2(n_57),
.B1(n_45),
.B2(n_55),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_90),
.A2(n_94),
.B1(n_97),
.B2(n_105),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_57),
.C(n_50),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_93),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_53),
.B1(n_58),
.B2(n_45),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_92),
.A2(n_100),
.B1(n_106),
.B2(n_107),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_50),
.C(n_66),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_69),
.A2(n_55),
.B1(n_46),
.B2(n_56),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_69),
.A2(n_46),
.B1(n_61),
.B2(n_48),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_43),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_109),
.Y(n_125)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_75),
.Y(n_112)
);

BUFx8_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_85),
.A2(n_46),
.B1(n_61),
.B2(n_51),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_76),
.A2(n_48),
.B1(n_51),
.B2(n_60),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_72),
.A2(n_48),
.B1(n_51),
.B2(n_60),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_80),
.A2(n_84),
.B1(n_75),
.B2(n_67),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_108),
.A2(n_109),
.B1(n_65),
.B2(n_59),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_67),
.A2(n_58),
.B1(n_43),
.B2(n_44),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_88),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_111),
.B(n_113),
.Y(n_149)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_119),
.B1(n_121),
.B2(n_129),
.Y(n_145)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_120),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_82),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_117),
.A2(n_18),
.B(n_42),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_90),
.A2(n_82),
.B1(n_86),
.B2(n_73),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_124),
.Y(n_151)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_125),
.B(n_127),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_73),
.Y(n_126)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_91),
.A2(n_79),
.B(n_71),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_130),
.B(n_133),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_92),
.A2(n_71),
.B1(n_68),
.B2(n_70),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_100),
.A2(n_79),
.B(n_26),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_88),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_131),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_99),
.A2(n_77),
.B1(n_42),
.B2(n_47),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_132),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_102),
.A2(n_47),
.B(n_18),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_121),
.Y(n_137)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

INVx4_ASAP7_75t_SL g138 ( 
.A(n_118),
.Y(n_138)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

NOR4xp25_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_100),
.C(n_108),
.D(n_101),
.Y(n_139)
);

A2O1A1O1Ixp25_ASAP7_75t_L g174 ( 
.A1(n_139),
.A2(n_130),
.B(n_117),
.C(n_115),
.D(n_121),
.Y(n_174)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_144),
.Y(n_169)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_120),
.B(n_101),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_148),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_123),
.B(n_105),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_150),
.A2(n_116),
.B(n_113),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_111),
.B(n_103),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_152),
.A2(n_154),
.B(n_155),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_83),
.C(n_62),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_127),
.C(n_131),
.Y(n_162)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_128),
.A2(n_18),
.B(n_62),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_157),
.A2(n_147),
.B1(n_146),
.B2(n_140),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_122),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_162),
.C(n_163),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_125),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_156),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_171),
.C(n_177),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_165),
.B(n_167),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_110),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_172),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_175),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_135),
.B(n_110),
.C(n_117),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_174),
.A2(n_178),
.B(n_151),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_149),
.Y(n_175)
);

OAI32xp33_ASAP7_75t_L g176 ( 
.A1(n_155),
.A2(n_124),
.A3(n_114),
.B1(n_133),
.B2(n_22),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_154),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_114),
.C(n_95),
.Y(n_177)
);

XNOR2x2_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_18),
.Y(n_178)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_141),
.Y(n_185)
);

AOI22x1_ASAP7_75t_L g182 ( 
.A1(n_178),
.A2(n_157),
.B1(n_145),
.B2(n_147),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_182),
.A2(n_183),
.B1(n_187),
.B2(n_167),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_179),
.A2(n_144),
.B1(n_141),
.B2(n_142),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_199),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_185),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_152),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_188),
.A2(n_191),
.B1(n_194),
.B2(n_202),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_158),
.A2(n_136),
.B(n_149),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_190),
.B(n_200),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_171),
.A2(n_145),
.B1(n_150),
.B2(n_134),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_134),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_193),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_169),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_168),
.A2(n_148),
.B1(n_137),
.B2(n_77),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_95),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_201),
.Y(n_216)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_170),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_158),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_95),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_180),
.A2(n_77),
.B1(n_104),
.B2(n_22),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_164),
.B(n_104),
.C(n_22),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_162),
.C(n_177),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_212),
.C(n_219),
.Y(n_229)
);

NAND2x1_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_174),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_206),
.A2(n_11),
.B1(n_10),
.B2(n_8),
.Y(n_236)
);

INVxp33_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_208),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_191),
.A2(n_181),
.B1(n_176),
.B2(n_173),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_210),
.A2(n_217),
.B1(n_0),
.B2(n_1),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_181),
.C(n_160),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_218),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_194),
.B(n_11),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_214),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_104),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_220),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_188),
.A2(n_22),
.B1(n_20),
.B2(n_19),
.Y(n_217)
);

INVxp33_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_218),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_20),
.C(n_1),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_20),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_211),
.B(n_190),
.Y(n_224)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_224),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_205),
.A2(n_196),
.B1(n_184),
.B2(n_189),
.Y(n_225)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_225),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_221),
.A2(n_198),
.B(n_203),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_227),
.A2(n_212),
.B(n_219),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_228),
.A2(n_230),
.B(n_232),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_206),
.A2(n_183),
.B(n_198),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_205),
.A2(n_195),
.B1(n_20),
.B2(n_2),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_210),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_0),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_220),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_209),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_236),
.A2(n_10),
.B(n_11),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_238),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_217),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_241),
.A2(n_243),
.B(n_246),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_204),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_242),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_229),
.C(n_233),
.Y(n_253)
);

NAND3xp33_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_215),
.C(n_216),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_223),
.A2(n_10),
.B(n_8),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_247),
.A2(n_235),
.B1(n_223),
.B2(n_226),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_232),
.Y(n_248)
);

AOI21xp33_ASAP7_75t_L g251 ( 
.A1(n_248),
.A2(n_247),
.B(n_246),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_250),
.B(n_242),
.Y(n_261)
);

NOR2x1_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_257),
.Y(n_258)
);

AOI21x1_ASAP7_75t_L g252 ( 
.A1(n_238),
.A2(n_227),
.B(n_234),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_253),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_245),
.A2(n_229),
.B1(n_4),
.B2(n_5),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_239),
.B(n_4),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_256),
.B(n_240),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_259),
.A2(n_255),
.B(n_253),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_261),
.B(n_6),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_5),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_262),
.B(n_5),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_265),
.Y(n_268)
);

AOI21xp33_ASAP7_75t_L g264 ( 
.A1(n_258),
.A2(n_254),
.B(n_257),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_266),
.C(n_267),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_6),
.C(n_7),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_6),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_270),
.A2(n_268),
.B(n_7),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_7),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_7),
.Y(n_273)
);


endmodule