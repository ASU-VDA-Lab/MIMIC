module real_jpeg_32978_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_325;
wire n_594;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_604;
wire n_420;
wire n_431;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_588;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_0),
.Y(n_146)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_0),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_0),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_0),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_1),
.B(n_47),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_1),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_1),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_1),
.B(n_175),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_1),
.B(n_376),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_1),
.B(n_388),
.Y(n_387)
);

NAND2x1_ASAP7_75t_L g488 ( 
.A(n_1),
.B(n_489),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_1),
.B(n_494),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_2),
.B(n_62),
.Y(n_61)
);

AND2x4_ASAP7_75t_SL g79 ( 
.A(n_2),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_2),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_2),
.B(n_119),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_2),
.B(n_401),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_2),
.B(n_146),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_2),
.B(n_472),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_2),
.B(n_484),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_3),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_4),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_4),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_4),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_4),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_4),
.B(n_364),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_4),
.B(n_393),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_4),
.B(n_460),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_4),
.Y(n_478)
);

AND2x2_ASAP7_75t_SL g194 ( 
.A(n_5),
.B(n_195),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_5),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_5),
.B(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_5),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_5),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_5),
.B(n_379),
.Y(n_378)
);

AND2x2_ASAP7_75t_SL g390 ( 
.A(n_5),
.B(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_5),
.B(n_49),
.Y(n_463)
);

NAND2xp33_ASAP7_75t_R g161 ( 
.A(n_6),
.B(n_162),
.Y(n_161)
);

AO22x1_ASAP7_75t_L g171 ( 
.A1(n_6),
.A2(n_12),
.B1(n_162),
.B2(n_172),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_6),
.B(n_217),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_6),
.B(n_233),
.Y(n_232)
);

NAND2x1_ASAP7_75t_L g271 ( 
.A(n_6),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_6),
.B(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_6),
.B(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_6),
.B(n_98),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_6),
.B(n_398),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_7),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_8),
.Y(n_238)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_9),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_9),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_9),
.Y(n_285)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_10),
.Y(n_103)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_10),
.Y(n_189)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_10),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_11),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_11),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_11),
.B(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_11),
.B(n_101),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_11),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_11),
.B(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_11),
.B(n_500),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_12),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_12),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_12),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_12),
.B(n_167),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_12),
.B(n_256),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_12),
.B(n_418),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_12),
.B(n_474),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_12),
.B(n_43),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_13),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_13),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_13),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_13),
.B(n_195),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_13),
.B(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_13),
.Y(n_332)
);

NAND2x1_ASAP7_75t_L g147 ( 
.A(n_14),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_14),
.B(n_182),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_14),
.B(n_222),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_14),
.B(n_146),
.Y(n_258)
);

AND2x4_ASAP7_75t_SL g367 ( 
.A(n_14),
.B(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_14),
.B(n_420),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_14),
.B(n_157),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_14),
.B(n_515),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g20 ( 
.A1(n_15),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_20)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_16),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_16),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_16),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_17),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_17),
.B(n_199),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_17),
.B(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_17),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_17),
.B(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_17),
.B(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_17),
.B(n_78),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_18),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_135),
.B(n_603),
.Y(n_22)
);

OAI21xp33_ASAP7_75t_L g603 ( 
.A1(n_23),
.A2(n_604),
.B(n_607),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_134),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_108),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_25),
.B(n_108),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_67),
.C(n_88),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_27),
.B(n_67),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_53),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_33),
.B1(n_51),
.B2(n_52),
.Y(n_28)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_29),
.B(n_110),
.C(n_111),
.Y(n_109)
);

BUFx4f_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g398 ( 
.A(n_31),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_41),
.C(n_46),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_35),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_34),
.Y(n_116)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_36),
.A2(n_41),
.B1(n_42),
.B2(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_36),
.Y(n_107)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_39),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_40),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_40),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_40),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_40),
.Y(n_490)
);

AOI22xp33_ASAP7_75t_SL g559 ( 
.A1(n_41),
.A2(n_42),
.B1(n_99),
.B2(n_100),
.Y(n_559)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_42),
.B(n_93),
.C(n_99),
.Y(n_92)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_46),
.B(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_50),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_61),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_55),
.B(n_115),
.C(n_116),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_55),
.A2(n_125),
.B1(n_126),
.B2(n_132),
.Y(n_124)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_55),
.Y(n_132)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_60),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_66),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_66),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_81),
.C(n_84),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_76),
.C(n_79),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g570 ( 
.A1(n_69),
.A2(n_70),
.B1(n_79),
.B2(n_571),
.Y(n_570)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_74),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_75),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g421 ( 
.A(n_75),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_76),
.B(n_570),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g571 ( 
.A(n_79),
.Y(n_571)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_80),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_84),
.Y(n_91)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_87),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_88),
.B(n_580),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.C(n_104),
.Y(n_88)
);

INVxp67_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_90),
.B(n_588),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_92),
.B(n_105),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_93),
.B(n_559),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_99),
.B(n_498),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_99),
.B(n_493),
.C(n_498),
.Y(n_561)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_103),
.Y(n_335)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_103),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_133),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_117),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_124),
.Y(n_117)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_131),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI21xp33_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_545),
.B(n_594),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_137),
.Y(n_606)
);

OAI21x1_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_449),
.B(n_542),
.Y(n_137)
);

AOI21x1_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_355),
.B(n_446),
.Y(n_138)
);

AO21x2_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_259),
.B(n_354),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_240),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_141),
.B(n_240),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_191),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_142),
.B(n_444),
.C(n_445),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_159),
.Y(n_142)
);

MAJx2_ASAP7_75t_L g438 ( 
.A(n_143),
.B(n_160),
.C(n_176),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_151),
.C(n_155),
.Y(n_143)
);

XNOR2x2_ASAP7_75t_L g244 ( 
.A(n_144),
.B(n_245),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_145),
.B(n_147),
.Y(n_247)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_150),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_150),
.Y(n_319)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_150),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_151),
.B(n_156),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_154),
.Y(n_382)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_176),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_166),
.B(n_171),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_165),
.Y(n_496)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_170),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_171),
.B(n_406),
.C(n_411),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_171),
.A2(n_411),
.B1(n_412),
.B2(n_437),
.Y(n_436)
);

INVxp67_ASAP7_75t_SL g437 ( 
.A(n_171),
.Y(n_437)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_175),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_175),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_180),
.Y(n_176)
);

MAJx2_ASAP7_75t_L g383 ( 
.A(n_177),
.B(n_185),
.C(n_190),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_179),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_185),
.B1(n_186),
.B2(n_190),
.Y(n_180)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_181),
.Y(n_190)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_183),
.Y(n_220)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_183),
.Y(n_472)
);

BUFx5_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_188),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_188),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_189),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_225),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_192),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_206),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_193),
.B(n_207),
.C(n_360),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_194),
.B(n_200),
.C(n_204),
.Y(n_412)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_200),
.B1(n_204),
.B2(n_205),
.Y(n_197)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_198),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_200),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_203),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_215),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_213),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_208),
.A2(n_209),
.B1(n_213),
.B2(n_214),
.Y(n_239)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_215),
.Y(n_360)
);

MAJx2_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_219),
.C(n_221),
.Y(n_215)
);

XNOR2x1_ASAP7_75t_SL g227 ( 
.A(n_216),
.B(n_219),
.Y(n_227)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_225),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.C(n_239),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_239),
.Y(n_243)
);

MAJx2_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_232),
.C(n_235),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_229),
.A2(n_230),
.B1(n_235),
.B2(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_232),
.B(n_295),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_234),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_234),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_235),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_244),
.C(n_246),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_242),
.B(n_352),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_244),
.B(n_246),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.C(n_253),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_247),
.B(n_248),
.Y(n_298)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_251),
.Y(n_273)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx6_ASAP7_75t_L g418 ( 
.A(n_252),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_253),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_258),
.Y(n_253)
);

AO22x1_ASAP7_75t_SL g279 ( 
.A1(n_254),
.A2(n_255),
.B1(n_258),
.B2(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_258),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_348),
.B(n_353),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_299),
.B(n_347),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_291),
.Y(n_261)
);

NOR2xp67_ASAP7_75t_L g347 ( 
.A(n_262),
.B(n_291),
.Y(n_347)
);

OAI21x1_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_277),
.B(n_290),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_264),
.B(n_311),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_270),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_265),
.B(n_274),
.C(n_276),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_267),
.Y(n_309)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_274),
.B1(n_275),
.B2(n_276),
.Y(n_270)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_271),
.Y(n_276)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_281),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_281),
.Y(n_290)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_279),
.B(n_281),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_286),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_282),
.A2(n_283),
.B1(n_286),
.B2(n_287),
.Y(n_303)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_285),
.Y(n_500)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

BUFx4f_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_297),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_293),
.B(n_297),
.C(n_350),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_294),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_312),
.B(n_346),
.Y(n_299)
);

NOR2xp67_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_310),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_301),
.B(n_310),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_304),
.C(n_308),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_302),
.A2(n_303),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

NAND2xp33_ASAP7_75t_L g345 ( 
.A(n_302),
.B(n_328),
.Y(n_345)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_303),
.B(n_327),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_305),
.B(n_308),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_329),
.B(n_343),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_326),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_314),
.A2(n_344),
.B(n_345),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_320),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_315),
.A2(n_316),
.B1(n_320),
.B2(n_321),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_315),
.B(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_337),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_336),
.Y(n_330)
);

OAI21xp33_ASAP7_75t_L g337 ( 
.A1(n_331),
.A2(n_336),
.B(n_338),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_332),
.B(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx8_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_351),
.Y(n_348)
);

NAND2xp33_ASAP7_75t_SL g353 ( 
.A(n_349),
.B(n_351),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_431),
.B(n_439),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_356),
.B(n_431),
.C(n_447),
.Y(n_446)
);

XNOR2x1_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_384),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_357),
.B(n_385),
.C(n_539),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_361),
.C(n_372),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

XOR2x2_ASAP7_75t_L g432 ( 
.A(n_359),
.B(n_433),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_362),
.A2(n_372),
.B1(n_373),
.B2(n_434),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_362),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_365),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_363),
.B(n_366),
.C(n_370),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_366),
.A2(n_367),
.B1(n_370),
.B2(n_371),
.Y(n_365)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_366),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_367),
.Y(n_370)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

XOR2x2_ASAP7_75t_SL g373 ( 
.A(n_374),
.B(n_383),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_378),
.Y(n_374)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_375),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_378),
.Y(n_427)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_383),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_404),
.Y(n_384)
);

XOR2x2_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_394),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_386),
.B(n_395),
.C(n_396),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_389),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_387),
.B(n_390),
.C(n_392),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_387),
.B(n_390),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_387),
.B(n_390),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_392),
.Y(n_389)
);

AO21x1_ASAP7_75t_L g518 ( 
.A1(n_392),
.A2(n_458),
.B(n_463),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_396),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_399),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_397),
.B(n_400),
.C(n_402),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_402),
.Y(n_399)
);

XNOR2x1_ASAP7_75t_L g509 ( 
.A(n_402),
.B(n_498),
.Y(n_509)
);

MAJx2_ASAP7_75t_L g516 ( 
.A(n_402),
.B(n_499),
.C(n_508),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_404),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_413),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_405),
.Y(n_532)
);

XOR2x2_ASAP7_75t_L g435 ( 
.A(n_406),
.B(n_436),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_SL g406 ( 
.A(n_407),
.B(n_410),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_409),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_408),
.B(n_409),
.C(n_410),
.Y(n_415)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_422),
.B1(n_423),
.B2(n_430),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g430 ( 
.A(n_414),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_414),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_416),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_415),
.B(n_417),
.C(n_465),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_419),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_419),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_423),
.Y(n_533)
);

A2O1A1Ixp33_ASAP7_75t_L g423 ( 
.A1(n_424),
.A2(n_426),
.B(n_428),
.C(n_429),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_425),
.B(n_427),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_435),
.C(n_438),
.Y(n_431)
);

AOI221xp5_ASAP7_75t_L g439 ( 
.A1(n_432),
.A2(n_440),
.B1(n_441),
.B2(n_442),
.C(n_443),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_432),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_432),
.B(n_440),
.Y(n_448)
);

XNOR2x1_ASAP7_75t_L g440 ( 
.A(n_435),
.B(n_438),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_440),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_443),
.B(n_448),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_537),
.Y(n_449)
);

AOI21x1_ASAP7_75t_L g542 ( 
.A1(n_450),
.A2(n_543),
.B(n_544),
.Y(n_542)
);

OR2x2_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_526),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_451),
.B(n_526),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_466),
.Y(n_451)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_452),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_455),
.C(n_464),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_453),
.A2(n_454),
.B1(n_529),
.B2(n_530),
.Y(n_528)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_455),
.B(n_464),
.Y(n_529)
);

XNOR2x1_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_457),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_458),
.A2(n_459),
.B1(n_462),
.B2(n_463),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_458),
.A2(n_459),
.B1(n_513),
.B2(n_514),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_458),
.B(n_463),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_458),
.B(n_463),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_458),
.B(n_514),
.C(n_516),
.Y(n_568)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx3_ASAP7_75t_SL g460 ( 
.A(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_467),
.A2(n_501),
.B1(n_524),
.B2(n_525),
.Y(n_466)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_467),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_467),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_491),
.Y(n_467)
);

XNOR2x1_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_482),
.Y(n_468)
);

MAJx2_ASAP7_75t_L g572 ( 
.A(n_469),
.B(n_482),
.C(n_492),
.Y(n_572)
);

XNOR2x2_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_477),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_473),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_471),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_473),
.Y(n_564)
);

INVx5_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx5_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_477),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_479),
.Y(n_477)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_486),
.C(n_488),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_483),
.B(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_487),
.B(n_488),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_497),
.Y(n_492)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVxp67_ASAP7_75t_SL g495 ( 
.A(n_496),
.Y(n_495)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_501),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_510),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g553 ( 
.A(n_502),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_505),
.C(n_506),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_503),
.B(n_505),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_506),
.B(n_536),
.Y(n_535)
);

XNOR2x1_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_509),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_517),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_511),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_516),
.Y(n_511)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_514),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_517),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_518),
.A2(n_519),
.B(n_520),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_521),
.A2(n_522),
.B(n_523),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_525),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_527),
.B(n_531),
.C(n_535),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_528),
.B(n_535),
.Y(n_541)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_529),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_531),
.B(n_541),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_533),
.C(n_534),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_538),
.B(n_540),
.Y(n_537)
);

NOR2x1_ASAP7_75t_L g543 ( 
.A(n_538),
.B(n_540),
.Y(n_543)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_546),
.Y(n_605)
);

NOR3x1_ASAP7_75t_L g546 ( 
.A(n_547),
.B(n_577),
.C(n_589),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_549),
.B(n_573),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_549),
.B(n_573),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_550),
.B(n_556),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_552),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_552),
.B(n_557),
.C(n_566),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_553),
.B(n_554),
.C(n_555),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_557),
.B(n_566),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_558),
.B(n_560),
.Y(n_557)
);

MAJx2_ASAP7_75t_L g585 ( 
.A(n_558),
.B(n_561),
.C(n_562),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_561),
.B(n_562),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_563),
.B(n_564),
.C(n_565),
.Y(n_562)
);

XNOR2x1_ASAP7_75t_L g566 ( 
.A(n_567),
.B(n_572),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_568),
.B(n_569),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_568),
.B(n_572),
.C(n_583),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_569),
.Y(n_583)
);

MAJx2_ASAP7_75t_L g573 ( 
.A(n_574),
.B(n_575),
.C(n_576),
.Y(n_573)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_577),
.Y(n_597)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_578),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_SL g578 ( 
.A(n_579),
.B(n_581),
.Y(n_578)
);

NAND2xp33_ASAP7_75t_SL g602 ( 
.A(n_579),
.B(n_581),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_582),
.B(n_584),
.C(n_586),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g592 ( 
.A(n_582),
.B(n_593),
.Y(n_592)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_585),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_585),
.B(n_587),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_590),
.Y(n_589)
);

OAI21x1_ASAP7_75t_L g598 ( 
.A1(n_590),
.A2(n_599),
.B(n_600),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_591),
.B(n_592),
.Y(n_590)
);

OR2x2_ASAP7_75t_L g600 ( 
.A(n_591),
.B(n_592),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_595),
.B(n_601),
.Y(n_594)
);

INVxp33_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_597),
.B(n_598),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_597),
.B(n_598),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_601),
.Y(n_610)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_602),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_605),
.B(n_606),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_608),
.B(n_610),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_609),
.Y(n_608)
);


endmodule