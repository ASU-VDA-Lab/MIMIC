module fake_jpeg_9786_n_336 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_0),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_25),
.Y(n_68)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_17),
.B1(n_28),
.B2(n_20),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_50),
.A2(n_55),
.B1(n_64),
.B2(n_66),
.Y(n_96)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_54),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_17),
.B1(n_28),
.B2(n_20),
.Y(n_55)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_68),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_40),
.A2(n_28),
.B1(n_20),
.B2(n_21),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_21),
.B1(n_29),
.B2(n_33),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_68),
.B(n_33),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_71),
.B(n_93),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_58),
.A2(n_25),
.B1(n_27),
.B2(n_29),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_72),
.A2(n_94),
.B1(n_97),
.B2(n_33),
.Y(n_102)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_75),
.B(n_80),
.Y(n_105)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_78),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_56),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_82),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_35),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_56),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_46),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_95),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_54),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_88),
.Y(n_119)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

AO22x2_ASAP7_75t_L g86 ( 
.A1(n_62),
.A2(n_37),
.B1(n_45),
.B2(n_46),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_86),
.A2(n_49),
.B1(n_51),
.B2(n_60),
.Y(n_112)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_91),
.Y(n_121)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_62),
.A2(n_30),
.B1(n_29),
.B2(n_27),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_46),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_49),
.A2(n_43),
.B1(n_27),
.B2(n_25),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g134 ( 
.A(n_98),
.Y(n_134)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_99),
.B(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

OA22x2_ASAP7_75t_L g133 ( 
.A1(n_102),
.A2(n_122),
.B1(n_123),
.B2(n_81),
.Y(n_133)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_106),
.Y(n_132)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_107),
.Y(n_137)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_108),
.Y(n_142)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_110),
.Y(n_135)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_112),
.A2(n_120),
.B1(n_74),
.B2(n_51),
.Y(n_130)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_113),
.Y(n_140)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_75),
.A2(n_36),
.B1(n_39),
.B2(n_41),
.Y(n_120)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_125),
.A2(n_124),
.B1(n_114),
.B2(n_92),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_61),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_126),
.A2(n_48),
.B(n_67),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_111),
.A2(n_96),
.B1(n_71),
.B2(n_61),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_127),
.A2(n_130),
.B1(n_131),
.B2(n_153),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_99),
.A2(n_36),
.B1(n_39),
.B2(n_44),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_129),
.A2(n_138),
.B1(n_145),
.B2(n_148),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_112),
.A2(n_41),
.B1(n_44),
.B2(n_92),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_133),
.A2(n_136),
.B1(n_116),
.B2(n_67),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_100),
.A2(n_53),
.B1(n_59),
.B2(n_70),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_109),
.B(n_80),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_141),
.A2(n_119),
.B(n_103),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_110),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_109),
.A2(n_70),
.B1(n_81),
.B2(n_30),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_104),
.A2(n_30),
.B1(n_35),
.B2(n_23),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_104),
.B(n_45),
.C(n_38),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_69),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_105),
.A2(n_120),
.B1(n_124),
.B2(n_106),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_150),
.A2(n_151),
.B1(n_154),
.B2(n_24),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_117),
.A2(n_23),
.B1(n_32),
.B2(n_19),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_1),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_152),
.A2(n_34),
.B(n_22),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_121),
.A2(n_32),
.B1(n_19),
.B2(n_48),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_123),
.A2(n_34),
.B1(n_24),
.B2(n_18),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_155),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_156),
.A2(n_159),
.B(n_177),
.Y(n_196)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_157),
.B(n_160),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_141),
.B(n_148),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_158),
.B(n_137),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_146),
.A2(n_34),
.B(n_22),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_122),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_162),
.Y(n_191)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_163),
.A2(n_167),
.B1(n_169),
.B2(n_170),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_113),
.Y(n_164)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_164),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_115),
.Y(n_165)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_165),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_139),
.A2(n_116),
.B1(n_114),
.B2(n_98),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_166),
.A2(n_184),
.B1(n_132),
.B2(n_140),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_147),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_168),
.Y(n_190)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

OA21x2_ASAP7_75t_L g189 ( 
.A1(n_172),
.A2(n_183),
.B(n_133),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_145),
.Y(n_173)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_173),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_127),
.B(n_139),
.Y(n_174)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_143),
.C(n_130),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_147),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_176),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_133),
.A2(n_31),
.B1(n_24),
.B2(n_18),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_150),
.A2(n_22),
.B(n_24),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_162),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_152),
.Y(n_180)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_22),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_154),
.Y(n_194)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_138),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_169),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_1),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_186),
.B(n_198),
.C(n_212),
.Y(n_227)
);

OAI32xp33_ASAP7_75t_L g187 ( 
.A1(n_174),
.A2(n_133),
.A3(n_131),
.B1(n_137),
.B2(n_153),
.Y(n_187)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_188),
.B(n_203),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_197),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_192),
.A2(n_159),
.B(n_178),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_202),
.Y(n_221)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_155),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_132),
.C(n_140),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_199),
.A2(n_209),
.B(n_181),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_165),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_160),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_157),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_207),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_170),
.A2(n_135),
.B1(n_31),
.B2(n_24),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_173),
.B(n_78),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_156),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_213),
.B(n_195),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_204),
.A2(n_182),
.B1(n_179),
.B2(n_184),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_215),
.A2(n_239),
.B1(n_10),
.B2(n_16),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_206),
.A2(n_171),
.B1(n_177),
.B2(n_180),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_217),
.A2(n_233),
.B1(n_189),
.B2(n_190),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_218),
.A2(n_231),
.B(n_209),
.Y(n_247)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_222),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_197),
.Y(n_223)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_158),
.Y(n_224)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_224),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_185),
.A2(n_171),
.B1(n_179),
.B2(n_163),
.Y(n_225)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_225),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_188),
.B(n_183),
.Y(n_226)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_226),
.Y(n_260)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_229),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_183),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_235),
.C(n_193),
.Y(n_251)
);

XOR2x2_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_176),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_208),
.B(n_168),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_232),
.B(n_234),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_186),
.A2(n_135),
.B1(n_161),
.B2(n_144),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_200),
.B(n_201),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_194),
.B(n_191),
.C(n_196),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_192),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_238),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_161),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_189),
.A2(n_13),
.B1(n_16),
.B2(n_15),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_240),
.A2(n_244),
.B1(n_262),
.B2(n_1),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_214),
.A2(n_192),
.B1(n_211),
.B2(n_187),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_196),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_249),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_247),
.B(n_253),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_231),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_226),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_256),
.Y(n_272)
);

MAJx2_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_221),
.C(n_218),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_255),
.A2(n_215),
.B1(n_9),
.B2(n_10),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_78),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_221),
.B(n_89),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_261),
.C(n_233),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_230),
.B(n_24),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_219),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_144),
.C(n_76),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_216),
.A2(n_18),
.B1(n_8),
.B2(n_9),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_279),
.Y(n_282)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_241),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_266),
.Y(n_286)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_252),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_273),
.C(n_261),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_242),
.A2(n_238),
.B(n_229),
.Y(n_268)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_268),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_224),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_278),
.C(n_253),
.Y(n_292)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_246),
.Y(n_271)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_271),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_237),
.C(n_217),
.Y(n_273)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_274),
.Y(n_295)
);

OAI21xp33_ASAP7_75t_L g275 ( 
.A1(n_254),
.A2(n_220),
.B(n_239),
.Y(n_275)
);

MAJx2_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_243),
.C(n_260),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_276),
.B(n_277),
.Y(n_284)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_244),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_248),
.B(n_18),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_240),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_259),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_293),
.C(n_272),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_283),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_256),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_290),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_282),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_249),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_245),
.C(n_257),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_294),
.C(n_7),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_292),
.B(n_6),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_7),
.C(n_15),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_270),
.B(n_6),
.C(n_14),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_296),
.B(n_300),
.C(n_302),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_295),
.B(n_272),
.Y(n_298)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_298),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_264),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_285),
.A2(n_264),
.B1(n_275),
.B2(n_263),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_5),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_286),
.C(n_289),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_306),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_304),
.B(n_305),
.Y(n_316)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_284),
.Y(n_305)
);

INVxp33_ASAP7_75t_L g306 ( 
.A(n_288),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_307),
.B(n_7),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_2),
.C(n_3),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_308),
.Y(n_313)
);

BUFx24_ASAP7_75t_SL g309 ( 
.A(n_299),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_309),
.B(n_311),
.Y(n_322)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_310),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_297),
.A2(n_306),
.B1(n_304),
.B2(n_307),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_14),
.C(n_16),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_300),
.B(n_5),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_318),
.B(n_308),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_319),
.Y(n_329)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_314),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_320),
.B(n_323),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_9),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_325),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_2),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_2),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_326),
.A2(n_316),
.B(n_321),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_330),
.A2(n_316),
.B(n_322),
.Y(n_331)
);

AOI321xp33_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_329),
.A3(n_320),
.B1(n_327),
.B2(n_319),
.C(n_328),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_332),
.A2(n_2),
.B(n_3),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_3),
.B(n_4),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_3),
.C(n_4),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_4),
.B(n_327),
.Y(n_336)
);


endmodule