module fake_jpeg_9141_n_38 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_38);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_38;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

INVx2_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_5),
.A2(n_14),
.B1(n_4),
.B2(n_3),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_1),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_3),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_22),
.B(n_19),
.Y(n_30)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx24_ASAP7_75t_SL g31 ( 
.A(n_25),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_20),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_10),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_33),
.C(n_21),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_13),
.B1(n_15),
.B2(n_27),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_24),
.B(n_11),
.Y(n_33)
);

NAND3xp33_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_35),
.C(n_31),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_28),
.B1(n_29),
.B2(n_22),
.Y(n_37)
);

BUFx24_ASAP7_75t_SL g38 ( 
.A(n_37),
.Y(n_38)
);


endmodule