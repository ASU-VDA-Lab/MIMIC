module fake_jpeg_18045_n_241 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_241);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_241;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_9),
.B(n_8),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx5_ASAP7_75t_SL g76 ( 
.A(n_41),
.Y(n_76)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_25),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_16),
.B(n_1),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_46),
.B(n_48),
.Y(n_79)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_16),
.B(n_2),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_27),
.B(n_2),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_51),
.B(n_52),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_27),
.B(n_2),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_28),
.B(n_4),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_28),
.B(n_5),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_58),
.Y(n_80)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_57),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

NOR3xp33_ASAP7_75t_L g59 ( 
.A(n_30),
.B(n_23),
.C(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_60),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_18),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_19),
.Y(n_95)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_43),
.A2(n_31),
.B1(n_22),
.B2(n_38),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_74),
.A2(n_86),
.B(n_89),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_42),
.A2(n_31),
.B(n_22),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_75),
.B(n_82),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_26),
.C(n_19),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_77),
.B(n_85),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_23),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_24),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_83),
.B(n_84),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_39),
.B(n_24),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_63),
.A2(n_36),
.B1(n_35),
.B2(n_34),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_49),
.A2(n_38),
.B1(n_35),
.B2(n_34),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_64),
.A2(n_33),
.B1(n_29),
.B2(n_26),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_47),
.B(n_33),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_90),
.B(n_94),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_5),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_103),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_97),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_7),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_100),
.B(n_104),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_14),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_41),
.B(n_7),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_57),
.B(n_7),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_106),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_41),
.B(n_8),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_40),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_107),
.A2(n_13),
.B1(n_67),
.B2(n_101),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_67),
.A2(n_75),
.B1(n_86),
.B2(n_74),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_108),
.A2(n_116),
.B1(n_134),
.B2(n_87),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_73),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_109),
.B(n_125),
.Y(n_155)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

AOI32xp33_ASAP7_75t_L g113 ( 
.A1(n_93),
.A2(n_44),
.A3(n_58),
.B1(n_66),
.B2(n_65),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_70),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_44),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_115),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_11),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_81),
.A2(n_13),
.B1(n_66),
.B2(n_98),
.Y(n_116)
);

INVx5_ASAP7_75t_SL g117 ( 
.A(n_68),
.Y(n_117)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_105),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_130),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_89),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_124),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_78),
.B(n_91),
.Y(n_125)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_68),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_132),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_71),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_68),
.Y(n_133)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_102),
.A2(n_70),
.B1(n_72),
.B2(n_76),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_69),
.B(n_97),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_69),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_139),
.Y(n_147)
);

INVx13_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_107),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_142),
.A2(n_134),
.B(n_126),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_148),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_112),
.B(n_72),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_112),
.B(n_114),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_121),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_131),
.Y(n_182)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

INVxp33_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_71),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_115),
.C(n_122),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_156),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_130),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_158),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_109),
.B(n_88),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_159),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_110),
.Y(n_160)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_160),
.Y(n_167)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_88),
.Y(n_163)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_163),
.Y(n_178)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_165),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_142),
.A2(n_128),
.B1(n_129),
.B2(n_126),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_166),
.A2(n_171),
.B1(n_181),
.B2(n_184),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_142),
.A2(n_128),
.B1(n_113),
.B2(n_129),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_173),
.Y(n_194)
);

MAJx2_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_172),
.C(n_182),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_165),
.A2(n_150),
.B1(n_158),
.B2(n_143),
.Y(n_171)
);

MAJx2_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_136),
.C(n_135),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_141),
.A2(n_111),
.B(n_138),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_185),
.Y(n_188)
);

OAI321xp33_ASAP7_75t_L g189 ( 
.A1(n_179),
.A2(n_140),
.A3(n_155),
.B1(n_145),
.B2(n_160),
.C(n_154),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_156),
.A2(n_127),
.B1(n_111),
.B2(n_117),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_143),
.B(n_133),
.C(n_139),
.Y(n_185)
);

A2O1A1O1Ixp25_ASAP7_75t_L g186 ( 
.A1(n_182),
.A2(n_148),
.B(n_149),
.C(n_140),
.D(n_155),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_SL g213 ( 
.A(n_186),
.B(n_187),
.C(n_189),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_144),
.Y(n_190)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_190),
.Y(n_210)
);

A2O1A1O1Ixp25_ASAP7_75t_L g191 ( 
.A1(n_168),
.A2(n_157),
.B(n_153),
.C(n_147),
.D(n_154),
.Y(n_191)
);

A2O1A1Ixp33_ASAP7_75t_L g203 ( 
.A1(n_191),
.A2(n_169),
.B(n_183),
.C(n_188),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_184),
.A2(n_157),
.B1(n_153),
.B2(n_144),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_192),
.A2(n_200),
.B1(n_183),
.B2(n_180),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_177),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_193),
.B(n_201),
.Y(n_205)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_195),
.Y(n_206)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_196),
.Y(n_208)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_198),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_180),
.A2(n_161),
.B1(n_151),
.B2(n_164),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_178),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_181),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_199),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_191),
.A2(n_162),
.B1(n_164),
.B2(n_176),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_204),
.A2(n_207),
.B1(n_187),
.B2(n_192),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_188),
.A2(n_175),
.B1(n_166),
.B2(n_185),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_190),
.A2(n_179),
.B(n_171),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_211),
.A2(n_194),
.B(n_199),
.Y(n_219)
);

NOR3xp33_ASAP7_75t_SL g214 ( 
.A(n_213),
.B(n_186),
.C(n_172),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_214),
.A2(n_219),
.B(n_172),
.Y(n_226)
);

A2O1A1Ixp33_ASAP7_75t_SL g223 ( 
.A1(n_215),
.A2(n_216),
.B(n_207),
.C(n_202),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_210),
.A2(n_211),
.B1(n_194),
.B2(n_203),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_174),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_217),
.B(n_220),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_200),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_209),
.B(n_173),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_221),
.B(n_210),
.Y(n_224)
);

AO21x1_ASAP7_75t_L g232 ( 
.A1(n_223),
.A2(n_225),
.B(n_226),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_227),
.Y(n_231)
);

NOR2xp67_ASAP7_75t_SL g225 ( 
.A(n_219),
.B(n_213),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_216),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_215),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_229),
.B(n_233),
.C(n_212),
.Y(n_234)
);

NOR3xp33_ASAP7_75t_SL g230 ( 
.A(n_222),
.B(n_214),
.C(n_218),
.Y(n_230)
);

AOI31xp33_ASAP7_75t_SL g237 ( 
.A1(n_230),
.A2(n_133),
.A3(n_161),
.B(n_232),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_206),
.C(n_208),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_234),
.B(n_235),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_170),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_232),
.B(n_146),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_236),
.A2(n_237),
.B(n_230),
.Y(n_239)
);

BUFx24_ASAP7_75t_SL g240 ( 
.A(n_239),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_240),
.B(n_238),
.Y(n_241)
);


endmodule