module fake_jpeg_16514_n_293 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_293);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_293;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_272;
wire n_265;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_4),
.B(n_8),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx4_ASAP7_75t_SL g33 ( 
.A(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_8),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_42),
.Y(n_45)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_32),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_34),
.A2(n_24),
.B1(n_22),
.B2(n_28),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_33),
.B1(n_23),
.B2(n_27),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_30),
.Y(n_51)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_25),
.Y(n_52)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_24),
.B1(n_28),
.B2(n_22),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_54),
.A2(n_25),
.B1(n_23),
.B2(n_27),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_30),
.Y(n_56)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_25),
.Y(n_59)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_37),
.A2(n_24),
.B1(n_28),
.B2(n_22),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_61),
.A2(n_22),
.B1(n_24),
.B2(n_28),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_75),
.B1(n_23),
.B2(n_43),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_21),
.Y(n_63)
);

OAI32xp33_ASAP7_75t_L g99 ( 
.A1(n_63),
.A2(n_45),
.A3(n_56),
.B1(n_51),
.B2(n_48),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_65),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_69),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_58),
.Y(n_72)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_52),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_73),
.B(n_76),
.Y(n_109)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_57),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_77),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_54),
.A2(n_36),
.B1(n_20),
.B2(n_26),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_78),
.A2(n_79),
.B1(n_61),
.B2(n_27),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_82),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_58),
.Y(n_83)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_84),
.Y(n_113)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_85),
.Y(n_96)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_90),
.B1(n_112),
.B2(n_81),
.Y(n_116)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_67),
.A2(n_26),
.B1(n_20),
.B2(n_47),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_63),
.Y(n_119)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_73),
.B(n_64),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_103),
.A2(n_111),
.B(n_21),
.Y(n_140)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_70),
.A2(n_47),
.B1(n_55),
.B2(n_49),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_108),
.A2(n_33),
.B1(n_39),
.B2(n_46),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_72),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_72),
.Y(n_121)
);

NOR2x1_ASAP7_75t_R g111 ( 
.A(n_70),
.B(n_21),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_67),
.A2(n_71),
.B1(n_81),
.B2(n_80),
.Y(n_112)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_116),
.A2(n_126),
.B1(n_136),
.B2(n_137),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_119),
.B(n_95),
.Y(n_164)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_71),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_122),
.B(n_132),
.Y(n_166)
);

OA22x2_ASAP7_75t_L g123 ( 
.A1(n_111),
.A2(n_83),
.B1(n_85),
.B2(n_68),
.Y(n_123)
);

OA21x2_ASAP7_75t_L g155 ( 
.A1(n_123),
.A2(n_95),
.B(n_21),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_68),
.C(n_62),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_108),
.C(n_101),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_99),
.A2(n_55),
.B1(n_83),
.B2(n_49),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_91),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_130),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_94),
.A2(n_79),
.B(n_21),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_128),
.A2(n_140),
.B(n_96),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_115),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_55),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_77),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_135),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_60),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_90),
.A2(n_60),
.B1(n_40),
.B2(n_38),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_89),
.A2(n_60),
.B1(n_40),
.B2(n_38),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_46),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_138),
.B(n_139),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_144),
.C(n_147),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_97),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_143),
.A2(n_155),
.B(n_165),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_124),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_106),
.C(n_97),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_133),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_149),
.B(n_156),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_126),
.A2(n_101),
.B1(n_107),
.B2(n_110),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_150),
.A2(n_154),
.B1(n_161),
.B2(n_33),
.Y(n_194)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_117),
.Y(n_151)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_152),
.Y(n_176)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_125),
.A2(n_110),
.B1(n_105),
.B2(n_100),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_117),
.Y(n_156)
);

INVx13_ASAP7_75t_L g157 ( 
.A(n_118),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

AND2x2_ASAP7_75t_SL g159 ( 
.A(n_132),
.B(n_123),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_159),
.A2(n_131),
.B1(n_120),
.B2(n_136),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_118),
.B(n_106),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_162),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_125),
.A2(n_105),
.B1(n_100),
.B2(n_92),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_129),
.Y(n_162)
);

INVx13_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_122),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_128),
.A2(n_92),
.B(n_2),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_168),
.A2(n_123),
.B(n_121),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_120),
.B(n_88),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_169),
.B(n_131),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_179),
.C(n_181),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_172),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_173),
.A2(n_174),
.B(n_191),
.Y(n_220)
);

FAx1_ASAP7_75t_SL g177 ( 
.A(n_144),
.B(n_137),
.CI(n_139),
.CON(n_177),
.SN(n_177)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_177),
.B(n_180),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_102),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_145),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_142),
.B(n_129),
.C(n_65),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_166),
.B(n_26),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_183),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_20),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_40),
.C(n_32),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_187),
.C(n_189),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_143),
.A2(n_16),
.B(n_19),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_186),
.A2(n_141),
.B(n_149),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_166),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_152),
.B(n_32),
.C(n_38),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_168),
.A2(n_16),
.B(n_19),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_153),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_193),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_158),
.B(n_16),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_194),
.A2(n_156),
.B1(n_162),
.B2(n_146),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_143),
.B(n_21),
.Y(n_195)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_195),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_46),
.C(n_31),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_154),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_159),
.A2(n_46),
.B1(n_29),
.B2(n_19),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_197),
.A2(n_198),
.B1(n_29),
.B2(n_148),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_148),
.A2(n_29),
.B1(n_2),
.B2(n_3),
.Y(n_198)
);

O2A1O1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_173),
.A2(n_155),
.B(n_167),
.C(n_141),
.Y(n_200)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_200),
.Y(n_223)
);

OA21x2_ASAP7_75t_L g201 ( 
.A1(n_170),
.A2(n_155),
.B(n_150),
.Y(n_201)
);

OA22x2_ASAP7_75t_L g231 ( 
.A1(n_201),
.A2(n_195),
.B1(n_21),
.B2(n_15),
.Y(n_231)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_188),
.Y(n_203)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_203),
.Y(n_224)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_190),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_206),
.B(n_198),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_185),
.B(n_167),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_207),
.B(n_213),
.Y(n_222)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_175),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_217),
.Y(n_238)
);

BUFx12_ASAP7_75t_L g213 ( 
.A(n_181),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_31),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_177),
.A2(n_146),
.B1(n_161),
.B2(n_157),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_215),
.A2(n_218),
.B1(n_219),
.B2(n_39),
.Y(n_237)
);

AOI322xp5_ASAP7_75t_SL g217 ( 
.A1(n_187),
.A2(n_171),
.A3(n_191),
.B1(n_179),
.B2(n_178),
.C1(n_170),
.C2(n_186),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_177),
.A2(n_163),
.B1(n_151),
.B2(n_3),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_174),
.A2(n_163),
.B(n_2),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_225),
.B(n_207),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_178),
.C(n_184),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_233),
.C(n_239),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_211),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_236),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_214),
.A2(n_176),
.B1(n_196),
.B2(n_189),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_228),
.A2(n_232),
.B1(n_234),
.B2(n_223),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_199),
.B(n_197),
.Y(n_230)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_230),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_231),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_203),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_215),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_202),
.A2(n_10),
.B1(n_14),
.B2(n_13),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_235),
.A2(n_204),
.B1(n_212),
.B2(n_201),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_220),
.B(n_10),
.Y(n_236)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_237),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_31),
.C(n_4),
.Y(n_239)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_240),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_221),
.C(n_213),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_246),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_253),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_213),
.C(n_218),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_238),
.A2(n_219),
.B(n_208),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_247),
.A2(n_224),
.B(n_229),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_220),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_241),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_222),
.B(n_216),
.Y(n_251)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_251),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_206),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_252),
.B(n_234),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_255),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_244),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_253),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_259),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_249),
.A2(n_210),
.B1(n_231),
.B2(n_233),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_262),
.A2(n_239),
.B1(n_245),
.B2(n_241),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_250),
.C(n_231),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_260),
.A2(n_244),
.B(n_248),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_264),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_266),
.A2(n_269),
.B(n_273),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_242),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_267),
.B(n_272),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_270),
.C(n_265),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_258),
.A2(n_9),
.B(n_14),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_31),
.C(n_5),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_261),
.B(n_9),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_259),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_274),
.B(n_275),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_31),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_12),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_277),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_12),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_273),
.B(n_13),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_279),
.B(n_6),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_285),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_280),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_275),
.A2(n_7),
.B(n_281),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_286),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_282),
.Y(n_289)
);

BUFx24_ASAP7_75t_SL g290 ( 
.A(n_289),
.Y(n_290)
);

XNOR2x2_ASAP7_75t_SL g291 ( 
.A(n_290),
.B(n_282),
.Y(n_291)
);

AOI21x1_ASAP7_75t_L g292 ( 
.A1(n_291),
.A2(n_287),
.B(n_284),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_288),
.Y(n_293)
);


endmodule