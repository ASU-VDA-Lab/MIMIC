module fake_jpeg_16087_n_245 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_245);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_245;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVxp33_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_42),
.Y(n_55)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_23),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_19),
.B(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_18),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx5_ASAP7_75t_SL g58 ( 
.A(n_44),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_24),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_38),
.A2(n_29),
.B1(n_23),
.B2(n_17),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_56),
.B1(n_33),
.B2(n_32),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_27),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_47),
.B(n_60),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_49),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_17),
.B1(n_29),
.B2(n_25),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_51),
.A2(n_61),
.B1(n_39),
.B2(n_37),
.Y(n_74)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_36),
.A2(n_25),
.B1(n_22),
.B2(n_30),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_57),
.B(n_62),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_28),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_36),
.A2(n_22),
.B1(n_18),
.B2(n_33),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_26),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_39),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_76),
.Y(n_102)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_55),
.B(n_26),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_71),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_45),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_72),
.B(n_81),
.Y(n_119)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_74),
.A2(n_53),
.B1(n_59),
.B2(n_50),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_0),
.Y(n_75)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_1),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_37),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_83),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_46),
.A2(n_35),
.B1(n_32),
.B2(n_21),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_79),
.A2(n_88),
.B1(n_94),
.B2(n_10),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_51),
.A2(n_24),
.B1(n_34),
.B2(n_3),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_82),
.B1(n_7),
.B2(n_9),
.Y(n_97)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_34),
.B1(n_2),
.B2(n_4),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_47),
.B(n_1),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_58),
.A2(n_48),
.B1(n_52),
.B2(n_53),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_85),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_1),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_86),
.A2(n_7),
.B(n_9),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_60),
.B(n_2),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_89),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_48),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_5),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_58),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_91),
.A2(n_58),
.B(n_49),
.Y(n_95)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_15),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_52),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_95),
.B(n_73),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_96),
.B(n_88),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_97),
.A2(n_99),
.B1(n_108),
.B2(n_91),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_52),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_100),
.C(n_70),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_90),
.A2(n_49),
.B(n_59),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_59),
.B1(n_11),
.B2(n_12),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_105),
.A2(n_111),
.B1(n_76),
.B2(n_83),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_75),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_109),
.A2(n_80),
.B1(n_89),
.B2(n_16),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_64),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_90),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_65),
.B(n_15),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_86),
.Y(n_132)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_121),
.B(n_132),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_114),
.A2(n_81),
.B1(n_69),
.B2(n_82),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_133),
.B1(n_105),
.B2(n_97),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_119),
.B(n_107),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_127),
.Y(n_150)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_107),
.B(n_68),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_139),
.Y(n_151)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_113),
.A2(n_79),
.B1(n_86),
.B2(n_71),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_134),
.A2(n_144),
.B(n_101),
.Y(n_169)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_136),
.A2(n_145),
.B1(n_118),
.B2(n_116),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_142),
.Y(n_157)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_117),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_146),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_98),
.B(n_87),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_143),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_68),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_106),
.B(n_93),
.C(n_92),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_113),
.A2(n_77),
.B1(n_85),
.B2(n_66),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_155),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_122),
.A2(n_120),
.B1(n_100),
.B2(n_102),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_158),
.A2(n_170),
.B(n_95),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_163),
.B(n_168),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_133),
.A2(n_120),
.B1(n_102),
.B2(n_108),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_164),
.A2(n_169),
.B1(n_156),
.B2(n_153),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_93),
.Y(n_165)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_165),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_103),
.Y(n_166)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_123),
.B(n_103),
.Y(n_167)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_167),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_135),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_169),
.B(n_121),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_138),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_142),
.Y(n_171)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_137),
.C(n_141),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_172),
.B(n_176),
.Y(n_194)
);

OAI21xp33_ASAP7_75t_L g173 ( 
.A1(n_154),
.A2(n_101),
.B(n_132),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_173),
.A2(n_179),
.B(n_180),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_149),
.A2(n_124),
.B1(n_123),
.B2(n_144),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_186),
.B1(n_162),
.B2(n_161),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_149),
.A2(n_99),
.B(n_130),
.Y(n_179)
);

OAI322xp33_ASAP7_75t_L g181 ( 
.A1(n_156),
.A2(n_96),
.A3(n_111),
.B1(n_126),
.B2(n_129),
.C1(n_112),
.C2(n_109),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_181),
.B(n_189),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_67),
.Y(n_183)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_183),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_184),
.A2(n_148),
.B1(n_152),
.B2(n_159),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_158),
.A2(n_164),
.B1(n_168),
.B2(n_163),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_147),
.C(n_148),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_147),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_162),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_188),
.B(n_160),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_150),
.B(n_151),
.Y(n_189)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_193),
.B(n_175),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_189),
.C(n_175),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_188),
.B(n_178),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_198),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_197),
.A2(n_201),
.B1(n_190),
.B2(n_203),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_185),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_152),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_200),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_183),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_174),
.A2(n_155),
.B1(n_159),
.B2(n_179),
.Y(n_201)
);

INVxp67_ASAP7_75t_SL g202 ( 
.A(n_177),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_202),
.B(n_186),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_185),
.Y(n_205)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_205),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_187),
.C(n_172),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_208),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_182),
.Y(n_210)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_210),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_184),
.C(n_180),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_204),
.Y(n_225)
);

INVxp33_ASAP7_75t_SL g213 ( 
.A(n_200),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_213),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_215),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_216),
.A2(n_199),
.B1(n_196),
.B2(n_203),
.Y(n_217)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_209),
.B(n_191),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_222),
.B(n_218),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_204),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_225),
.Y(n_231)
);

NOR3xp33_ASAP7_75t_SL g226 ( 
.A(n_223),
.B(n_181),
.C(n_176),
.Y(n_226)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_226),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_207),
.C(n_213),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_230),
.Y(n_235)
);

OAI321xp33_ASAP7_75t_L g233 ( 
.A1(n_228),
.A2(n_229),
.A3(n_217),
.B1(n_219),
.B2(n_224),
.C(n_182),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_218),
.A2(n_212),
.B1(n_206),
.B2(n_192),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_192),
.C(n_171),
.Y(n_230)
);

AO21x1_ASAP7_75t_L g238 ( 
.A1(n_233),
.A2(n_237),
.B(n_236),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_231),
.A2(n_225),
.B(n_232),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_231),
.Y(n_240)
);

NOR2xp67_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_227),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_238),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_230),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_239),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_242),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_243),
.B(n_241),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_244),
.B(n_240),
.Y(n_245)
);


endmodule