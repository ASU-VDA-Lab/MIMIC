module real_aes_9468_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_900, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_900;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_887;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_892;
wire n_528;
wire n_372;
wire n_202;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_875;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_733;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_880;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_869;
wire n_613;
wire n_642;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_898;
wire n_115;
wire n_604;
wire n_110;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_0), .A2(n_84), .B1(n_532), .B2(n_533), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_1), .B(n_202), .Y(n_584) );
AOI22x1_ASAP7_75t_SL g866 ( .A1(n_2), .A2(n_72), .B1(n_867), .B2(n_868), .Y(n_866) );
INVx1_ASAP7_75t_L g867 ( .A(n_2), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_3), .A2(n_102), .B1(n_887), .B2(n_898), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_4), .B(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_5), .B(n_143), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g588 ( .A(n_6), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_7), .A2(n_39), .B1(n_174), .B2(n_530), .Y(n_645) );
NOR2xp67_ASAP7_75t_L g112 ( .A(n_8), .B(n_86), .Y(n_112) );
INVx1_ASAP7_75t_L g892 ( .A(n_8), .Y(n_892) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_9), .B(n_154), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_10), .B(n_135), .Y(n_162) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_11), .A2(n_62), .B1(n_174), .B2(n_213), .Y(n_543) );
NAND3xp33_ASAP7_75t_L g605 ( .A(n_12), .B(n_157), .C(n_174), .Y(n_605) );
NAND2x1p5_ASAP7_75t_L g238 ( .A(n_13), .B(n_135), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_14), .B(n_193), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g582 ( .A(n_15), .Y(n_582) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_16), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_17), .B(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_18), .B(n_147), .Y(n_569) );
AND2x2_ASAP7_75t_L g212 ( .A(n_19), .B(n_213), .Y(n_212) );
NAND3xp33_ASAP7_75t_L g602 ( .A(n_20), .B(n_150), .C(n_154), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_21), .A2(n_28), .B1(n_154), .B2(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_22), .B(n_571), .Y(n_619) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_23), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_24), .B(n_275), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_25), .B(n_201), .Y(n_200) );
NAND2xp33_ASAP7_75t_L g231 ( .A(n_26), .B(n_142), .Y(n_231) );
NAND2xp33_ASAP7_75t_L g155 ( .A(n_27), .B(n_142), .Y(n_155) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_29), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_30), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_31), .B(n_561), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g120 ( .A1(n_32), .A2(n_81), .B1(n_121), .B2(n_122), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_32), .Y(n_121) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_33), .A2(n_52), .B1(n_142), .B2(n_213), .Y(n_646) );
NAND2xp5_ASAP7_75t_SL g600 ( .A(n_34), .B(n_150), .Y(n_600) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_35), .B(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g111 ( .A(n_36), .Y(n_111) );
OAI21x1_ASAP7_75t_L g137 ( .A1(n_37), .A2(n_65), .B(n_138), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_38), .A2(n_176), .B(n_218), .C(n_219), .Y(n_217) );
NAND2xp33_ASAP7_75t_L g272 ( .A(n_40), .B(n_180), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g289 ( .A(n_41), .B(n_174), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_42), .Y(n_291) );
AND2x6_ASAP7_75t_L g160 ( .A(n_43), .B(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_L g545 ( .A(n_44), .B(n_275), .Y(n_545) );
NAND2x1p5_ASAP7_75t_L g606 ( .A(n_45), .B(n_275), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_46), .B(n_173), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_47), .B(n_153), .Y(n_152) );
NAND2xp33_ASAP7_75t_L g198 ( .A(n_48), .B(n_180), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_49), .B(n_147), .Y(n_621) );
INVx1_ASAP7_75t_L g161 ( .A(n_50), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_51), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_53), .B(n_180), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_54), .B(n_275), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_55), .B(n_154), .Y(n_576) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_56), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_57), .B(n_154), .Y(n_559) );
NAND2x1_ASAP7_75t_L g625 ( .A(n_58), .B(n_275), .Y(n_625) );
AND2x2_ASAP7_75t_L g221 ( .A(n_59), .B(n_201), .Y(n_221) );
AND2x2_ASAP7_75t_L g895 ( .A(n_60), .B(n_896), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_61), .B(n_157), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_63), .B(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_64), .B(n_553), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_66), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g556 ( .A(n_67), .Y(n_556) );
NAND2xp33_ASAP7_75t_L g254 ( .A(n_68), .B(n_147), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_69), .B(n_157), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_70), .A2(n_75), .B1(n_154), .B2(n_530), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_71), .B(n_230), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g868 ( .A(n_72), .Y(n_868) );
CKINVDCx5p33_ASAP7_75t_R g592 ( .A(n_73), .Y(n_592) );
BUFx10_ASAP7_75t_L g115 ( .A(n_74), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_76), .B(n_146), .Y(n_145) );
INVx1_ASAP7_75t_SL g536 ( .A(n_77), .Y(n_536) );
NAND2xp33_ASAP7_75t_L g259 ( .A(n_78), .B(n_154), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g882 ( .A(n_79), .Y(n_882) );
CKINVDCx5p33_ASAP7_75t_R g648 ( .A(n_80), .Y(n_648) );
INVx1_ASAP7_75t_L g122 ( .A(n_81), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_82), .B(n_142), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g624 ( .A(n_83), .Y(n_624) );
CKINVDCx5p33_ASAP7_75t_R g220 ( .A(n_85), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g891 ( .A(n_86), .B(n_892), .Y(n_891) );
INVx2_ASAP7_75t_L g138 ( .A(n_87), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_88), .B(n_157), .Y(n_604) );
OR2x2_ASAP7_75t_L g108 ( .A(n_89), .B(n_109), .Y(n_108) );
BUFx2_ASAP7_75t_L g875 ( .A(n_89), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_89), .B(n_110), .Y(n_886) );
INVx1_ASAP7_75t_L g897 ( .A(n_89), .Y(n_897) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_90), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_91), .B(n_180), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_92), .B(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_93), .B(n_237), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_94), .Y(n_191) );
INVx1_ASAP7_75t_L g896 ( .A(n_95), .Y(n_896) );
INVx1_ASAP7_75t_L g211 ( .A(n_96), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_97), .Y(n_172) );
AND2x2_ASAP7_75t_L g185 ( .A(n_98), .B(n_135), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_99), .B(n_183), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_100), .B(n_201), .Y(n_260) );
OR2x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_113), .Y(n_102) );
AOI21xp33_ASAP7_75t_L g116 ( .A1(n_103), .A2(n_117), .B(n_513), .Y(n_116) );
NOR2x1_ASAP7_75t_R g103 ( .A(n_104), .B(n_105), .Y(n_103) );
INVx5_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx4_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx5_ASAP7_75t_L g516 ( .A(n_107), .Y(n_516) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g874 ( .A(n_109), .B(n_875), .Y(n_874) );
AND2x4_ASAP7_75t_L g879 ( .A(n_109), .B(n_880), .Y(n_879) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x4_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
NOR3xp33_ASAP7_75t_L g893 ( .A(n_111), .B(n_894), .C(n_897), .Y(n_893) );
OAI21xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_116), .B(n_517), .Y(n_113) );
BUFx12f_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx6_ASAP7_75t_L g873 ( .A(n_115), .Y(n_873) );
INVx2_ASAP7_75t_SL g885 ( .A(n_115), .Y(n_885) );
OAI21xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_123), .B(n_511), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_120), .B(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
BUFx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g512 ( .A(n_125), .Y(n_512) );
NAND2x1p5_ASAP7_75t_L g125 ( .A(n_126), .B(n_428), .Y(n_125) );
AND5x1_ASAP7_75t_L g126 ( .A(n_127), .B(n_331), .C(n_370), .D(n_396), .E(n_411), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_128), .B(n_298), .Y(n_127) );
OAI221xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_222), .B1(n_239), .B2(n_249), .C(n_277), .Y(n_128) );
OR2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_163), .Y(n_129) );
INVx1_ASAP7_75t_L g395 ( .A(n_130), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_130), .B(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_130), .B(n_280), .Y(n_479) );
AOI322xp5_ASAP7_75t_L g492 ( .A1(n_130), .A2(n_361), .A3(n_414), .B1(n_493), .B2(n_495), .C1(n_496), .C2(n_499), .Y(n_492) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_L g380 ( .A(n_131), .B(n_247), .Y(n_380) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_132), .Y(n_248) );
INVx1_ASAP7_75t_L g315 ( .A(n_132), .Y(n_315) );
AND2x2_ASAP7_75t_L g320 ( .A(n_132), .B(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g330 ( .A(n_132), .B(n_244), .Y(n_330) );
AND2x2_ASAP7_75t_L g338 ( .A(n_132), .B(n_186), .Y(n_338) );
INVx1_ASAP7_75t_L g352 ( .A(n_132), .Y(n_352) );
OAI21x1_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_139), .B(n_162), .Y(n_132) );
OAI21x1_ASAP7_75t_L g265 ( .A1(n_133), .A2(n_266), .B(n_274), .Y(n_265) );
OAI21xp5_ASAP7_75t_L g294 ( .A1(n_133), .A2(n_266), .B(n_274), .Y(n_294) );
OAI21x1_ASAP7_75t_L g597 ( .A1(n_133), .A2(n_598), .B(n_606), .Y(n_597) );
OAI21x1_ASAP7_75t_L g656 ( .A1(n_133), .A2(n_598), .B(n_606), .Y(n_656) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g643 ( .A(n_134), .B(n_158), .Y(n_643) );
INVx3_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx4_ASAP7_75t_L g166 ( .A(n_135), .Y(n_166) );
BUFx4f_ASAP7_75t_L g188 ( .A(n_135), .Y(n_188) );
OA21x2_ASAP7_75t_L g251 ( .A1(n_135), .A2(n_252), .B(n_260), .Y(n_251) );
OA21x2_ASAP7_75t_L g297 ( .A1(n_135), .A2(n_252), .B(n_260), .Y(n_297) );
OA21x2_ASAP7_75t_L g302 ( .A1(n_135), .A2(n_252), .B(n_260), .Y(n_302) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_135), .Y(n_609) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g276 ( .A(n_136), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_136), .B(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g202 ( .A(n_137), .Y(n_202) );
OAI21x1_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_151), .B(n_158), .Y(n_139) );
AOI21xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_145), .B(n_148), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_142), .B(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g180 ( .A(n_143), .Y(n_180) );
INVx1_ASAP7_75t_L g237 ( .A(n_143), .Y(n_237) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_144), .Y(n_147) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_144), .Y(n_154) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_144), .Y(n_174) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_144), .Y(n_183) );
INVx1_ASAP7_75t_L g215 ( .A(n_144), .Y(n_215) );
INVx1_ASAP7_75t_L g288 ( .A(n_146), .Y(n_288) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g193 ( .A(n_147), .Y(n_193) );
INVx2_ASAP7_75t_L g256 ( .A(n_147), .Y(n_256) );
INVx2_ASAP7_75t_L g532 ( .A(n_147), .Y(n_532) );
INVx1_ASAP7_75t_L g575 ( .A(n_147), .Y(n_575) );
INVx2_ASAP7_75t_L g590 ( .A(n_147), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_147), .B(n_592), .Y(n_591) );
OAI21xp33_ASAP7_75t_L g177 ( .A1(n_148), .A2(n_178), .B(n_181), .Y(n_177) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_148), .A2(n_199), .B1(n_645), .B2(n_646), .Y(n_644) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_149), .Y(n_148) );
INVx3_ASAP7_75t_L g195 ( .A(n_149), .Y(n_195) );
BUFx2_ASAP7_75t_L g216 ( .A(n_149), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_149), .A2(n_271), .B(n_272), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_149), .A2(n_559), .B(n_560), .Y(n_558) );
AOI21x1_ASAP7_75t_L g620 ( .A1(n_149), .A2(n_621), .B(n_622), .Y(n_620) );
BUFx12f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx5_ASAP7_75t_L g157 ( .A(n_150), .Y(n_157) );
INVx5_ASAP7_75t_L g176 ( .A(n_150), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_L g286 ( .A1(n_150), .A2(n_287), .B(n_288), .C(n_289), .Y(n_286) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_150), .A2(n_573), .B1(n_574), .B2(n_576), .Y(n_572) );
OAI321xp33_ASAP7_75t_L g581 ( .A1(n_150), .A2(n_154), .A3(n_532), .B1(n_582), .B2(n_583), .C(n_584), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_155), .B(n_156), .Y(n_151) );
INVx2_ASAP7_75t_L g218 ( .A(n_153), .Y(n_218) );
INVx2_ASAP7_75t_SL g153 ( .A(n_154), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_154), .B(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g230 ( .A(n_154), .Y(n_230) );
INVx2_ASAP7_75t_L g235 ( .A(n_154), .Y(n_235) );
O2A1O1Ixp33_ASAP7_75t_L g555 ( .A1(n_154), .A2(n_157), .B(n_556), .C(n_557), .Y(n_555) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_157), .A2(n_258), .B(n_259), .Y(n_257) );
AOI21x1_ASAP7_75t_L g267 ( .A1(n_157), .A2(n_268), .B(n_269), .Y(n_267) );
OAI21xp5_ASAP7_75t_L g189 ( .A1(n_158), .A2(n_190), .B(n_196), .Y(n_189) );
OAI21x1_ASAP7_75t_L g227 ( .A1(n_158), .A2(n_228), .B(n_232), .Y(n_227) );
OAI21x1_ASAP7_75t_L g252 ( .A1(n_158), .A2(n_253), .B(n_257), .Y(n_252) );
OAI21x1_ASAP7_75t_L g285 ( .A1(n_158), .A2(n_286), .B(n_290), .Y(n_285) );
AO31x2_ASAP7_75t_L g527 ( .A1(n_158), .A2(n_166), .A3(n_528), .B(n_534), .Y(n_527) );
INVx8_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_159), .A2(n_168), .B(n_177), .Y(n_167) );
NOR2xp67_ASAP7_75t_L g206 ( .A(n_159), .B(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g540 ( .A(n_159), .Y(n_540) );
OAI21xp5_ASAP7_75t_L g593 ( .A1(n_159), .A2(n_584), .B(n_594), .Y(n_593) );
INVx8_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
BUFx2_ASAP7_75t_L g273 ( .A(n_160), .Y(n_273) );
INVx1_ASAP7_75t_L g563 ( .A(n_160), .Y(n_563) );
OAI21x1_ASAP7_75t_L g567 ( .A1(n_160), .A2(n_568), .B(n_572), .Y(n_567) );
OAI21x1_ASAP7_75t_L g598 ( .A1(n_160), .A2(n_599), .B(n_603), .Y(n_598) );
INVx1_ASAP7_75t_L g481 ( .A(n_163), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_164), .B(n_203), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_165), .B(n_186), .Y(n_164) );
INVx1_ASAP7_75t_L g319 ( .A(n_165), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_165), .B(n_352), .Y(n_351) );
INVx2_ASAP7_75t_SL g363 ( .A(n_165), .Y(n_363) );
AO21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_185), .Y(n_165) );
INVx3_ASAP7_75t_L g207 ( .A(n_166), .Y(n_207) );
AO21x2_ASAP7_75t_L g244 ( .A1(n_166), .A2(n_167), .B(n_185), .Y(n_244) );
OAI21xp5_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_171), .B(n_175), .Y(n_168) );
NOR2xp67_ASAP7_75t_L g171 ( .A(n_172), .B(n_173), .Y(n_171) );
INVx5_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_SL g175 ( .A(n_176), .Y(n_175) );
CKINVDCx6p67_ASAP7_75t_R g199 ( .A(n_176), .Y(n_199) );
AOI21x1_ASAP7_75t_L g568 ( .A1(n_176), .A2(n_569), .B(n_570), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_176), .A2(n_586), .B(n_591), .Y(n_585) );
AOI21x1_ASAP7_75t_L g617 ( .A1(n_176), .A2(n_618), .B(n_619), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
NOR2xp33_ASAP7_75t_SL g181 ( .A(n_182), .B(n_184), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_182), .B(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g530 ( .A(n_183), .Y(n_530) );
INVx2_ASAP7_75t_L g561 ( .A(n_183), .Y(n_561) );
INVx2_ASAP7_75t_L g571 ( .A(n_183), .Y(n_571) );
OR2x2_ASAP7_75t_L g314 ( .A(n_186), .B(n_315), .Y(n_314) );
BUFx3_ASAP7_75t_L g368 ( .A(n_186), .Y(n_368) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g247 ( .A(n_187), .Y(n_247) );
AND2x2_ASAP7_75t_L g345 ( .A(n_187), .B(n_244), .Y(n_345) );
OA21x2_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_200), .Y(n_187) );
OAI21x1_ASAP7_75t_L g226 ( .A1(n_188), .A2(n_227), .B(n_238), .Y(n_226) );
OAI21x1_ASAP7_75t_L g284 ( .A1(n_188), .A2(n_285), .B(n_293), .Y(n_284) );
OAI21x1_ASAP7_75t_L g307 ( .A1(n_188), .A2(n_285), .B(n_293), .Y(n_307) );
OA21x2_ASAP7_75t_L g326 ( .A1(n_188), .A2(n_227), .B(n_238), .Y(n_326) );
O2A1O1Ixp5_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_194), .C(n_195), .Y(n_190) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
O2A1O1Ixp5_ASAP7_75t_L g232 ( .A1(n_195), .A2(n_233), .B(n_234), .C(n_236), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g290 ( .A1(n_195), .A2(n_234), .B(n_291), .C(n_292), .Y(n_290) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_195), .A2(n_199), .B1(n_529), .B2(n_531), .Y(n_528) );
OA22x2_ASAP7_75t_L g541 ( .A1(n_195), .A2(n_199), .B1(n_542), .B2(n_543), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B(n_199), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_199), .A2(n_229), .B(n_231), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_199), .A2(n_254), .B(n_255), .Y(n_253) );
INVx2_ASAP7_75t_L g539 ( .A(n_201), .Y(n_539) );
BUFx5_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g535 ( .A(n_202), .Y(n_535) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_202), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_203), .B(n_247), .Y(n_508) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVxp67_ASAP7_75t_SL g312 ( .A(n_204), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_204), .B(n_247), .Y(n_353) );
INVx1_ASAP7_75t_L g378 ( .A(n_204), .Y(n_378) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx2_ASAP7_75t_L g243 ( .A(n_205), .Y(n_243) );
AOI21x1_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_208), .B(n_221), .Y(n_205) );
OAI21x1_ASAP7_75t_L g566 ( .A1(n_207), .A2(n_567), .B(n_577), .Y(n_566) );
OAI21x1_ASAP7_75t_L g615 ( .A1(n_207), .A2(n_616), .B(n_625), .Y(n_615) );
OAI21x1_ASAP7_75t_L g672 ( .A1(n_207), .A2(n_616), .B(n_625), .Y(n_672) );
OAI21x1_ASAP7_75t_L g707 ( .A1(n_207), .A2(n_567), .B(n_577), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_209), .B(n_217), .Y(n_208) );
OAI21x1_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_212), .B(n_216), .Y(n_209) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g533 ( .A(n_215), .Y(n_533) );
OAI21xp5_ASAP7_75t_L g603 ( .A1(n_218), .A2(n_604), .B(n_605), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_222), .A2(n_465), .B1(n_468), .B2(n_469), .Y(n_464) );
INVx1_ASAP7_75t_L g468 ( .A(n_222), .Y(n_468) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
NAND2x1_ASAP7_75t_L g348 ( .A(n_223), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
OR2x2_ASAP7_75t_L g296 ( .A(n_224), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g336 ( .A(n_224), .B(n_297), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_224), .B(n_325), .Y(n_374) );
OR2x2_ASAP7_75t_L g426 ( .A(n_224), .B(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g308 ( .A(n_225), .B(n_264), .Y(n_308) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g263 ( .A(n_226), .B(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x4_ASAP7_75t_L g240 ( .A(n_241), .B(n_245), .Y(n_240) );
INVx1_ASAP7_75t_L g420 ( .A(n_241), .Y(n_420) );
NAND2xp67_ASAP7_75t_L g451 ( .A(n_241), .B(n_338), .Y(n_451) );
INVx1_ASAP7_75t_L g494 ( .A(n_241), .Y(n_494) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_244), .Y(n_241) );
INVx1_ASAP7_75t_L g329 ( .A(n_242), .Y(n_329) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g280 ( .A(n_243), .B(n_244), .Y(n_280) );
INVx1_ASAP7_75t_L g321 ( .A(n_243), .Y(n_321) );
AND2x2_ASAP7_75t_L g362 ( .A(n_243), .B(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g382 ( .A(n_246), .B(n_279), .Y(n_382) );
OR2x2_ASAP7_75t_L g410 ( .A(n_246), .B(n_311), .Y(n_410) );
OR2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
INVx2_ASAP7_75t_L g387 ( .A(n_247), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_247), .B(n_319), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_261), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_250), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g367 ( .A(n_250), .B(n_368), .Y(n_367) );
NAND4xp25_ASAP7_75t_L g394 ( .A(n_250), .B(n_311), .C(n_317), .D(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g412 ( .A(n_250), .B(n_304), .Y(n_412) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g323 ( .A(n_251), .Y(n_323) );
AND2x2_ASAP7_75t_L g504 ( .A(n_251), .B(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g448 ( .A(n_261), .Y(n_448) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g317 ( .A(n_263), .B(n_305), .Y(n_317) );
BUFx2_ASAP7_75t_L g342 ( .A(n_263), .Y(n_342) );
AND2x2_ASAP7_75t_SL g443 ( .A(n_263), .B(n_403), .Y(n_443) );
INVx2_ASAP7_75t_L g325 ( .A(n_264), .Y(n_325) );
OR2x2_ASAP7_75t_L g439 ( .A(n_264), .B(n_284), .Y(n_439) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
OAI21x1_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_270), .B(n_273), .Y(n_266) );
OAI21x1_ASAP7_75t_L g616 ( .A1(n_273), .A2(n_617), .B(n_620), .Y(n_616) );
INVx3_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_281), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_278), .B(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_280), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g397 ( .A(n_280), .B(n_313), .Y(n_397) );
AND2x2_ASAP7_75t_L g490 ( .A(n_280), .B(n_466), .Y(n_490) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_295), .Y(n_281) );
INVx2_ASAP7_75t_L g497 ( .A(n_282), .Y(n_497) );
BUFx3_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_283), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_294), .Y(n_283) );
INVx1_ASAP7_75t_L g341 ( .A(n_284), .Y(n_341) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp33_ASAP7_75t_R g385 ( .A(n_296), .B(n_340), .Y(n_385) );
INVx1_ASAP7_75t_L g484 ( .A(n_296), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_297), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g391 ( .A(n_297), .Y(n_391) );
OAI21xp33_ASAP7_75t_SL g298 ( .A1(n_299), .A2(n_309), .B(n_316), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
O2A1O1Ixp5_ASAP7_75t_L g370 ( .A1(n_300), .A2(n_371), .B(n_375), .C(n_381), .Y(n_370) );
NOR2x1p5_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
INVx1_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g347 ( .A(n_302), .Y(n_347) );
BUFx2_ASAP7_75t_L g358 ( .A(n_302), .Y(n_358) );
INVx2_ASAP7_75t_SL g427 ( .A(n_302), .Y(n_427) );
INVx3_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_305), .B(n_308), .Y(n_304) );
AND2x4_ASAP7_75t_L g333 ( .A(n_305), .B(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g349 ( .A(n_307), .Y(n_349) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_307), .Y(n_373) );
AND2x2_ASAP7_75t_L g356 ( .A(n_308), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g503 ( .A(n_308), .Y(n_503) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_313), .Y(n_310) );
INVx1_ASAP7_75t_L g486 ( .A(n_311), .Y(n_486) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g407 ( .A(n_314), .Y(n_407) );
INVx1_ASAP7_75t_SL g417 ( .A(n_314), .Y(n_417) );
OR2x2_ASAP7_75t_L g453 ( .A(n_314), .B(n_377), .Y(n_453) );
OR2x2_ASAP7_75t_L g475 ( .A(n_314), .B(n_463), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_318), .B1(n_322), .B2(n_327), .Y(n_316) );
INVx2_ASAP7_75t_L g409 ( .A(n_317), .Y(n_409) );
INVx1_ASAP7_75t_L g359 ( .A(n_318), .Y(n_359) );
AND2x4_ASAP7_75t_L g441 ( .A(n_318), .B(n_387), .Y(n_441) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
BUFx2_ASAP7_75t_SL g470 ( .A(n_319), .Y(n_470) );
AND2x4_ASAP7_75t_L g344 ( .A(n_320), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g435 ( .A(n_320), .Y(n_435) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
OR2x6_ASAP7_75t_SL g438 ( .A(n_323), .B(n_439), .Y(n_438) );
OAI211xp5_ASAP7_75t_L g488 ( .A1(n_323), .A2(n_489), .B(n_492), .C(n_500), .Y(n_488) );
AND2x2_ASAP7_75t_L g495 ( .A(n_323), .B(n_443), .Y(n_495) );
INVx2_ASAP7_75t_L g404 ( .A(n_324), .Y(n_404) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVx2_ASAP7_75t_L g334 ( .A(n_325), .Y(n_334) );
INVx2_ASAP7_75t_L g392 ( .A(n_326), .Y(n_392) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx2_ASAP7_75t_L g413 ( .A(n_329), .Y(n_413) );
INVxp67_ASAP7_75t_SL g369 ( .A(n_330), .Y(n_369) );
INVx2_ASAP7_75t_L g388 ( .A(n_330), .Y(n_388) );
OR2x2_ASAP7_75t_L g445 ( .A(n_330), .B(n_378), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_332), .B(n_354), .Y(n_331) );
OAI332xp33_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_335), .A3(n_337), .B1(n_339), .B2(n_342), .B3(n_343), .C1(n_346), .C2(n_350), .Y(n_332) );
INVx2_ASAP7_75t_L g405 ( .A(n_333), .Y(n_405) );
AND2x4_ASAP7_75t_SL g365 ( .A(n_334), .B(n_349), .Y(n_365) );
BUFx2_ASAP7_75t_L g472 ( .A(n_334), .Y(n_472) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OAI311xp33_ASAP7_75t_L g381 ( .A1(n_336), .A2(n_382), .A3(n_383), .B1(n_384), .C1(n_394), .Y(n_381) );
AND2x2_ASAP7_75t_L g398 ( .A(n_336), .B(n_399), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_337), .A2(n_401), .B1(n_405), .B2(n_406), .Y(n_400) );
AND2x4_ASAP7_75t_L g361 ( .A(n_338), .B(n_362), .Y(n_361) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
BUFx2_ASAP7_75t_L g403 ( .A(n_341), .Y(n_403) );
NAND3xp33_ASAP7_75t_L g366 ( .A(n_342), .B(n_367), .C(n_369), .Y(n_366) );
AOI22xp33_ASAP7_75t_SL g442 ( .A1(n_342), .A2(n_393), .B1(n_443), .B2(n_444), .Y(n_442) );
INVx2_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
OR2x2_ASAP7_75t_L g437 ( .A(n_347), .B(n_404), .Y(n_437) );
BUFx2_ASAP7_75t_L g383 ( .A(n_349), .Y(n_383) );
INVx1_ASAP7_75t_L g399 ( .A(n_349), .Y(n_399) );
OR2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
OR2x2_ASAP7_75t_L g510 ( .A(n_351), .B(n_508), .Y(n_510) );
INVx1_ASAP7_75t_L g467 ( .A(n_352), .Y(n_467) );
INVx1_ASAP7_75t_L g423 ( .A(n_353), .Y(n_423) );
OAI221xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_359), .B1(n_360), .B2(n_364), .C(n_366), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g393 ( .A(n_362), .B(n_368), .Y(n_393) );
AND2x2_ASAP7_75t_L g416 ( .A(n_362), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g476 ( .A(n_362), .Y(n_476) );
INVx2_ASAP7_75t_L g449 ( .A(n_365), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_365), .A2(n_472), .B1(n_490), .B2(n_491), .Y(n_489) );
AND2x2_ASAP7_75t_L g506 ( .A(n_369), .B(n_507), .Y(n_506) );
INVx2_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
INVxp67_ASAP7_75t_SL g425 ( .A(n_373), .Y(n_425) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_373), .Y(n_483) );
INVx1_ASAP7_75t_L g505 ( .A(n_374), .Y(n_505) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_379), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_386), .B1(n_389), .B2(n_393), .Y(n_384) );
INVx3_ASAP7_75t_L g487 ( .A(n_386), .Y(n_487) );
AND2x4_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
AOI321xp33_ASAP7_75t_L g411 ( .A1(n_387), .A2(n_412), .A3(n_413), .B1(n_414), .B2(n_416), .C(n_418), .Y(n_411) );
OR2x2_ASAP7_75t_L g419 ( .A(n_387), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g460 ( .A(n_387), .B(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g422 ( .A(n_388), .B(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g415 ( .A(n_390), .Y(n_415) );
INVxp67_ASAP7_75t_SL g458 ( .A(n_390), .Y(n_458) );
NAND2x1p5_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
AOI211xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_398), .B(n_400), .C(n_408), .Y(n_396) );
AOI222xp33_ASAP7_75t_L g500 ( .A1(n_397), .A2(n_501), .B1(n_504), .B2(n_506), .C1(n_509), .C2(n_900), .Y(n_500) );
NAND2x1_ASAP7_75t_L g440 ( .A(n_398), .B(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g414 ( .A(n_399), .B(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_404), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OAI32xp33_ASAP7_75t_L g485 ( .A1(n_404), .A2(n_439), .A3(n_475), .B1(n_486), .B2(n_487), .Y(n_485) );
NOR2xp67_ASAP7_75t_SL g408 ( .A(n_409), .B(n_410), .Y(n_408) );
INVx1_ASAP7_75t_L g499 ( .A(n_410), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_413), .B(n_466), .Y(n_465) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_415), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_421), .B(n_424), .Y(n_418) );
INVx1_ASAP7_75t_L g491 ( .A(n_419), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g452 ( .A1(n_421), .A2(n_453), .B1(n_454), .B2(n_457), .Y(n_452) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OR2x2_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
INVx1_ASAP7_75t_L g456 ( .A(n_426), .Y(n_456) );
INVx1_ASAP7_75t_L g463 ( .A(n_427), .Y(n_463) );
NOR2x1_ASAP7_75t_L g428 ( .A(n_429), .B(n_488), .Y(n_428) );
NAND4xp75_ASAP7_75t_L g429 ( .A(n_430), .B(n_446), .C(n_459), .D(n_477), .Y(n_429) );
AND3x1_ASAP7_75t_L g430 ( .A(n_431), .B(n_440), .C(n_442), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_436), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
NAND2xp33_ASAP7_75t_SL g436 ( .A(n_437), .B(n_438), .Y(n_436) );
INVx2_ASAP7_75t_L g455 ( .A(n_439), .Y(n_455) );
OR2x2_ASAP7_75t_L g462 ( .A(n_439), .B(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_450), .B(n_452), .Y(n_446) );
NAND2xp33_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NAND2x1_ASAP7_75t_SL g454 ( .A(n_455), .B(n_456), .Y(n_454) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AOI21x1_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_464), .B(n_471), .Y(n_459) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NOR2x1_ASAP7_75t_L g471 ( .A(n_472), .B(n_473), .Y(n_471) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NOR2x1_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_482), .B(n_485), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AND2x4_ASAP7_75t_L g482 ( .A(n_483), .B(n_484), .Y(n_482) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
BUFx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
XNOR2xp5_ASAP7_75t_L g877 ( .A(n_512), .B(n_866), .Y(n_877) );
BUFx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
BUFx3_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx6_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AOI221xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_869), .B1(n_876), .B2(n_878), .C(n_881), .Y(n_517) );
XNOR2x1_ASAP7_75t_L g518 ( .A(n_519), .B(n_866), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
NOR2x1_ASAP7_75t_L g520 ( .A(n_521), .B(n_771), .Y(n_520) );
NAND4xp25_ASAP7_75t_L g521 ( .A(n_522), .B(n_675), .C(n_722), .D(n_759), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_612), .B(n_626), .Y(n_522) );
AO22x1_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_564), .B1(n_595), .B2(n_611), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_546), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_525), .B(n_547), .Y(n_688) );
AND2x2_ASAP7_75t_L g791 ( .A(n_525), .B(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g742 ( .A(n_526), .B(n_743), .Y(n_742) );
INVxp67_ASAP7_75t_L g827 ( .A(n_526), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_537), .Y(n_526) );
AND2x2_ASAP7_75t_L g607 ( .A(n_527), .B(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g633 ( .A(n_527), .Y(n_633) );
INVx1_ASAP7_75t_L g654 ( .A(n_527), .Y(n_654) );
INVx1_ASAP7_75t_L g684 ( .A(n_527), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
INVx1_ASAP7_75t_L g553 ( .A(n_535), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_535), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g682 ( .A(n_537), .Y(n_682) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_537), .Y(n_700) );
INVx1_ASAP7_75t_L g727 ( .A(n_537), .Y(n_727) );
INVxp67_ASAP7_75t_SL g757 ( .A(n_537), .Y(n_757) );
INVx1_ASAP7_75t_L g806 ( .A(n_537), .Y(n_806) );
OAI21x1_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_541), .B(n_544), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
OA21x2_ASAP7_75t_L g608 ( .A1(n_541), .A2(n_609), .B(n_610), .Y(n_608) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVxp67_ASAP7_75t_L g610 ( .A(n_545), .Y(n_610) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g822 ( .A(n_547), .B(n_607), .Y(n_822) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
NOR2xp67_ASAP7_75t_L g653 ( .A(n_548), .B(n_654), .Y(n_653) );
NAND3xp33_ASAP7_75t_L g801 ( .A(n_548), .B(n_726), .C(n_802), .Y(n_801) );
AND2x2_ASAP7_75t_L g805 ( .A(n_548), .B(n_806), .Y(n_805) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g629 ( .A(n_549), .B(n_608), .Y(n_629) );
AND2x2_ASAP7_75t_L g728 ( .A(n_549), .B(n_692), .Y(n_728) );
AND2x2_ASAP7_75t_L g736 ( .A(n_549), .B(n_654), .Y(n_736) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g686 ( .A(n_550), .B(n_597), .Y(n_686) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g660 ( .A(n_551), .Y(n_660) );
AND2x2_ASAP7_75t_L g770 ( .A(n_551), .B(n_597), .Y(n_770) );
NAND2x1p5_ASAP7_75t_L g551 ( .A(n_552), .B(n_554), .Y(n_551) );
OAI21x1_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_558), .B(n_562), .Y(n_554) );
AND2x2_ASAP7_75t_L g763 ( .A(n_564), .B(n_764), .Y(n_763) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_578), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_565), .B(n_673), .Y(n_678) );
INVx1_ASAP7_75t_L g746 ( .A(n_565), .Y(n_746) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g637 ( .A(n_566), .Y(n_637) );
INVxp67_ASAP7_75t_L g601 ( .A(n_571), .Y(n_601) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_575), .B(n_623), .Y(n_622) );
BUFx2_ASAP7_75t_L g611 ( .A(n_578), .Y(n_611) );
AND2x4_ASAP7_75t_L g788 ( .A(n_578), .B(n_733), .Y(n_788) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_579), .B(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g740 ( .A(n_579), .B(n_672), .Y(n_740) );
AND2x2_ASAP7_75t_L g854 ( .A(n_579), .B(n_749), .Y(n_854) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g640 ( .A(n_580), .B(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g651 ( .A(n_580), .Y(n_651) );
OAI21x1_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_585), .B(n_593), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AOI32xp33_ASAP7_75t_L g663 ( .A1(n_595), .A2(n_657), .A3(n_664), .B1(n_665), .B2(n_668), .Y(n_663) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_607), .Y(n_595) );
NOR2xp67_ASAP7_75t_L g630 ( .A(n_596), .B(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g658 ( .A(n_596), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_596), .B(n_684), .Y(n_721) );
OAI32xp33_ASAP7_75t_L g773 ( .A1(n_596), .A2(n_681), .A3(n_774), .B1(n_777), .B2(n_779), .Y(n_773) );
NOR3xp33_ASAP7_75t_L g808 ( .A(n_596), .B(n_674), .C(n_809), .Y(n_808) );
BUFx3_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OAI21xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_601), .B(n_602), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_607), .B(n_758), .Y(n_863) );
AND2x2_ASAP7_75t_L g655 ( .A(n_608), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g664 ( .A(n_611), .Y(n_664) );
INVx1_ASAP7_75t_L g832 ( .A(n_611), .Y(n_832) );
OR2x2_ASAP7_75t_L g859 ( .A(n_612), .B(n_775), .Y(n_859) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
OR2x2_ASAP7_75t_L g635 ( .A(n_613), .B(n_636), .Y(n_635) );
BUFx2_ASAP7_75t_L g679 ( .A(n_613), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_613), .B(n_636), .Y(n_776) );
AND2x2_ASAP7_75t_L g798 ( .A(n_613), .B(n_699), .Y(n_798) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g662 ( .A(n_614), .B(n_641), .Y(n_662) );
HB1xp67_ASAP7_75t_L g852 ( .A(n_614), .Y(n_852) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g714 ( .A(n_615), .Y(n_714) );
INVx4_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_663), .Y(n_626) );
AOI322xp5_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_634), .A3(n_638), .B1(n_649), .B2(n_652), .C1(n_657), .C2(n_661), .Y(n_627) );
AND2x4_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
INVx2_ASAP7_75t_L g720 ( .A(n_629), .Y(n_720) );
AND2x2_ASAP7_75t_L g847 ( .A(n_629), .B(n_691), .Y(n_847) );
INVxp67_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g836 ( .A(n_632), .B(n_660), .Y(n_836) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AND2x4_ASAP7_75t_L g659 ( .A(n_633), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g691 ( .A(n_633), .B(n_692), .Y(n_691) );
INVx2_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_635), .B(n_662), .Y(n_661) );
OR2x2_ASAP7_75t_L g650 ( .A(n_636), .B(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g840 ( .A(n_636), .B(n_745), .Y(n_840) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_SL g674 ( .A(n_637), .Y(n_674) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_639), .B(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g732 ( .A(n_640), .B(n_733), .Y(n_732) );
BUFx3_ASAP7_75t_L g796 ( .A(n_640), .Y(n_796) );
AND2x2_ASAP7_75t_L g817 ( .A(n_640), .B(n_734), .Y(n_817) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_641), .Y(n_667) );
INVx2_ASAP7_75t_L g673 ( .A(n_641), .Y(n_673) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g749 ( .A(n_642), .Y(n_749) );
AOI21x1_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_644), .B(n_647), .Y(n_642) );
AND2x2_ASAP7_75t_L g706 ( .A(n_651), .B(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g717 ( .A(n_651), .B(n_718), .Y(n_717) );
OR2x2_ASAP7_75t_L g775 ( .A(n_651), .B(n_749), .Y(n_775) );
INVxp67_ASAP7_75t_SL g790 ( .A(n_651), .Y(n_790) );
AND2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_655), .Y(n_652) );
INVx1_ASAP7_75t_L g767 ( .A(n_654), .Y(n_767) );
AND2x4_ASAP7_75t_L g835 ( .A(n_655), .B(n_836), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_655), .B(n_856), .Y(n_855) );
INVx2_ASAP7_75t_L g692 ( .A(n_656), .Y(n_692) );
AND2x4_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx2_ASAP7_75t_L g701 ( .A(n_659), .Y(n_701) );
AND2x2_ASAP7_75t_L g737 ( .A(n_659), .B(n_727), .Y(n_737) );
BUFx2_ASAP7_75t_L g800 ( .A(n_659), .Y(n_800) );
INVx1_ASAP7_75t_L g857 ( .A(n_659), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_660), .B(n_692), .Y(n_743) );
INVx2_ASAP7_75t_L g694 ( .A(n_662), .Y(n_694) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OAI221xp5_ASAP7_75t_L g804 ( .A1(n_666), .A2(n_736), .B1(n_805), .B2(n_807), .C(n_808), .Y(n_804) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_667), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g807 ( .A(n_667), .Y(n_807) );
INVx1_ASAP7_75t_L g696 ( .A(n_668), .Y(n_696) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_670), .B(n_674), .Y(n_669) );
INVx2_ASAP7_75t_L g781 ( .A(n_670), .Y(n_781) );
AND2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_673), .Y(n_670) );
INVx2_ASAP7_75t_L g709 ( .A(n_671), .Y(n_709) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g710 ( .A(n_673), .Y(n_710) );
HB1xp67_ASAP7_75t_L g739 ( .A(n_673), .Y(n_739) );
AND2x2_ASAP7_75t_L g693 ( .A(n_674), .B(n_694), .Y(n_693) );
AND2x4_ASAP7_75t_L g729 ( .A(n_674), .B(n_708), .Y(n_729) );
AND2x2_ASAP7_75t_L g813 ( .A(n_674), .B(n_716), .Y(n_813) );
AOI221xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_680), .B1(n_687), .B2(n_693), .C(n_695), .Y(n_675) );
INVx2_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
OR2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g789 ( .A(n_678), .B(n_790), .Y(n_789) );
AND2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_683), .Y(n_680) );
OR2x2_ASAP7_75t_L g689 ( .A(n_681), .B(n_690), .Y(n_689) );
OR2x2_ASAP7_75t_L g777 ( .A(n_681), .B(n_778), .Y(n_777) );
INVx2_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g735 ( .A(n_682), .B(n_736), .Y(n_735) );
NOR2x1_ASAP7_75t_L g831 ( .A(n_682), .B(n_767), .Y(n_831) );
NOR2x1_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
INVx1_ASAP7_75t_L g703 ( .A(n_684), .Y(n_703) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_684), .Y(n_724) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g750 ( .A(n_686), .B(n_727), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
NOR2x1p5_ASAP7_75t_L g837 ( .A(n_690), .B(n_838), .Y(n_837) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g699 ( .A(n_692), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_694), .B(n_706), .Y(n_825) );
OAI221xp5_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_697), .B1(n_702), .B2(n_704), .C(n_711), .Y(n_695) );
OAI222xp33_ASAP7_75t_L g860 ( .A1(n_697), .A2(n_762), .B1(n_861), .B2(n_862), .C1(n_863), .C2(n_864), .Y(n_860) );
OR2x2_ASAP7_75t_L g697 ( .A(n_698), .B(n_701), .Y(n_697) );
OR2x2_ASAP7_75t_L g702 ( .A(n_698), .B(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
OR2x6_ASAP7_75t_L g845 ( .A(n_701), .B(n_806), .Y(n_845) );
INVx2_ASAP7_75t_L g818 ( .A(n_702), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_705), .B(n_708), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g760 ( .A(n_705), .B(n_761), .Y(n_760) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g718 ( .A(n_707), .Y(n_718) );
INVx2_ASAP7_75t_L g734 ( .A(n_707), .Y(n_734) );
INVx1_ASAP7_75t_L g762 ( .A(n_708), .Y(n_762) );
AND2x2_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
INVx2_ASAP7_75t_L g716 ( .A(n_709), .Y(n_716) );
HB1xp67_ASAP7_75t_L g764 ( .A(n_709), .Y(n_764) );
AND2x2_ASAP7_75t_L g829 ( .A(n_709), .B(n_728), .Y(n_829) );
AND2x2_ASAP7_75t_L g745 ( .A(n_710), .B(n_714), .Y(n_745) );
OAI21xp33_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_715), .B(n_719), .Y(n_711) );
BUFx2_ASAP7_75t_L g803 ( .A(n_714), .Y(n_803) );
INVxp67_ASAP7_75t_SL g865 ( .A(n_714), .Y(n_865) );
AND2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
AND2x2_ASAP7_75t_L g747 ( .A(n_717), .B(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g780 ( .A(n_717), .Y(n_780) );
NOR2x1p5_ASAP7_75t_SL g719 ( .A(n_720), .B(n_721), .Y(n_719) );
AOI211xp5_ASAP7_75t_SL g722 ( .A1(n_723), .A2(n_729), .B(n_730), .C(n_751), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
INVx2_ASAP7_75t_L g816 ( .A(n_725), .Y(n_816) );
AND2x2_ASAP7_75t_L g725 ( .A(n_726), .B(n_728), .Y(n_725) );
AO22x1_ASAP7_75t_L g830 ( .A1(n_726), .A2(n_831), .B1(n_832), .B2(n_833), .Y(n_830) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g778 ( .A(n_728), .Y(n_778) );
AND2x2_ASAP7_75t_L g841 ( .A(n_728), .B(n_827), .Y(n_841) );
INVx1_ASAP7_75t_L g753 ( .A(n_729), .Y(n_753) );
NAND2xp33_ASAP7_75t_L g730 ( .A(n_731), .B(n_741), .Y(n_730) );
AOI22xp5_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_735), .B1(n_737), .B2(n_738), .Y(n_731) );
INVx2_ASAP7_75t_SL g752 ( .A(n_732), .Y(n_752) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g858 ( .A(n_735), .Y(n_858) );
AND2x2_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
INVx1_ASAP7_75t_L g809 ( .A(n_740), .Y(n_809) );
AOI32xp33_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_744), .A3(n_746), .B1(n_747), .B2(n_750), .Y(n_741) );
INVx1_ASAP7_75t_L g758 ( .A(n_743), .Y(n_758) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
BUFx2_ASAP7_75t_L g784 ( .A(n_745), .Y(n_784) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g815 ( .A(n_750), .Y(n_815) );
AOI21xp33_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_753), .B(n_754), .Y(n_751) );
OAI321xp33_ASAP7_75t_L g794 ( .A1(n_752), .A2(n_795), .A3(n_797), .B1(n_799), .B2(n_801), .C(n_804), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_755), .B(n_758), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
NAND2x1p5_ASAP7_75t_L g769 ( .A(n_756), .B(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
OAI21xp33_ASAP7_75t_L g759 ( .A1(n_760), .A2(n_763), .B(n_765), .Y(n_759) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
AND2x4_ASAP7_75t_L g765 ( .A(n_766), .B(n_768), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx2_ASAP7_75t_L g793 ( .A(n_770), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_772), .B(n_819), .Y(n_771) );
NOR4xp25_ASAP7_75t_L g772 ( .A(n_773), .B(n_782), .C(n_794), .D(n_810), .Y(n_772) );
OR2x2_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
INVx2_ASAP7_75t_L g812 ( .A(n_775), .Y(n_812) );
OR2x2_ASAP7_75t_L g779 ( .A(n_780), .B(n_781), .Y(n_779) );
INVx2_ASAP7_75t_L g833 ( .A(n_780), .Y(n_833) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
A2O1A1Ixp33_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_785), .B(n_789), .C(n_791), .Y(n_783) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
OAI21xp33_ASAP7_75t_L g839 ( .A1(n_786), .A2(n_840), .B(n_841), .Y(n_839) );
INVx2_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx4_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
OAI21xp33_ASAP7_75t_L g844 ( .A1(n_795), .A2(n_845), .B(n_846), .Y(n_844) );
INVx2_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_796), .B(n_865), .Y(n_864) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
AND2x2_ASAP7_75t_L g823 ( .A(n_802), .B(n_817), .Y(n_823) );
INVxp67_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx2_ASAP7_75t_L g838 ( .A(n_805), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_807), .A2(n_812), .B1(n_835), .B2(n_837), .Y(n_834) );
AO22x1_ASAP7_75t_L g810 ( .A1(n_811), .A2(n_814), .B1(n_817), .B2(n_818), .Y(n_810) );
AND2x2_ASAP7_75t_L g811 ( .A(n_812), .B(n_813), .Y(n_811) );
INVx1_ASAP7_75t_L g862 ( .A(n_812), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_815), .B(n_816), .Y(n_814) );
NOR3xp33_ASAP7_75t_L g819 ( .A(n_820), .B(n_842), .C(n_860), .Y(n_819) );
NAND4xp25_ASAP7_75t_L g820 ( .A(n_821), .B(n_828), .C(n_834), .D(n_839), .Y(n_820) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_822), .A2(n_823), .B1(n_824), .B2(n_826), .Y(n_821) );
INVxp67_ASAP7_75t_SL g824 ( .A(n_825), .Y(n_824) );
BUFx2_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_829), .B(n_830), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_840), .B(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g861 ( .A(n_841), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_843), .B(n_848), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
OAI22xp33_ASAP7_75t_L g849 ( .A1(n_850), .A2(n_855), .B1(n_858), .B2(n_859), .Y(n_849) );
OR2x2_ASAP7_75t_L g850 ( .A(n_851), .B(n_853), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx2_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx4_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx3_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
AND2x6_ASAP7_75t_L g871 ( .A(n_872), .B(n_874), .Y(n_871) );
AND2x2_ASAP7_75t_SL g878 ( .A(n_872), .B(n_879), .Y(n_878) );
INVx1_ASAP7_75t_SL g872 ( .A(n_873), .Y(n_872) );
CKINVDCx5p33_ASAP7_75t_R g880 ( .A(n_875), .Y(n_880) );
INVx1_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
NOR2xp33_ASAP7_75t_L g881 ( .A(n_882), .B(n_883), .Y(n_881) );
BUFx12f_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
OR2x2_ASAP7_75t_L g884 ( .A(n_885), .B(n_886), .Y(n_884) );
CKINVDCx14_ASAP7_75t_R g887 ( .A(n_888), .Y(n_887) );
CKINVDCx11_ASAP7_75t_R g888 ( .A(n_889), .Y(n_888) );
BUFx6f_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
INVx6_ASAP7_75t_SL g898 ( .A(n_890), .Y(n_898) );
AND2x4_ASAP7_75t_L g890 ( .A(n_891), .B(n_893), .Y(n_890) );
INVx4_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
endmodule