module fake_jpeg_20849_n_239 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_239);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_239;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_14),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_14),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_26),
.Y(n_63)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_26),
.B1(n_32),
.B2(n_17),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_17),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_53),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_48),
.B(n_49),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_42),
.B(n_16),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_26),
.B1(n_32),
.B2(n_29),
.Y(n_50)
);

AO22x1_ASAP7_75t_SL g91 ( 
.A1(n_50),
.A2(n_75),
.B1(n_79),
.B2(n_63),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_27),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_27),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_57),
.B(n_60),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_15),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_15),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_61),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_29),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_70),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_77),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_32),
.B1(n_28),
.B2(n_21),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_65),
.A2(n_79),
.B1(n_25),
.B2(n_2),
.Y(n_99)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_34),
.B(n_28),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_68),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_34),
.B(n_21),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_69),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_29),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_34),
.B(n_19),
.C(n_29),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_40),
.C(n_23),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_38),
.A2(n_23),
.B1(n_29),
.B2(n_18),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_72),
.A2(n_74),
.B1(n_41),
.B2(n_40),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_38),
.A2(n_23),
.B1(n_29),
.B2(n_18),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_34),
.B(n_19),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_76),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_40),
.B(n_30),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_41),
.A2(n_30),
.B1(n_25),
.B2(n_18),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_84),
.B(n_88),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_62),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_94),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_91),
.A2(n_99),
.B1(n_75),
.B2(n_73),
.Y(n_115)
);

BUFx4f_ASAP7_75t_SL g92 ( 
.A(n_78),
.Y(n_92)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_50),
.A2(n_25),
.B1(n_31),
.B2(n_24),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_95),
.B1(n_80),
.B2(n_55),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_40),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_63),
.A2(n_25),
.B1(n_31),
.B2(n_24),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_31),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_101),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_49),
.B(n_24),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_50),
.A2(n_19),
.B(n_3),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_102),
.A2(n_4),
.B(n_6),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_1),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_54),
.Y(n_121)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_50),
.B(n_1),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_105),
.A2(n_71),
.B1(n_66),
.B2(n_77),
.Y(n_110)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_52),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_88),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_91),
.A2(n_73),
.B1(n_65),
.B2(n_58),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_112),
.A2(n_115),
.B1(n_129),
.B2(n_132),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_48),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_116),
.B(n_121),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_96),
.A2(n_51),
.B1(n_75),
.B2(n_58),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_117),
.A2(n_133),
.B(n_134),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_90),
.A2(n_64),
.B(n_55),
.C(n_78),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_122),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_120),
.A2(n_126),
.B1(n_96),
.B2(n_91),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_67),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_67),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_124),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_67),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_86),
.B(n_56),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_125),
.B(n_127),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_51),
.B1(n_56),
.B2(n_78),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_87),
.B(n_94),
.Y(n_127)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

OAI32xp33_ASAP7_75t_L g129 ( 
.A1(n_95),
.A2(n_3),
.A3(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_54),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_136),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_99),
.A2(n_52),
.B1(n_54),
.B2(n_7),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_84),
.B(n_54),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_86),
.B(n_7),
.Y(n_135)
);

BUFx24_ASAP7_75t_SL g152 ( 
.A(n_135),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_87),
.B(n_8),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_8),
.C(n_9),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_101),
.C(n_82),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_97),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_145),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_154),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_147),
.A2(n_155),
.B1(n_131),
.B2(n_133),
.Y(n_170)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_97),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

NAND3xp33_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_98),
.C(n_102),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_115),
.A2(n_105),
.B1(n_88),
.B2(n_109),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_111),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_157),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_124),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_83),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_160),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_83),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_106),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_119),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_113),
.Y(n_163)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_163),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_170),
.A2(n_161),
.B1(n_155),
.B2(n_147),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_131),
.C(n_133),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_173),
.B(n_161),
.C(n_145),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_178),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_159),
.A2(n_131),
.B(n_127),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_176),
.B(n_141),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_159),
.A2(n_126),
.B(n_120),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_139),
.A2(n_134),
.B1(n_129),
.B2(n_118),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_177),
.A2(n_179),
.B1(n_141),
.B2(n_140),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_118),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_139),
.A2(n_110),
.B1(n_132),
.B2(n_88),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_150),
.B(n_107),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_162),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_189),
.C(n_181),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_195),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_153),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_186),
.Y(n_205)
);

AO21x1_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_145),
.B(n_150),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_172),
.B(n_156),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_187),
.B(n_188),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_142),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_151),
.C(n_157),
.Y(n_189)
);

AOI322xp5_ASAP7_75t_L g202 ( 
.A1(n_190),
.A2(n_165),
.A3(n_144),
.B1(n_146),
.B2(n_85),
.C1(n_92),
.C2(n_163),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_191),
.A2(n_170),
.B1(n_176),
.B2(n_175),
.Y(n_197)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_192),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_142),
.Y(n_193)
);

NOR3xp33_ASAP7_75t_SL g207 ( 
.A(n_193),
.B(n_196),
.C(n_163),
.Y(n_207)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_171),
.Y(n_194)
);

OAI322xp33_ASAP7_75t_L g201 ( 
.A1(n_194),
.A2(n_144),
.A3(n_180),
.B1(n_85),
.B2(n_152),
.C1(n_116),
.C2(n_171),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_167),
.B(n_169),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_104),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_192),
.C(n_184),
.Y(n_210)
);

OAI321xp33_ASAP7_75t_L g200 ( 
.A1(n_182),
.A2(n_180),
.A3(n_172),
.B1(n_179),
.B2(n_169),
.C(n_164),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_200),
.A2(n_202),
.B1(n_9),
.B2(n_10),
.Y(n_217)
);

AOI31xp67_ASAP7_75t_L g216 ( 
.A1(n_201),
.A2(n_81),
.A3(n_10),
.B(n_11),
.Y(n_216)
);

A2O1A1Ixp33_ASAP7_75t_L g203 ( 
.A1(n_186),
.A2(n_182),
.B(n_195),
.C(n_185),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_191),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_165),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_189),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_198),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_213),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_212),
.B(n_216),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_92),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_113),
.C(n_108),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_217),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_215),
.A2(n_203),
.B(n_206),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_213),
.A2(n_197),
.B1(n_205),
.B2(n_198),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_220),
.A2(n_223),
.B1(n_224),
.B2(n_208),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_210),
.C(n_11),
.Y(n_228)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_211),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_225),
.B(n_226),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_222),
.A2(n_205),
.B(n_209),
.Y(n_226)
);

OAI21x1_ASAP7_75t_L g227 ( 
.A1(n_220),
.A2(n_207),
.B(n_214),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_229),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_219),
.C(n_221),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_218),
.A2(n_10),
.B(n_12),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_228),
.B(n_219),
.Y(n_230)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_230),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_12),
.C(n_13),
.Y(n_236)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_231),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_235),
.B(n_236),
.Y(n_237)
);

AO21x1_ASAP7_75t_L g238 ( 
.A1(n_234),
.A2(n_232),
.B(n_13),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_238),
.B(n_237),
.Y(n_239)
);


endmodule