module fake_jpeg_5481_n_104 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_104);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_9),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx4f_ASAP7_75t_SL g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_21),
.B(n_0),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_12),
.Y(n_45)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_31),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_30),
.A2(n_11),
.B1(n_20),
.B2(n_22),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_41),
.B1(n_22),
.B2(n_18),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_0),
.B1(n_1),
.B2(n_21),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_45),
.B(n_14),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_47),
.Y(n_72)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

INVxp67_ASAP7_75t_SL g68 ( 
.A(n_48),
.Y(n_68)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_53),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_50),
.A2(n_55),
.B1(n_58),
.B2(n_59),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_45),
.B(n_26),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_54),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_15),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_24),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_56),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_40),
.A2(n_27),
.B1(n_24),
.B2(n_12),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_57),
.A2(n_42),
.B1(n_44),
.B2(n_38),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_41),
.B(n_13),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_37),
.B(n_2),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_42),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_61),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_31),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_63),
.A2(n_25),
.B1(n_29),
.B2(n_31),
.Y(n_78)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

AND2x6_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_25),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_4),
.C(n_6),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_70),
.A2(n_58),
.B1(n_55),
.B2(n_53),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_73),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_69),
.A2(n_51),
.B1(n_49),
.B2(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_78),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_54),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_79),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_52),
.B1(n_38),
.B2(n_25),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_77),
.B(n_65),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_29),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_29),
.B1(n_6),
.B2(n_7),
.Y(n_80)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_81),
.A2(n_62),
.B(n_66),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_83),
.A2(n_66),
.B1(n_72),
.B2(n_78),
.Y(n_91)
);

AO21x1_ASAP7_75t_L g90 ( 
.A1(n_85),
.A2(n_64),
.B(n_72),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_74),
.B(n_79),
.C(n_68),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_88),
.B(n_86),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_87),
.A2(n_81),
.B1(n_76),
.B2(n_80),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_90),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_92),
.Y(n_94)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

XOR2x2_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_88),
.Y(n_98)
);

XNOR2x1_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_84),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_96),
.A2(n_89),
.B1(n_75),
.B2(n_67),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_85),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_98),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_93),
.C(n_8),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_100),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_9),
.Y(n_104)
);


endmodule