module fake_ariane_1089_n_796 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_796);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_796;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_784;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_166;
wire n_561;
wire n_770;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_780;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_617;
wire n_658;
wire n_616;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_742;
wire n_716;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_769;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_793;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_542;
wire n_548;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_791;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_531;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g158 ( 
.A(n_98),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_118),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_8),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_12),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_32),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_148),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_134),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_22),
.Y(n_166)
);

BUFx2_ASAP7_75t_SL g167 ( 
.A(n_82),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_52),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_85),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_39),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_88),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_142),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_33),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_35),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_155),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_67),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_153),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_12),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_116),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_79),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_47),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_133),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_77),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_126),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_110),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_10),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_101),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_119),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_121),
.Y(n_191)
);

BUFx8_ASAP7_75t_SL g192 ( 
.A(n_58),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_5),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_38),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_135),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_140),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_75),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_157),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_62),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_53),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_42),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_59),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_130),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_149),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_95),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_50),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_74),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_87),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_113),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_8),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_154),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_2),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_19),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_177),
.Y(n_214)
);

NOR2xp67_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_0),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_162),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_158),
.B(n_0),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g218 ( 
.A(n_160),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_192),
.Y(n_219)
);

OAI22x1_ASAP7_75t_R g220 ( 
.A1(n_193),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_182),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_177),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_172),
.B(n_1),
.Y(n_223)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_182),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_161),
.B(n_3),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_182),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g227 ( 
.A(n_159),
.Y(n_227)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_182),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_169),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_207),
.Y(n_231)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_178),
.Y(n_232)
);

AND2x4_ASAP7_75t_L g233 ( 
.A(n_180),
.B(n_4),
.Y(n_233)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_172),
.Y(n_234)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_164),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_188),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_206),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_170),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_189),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_186),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_168),
.Y(n_242)
);

CKINVDCx11_ASAP7_75t_R g243 ( 
.A(n_163),
.Y(n_243)
);

BUFx8_ASAP7_75t_L g244 ( 
.A(n_168),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_173),
.Y(n_245)
);

OA21x2_ASAP7_75t_L g246 ( 
.A1(n_196),
.A2(n_6),
.B(n_7),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_173),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_187),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_202),
.B(n_7),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_208),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_213),
.Y(n_251)
);

INVx5_ASAP7_75t_L g252 ( 
.A(n_187),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_186),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_198),
.Y(n_254)
);

BUFx12f_ASAP7_75t_L g255 ( 
.A(n_165),
.Y(n_255)
);

BUFx8_ASAP7_75t_SL g256 ( 
.A(n_198),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_R g257 ( 
.A(n_219),
.B(n_241),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_216),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_230),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_230),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_R g261 ( 
.A(n_253),
.B(n_234),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_243),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_230),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_221),
.Y(n_264)
);

NAND2xp33_ASAP7_75t_R g265 ( 
.A(n_237),
.B(n_166),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_221),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_243),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_229),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_229),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_227),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_236),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_R g272 ( 
.A(n_234),
.B(n_171),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_254),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_230),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_255),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_242),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_218),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_R g278 ( 
.A(n_234),
.B(n_211),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_221),
.Y(n_279)
);

OAI21x1_ASAP7_75t_L g280 ( 
.A1(n_250),
.A2(n_167),
.B(n_179),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_242),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_232),
.B(n_174),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_226),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_256),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_256),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_232),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_226),
.Y(n_287)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_224),
.Y(n_288)
);

BUFx10_ASAP7_75t_L g289 ( 
.A(n_233),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_223),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_235),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_232),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_242),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_242),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_214),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_235),
.Y(n_296)
);

NAND2xp33_ASAP7_75t_R g297 ( 
.A(n_246),
.B(n_175),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_232),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_245),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_222),
.B(n_176),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_244),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_244),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_245),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_239),
.B(n_181),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_245),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_265),
.A2(n_215),
.B1(n_249),
.B2(n_217),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_276),
.B(n_252),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g308 ( 
.A(n_289),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_258),
.A2(n_233),
.B1(n_254),
.B2(n_217),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_295),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_281),
.Y(n_311)
);

INVx2_ASAP7_75t_SL g312 ( 
.A(n_289),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_303),
.Y(n_313)
);

BUFx2_ASAP7_75t_R g314 ( 
.A(n_262),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_291),
.B(n_231),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_296),
.B(n_231),
.Y(n_316)
);

NOR3xp33_ASAP7_75t_L g317 ( 
.A(n_271),
.B(n_225),
.C(n_249),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_271),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_259),
.Y(n_319)
);

NOR2xp67_ASAP7_75t_L g320 ( 
.A(n_270),
.B(n_275),
.Y(n_320)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_266),
.Y(n_321)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_279),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_293),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_273),
.B(n_240),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_294),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_299),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_268),
.B(n_238),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_273),
.B(n_251),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_298),
.B(n_225),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_290),
.B(n_261),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_305),
.B(n_252),
.Y(n_331)
);

AO21x2_ASAP7_75t_L g332 ( 
.A1(n_280),
.A2(n_236),
.B(n_246),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_257),
.B(n_247),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_260),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_264),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_300),
.B(n_252),
.Y(n_336)
);

AO221x1_ASAP7_75t_L g337 ( 
.A1(n_263),
.A2(n_220),
.B1(n_247),
.B2(n_248),
.C(n_245),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_301),
.B(n_231),
.Y(n_338)
);

NOR2xp67_ASAP7_75t_L g339 ( 
.A(n_277),
.B(n_231),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_274),
.Y(n_340)
);

INVx8_ASAP7_75t_L g341 ( 
.A(n_286),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_282),
.B(n_252),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_300),
.B(n_248),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_272),
.B(n_183),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_292),
.B(n_248),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_264),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_304),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_304),
.B(n_248),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_264),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_288),
.B(n_224),
.Y(n_350)
);

NOR3xp33_ASAP7_75t_L g351 ( 
.A(n_269),
.B(n_201),
.C(n_185),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_283),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_278),
.B(n_184),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_283),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_288),
.B(n_224),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_283),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_302),
.B(n_224),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_L g358 ( 
.A1(n_297),
.A2(n_226),
.B1(n_200),
.B2(n_209),
.Y(n_358)
);

INVxp33_ASAP7_75t_L g359 ( 
.A(n_267),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_287),
.B(n_228),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_287),
.B(n_228),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_287),
.Y(n_362)
);

INVxp33_ASAP7_75t_L g363 ( 
.A(n_284),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_285),
.B(n_228),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_276),
.B(n_228),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_273),
.B(n_190),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_265),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_295),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_295),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_265),
.A2(n_199),
.B1(n_205),
.B2(n_204),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_303),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g372 ( 
.A(n_333),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_347),
.B(n_191),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_335),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_367),
.B(n_194),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_311),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_L g377 ( 
.A1(n_317),
.A2(n_226),
.B1(n_203),
.B2(n_197),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_306),
.A2(n_195),
.B1(n_10),
.B2(n_11),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_341),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_329),
.B(n_9),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_313),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_335),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_341),
.Y(n_383)
);

AND2x4_ASAP7_75t_L g384 ( 
.A(n_308),
.B(n_9),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g385 ( 
.A(n_312),
.B(n_11),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_318),
.B(n_13),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_330),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_370),
.B(n_13),
.Y(n_388)
);

AND2x4_ASAP7_75t_L g389 ( 
.A(n_339),
.B(n_14),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_323),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_L g391 ( 
.A1(n_309),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_324),
.B(n_15),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_325),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_371),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_366),
.B(n_17),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_341),
.Y(n_396)
);

HB1xp67_ASAP7_75t_SL g397 ( 
.A(n_314),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_319),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_328),
.B(n_18),
.Y(n_399)
);

NAND2x1p5_ASAP7_75t_L g400 ( 
.A(n_310),
.B(n_20),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_345),
.B(n_21),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_348),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_348),
.A2(n_23),
.B(n_24),
.Y(n_403)
);

BUFx8_ASAP7_75t_L g404 ( 
.A(n_338),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_343),
.B(n_25),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_L g406 ( 
.A1(n_358),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_320),
.B(n_29),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_334),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_326),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_335),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_340),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_346),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_346),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_368),
.B(n_30),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_369),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_321),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_321),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_364),
.B(n_31),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_322),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_346),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_322),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_349),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_364),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_332),
.B(n_336),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_351),
.B(n_34),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_359),
.B(n_36),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_354),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_356),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_L g429 ( 
.A1(n_337),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_327),
.B(n_43),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_344),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_332),
.B(n_48),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_336),
.A2(n_156),
.B(n_51),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_357),
.B(n_49),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_315),
.B(n_54),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_316),
.B(n_55),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_352),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_356),
.B(n_56),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_362),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_353),
.B(n_57),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_376),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_398),
.Y(n_442)
);

AND2x4_ASAP7_75t_L g443 ( 
.A(n_383),
.B(n_307),
.Y(n_443)
);

NAND3xp33_ASAP7_75t_L g444 ( 
.A(n_391),
.B(n_378),
.C(n_377),
.Y(n_444)
);

AOI21x1_ASAP7_75t_L g445 ( 
.A1(n_424),
.A2(n_342),
.B(n_365),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_396),
.Y(n_446)
);

AOI21x1_ASAP7_75t_L g447 ( 
.A1(n_424),
.A2(n_365),
.B(n_331),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_379),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_405),
.A2(n_355),
.B(n_350),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_408),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_395),
.A2(n_363),
.B1(n_355),
.B2(n_350),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_387),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_405),
.A2(n_331),
.B(n_307),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_374),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_R g455 ( 
.A(n_423),
.B(n_60),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_387),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_402),
.B(n_361),
.Y(n_457)
);

OAI22x1_ASAP7_75t_L g458 ( 
.A1(n_384),
.A2(n_360),
.B1(n_63),
.B2(n_64),
.Y(n_458)
);

A2O1A1Ixp33_ASAP7_75t_L g459 ( 
.A1(n_392),
.A2(n_61),
.B(n_65),
.C(n_66),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_384),
.B(n_68),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_R g461 ( 
.A(n_397),
.B(n_69),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_374),
.Y(n_462)
);

OAI21x1_ASAP7_75t_L g463 ( 
.A1(n_432),
.A2(n_70),
.B(n_71),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_381),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_374),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_385),
.B(n_72),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_402),
.A2(n_73),
.B(n_76),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_373),
.B(n_78),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_372),
.B(n_80),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_373),
.B(n_81),
.Y(n_470)
);

NOR2x1_ASAP7_75t_R g471 ( 
.A(n_385),
.B(n_83),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_430),
.B(n_84),
.Y(n_472)
);

O2A1O1Ixp33_ASAP7_75t_L g473 ( 
.A1(n_392),
.A2(n_86),
.B(n_89),
.C(n_90),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_399),
.B(n_91),
.Y(n_474)
);

AO21x1_ASAP7_75t_L g475 ( 
.A1(n_432),
.A2(n_92),
.B(n_93),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_415),
.B(n_94),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_390),
.B(n_96),
.Y(n_477)
);

A2O1A1Ixp33_ASAP7_75t_L g478 ( 
.A1(n_391),
.A2(n_97),
.B(n_99),
.C(n_100),
.Y(n_478)
);

A2O1A1Ixp33_ASAP7_75t_L g479 ( 
.A1(n_386),
.A2(n_102),
.B(n_103),
.C(n_104),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_393),
.B(n_105),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_428),
.A2(n_106),
.B(n_107),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_409),
.B(n_108),
.Y(n_482)
);

O2A1O1Ixp33_ASAP7_75t_L g483 ( 
.A1(n_380),
.A2(n_109),
.B(n_111),
.C(n_112),
.Y(n_483)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_416),
.B(n_114),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_411),
.B(n_115),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_404),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_382),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_428),
.A2(n_117),
.B(n_120),
.Y(n_488)
);

O2A1O1Ixp33_ASAP7_75t_L g489 ( 
.A1(n_388),
.A2(n_123),
.B(n_124),
.C(n_125),
.Y(n_489)
);

O2A1O1Ixp33_ASAP7_75t_L g490 ( 
.A1(n_425),
.A2(n_127),
.B(n_128),
.C(n_129),
.Y(n_490)
);

INVx1_ASAP7_75t_SL g491 ( 
.A(n_389),
.Y(n_491)
);

CKINVDCx8_ASAP7_75t_R g492 ( 
.A(n_397),
.Y(n_492)
);

O2A1O1Ixp33_ASAP7_75t_L g493 ( 
.A1(n_377),
.A2(n_131),
.B(n_132),
.C(n_137),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_394),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_422),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_R g496 ( 
.A(n_404),
.B(n_138),
.Y(n_496)
);

O2A1O1Ixp33_ASAP7_75t_L g497 ( 
.A1(n_375),
.A2(n_139),
.B(n_141),
.C(n_143),
.Y(n_497)
);

INVx4_ASAP7_75t_L g498 ( 
.A(n_446),
.Y(n_498)
);

AO21x2_ASAP7_75t_L g499 ( 
.A1(n_445),
.A2(n_401),
.B(n_438),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_441),
.B(n_426),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_444),
.B(n_417),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_486),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_491),
.B(n_414),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_441),
.B(n_472),
.Y(n_504)
);

BUFx2_ASAP7_75t_SL g505 ( 
.A(n_492),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_495),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_468),
.A2(n_427),
.B(n_438),
.Y(n_507)
);

AO21x2_ASAP7_75t_L g508 ( 
.A1(n_447),
.A2(n_453),
.B(n_449),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_450),
.Y(n_509)
);

INVx5_ASAP7_75t_L g510 ( 
.A(n_454),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_448),
.B(n_414),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_442),
.Y(n_512)
);

OAI21x1_ASAP7_75t_L g513 ( 
.A1(n_463),
.A2(n_403),
.B(n_433),
.Y(n_513)
);

BUFx2_ASAP7_75t_R g514 ( 
.A(n_460),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_464),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_452),
.B(n_389),
.Y(n_516)
);

AO21x2_ASAP7_75t_L g517 ( 
.A1(n_470),
.A2(n_474),
.B(n_477),
.Y(n_517)
);

NAND2x1p5_ASAP7_75t_L g518 ( 
.A(n_454),
.B(n_420),
.Y(n_518)
);

AOI22x1_ASAP7_75t_L g519 ( 
.A1(n_467),
.A2(n_407),
.B1(n_403),
.B2(n_433),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_454),
.Y(n_520)
);

AND2x6_ASAP7_75t_L g521 ( 
.A(n_462),
.B(n_487),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_456),
.B(n_457),
.Y(n_522)
);

OA21x2_ASAP7_75t_L g523 ( 
.A1(n_475),
.A2(n_436),
.B(n_435),
.Y(n_523)
);

BUFx12f_ASAP7_75t_L g524 ( 
.A(n_484),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_494),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_480),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_482),
.Y(n_527)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_455),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_443),
.B(n_410),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_485),
.Y(n_530)
);

OAI21x1_ASAP7_75t_L g531 ( 
.A1(n_481),
.A2(n_400),
.B(n_418),
.Y(n_531)
);

INVx5_ASAP7_75t_L g532 ( 
.A(n_462),
.Y(n_532)
);

CKINVDCx16_ASAP7_75t_R g533 ( 
.A(n_496),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_461),
.Y(n_534)
);

INVx2_ASAP7_75t_SL g535 ( 
.A(n_443),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_462),
.Y(n_536)
);

BUFx2_ASAP7_75t_L g537 ( 
.A(n_465),
.Y(n_537)
);

AOI22x1_ASAP7_75t_L g538 ( 
.A1(n_458),
.A2(n_400),
.B1(n_434),
.B2(n_421),
.Y(n_538)
);

BUFx12f_ASAP7_75t_L g539 ( 
.A(n_465),
.Y(n_539)
);

BUFx12f_ASAP7_75t_L g540 ( 
.A(n_465),
.Y(n_540)
);

AO21x1_ASAP7_75t_L g541 ( 
.A1(n_493),
.A2(n_440),
.B(n_431),
.Y(n_541)
);

BUFx12f_ASAP7_75t_L g542 ( 
.A(n_487),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_476),
.B(n_429),
.Y(n_543)
);

INVxp67_ASAP7_75t_SL g544 ( 
.A(n_487),
.Y(n_544)
);

OAI21x1_ASAP7_75t_L g545 ( 
.A1(n_488),
.A2(n_410),
.B(n_420),
.Y(n_545)
);

BUFx4f_ASAP7_75t_SL g546 ( 
.A(n_466),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_469),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_512),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_506),
.Y(n_549)
);

AOI21x1_ASAP7_75t_L g550 ( 
.A1(n_543),
.A2(n_451),
.B(n_439),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_512),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_501),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_501),
.B(n_429),
.Y(n_553)
);

NAND2x1_ASAP7_75t_L g554 ( 
.A(n_526),
.B(n_527),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_543),
.A2(n_419),
.B1(n_437),
.B2(n_434),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_503),
.A2(n_406),
.B1(n_471),
.B2(n_412),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_515),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_533),
.Y(n_558)
);

CKINVDCx11_ASAP7_75t_R g559 ( 
.A(n_502),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_510),
.Y(n_560)
);

NAND2x1p5_ASAP7_75t_L g561 ( 
.A(n_510),
.B(n_413),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_515),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_516),
.Y(n_563)
);

BUFx2_ASAP7_75t_R g564 ( 
.A(n_505),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_503),
.A2(n_413),
.B1(n_412),
.B2(n_382),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_509),
.Y(n_566)
);

NAND2x1p5_ASAP7_75t_L g567 ( 
.A(n_510),
.B(n_413),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_539),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_529),
.B(n_412),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_525),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_503),
.B(n_478),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_524),
.A2(n_382),
.B1(n_489),
.B2(n_483),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_522),
.Y(n_573)
);

OAI21x1_ASAP7_75t_L g574 ( 
.A1(n_513),
.A2(n_473),
.B(n_497),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_535),
.Y(n_575)
);

AO21x2_ASAP7_75t_L g576 ( 
.A1(n_507),
.A2(n_459),
.B(n_479),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_539),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_SL g578 ( 
.A1(n_538),
.A2(n_490),
.B1(n_145),
.B2(n_146),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_537),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_521),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_526),
.Y(n_581)
);

OAI21x1_ASAP7_75t_L g582 ( 
.A1(n_513),
.A2(n_144),
.B(n_147),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_524),
.A2(n_150),
.B1(n_151),
.B2(n_546),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_508),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_508),
.Y(n_585)
);

OR2x6_ASAP7_75t_L g586 ( 
.A(n_511),
.B(n_504),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_500),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_545),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_545),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_499),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_559),
.Y(n_591)
);

CKINVDCx16_ASAP7_75t_R g592 ( 
.A(n_558),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_558),
.B(n_534),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_552),
.B(n_544),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_566),
.Y(n_595)
);

NAND3xp33_ASAP7_75t_L g596 ( 
.A(n_553),
.B(n_530),
.C(n_519),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_563),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_553),
.A2(n_546),
.B1(n_514),
.B2(n_511),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_566),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_564),
.Y(n_600)
);

INVxp33_ASAP7_75t_SL g601 ( 
.A(n_577),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_568),
.Y(n_602)
);

OR2x2_ASAP7_75t_SL g603 ( 
.A(n_573),
.B(n_547),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_552),
.B(n_511),
.Y(n_604)
);

OR2x6_ASAP7_75t_L g605 ( 
.A(n_586),
.B(n_571),
.Y(n_605)
);

AND2x6_ASAP7_75t_L g606 ( 
.A(n_580),
.B(n_529),
.Y(n_606)
);

CKINVDCx16_ASAP7_75t_R g607 ( 
.A(n_568),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_570),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_579),
.B(n_528),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_569),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_586),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_586),
.B(n_529),
.Y(n_612)
);

OR2x2_ASAP7_75t_SL g613 ( 
.A(n_549),
.B(n_534),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_586),
.Y(n_614)
);

OAI21xp5_ASAP7_75t_SL g615 ( 
.A1(n_578),
.A2(n_541),
.B(n_518),
.Y(n_615)
);

CKINVDCx16_ASAP7_75t_R g616 ( 
.A(n_569),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_549),
.B(n_502),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_571),
.A2(n_517),
.B1(n_523),
.B2(n_540),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_587),
.B(n_581),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_SL g620 ( 
.A(n_580),
.B(n_498),
.Y(n_620)
);

OR2x6_ASAP7_75t_L g621 ( 
.A(n_554),
.B(n_542),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_581),
.A2(n_570),
.B1(n_556),
.B2(n_555),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_548),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_569),
.B(n_536),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_575),
.B(n_536),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_561),
.Y(n_626)
);

NAND2xp33_ASAP7_75t_R g627 ( 
.A(n_580),
.B(n_523),
.Y(n_627)
);

AND2x2_ASAP7_75t_SL g628 ( 
.A(n_583),
.B(n_498),
.Y(n_628)
);

OR2x6_ASAP7_75t_L g629 ( 
.A(n_554),
.B(n_542),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_560),
.Y(n_630)
);

NAND2xp33_ASAP7_75t_R g631 ( 
.A(n_548),
.B(n_523),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_R g632 ( 
.A(n_550),
.B(n_540),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_561),
.B(n_520),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_551),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_561),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_551),
.A2(n_517),
.B1(n_499),
.B2(n_521),
.Y(n_636)
);

AO21x1_ASAP7_75t_L g637 ( 
.A1(n_550),
.A2(n_584),
.B(n_585),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_567),
.B(n_510),
.Y(n_638)
);

BUFx2_ASAP7_75t_L g639 ( 
.A(n_567),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_567),
.Y(n_640)
);

HB1xp67_ASAP7_75t_L g641 ( 
.A(n_597),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_605),
.B(n_584),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_605),
.Y(n_643)
);

AOI21xp33_ASAP7_75t_L g644 ( 
.A1(n_631),
.A2(n_576),
.B(n_572),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_617),
.B(n_557),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_623),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_619),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_604),
.B(n_562),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_594),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_599),
.B(n_589),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_619),
.Y(n_651)
);

INVx1_ASAP7_75t_SL g652 ( 
.A(n_602),
.Y(n_652)
);

INVx1_ASAP7_75t_SL g653 ( 
.A(n_609),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_SL g654 ( 
.A(n_600),
.B(n_592),
.Y(n_654)
);

INVxp33_ASAP7_75t_L g655 ( 
.A(n_593),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_594),
.B(n_590),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_608),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_612),
.B(n_588),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_634),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_595),
.B(n_589),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_618),
.B(n_588),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_637),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_603),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_630),
.Y(n_664)
);

INVx1_ASAP7_75t_SL g665 ( 
.A(n_601),
.Y(n_665)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_625),
.Y(n_666)
);

OR2x2_ASAP7_75t_L g667 ( 
.A(n_613),
.B(n_596),
.Y(n_667)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_596),
.B(n_576),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_636),
.Y(n_669)
);

HB1xp67_ASAP7_75t_L g670 ( 
.A(n_621),
.Y(n_670)
);

BUFx2_ASAP7_75t_L g671 ( 
.A(n_621),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_611),
.Y(n_672)
);

AO21x2_ASAP7_75t_L g673 ( 
.A1(n_632),
.A2(n_574),
.B(n_582),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_621),
.Y(n_674)
);

AOI21x1_ASAP7_75t_L g675 ( 
.A1(n_629),
.A2(n_574),
.B(n_582),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_629),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_653),
.B(n_607),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_657),
.Y(n_678)
);

AND2x4_ASAP7_75t_SL g679 ( 
.A(n_641),
.B(n_629),
.Y(n_679)
);

INVxp67_ASAP7_75t_SL g680 ( 
.A(n_649),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g681 ( 
.A(n_666),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_643),
.B(n_610),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_643),
.B(n_633),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_664),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_658),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_657),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_647),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_643),
.B(n_614),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_647),
.B(n_628),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_651),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_667),
.B(n_598),
.Y(n_691)
);

HB1xp67_ASAP7_75t_L g692 ( 
.A(n_651),
.Y(n_692)
);

NOR3xp33_ASAP7_75t_L g693 ( 
.A(n_667),
.B(n_598),
.C(n_615),
.Y(n_693)
);

AND2x4_ASAP7_75t_SL g694 ( 
.A(n_670),
.B(n_638),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_646),
.Y(n_695)
);

INVx1_ASAP7_75t_SL g696 ( 
.A(n_665),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_658),
.B(n_650),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_650),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_663),
.B(n_615),
.Y(n_699)
);

AND2x4_ASAP7_75t_SL g700 ( 
.A(n_676),
.B(n_624),
.Y(n_700)
);

OR2x2_ASAP7_75t_L g701 ( 
.A(n_645),
.B(n_616),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_646),
.Y(n_702)
);

AOI221xp5_ASAP7_75t_L g703 ( 
.A1(n_644),
.A2(n_622),
.B1(n_591),
.B2(n_620),
.C(n_565),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_660),
.Y(n_704)
);

OR2x2_ASAP7_75t_L g705 ( 
.A(n_658),
.B(n_639),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_661),
.B(n_640),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_668),
.B(n_640),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_661),
.B(n_635),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_680),
.B(n_668),
.Y(n_709)
);

AND2x2_ASAP7_75t_SL g710 ( 
.A(n_693),
.B(n_663),
.Y(n_710)
);

HB1xp67_ASAP7_75t_L g711 ( 
.A(n_681),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_692),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_697),
.B(n_664),
.Y(n_713)
);

AND2x4_ASAP7_75t_SL g714 ( 
.A(n_688),
.B(n_672),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_697),
.B(n_652),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_685),
.B(n_654),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_686),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_685),
.B(n_671),
.Y(n_718)
);

OR2x2_ASAP7_75t_L g719 ( 
.A(n_704),
.B(n_656),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_685),
.B(n_671),
.Y(n_720)
);

OR2x2_ASAP7_75t_L g721 ( 
.A(n_698),
.B(n_656),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_677),
.B(n_642),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_687),
.B(n_660),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_691),
.A2(n_642),
.B1(n_627),
.B2(n_669),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_684),
.B(n_655),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_717),
.Y(n_726)
);

NAND2x2_ASAP7_75t_L g727 ( 
.A(n_709),
.B(n_684),
.Y(n_727)
);

NAND2x1p5_ASAP7_75t_L g728 ( 
.A(n_725),
.B(n_696),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_712),
.Y(n_729)
);

XNOR2xp5_ASAP7_75t_L g730 ( 
.A(n_710),
.B(n_691),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_711),
.B(n_690),
.Y(n_731)
);

OAI22xp5_ASAP7_75t_SL g732 ( 
.A1(n_710),
.A2(n_699),
.B1(n_689),
.B2(n_688),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_711),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_717),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_723),
.Y(n_735)
);

INVxp67_ASAP7_75t_L g736 ( 
.A(n_729),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_730),
.A2(n_699),
.B1(n_724),
.B2(n_669),
.Y(n_737)
);

INVxp67_ASAP7_75t_L g738 ( 
.A(n_731),
.Y(n_738)
);

AOI21xp33_ASAP7_75t_SL g739 ( 
.A1(n_728),
.A2(n_732),
.B(n_733),
.Y(n_739)
);

OR2x2_ASAP7_75t_L g740 ( 
.A(n_735),
.B(n_709),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_736),
.Y(n_741)
);

OR2x2_ASAP7_75t_L g742 ( 
.A(n_738),
.B(n_740),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_737),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_739),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_741),
.Y(n_745)
);

NOR3xp33_ASAP7_75t_SL g746 ( 
.A(n_744),
.B(n_703),
.C(n_727),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_742),
.Y(n_747)
);

AOI211xp5_ASAP7_75t_L g748 ( 
.A1(n_743),
.A2(n_716),
.B(n_713),
.C(n_723),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_747),
.Y(n_749)
);

OA22x2_ASAP7_75t_L g750 ( 
.A1(n_745),
.A2(n_714),
.B1(n_715),
.B2(n_679),
.Y(n_750)
);

AOI221xp5_ASAP7_75t_L g751 ( 
.A1(n_749),
.A2(n_746),
.B1(n_748),
.B2(n_726),
.C(n_678),
.Y(n_751)
);

OAI211xp5_ASAP7_75t_L g752 ( 
.A1(n_750),
.A2(n_675),
.B(n_718),
.C(n_720),
.Y(n_752)
);

NOR3xp33_ASAP7_75t_L g753 ( 
.A(n_749),
.B(n_707),
.C(n_674),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_753),
.Y(n_754)
);

NOR2x1_ASAP7_75t_L g755 ( 
.A(n_752),
.B(n_751),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_753),
.Y(n_756)
);

INVxp33_ASAP7_75t_SL g757 ( 
.A(n_751),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_751),
.A2(n_679),
.B1(n_714),
.B2(n_700),
.Y(n_758)
);

INVxp33_ASAP7_75t_SL g759 ( 
.A(n_751),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_754),
.Y(n_760)
);

OR2x6_ASAP7_75t_L g761 ( 
.A(n_756),
.B(n_722),
.Y(n_761)
);

NAND3xp33_ASAP7_75t_L g762 ( 
.A(n_755),
.B(n_532),
.C(n_662),
.Y(n_762)
);

NAND4xp25_ASAP7_75t_L g763 ( 
.A(n_757),
.B(n_688),
.C(n_705),
.D(n_721),
.Y(n_763)
);

NAND4xp75_ASAP7_75t_L g764 ( 
.A(n_758),
.B(n_674),
.C(n_707),
.D(n_708),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_759),
.Y(n_765)
);

NAND4xp75_ASAP7_75t_L g766 ( 
.A(n_755),
.B(n_708),
.C(n_662),
.D(n_706),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_761),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_765),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_760),
.Y(n_769)
);

INVx1_ASAP7_75t_SL g770 ( 
.A(n_762),
.Y(n_770)
);

BUFx2_ASAP7_75t_L g771 ( 
.A(n_763),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_768),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_767),
.Y(n_773)
);

HB1xp67_ASAP7_75t_L g774 ( 
.A(n_769),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_769),
.Y(n_775)
);

INVxp67_ASAP7_75t_SL g776 ( 
.A(n_771),
.Y(n_776)
);

INVxp67_ASAP7_75t_L g777 ( 
.A(n_770),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_768),
.Y(n_778)
);

AOI31xp33_ASAP7_75t_L g779 ( 
.A1(n_776),
.A2(n_766),
.A3(n_764),
.B(n_518),
.Y(n_779)
);

OAI31xp33_ASAP7_75t_SL g780 ( 
.A1(n_775),
.A2(n_726),
.A3(n_531),
.B(n_682),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_774),
.B(n_734),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_773),
.Y(n_782)
);

A2O1A1Ixp33_ASAP7_75t_SL g783 ( 
.A1(n_772),
.A2(n_686),
.B(n_706),
.C(n_532),
.Y(n_783)
);

AOI22xp5_ASAP7_75t_L g784 ( 
.A1(n_777),
.A2(n_673),
.B1(n_700),
.B2(n_606),
.Y(n_784)
);

OAI22xp5_ASAP7_75t_L g785 ( 
.A1(n_782),
.A2(n_777),
.B1(n_778),
.B2(n_719),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_781),
.B(n_673),
.Y(n_786)
);

BUFx2_ASAP7_75t_L g787 ( 
.A(n_784),
.Y(n_787)
);

OAI22xp5_ASAP7_75t_L g788 ( 
.A1(n_779),
.A2(n_675),
.B1(n_701),
.B2(n_694),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_785),
.A2(n_780),
.B1(n_783),
.B2(n_673),
.Y(n_789)
);

CKINVDCx20_ASAP7_75t_R g790 ( 
.A(n_787),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_SL g791 ( 
.A1(n_788),
.A2(n_532),
.B1(n_626),
.B2(n_682),
.Y(n_791)
);

OAI21xp5_ASAP7_75t_L g792 ( 
.A1(n_790),
.A2(n_786),
.B(n_532),
.Y(n_792)
);

AOI21xp33_ASAP7_75t_L g793 ( 
.A1(n_789),
.A2(n_702),
.B(n_695),
.Y(n_793)
);

AOI322xp5_ASAP7_75t_L g794 ( 
.A1(n_793),
.A2(n_791),
.A3(n_683),
.B1(n_682),
.B2(n_702),
.C1(n_695),
.C2(n_648),
.Y(n_794)
);

AOI221xp5_ASAP7_75t_L g795 ( 
.A1(n_794),
.A2(n_792),
.B1(n_694),
.B2(n_683),
.C(n_659),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_795),
.A2(n_521),
.B1(n_606),
.B2(n_659),
.Y(n_796)
);


endmodule