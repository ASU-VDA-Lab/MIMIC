module real_jpeg_33109_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_0),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_0),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_1),
.A2(n_19),
.B(n_452),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_1),
.B(n_453),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_2),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_3),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_4),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_4),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_4),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_4),
.B(n_198),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_4),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_4),
.B(n_306),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_4),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_4),
.B(n_360),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_5),
.Y(n_304)
);

NAND2x1_ASAP7_75t_SL g38 ( 
.A(n_6),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_6),
.B(n_49),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_6),
.B(n_107),
.Y(n_106)
);

NAND2xp33_ASAP7_75t_SL g173 ( 
.A(n_6),
.B(n_96),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_6),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_6),
.B(n_439),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_7),
.Y(n_81)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_7),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_7),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_8),
.B(n_54),
.Y(n_53)
);

NAND2xp67_ASAP7_75t_SL g73 ( 
.A(n_8),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_8),
.B(n_94),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_8),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_8),
.B(n_203),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_8),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_8),
.B(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_8),
.B(n_329),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_9),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_9),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_9),
.B(n_29),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_9),
.B(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_9),
.B(n_135),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_9),
.B(n_176),
.Y(n_175)
);

AND2x2_ASAP7_75t_SL g206 ( 
.A(n_9),
.B(n_207),
.Y(n_206)
);

AND2x2_ASAP7_75t_SL g432 ( 
.A(n_9),
.B(n_127),
.Y(n_432)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_10),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_10),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_11),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_11),
.B(n_191),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_11),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_11),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_11),
.B(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_11),
.B(n_365),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_11),
.B(n_369),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_13),
.Y(n_91)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_13),
.Y(n_343)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_14),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_14),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_14),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_15),
.B(n_29),
.Y(n_62)
);

NAND2x1_ASAP7_75t_L g72 ( 
.A(n_15),
.B(n_49),
.Y(n_72)
);

NAND2x1p5_ASAP7_75t_L g87 ( 
.A(n_15),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_15),
.B(n_143),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_15),
.B(n_158),
.Y(n_157)
);

BUFx24_ASAP7_75t_L g163 ( 
.A(n_15),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_16),
.B(n_29),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_16),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_16),
.B(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_16),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_16),
.B(n_423),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_17),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_17),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_17),
.B(n_235),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_17),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_17),
.B(n_295),
.Y(n_294)
);

AND2x2_ASAP7_75t_SL g340 ( 
.A(n_17),
.B(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_17),
.B(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_17),
.B(n_374),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_409),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_223),
.B(n_407),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_179),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_24),
.B(n_180),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_111),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_25),
.B(n_112),
.C(n_177),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_45),
.C(n_68),
.Y(n_25)
);

XOR2x1_ASAP7_75t_L g183 ( 
.A(n_26),
.B(n_46),
.Y(n_183)
);

MAJx2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_34),
.C(n_38),
.Y(n_26)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_27),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

OA21x2_ASAP7_75t_L g229 ( 
.A1(n_28),
.A2(n_30),
.B(n_217),
.Y(n_229)
);

INVx4_ASAP7_75t_SL g312 ( 
.A(n_29),
.Y(n_312)
);

INVx8_ASAP7_75t_L g375 ( 
.A(n_29),
.Y(n_375)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_33),
.Y(n_176)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_33),
.Y(n_194)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_33),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_34),
.B(n_38),
.Y(n_216)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_42),
.Y(n_366)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_44),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_44),
.Y(n_208)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_44),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_56),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_52),
.B1(n_53),
.B2(n_55),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_48),
.Y(n_55)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_50),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_52),
.B(n_55),
.C(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_61),
.C(n_63),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_57),
.B(n_61),
.C(n_63),
.Y(n_168)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_58),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_58),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_60),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_60),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_61),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_211)
);

AO22x1_ASAP7_75t_SL g333 ( 
.A1(n_61),
.A2(n_62),
.B1(n_134),
.B2(n_248),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_62),
.B(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVxp67_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

XNOR2x1_ASAP7_75t_L g182 ( 
.A(n_69),
.B(n_183),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_82),
.C(n_97),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_70),
.B(n_82),
.Y(n_275)
);

XOR2x2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_77),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_72),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_72),
.A2(n_153),
.B1(n_422),
.B2(n_424),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_73),
.B(n_151),
.C(n_152),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_75),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_76),
.Y(n_144)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_77),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_79),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_81),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.C(n_92),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_83),
.B(n_231),
.Y(n_230)
);

BUFx4f_ASAP7_75t_SL g84 ( 
.A(n_85),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_86),
.B(n_93),
.Y(n_231)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XNOR2x1_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_87),
.B(n_116),
.C(n_118),
.Y(n_443)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_91),
.Y(n_331)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_97),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_103),
.C(n_106),
.Y(n_97)
);

XNOR2x1_ASAP7_75t_SL g187 ( 
.A(n_98),
.B(n_103),
.Y(n_187)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_102),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_106),
.B(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_106),
.B(n_187),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_109),
.Y(n_316)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_110),
.Y(n_358)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_110),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_145),
.B1(n_177),
.B2(n_178),
.Y(n_111)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_112),
.Y(n_178)
);

XNOR2x1_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_120),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_113),
.B(n_121),
.C(n_132),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_118),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_118),
.A2(n_119),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

MAJx2_ASAP7_75t_L g170 ( 
.A(n_118),
.B(n_157),
.C(n_162),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_118),
.B(n_318),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_119),
.B(n_318),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_132),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_125),
.C(n_129),
.Y(n_121)
);

XOR2x2_ASAP7_75t_SL g147 ( 
.A(n_122),
.B(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2x1_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_129),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_137),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_133),
.A2(n_247),
.B1(n_431),
.B2(n_432),
.Y(n_430)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_134),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_142),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_138),
.B(n_247),
.C(n_418),
.Y(n_417)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_141),
.Y(n_346)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_142),
.Y(n_418)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_166),
.Y(n_145)
);

INVxp67_ASAP7_75t_SL g448 ( 
.A(n_146),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.C(n_154),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_147),
.A2(n_149),
.B1(n_150),
.B2(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_147),
.Y(n_222)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_154),
.Y(n_220)
);

XNOR2x1_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_160),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_159),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_161),
.A2(n_162),
.B1(n_190),
.B2(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_162),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

AND2x2_ASAP7_75t_SL g425 ( 
.A(n_163),
.B(n_426),
.Y(n_425)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_167),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_169),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_170),
.B(n_172),
.C(n_174),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_175),
.B(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_184),
.C(n_218),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_182),
.B(n_219),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_184),
.B(n_285),
.Y(n_284)
);

MAJx2_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_209),
.C(n_214),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_185),
.B(n_278),
.Y(n_277)
);

MAJx2_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_188),
.C(n_195),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_188),
.A2(n_189),
.B1(n_195),
.B2(n_196),
.Y(n_270)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_190),
.Y(n_266)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_196),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_202),
.C(n_205),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_197),
.A2(n_205),
.B1(n_206),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_197),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_201),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_202),
.B(n_252),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_205),
.A2(n_206),
.B1(n_430),
.B2(n_433),
.Y(n_429)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_209),
.A2(n_210),
.B1(n_215),
.B2(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_211),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_215),
.Y(n_279)
);

XNOR2x1_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_286),
.B(n_404),
.Y(n_223)
);

NOR2x1_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_280),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_271),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g405 ( 
.A(n_226),
.B(n_271),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_249),
.C(n_267),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_227),
.B(n_402),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_232),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_229),
.B(n_230),
.C(n_232),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_240),
.C(n_246),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_233),
.A2(n_234),
.B1(n_240),
.B2(n_241),
.Y(n_393)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_246),
.B(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_250),
.B(n_268),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_254),
.C(n_264),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_251),
.B(n_395),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_254),
.A2(n_264),
.B1(n_265),
.B2(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_254),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_258),
.C(n_262),
.Y(n_254)
);

XNOR2x1_ASAP7_75t_SL g324 ( 
.A(n_255),
.B(n_262),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XNOR2x1_ASAP7_75t_SL g323 ( 
.A(n_258),
.B(n_324),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_261),
.Y(n_298)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_277),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_276),
.Y(n_272)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_273),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_282),
.C(n_283),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_277),
.Y(n_282)
);

OAI21x1_ASAP7_75t_L g404 ( 
.A1(n_280),
.A2(n_405),
.B(n_406),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_284),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_281),
.B(n_284),
.Y(n_406)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OA21x2_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_399),
.B(n_403),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_289),
.A2(n_386),
.B(n_398),
.Y(n_288)
);

OAI21x1_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_335),
.B(n_385),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_320),
.Y(n_290)
);

OR2x2_ASAP7_75t_L g385 ( 
.A(n_291),
.B(n_320),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_309),
.C(n_317),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_293),
.B(n_348),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_299),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_294),
.B(n_300),
.C(n_305),
.Y(n_322)
);

INVx2_ASAP7_75t_SL g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_305),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_309),
.A2(n_310),
.B1(n_317),
.B2(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_314),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_311),
.B(n_314),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_317),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_325),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_322),
.B(n_323),
.C(n_325),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_334),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_328),
.B1(n_332),
.B2(n_333),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_327),
.B(n_333),
.C(n_334),
.Y(n_390)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_350),
.B(n_384),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_347),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_337),
.B(n_347),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_340),
.C(n_344),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_338),
.A2(n_339),
.B1(n_380),
.B2(n_381),
.Y(n_379)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_340),
.A2(n_344),
.B1(n_345),
.B2(n_382),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_340),
.Y(n_382)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_377),
.B(n_383),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_352),
.A2(n_367),
.B(n_376),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_353),
.B(n_364),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_353),
.B(n_364),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_359),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_354),
.B(n_359),
.Y(n_378)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx3_ASAP7_75t_SL g360 ( 
.A(n_361),
.Y(n_360)
);

INVx8_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_373),
.Y(n_367)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx5_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_379),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_378),
.B(n_379),
.Y(n_383)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_387),
.B(n_397),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_387),
.B(n_397),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_394),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_389),
.A2(n_390),
.B1(n_391),
.B2(n_392),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_390),
.B(n_391),
.C(n_394),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_392),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_401),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_400),
.B(n_401),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_410),
.B(n_451),
.Y(n_409)
);

INVxp33_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

OR2x2_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_413),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_412),
.B(n_413),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_447),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_434),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_429),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_417),
.A2(n_419),
.B1(n_420),
.B2(n_428),
.Y(n_416)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_417),
.Y(n_428)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

XOR2x2_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_425),
.Y(n_420)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_422),
.Y(n_424)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_430),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_432),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_446),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_445),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_437),
.A2(n_442),
.B1(n_443),
.B2(n_444),
.Y(n_436)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_437),
.Y(n_444)
);

INVx5_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx8_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g442 ( 
.A(n_443),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_449),
.C(n_450),
.Y(n_447)
);


endmodule