module fake_jpeg_9712_n_197 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_197);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_197;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_35),
.Y(n_50)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_30),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_36),
.B(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_30),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_23),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_27),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_60),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_17),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_46),
.B(n_53),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_51),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_16),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_34),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_28),
.C(n_22),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_58),
.C(n_28),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_16),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_19),
.B1(n_23),
.B2(n_16),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_19),
.B1(n_23),
.B2(n_38),
.Y(n_69)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_61),
.B(n_65),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_57),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_67),
.Y(n_82)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_57),
.Y(n_67)
);

O2A1O1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_53),
.B(n_59),
.C(n_58),
.Y(n_86)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

NAND2x1_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_39),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_75),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_21),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_46),
.Y(n_80)
);

INVx6_ASAP7_75t_SL g74 ( 
.A(n_51),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_74),
.Y(n_84)
);

OAI32xp33_ASAP7_75t_L g76 ( 
.A1(n_42),
.A2(n_15),
.A3(n_25),
.B1(n_18),
.B2(n_31),
.Y(n_76)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

OR2x2_ASAP7_75t_SL g77 ( 
.A(n_44),
.B(n_19),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_55),
.Y(n_85)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_49),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_80),
.B(n_77),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_64),
.A2(n_45),
.B1(n_48),
.B2(n_54),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_81),
.A2(n_31),
.B(n_69),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_85),
.B(n_72),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_86),
.A2(n_64),
.B1(n_68),
.B2(n_34),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_61),
.A2(n_45),
.B1(n_48),
.B2(n_54),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_87),
.A2(n_64),
.B1(n_68),
.B2(n_72),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_31),
.C(n_39),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_94),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_89),
.B(n_91),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_29),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_29),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_96),
.Y(n_108)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_97),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_16),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_100),
.B(n_17),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_95),
.A2(n_75),
.B(n_76),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_102),
.A2(n_107),
.B(n_67),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_82),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_109),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_88),
.C(n_112),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_106),
.A2(n_95),
.B1(n_97),
.B2(n_89),
.Y(n_119)
);

CKINVDCx12_ASAP7_75t_R g109 ( 
.A(n_96),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_65),
.Y(n_110)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_98),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_111),
.A2(n_79),
.B1(n_93),
.B2(n_70),
.Y(n_135)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_114),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_73),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_116),
.Y(n_132)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_117),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_119),
.A2(n_133),
.B(n_134),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_122),
.C(n_129),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_116),
.A2(n_85),
.B(n_83),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_121),
.A2(n_130),
.B(n_100),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_83),
.C(n_85),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_113),
.A2(n_83),
.B1(n_84),
.B2(n_80),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_70),
.B1(n_25),
.B2(n_26),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_104),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_128),
.Y(n_150)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_102),
.C(n_115),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_111),
.A2(n_73),
.B(n_21),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_63),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_101),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_135),
.A2(n_106),
.B(n_107),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_126),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_140),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

INVxp67_ASAP7_75t_SL g162 ( 
.A(n_137),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g138 ( 
.A1(n_132),
.A2(n_99),
.B(n_103),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_138),
.B(n_145),
.Y(n_151)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_118),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_144),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_142),
.Y(n_159)
);

OAI32xp33_ASAP7_75t_L g143 ( 
.A1(n_118),
.A2(n_117),
.A3(n_101),
.B1(n_15),
.B2(n_25),
.Y(n_143)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

AOI322xp5_ASAP7_75t_L g147 ( 
.A1(n_134),
.A2(n_26),
.A3(n_22),
.B1(n_25),
.B2(n_43),
.C1(n_10),
.C2(n_14),
.Y(n_147)
);

OAI321xp33_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_143),
.A3(n_138),
.B1(n_145),
.B2(n_11),
.C(n_8),
.Y(n_161)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_130),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_127),
.A2(n_128),
.B1(n_121),
.B2(n_123),
.Y(n_149)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_120),
.C(n_122),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_155),
.C(n_144),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_150),
.B(n_129),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_154),
.B(n_0),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_131),
.C(n_119),
.Y(n_155)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_156),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_29),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_139),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_161),
.A2(n_141),
.B1(n_10),
.B2(n_8),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_170),
.C(n_173),
.Y(n_174)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_166),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_169),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_163),
.A2(n_137),
.B1(n_43),
.B2(n_2),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_168),
.A2(n_172),
.B1(n_162),
.B2(n_3),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_29),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_29),
.Y(n_170)
);

INVxp33_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

INVxp67_ASAP7_75t_SL g181 ( 
.A(n_171),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_1),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_171),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_176),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_164),
.A2(n_159),
.B1(n_158),
.B2(n_160),
.Y(n_176)
);

AND2x2_ASAP7_75t_SL g177 ( 
.A(n_166),
.B(n_159),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_177),
.A2(n_181),
.B(n_175),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_180),
.B(n_2),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_174),
.B(n_155),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_185),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_165),
.C(n_170),
.Y(n_183)
);

AO21x1_ASAP7_75t_L g186 ( 
.A1(n_179),
.A2(n_169),
.B(n_4),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_187),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_184),
.A2(n_181),
.B(n_177),
.Y(n_189)
);

INVxp33_ASAP7_75t_L g193 ( 
.A(n_189),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_5),
.C(n_6),
.Y(n_191)
);

AOI21x1_ASAP7_75t_L g192 ( 
.A1(n_191),
.A2(n_5),
.B(n_6),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_192),
.B(n_190),
.C(n_188),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_194),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_193),
.A2(n_5),
.B(n_6),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_195),
.Y(n_197)
);


endmodule