module fake_jpeg_24534_n_231 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_231);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_231;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_5),
.B(n_10),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_8),
.B(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_25),
.B(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_36),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_28),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_21),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_55),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_21),
.B1(n_24),
.B2(n_29),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_49),
.A2(n_54),
.B1(n_41),
.B2(n_19),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_50),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_34),
.A2(n_24),
.B1(n_31),
.B2(n_30),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_52),
.A2(n_19),
.B1(n_20),
.B2(n_16),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_20),
.B1(n_19),
.B2(n_30),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_41),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_34),
.A2(n_33),
.B1(n_28),
.B2(n_20),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_59),
.A2(n_23),
.B1(n_27),
.B2(n_25),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_45),
.B(n_35),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_60),
.B(n_63),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_39),
.C(n_35),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_65),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_45),
.B(n_37),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_79),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_39),
.C(n_20),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_67),
.A2(n_80),
.B1(n_83),
.B2(n_23),
.Y(n_93)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_32),
.Y(n_69)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVxp67_ASAP7_75t_SL g109 ( 
.A(n_70),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

OR2x4_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_39),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_72),
.A2(n_78),
.B1(n_85),
.B2(n_48),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_86),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_36),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_76),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_19),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_46),
.Y(n_79)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_82),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_58),
.B(n_37),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_46),
.A2(n_16),
.B(n_31),
.C(n_33),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_42),
.Y(n_108)
);

INVx3_ASAP7_75t_SL g85 ( 
.A(n_44),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_43),
.B(n_36),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_36),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_94),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_93),
.A2(n_110),
.B1(n_107),
.B2(n_91),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_36),
.Y(n_94)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_107),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_99),
.A2(n_78),
.B1(n_85),
.B2(n_79),
.Y(n_118)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_100),
.B(n_102),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_42),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_101),
.B(n_105),
.Y(n_113)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_42),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_106),
.B(n_110),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_83),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_108),
.Y(n_134)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_61),
.B(n_38),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_65),
.Y(n_130)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_112),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_114),
.B(n_120),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_115),
.A2(n_132),
.B1(n_98),
.B2(n_102),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_72),
.B(n_62),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_130),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_112),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_119),
.Y(n_143)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_122),
.B(n_127),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_73),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_125),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_80),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_136),
.C(n_89),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_79),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

NAND3xp33_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_27),
.C(n_1),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_129),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_109),
.Y(n_129)
);

NAND4xp25_ASAP7_75t_L g131 ( 
.A(n_90),
.B(n_84),
.C(n_85),
.D(n_70),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_131),
.A2(n_108),
.B1(n_106),
.B2(n_98),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_93),
.A2(n_74),
.B1(n_86),
.B2(n_38),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_101),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_89),
.B(n_38),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_142),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_147),
.B1(n_155),
.B2(n_134),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_153),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_119),
.B(n_91),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_100),
.Y(n_144)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_149),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_90),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_152),
.A2(n_113),
.B(n_127),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_90),
.C(n_88),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_116),
.B(n_88),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_154),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_115),
.A2(n_74),
.B1(n_95),
.B2(n_103),
.Y(n_155)
);

AOI322xp5_ASAP7_75t_L g156 ( 
.A1(n_117),
.A2(n_32),
.A3(n_70),
.B1(n_71),
.B2(n_22),
.C1(n_64),
.C2(n_97),
.Y(n_156)
);

OAI321xp33_ASAP7_75t_L g178 ( 
.A1(n_156),
.A2(n_71),
.A3(n_26),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_103),
.Y(n_157)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

XOR2x1_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_10),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_22),
.Y(n_176)
);

OAI21xp33_ASAP7_75t_L g182 ( 
.A1(n_163),
.A2(n_151),
.B(n_152),
.Y(n_182)
);

NAND3xp33_ASAP7_75t_SL g164 ( 
.A(n_147),
.B(n_131),
.C(n_133),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_167),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_165),
.A2(n_166),
.B1(n_173),
.B2(n_138),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_148),
.A2(n_118),
.B1(n_135),
.B2(n_122),
.Y(n_166)
);

NOR3xp33_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_120),
.C(n_114),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_143),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_176),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_148),
.A2(n_136),
.B(n_132),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_171),
.A2(n_150),
.B(n_159),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_146),
.A2(n_155),
.B1(n_144),
.B2(n_153),
.Y(n_173)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_162),
.Y(n_188)
);

OAI321xp33_ASAP7_75t_L g181 ( 
.A1(n_178),
.A2(n_142),
.A3(n_141),
.B1(n_137),
.B2(n_4),
.C(n_6),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_179),
.A2(n_184),
.B1(n_192),
.B2(n_161),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_180),
.A2(n_171),
.B(n_161),
.Y(n_194)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_181),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_182),
.A2(n_11),
.B1(n_6),
.B2(n_7),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_166),
.A2(n_152),
.B1(n_139),
.B2(n_158),
.Y(n_184)
);

INVx13_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_191),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_160),
.A2(n_149),
.B1(n_140),
.B2(n_158),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_186),
.A2(n_187),
.B1(n_168),
.B2(n_169),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_160),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_187)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_177),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_190),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_173),
.A2(n_0),
.B1(n_6),
.B2(n_7),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_172),
.C(n_163),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_197),
.C(n_202),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_203),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_172),
.C(n_176),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_179),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_200),
.A2(n_192),
.B1(n_185),
.B2(n_181),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_168),
.C(n_175),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_187),
.Y(n_204)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_204),
.Y(n_217)
);

NAND2xp67_ASAP7_75t_SL g205 ( 
.A(n_203),
.B(n_183),
.Y(n_205)
);

A2O1A1Ixp33_ASAP7_75t_SL g219 ( 
.A1(n_205),
.A2(n_211),
.B(n_208),
.C(n_9),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_188),
.C(n_189),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_197),
.Y(n_215)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_196),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_209),
.B(n_210),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_9),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_202),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_195),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_213),
.Y(n_224)
);

OAI321xp33_ASAP7_75t_L g223 ( 
.A1(n_214),
.A2(n_219),
.A3(n_12),
.B1(n_13),
.B2(n_15),
.C(n_217),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_206),
.Y(n_222)
);

AO21x1_ASAP7_75t_L g218 ( 
.A1(n_205),
.A2(n_201),
.B(n_199),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_218),
.A2(n_206),
.B(n_12),
.Y(n_221)
);

OA21x2_ASAP7_75t_SL g220 ( 
.A1(n_219),
.A2(n_207),
.B(n_208),
.Y(n_220)
);

AOI31xp67_ASAP7_75t_SL g225 ( 
.A1(n_220),
.A2(n_223),
.A3(n_12),
.B(n_13),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_222),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_225),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_224),
.A2(n_214),
.B(n_216),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_226),
.A2(n_0),
.B(n_227),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_229),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_230),
.B(n_228),
.Y(n_231)
);


endmodule