module fake_netlist_1_7155_n_760 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_760);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_760;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_724;
wire n_228;
wire n_599;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_751;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g83 ( .A(n_14), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_16), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_66), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_3), .Y(n_86) );
CKINVDCx20_ASAP7_75t_R g87 ( .A(n_70), .Y(n_87) );
INVx2_ASAP7_75t_L g88 ( .A(n_46), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_2), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_29), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_16), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_67), .Y(n_92) );
CKINVDCx20_ASAP7_75t_R g93 ( .A(n_64), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_9), .Y(n_94) );
INVxp67_ASAP7_75t_SL g95 ( .A(n_14), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_24), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_68), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_60), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_7), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_62), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_51), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_28), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_10), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_35), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_49), .Y(n_105) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_56), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_1), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_15), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_32), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_7), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_41), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_25), .Y(n_112) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_61), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_59), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_76), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_53), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_69), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_33), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_15), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_37), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_2), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_13), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_1), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_20), .Y(n_124) );
BUFx2_ASAP7_75t_L g125 ( .A(n_8), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_42), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_72), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_57), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_52), .Y(n_129) );
INVxp67_ASAP7_75t_L g130 ( .A(n_48), .Y(n_130) );
BUFx3_ASAP7_75t_L g131 ( .A(n_77), .Y(n_131) );
BUFx3_ASAP7_75t_L g132 ( .A(n_23), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_78), .Y(n_133) );
INVx3_ASAP7_75t_L g134 ( .A(n_133), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_96), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_88), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_96), .Y(n_137) );
BUFx3_ASAP7_75t_L g138 ( .A(n_131), .Y(n_138) );
AOI22xp5_ASAP7_75t_L g139 ( .A1(n_119), .A2(n_125), .B1(n_103), .B2(n_91), .Y(n_139) );
CKINVDCx16_ASAP7_75t_R g140 ( .A(n_106), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_88), .Y(n_141) );
OR2x2_ASAP7_75t_L g142 ( .A(n_119), .B(n_0), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_112), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_131), .Y(n_144) );
AND2x4_ASAP7_75t_L g145 ( .A(n_94), .B(n_0), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_98), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_98), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_112), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_101), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_115), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_101), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_132), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_133), .Y(n_153) );
BUFx8_ASAP7_75t_L g154 ( .A(n_125), .Y(n_154) );
BUFx3_ASAP7_75t_L g155 ( .A(n_132), .Y(n_155) );
BUFx3_ASAP7_75t_L g156 ( .A(n_115), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_120), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_92), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_120), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_94), .B(n_3), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_104), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_114), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_99), .B(n_4), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_113), .B(n_4), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_116), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_99), .B(n_5), .Y(n_166) );
NOR2xp33_ASAP7_75t_SL g167 ( .A(n_85), .B(n_39), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_128), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_83), .B(n_5), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_128), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_117), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_118), .Y(n_172) );
NAND2xp33_ASAP7_75t_L g173 ( .A(n_85), .B(n_40), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_84), .B(n_6), .Y(n_174) );
OAI22xp5_ASAP7_75t_L g175 ( .A1(n_84), .A2(n_6), .B1(n_8), .B2(n_9), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_126), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_86), .B(n_107), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_127), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_129), .Y(n_179) );
INVx2_ASAP7_75t_SL g180 ( .A(n_154), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_158), .B(n_103), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_145), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_140), .B(n_130), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_145), .Y(n_184) );
INVx2_ASAP7_75t_SL g185 ( .A(n_154), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_145), .Y(n_186) );
INVx2_ASAP7_75t_SL g187 ( .A(n_154), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_170), .Y(n_188) );
INVx3_ASAP7_75t_L g189 ( .A(n_145), .Y(n_189) );
NAND2xp33_ASAP7_75t_L g190 ( .A(n_135), .B(n_105), .Y(n_190) );
INVx1_ASAP7_75t_SL g191 ( .A(n_140), .Y(n_191) );
BUFx3_ASAP7_75t_L g192 ( .A(n_138), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_158), .B(n_91), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_161), .B(n_121), .Y(n_194) );
BUFx3_ASAP7_75t_L g195 ( .A(n_138), .Y(n_195) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_170), .Y(n_196) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_170), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_134), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g199 ( .A1(n_139), .A2(n_121), .B1(n_123), .B2(n_122), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_161), .B(n_100), .Y(n_200) );
INVx2_ASAP7_75t_SL g201 ( .A(n_154), .Y(n_201) );
OAI22xp33_ASAP7_75t_L g202 ( .A1(n_139), .A2(n_95), .B1(n_89), .B2(n_110), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_170), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_135), .B(n_108), .Y(n_204) );
CKINVDCx14_ASAP7_75t_R g205 ( .A(n_164), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_134), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_170), .Y(n_207) );
INVx4_ASAP7_75t_L g208 ( .A(n_138), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_170), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_162), .B(n_100), .Y(n_210) );
INVxp67_ASAP7_75t_SL g211 ( .A(n_142), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_134), .B(n_102), .Y(n_212) );
BUFx2_ASAP7_75t_L g213 ( .A(n_164), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_134), .B(n_102), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_162), .B(n_97), .Y(n_215) );
BUFx10_ASAP7_75t_L g216 ( .A(n_165), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_165), .B(n_97), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_146), .Y(n_218) );
BUFx10_ASAP7_75t_L g219 ( .A(n_178), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_178), .B(n_109), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_146), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_137), .B(n_109), .Y(n_222) );
NOR2x1p5_ASAP7_75t_L g223 ( .A(n_142), .B(n_105), .Y(n_223) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_170), .Y(n_224) );
BUFx10_ASAP7_75t_L g225 ( .A(n_179), .Y(n_225) );
INVx3_ASAP7_75t_L g226 ( .A(n_156), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_179), .B(n_90), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_146), .B(n_90), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_146), .B(n_124), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_147), .B(n_111), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_174), .B(n_93), .Y(n_231) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_152), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_147), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_137), .A2(n_87), .B1(n_11), .B2(n_12), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_147), .B(n_44), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_149), .B(n_43), .Y(n_236) );
NOR2x1p5_ASAP7_75t_L g237 ( .A(n_177), .B(n_10), .Y(n_237) );
BUFx3_ASAP7_75t_L g238 ( .A(n_155), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_174), .B(n_11), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_147), .Y(n_240) );
INVx3_ASAP7_75t_L g241 ( .A(n_156), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_156), .Y(n_242) );
AND2x4_ASAP7_75t_L g243 ( .A(n_149), .B(n_12), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_151), .B(n_13), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_151), .B(n_17), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_153), .B(n_17), .Y(n_246) );
BUFx10_ASAP7_75t_L g247 ( .A(n_153), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_152), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_152), .Y(n_249) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_211), .A2(n_167), .B1(n_173), .B2(n_175), .Y(n_250) );
AOI22xp5_ASAP7_75t_SL g251 ( .A1(n_231), .A2(n_175), .B1(n_163), .B2(n_166), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_247), .B(n_167), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_243), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_247), .B(n_176), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_243), .Y(n_255) );
OR2x2_ASAP7_75t_L g256 ( .A(n_191), .B(n_177), .Y(n_256) );
AOI22xp5_ASAP7_75t_L g257 ( .A1(n_223), .A2(n_169), .B1(n_160), .B2(n_166), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_247), .B(n_176), .Y(n_258) );
INVx4_ASAP7_75t_L g259 ( .A(n_216), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_216), .B(n_155), .Y(n_260) );
INVx8_ASAP7_75t_L g261 ( .A(n_222), .Y(n_261) );
AOI22xp5_ASAP7_75t_L g262 ( .A1(n_180), .A2(n_169), .B1(n_160), .B2(n_163), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_L g263 ( .A1(n_202), .A2(n_176), .B(n_172), .C(n_136), .Y(n_263) );
OAI21xp5_ASAP7_75t_L g264 ( .A1(n_182), .A2(n_172), .B(n_136), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_216), .B(n_219), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_219), .B(n_155), .Y(n_266) );
OAI22xp33_ASAP7_75t_L g267 ( .A1(n_199), .A2(n_172), .B1(n_157), .B2(n_168), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_219), .B(n_157), .Y(n_268) );
AND2x4_ASAP7_75t_L g269 ( .A(n_180), .B(n_157), .Y(n_269) );
AND2x4_ASAP7_75t_L g270 ( .A(n_185), .B(n_157), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_243), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_225), .B(n_168), .Y(n_272) );
INVxp67_ASAP7_75t_L g273 ( .A(n_231), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_225), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_225), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_210), .B(n_168), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_185), .B(n_171), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_222), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_183), .B(n_168), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_192), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_222), .B(n_171), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_215), .B(n_148), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_217), .B(n_148), .Y(n_283) );
AOI22xp33_ASAP7_75t_L g284 ( .A1(n_244), .A2(n_171), .B1(n_159), .B2(n_150), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_184), .B(n_171), .Y(n_285) );
OAI21xp5_ASAP7_75t_L g286 ( .A1(n_186), .A2(n_148), .B(n_159), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_226), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_226), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_192), .Y(n_289) );
NAND3xp33_ASAP7_75t_L g290 ( .A(n_190), .B(n_152), .C(n_144), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_220), .B(n_136), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_200), .B(n_159), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_187), .B(n_171), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_181), .B(n_171), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_227), .B(n_150), .Y(n_295) );
BUFx3_ASAP7_75t_L g296 ( .A(n_226), .Y(n_296) );
AND2x6_ASAP7_75t_SL g297 ( .A(n_193), .B(n_18), .Y(n_297) );
NAND2x1p5_ASAP7_75t_L g298 ( .A(n_187), .B(n_150), .Y(n_298) );
OAI21xp5_ASAP7_75t_L g299 ( .A1(n_198), .A2(n_143), .B(n_141), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_195), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_201), .Y(n_301) );
OAI22xp5_ASAP7_75t_SL g302 ( .A1(n_205), .A2(n_143), .B1(n_141), .B2(n_171), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_195), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_238), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_241), .Y(n_305) );
INVx2_ASAP7_75t_SL g306 ( .A(n_201), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_241), .Y(n_307) );
NAND2xp5_ASAP7_75t_SL g308 ( .A(n_204), .B(n_143), .Y(n_308) );
O2A1O1Ixp5_ASAP7_75t_L g309 ( .A1(n_212), .A2(n_141), .B(n_152), .C(n_144), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_213), .B(n_144), .Y(n_310) );
AOI22xp5_ASAP7_75t_L g311 ( .A1(n_190), .A2(n_144), .B1(n_152), .B2(n_18), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_238), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_189), .B(n_152), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_241), .Y(n_314) );
AOI22xp5_ASAP7_75t_L g315 ( .A1(n_205), .A2(n_144), .B1(n_21), .B2(n_22), .Y(n_315) );
O2A1O1Ixp33_ASAP7_75t_L g316 ( .A1(n_194), .A2(n_144), .B(n_26), .C(n_27), .Y(n_316) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_232), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_189), .B(n_19), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_229), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g320 ( .A1(n_239), .A2(n_30), .B1(n_31), .B2(n_34), .Y(n_320) );
NOR2x1p5_ASAP7_75t_L g321 ( .A(n_204), .B(n_36), .Y(n_321) );
NAND2x1p5_ASAP7_75t_L g322 ( .A(n_237), .B(n_38), .Y(n_322) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_232), .Y(n_323) );
AOI22xp5_ASAP7_75t_L g324 ( .A1(n_229), .A2(n_45), .B1(n_47), .B2(n_50), .Y(n_324) );
AOI21xp5_ASAP7_75t_L g325 ( .A1(n_254), .A2(n_189), .B(n_228), .Y(n_325) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_256), .B(n_230), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_259), .B(n_204), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_314), .Y(n_328) );
NAND2xp5_ASAP7_75t_SL g329 ( .A(n_259), .B(n_212), .Y(n_329) );
OR2x2_ASAP7_75t_L g330 ( .A(n_273), .B(n_230), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_310), .Y(n_331) );
INVx4_ASAP7_75t_L g332 ( .A(n_261), .Y(n_332) );
AOI21xp5_ASAP7_75t_L g333 ( .A1(n_254), .A2(n_228), .B(n_214), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_261), .B(n_214), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_261), .B(n_208), .Y(n_335) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_265), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_296), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_280), .Y(n_338) );
BUFx6f_ASAP7_75t_L g339 ( .A(n_298), .Y(n_339) );
NAND2xp33_ASAP7_75t_SL g340 ( .A(n_301), .B(n_234), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_262), .B(n_245), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_289), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_278), .B(n_208), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_258), .A2(n_208), .B(n_206), .Y(n_344) );
OR2x6_ASAP7_75t_L g345 ( .A(n_298), .B(n_246), .Y(n_345) );
INVx1_ASAP7_75t_SL g346 ( .A(n_258), .Y(n_346) );
NOR2xp67_ASAP7_75t_SL g347 ( .A(n_306), .B(n_235), .Y(n_347) );
AOI21xp5_ASAP7_75t_L g348 ( .A1(n_260), .A2(n_266), .B(n_313), .Y(n_348) );
O2A1O1Ixp33_ASAP7_75t_L g349 ( .A1(n_263), .A2(n_242), .B(n_218), .C(n_233), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_300), .Y(n_350) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_317), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_281), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_303), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_302), .A2(n_240), .B1(n_221), .B2(n_236), .Y(n_354) );
A2O1A1Ixp33_ASAP7_75t_L g355 ( .A1(n_253), .A2(n_235), .B(n_249), .C(n_248), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_257), .B(n_54), .Y(n_356) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_255), .A2(n_249), .B1(n_248), .B2(n_188), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_304), .Y(n_358) );
INVx2_ASAP7_75t_SL g359 ( .A(n_321), .Y(n_359) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_317), .Y(n_360) );
NOR3xp33_ASAP7_75t_L g361 ( .A(n_319), .B(n_209), .C(n_203), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_281), .Y(n_362) );
AOI21xp5_ASAP7_75t_L g363 ( .A1(n_313), .A2(n_318), .B(n_268), .Y(n_363) );
INVxp67_ASAP7_75t_L g364 ( .A(n_269), .Y(n_364) );
NAND2xp33_ASAP7_75t_L g365 ( .A(n_274), .B(n_232), .Y(n_365) );
O2A1O1Ixp33_ASAP7_75t_L g366 ( .A1(n_267), .A2(n_203), .B(n_188), .C(n_209), .Y(n_366) );
AOI21xp5_ASAP7_75t_L g367 ( .A1(n_318), .A2(n_232), .B(n_224), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_269), .B(n_224), .Y(n_368) );
AOI21xp5_ASAP7_75t_L g369 ( .A1(n_272), .A2(n_224), .B(n_207), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_312), .Y(n_370) );
NOR3xp33_ASAP7_75t_L g371 ( .A(n_250), .B(n_55), .C(n_58), .Y(n_371) );
NOR2xp33_ASAP7_75t_SL g372 ( .A(n_271), .B(n_224), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_279), .B(n_63), .Y(n_373) );
AOI21xp5_ASAP7_75t_L g374 ( .A1(n_285), .A2(n_207), .B(n_197), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_270), .B(n_207), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_275), .B(n_207), .Y(n_376) );
BUFx2_ASAP7_75t_L g377 ( .A(n_270), .Y(n_377) );
A2O1A1Ixp33_ASAP7_75t_SL g378 ( .A1(n_294), .A2(n_197), .B(n_196), .C(n_73), .Y(n_378) );
CKINVDCx20_ASAP7_75t_R g379 ( .A(n_251), .Y(n_379) );
AOI22xp33_ASAP7_75t_SL g380 ( .A1(n_322), .A2(n_197), .B1(n_196), .B2(n_74), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_308), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_285), .A2(n_197), .B(n_196), .Y(n_382) );
CKINVDCx8_ASAP7_75t_R g383 ( .A(n_297), .Y(n_383) );
NOR2xp33_ASAP7_75t_SL g384 ( .A(n_332), .B(n_322), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_331), .Y(n_385) );
A2O1A1Ixp33_ASAP7_75t_L g386 ( .A1(n_356), .A2(n_282), .B(n_283), .C(n_291), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_330), .B(n_326), .Y(n_387) );
OR2x6_ASAP7_75t_L g388 ( .A(n_332), .B(n_252), .Y(n_388) );
OAI21xp5_ASAP7_75t_L g389 ( .A1(n_325), .A2(n_309), .B(n_264), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_379), .A2(n_288), .B1(n_287), .B2(n_305), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_346), .B(n_276), .Y(n_391) );
AO31x2_ASAP7_75t_L g392 ( .A1(n_355), .A2(n_292), .A3(n_295), .B(n_307), .Y(n_392) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_351), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_340), .A2(n_264), .B1(n_286), .B2(n_299), .Y(n_394) );
AO31x2_ASAP7_75t_L g395 ( .A1(n_367), .A2(n_316), .A3(n_311), .B(n_286), .Y(n_395) );
CKINVDCx20_ASAP7_75t_R g396 ( .A(n_383), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g397 ( .A1(n_346), .A2(n_284), .B1(n_315), .B2(n_320), .Y(n_397) );
OAI22xp5_ASAP7_75t_SL g398 ( .A1(n_359), .A2(n_324), .B1(n_290), .B2(n_299), .Y(n_398) );
NOR2xp67_ASAP7_75t_L g399 ( .A(n_327), .B(n_293), .Y(n_399) );
BUFx3_ASAP7_75t_L g400 ( .A(n_336), .Y(n_400) );
CKINVDCx20_ASAP7_75t_R g401 ( .A(n_327), .Y(n_401) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_351), .Y(n_402) );
INVx4_ASAP7_75t_L g403 ( .A(n_339), .Y(n_403) );
O2A1O1Ixp5_ASAP7_75t_L g404 ( .A1(n_373), .A2(n_277), .B(n_317), .C(n_323), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_341), .B(n_323), .Y(n_405) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_336), .Y(n_406) );
NAND3xp33_ASAP7_75t_L g407 ( .A(n_371), .B(n_196), .C(n_323), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_381), .Y(n_408) );
INVx3_ASAP7_75t_SL g409 ( .A(n_345), .Y(n_409) );
A2O1A1Ixp33_ASAP7_75t_L g410 ( .A1(n_333), .A2(n_65), .B(n_71), .C(n_75), .Y(n_410) );
O2A1O1Ixp33_ASAP7_75t_SL g411 ( .A1(n_378), .A2(n_366), .B(n_376), .C(n_363), .Y(n_411) );
OAI221xp5_ASAP7_75t_L g412 ( .A1(n_364), .A2(n_377), .B1(n_354), .B2(n_334), .C(n_343), .Y(n_412) );
AOI21xp5_ASAP7_75t_L g413 ( .A1(n_376), .A2(n_79), .B(n_80), .Y(n_413) );
OAI21x1_ASAP7_75t_L g414 ( .A1(n_374), .A2(n_81), .B(n_82), .Y(n_414) );
CKINVDCx5p33_ASAP7_75t_R g415 ( .A(n_345), .Y(n_415) );
INVx5_ASAP7_75t_L g416 ( .A(n_339), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_352), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_337), .B(n_362), .Y(n_418) );
AOI21xp5_ASAP7_75t_L g419 ( .A1(n_369), .A2(n_348), .B(n_382), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_387), .B(n_336), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_417), .Y(n_421) );
AOI221xp5_ASAP7_75t_L g422 ( .A1(n_385), .A2(n_349), .B1(n_361), .B2(n_335), .C(n_357), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_401), .B(n_329), .Y(n_423) );
OAI21xp5_ASAP7_75t_L g424 ( .A1(n_386), .A2(n_344), .B(n_357), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_393), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_412), .A2(n_345), .B1(n_339), .B2(n_338), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_408), .Y(n_427) );
OA21x2_ASAP7_75t_L g428 ( .A1(n_419), .A2(n_368), .B(n_375), .Y(n_428) );
OAI21x1_ASAP7_75t_SL g429 ( .A1(n_403), .A2(n_328), .B(n_342), .Y(n_429) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_406), .Y(n_430) );
OAI21xp5_ASAP7_75t_L g431 ( .A1(n_394), .A2(n_389), .B(n_405), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_391), .Y(n_432) );
BUFx3_ASAP7_75t_L g433 ( .A(n_416), .Y(n_433) );
AND2x4_ASAP7_75t_L g434 ( .A(n_416), .B(n_350), .Y(n_434) );
AOI21xp5_ASAP7_75t_L g435 ( .A1(n_411), .A2(n_372), .B(n_351), .Y(n_435) );
AOI21xp5_ASAP7_75t_L g436 ( .A1(n_397), .A2(n_372), .B(n_360), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_418), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_409), .B(n_353), .Y(n_438) );
OAI21xp33_ASAP7_75t_SL g439 ( .A1(n_414), .A2(n_358), .B(n_370), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_390), .B(n_380), .Y(n_440) );
AOI21xp5_ASAP7_75t_L g441 ( .A1(n_398), .A2(n_360), .B(n_365), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_415), .B(n_347), .Y(n_442) );
AND2x4_ASAP7_75t_SL g443 ( .A(n_403), .B(n_360), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_416), .B(n_400), .Y(n_444) );
A2O1A1Ixp33_ASAP7_75t_L g445 ( .A1(n_384), .A2(n_407), .B(n_399), .C(n_413), .Y(n_445) );
OAI21x1_ASAP7_75t_L g446 ( .A1(n_404), .A2(n_392), .B(n_399), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_392), .Y(n_447) );
AO21x2_ASAP7_75t_L g448 ( .A1(n_410), .A2(n_392), .B(n_395), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_388), .B(n_398), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_393), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_428), .Y(n_451) );
INVx4_ASAP7_75t_L g452 ( .A(n_443), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_420), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_421), .Y(n_454) );
NAND4xp25_ASAP7_75t_L g455 ( .A(n_437), .B(n_396), .C(n_388), .D(n_395), .Y(n_455) );
INVxp67_ASAP7_75t_L g456 ( .A(n_432), .Y(n_456) );
BUFx3_ASAP7_75t_L g457 ( .A(n_433), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_421), .Y(n_458) );
AO21x2_ASAP7_75t_L g459 ( .A1(n_431), .A2(n_395), .B(n_393), .Y(n_459) );
OA21x2_ASAP7_75t_L g460 ( .A1(n_446), .A2(n_402), .B(n_388), .Y(n_460) );
AND2x4_ASAP7_75t_L g461 ( .A(n_425), .B(n_402), .Y(n_461) );
INVx3_ASAP7_75t_L g462 ( .A(n_443), .Y(n_462) );
OAI21xp5_ASAP7_75t_L g463 ( .A1(n_431), .A2(n_402), .B(n_424), .Y(n_463) );
OAI222xp33_ASAP7_75t_L g464 ( .A1(n_449), .A2(n_426), .B1(n_440), .B2(n_432), .C1(n_437), .C2(n_427), .Y(n_464) );
OR2x6_ASAP7_75t_L g465 ( .A(n_429), .B(n_441), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_423), .B(n_438), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_439), .A2(n_436), .B(n_435), .Y(n_467) );
BUFx3_ASAP7_75t_L g468 ( .A(n_433), .Y(n_468) );
OAI221xp5_ASAP7_75t_L g469 ( .A1(n_422), .A2(n_427), .B1(n_442), .B2(n_445), .C(n_447), .Y(n_469) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_430), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_447), .B(n_428), .Y(n_471) );
INVx3_ASAP7_75t_L g472 ( .A(n_443), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_444), .B(n_434), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_428), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_428), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_433), .B(n_448), .Y(n_476) );
AND2x4_ASAP7_75t_L g477 ( .A(n_425), .B(n_450), .Y(n_477) );
INVxp67_ASAP7_75t_SL g478 ( .A(n_446), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_434), .A2(n_444), .B1(n_448), .B2(n_429), .Y(n_479) );
INVx3_ASAP7_75t_L g480 ( .A(n_425), .Y(n_480) );
OAI21xp5_ASAP7_75t_L g481 ( .A1(n_439), .A2(n_450), .B(n_434), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_448), .Y(n_482) );
AND2x4_ASAP7_75t_L g483 ( .A(n_450), .B(n_434), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_432), .B(n_421), .Y(n_484) );
BUFx3_ASAP7_75t_L g485 ( .A(n_433), .Y(n_485) );
OAI22xp33_ASAP7_75t_L g486 ( .A1(n_449), .A2(n_401), .B1(n_379), .B2(n_384), .Y(n_486) );
OR2x6_ASAP7_75t_L g487 ( .A(n_449), .B(n_429), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_449), .A2(n_379), .B1(n_340), .B2(n_401), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_451), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_451), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_451), .Y(n_491) );
BUFx2_ASAP7_75t_L g492 ( .A(n_481), .Y(n_492) );
BUFx2_ASAP7_75t_L g493 ( .A(n_481), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_484), .B(n_454), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_455), .A2(n_486), .B1(n_488), .B2(n_456), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_464), .B(n_456), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_474), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_454), .Y(n_498) );
AOI221xp5_ASAP7_75t_L g499 ( .A1(n_464), .A2(n_455), .B1(n_484), .B2(n_469), .C(n_458), .Y(n_499) );
INVx2_ASAP7_75t_SL g500 ( .A(n_457), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_474), .B(n_475), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_458), .B(n_474), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_475), .B(n_473), .Y(n_503) );
BUFx2_ASAP7_75t_L g504 ( .A(n_487), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_471), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_471), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_473), .B(n_477), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_477), .B(n_459), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_476), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_477), .B(n_459), .Y(n_510) );
NAND3xp33_ASAP7_75t_SL g511 ( .A(n_466), .B(n_479), .C(n_469), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_482), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_477), .B(n_459), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_459), .B(n_480), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_453), .A2(n_470), .B1(n_452), .B2(n_487), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_476), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_480), .B(n_483), .Y(n_517) );
INVx3_ASAP7_75t_L g518 ( .A(n_465), .Y(n_518) );
BUFx2_ASAP7_75t_L g519 ( .A(n_487), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_480), .B(n_483), .Y(n_520) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_487), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_483), .B(n_480), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_482), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_487), .B(n_485), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_483), .B(n_463), .Y(n_525) );
BUFx2_ASAP7_75t_L g526 ( .A(n_465), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_463), .B(n_485), .Y(n_527) );
INVx3_ASAP7_75t_L g528 ( .A(n_465), .Y(n_528) );
NAND2x1_ASAP7_75t_L g529 ( .A(n_465), .B(n_460), .Y(n_529) );
INVx5_ASAP7_75t_SL g530 ( .A(n_465), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_457), .B(n_485), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_460), .Y(n_532) );
NOR2x1_ASAP7_75t_SL g533 ( .A(n_452), .B(n_457), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_460), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_460), .Y(n_535) );
AND2x4_ASAP7_75t_L g536 ( .A(n_478), .B(n_461), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_478), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_461), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_468), .B(n_461), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_468), .B(n_461), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_498), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_494), .B(n_468), .Y(n_542) );
NOR2x1_ASAP7_75t_L g543 ( .A(n_531), .B(n_452), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_503), .B(n_467), .Y(n_544) );
NOR2x1_ASAP7_75t_L g545 ( .A(n_531), .B(n_511), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_494), .B(n_452), .Y(n_546) );
NOR3xp33_ASAP7_75t_SL g547 ( .A(n_511), .B(n_467), .C(n_472), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_498), .Y(n_548) );
INVx2_ASAP7_75t_SL g549 ( .A(n_500), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_503), .B(n_462), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_502), .Y(n_551) );
AND2x4_ASAP7_75t_SL g552 ( .A(n_539), .B(n_462), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_502), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_508), .B(n_462), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_508), .B(n_462), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_510), .B(n_472), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_510), .B(n_513), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_513), .B(n_472), .Y(n_558) );
AND2x4_ASAP7_75t_L g559 ( .A(n_518), .B(n_472), .Y(n_559) );
AND2x4_ASAP7_75t_L g560 ( .A(n_518), .B(n_528), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_525), .B(n_501), .Y(n_561) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_500), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_525), .B(n_501), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_501), .B(n_516), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_505), .B(n_506), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_505), .B(n_506), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_509), .B(n_516), .Y(n_567) );
OAI21xp5_ASAP7_75t_L g568 ( .A1(n_499), .A2(n_496), .B(n_495), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_509), .B(n_514), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_524), .B(n_489), .Y(n_570) );
BUFx2_ASAP7_75t_L g571 ( .A(n_500), .Y(n_571) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_540), .Y(n_572) );
INVx1_ASAP7_75t_SL g573 ( .A(n_524), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_514), .B(n_520), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_517), .B(n_520), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_507), .B(n_495), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_517), .B(n_507), .Y(n_577) );
INVx1_ASAP7_75t_SL g578 ( .A(n_539), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_492), .B(n_493), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_523), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_492), .B(n_493), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_527), .B(n_489), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_496), .B(n_499), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_527), .B(n_489), .Y(n_584) );
INVx2_ASAP7_75t_SL g585 ( .A(n_540), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_523), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_490), .B(n_491), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_490), .B(n_491), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_490), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_491), .B(n_497), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_497), .B(n_538), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_497), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_538), .B(n_522), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_512), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_515), .B(n_533), .Y(n_595) );
INVxp67_ASAP7_75t_L g596 ( .A(n_533), .Y(n_596) );
AND2x4_ASAP7_75t_L g597 ( .A(n_518), .B(n_528), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_512), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_578), .B(n_522), .Y(n_599) );
AOI211xp5_ASAP7_75t_L g600 ( .A1(n_568), .A2(n_521), .B(n_526), .C(n_504), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_557), .B(n_536), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_583), .A2(n_515), .B1(n_504), .B2(n_519), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_578), .B(n_557), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_574), .B(n_536), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_541), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_574), .B(n_536), .Y(n_606) );
INVx3_ASAP7_75t_L g607 ( .A(n_560), .Y(n_607) );
NOR2xp33_ASAP7_75t_SL g608 ( .A(n_596), .B(n_519), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_569), .B(n_521), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_561), .B(n_536), .Y(n_610) );
NOR2xp33_ASAP7_75t_SL g611 ( .A(n_543), .B(n_526), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_561), .B(n_532), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_563), .B(n_532), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_541), .Y(n_614) );
NAND2xp5_ASAP7_75t_SL g615 ( .A(n_545), .B(n_530), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_548), .Y(n_616) );
AND2x4_ASAP7_75t_L g617 ( .A(n_560), .B(n_597), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_548), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_569), .B(n_538), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_583), .B(n_518), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_563), .B(n_534), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_564), .B(n_534), .Y(n_622) );
INVx1_ASAP7_75t_SL g623 ( .A(n_552), .Y(n_623) );
OR2x2_ASAP7_75t_L g624 ( .A(n_542), .B(n_537), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_582), .B(n_535), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_577), .B(n_528), .Y(n_626) );
NAND2xp33_ASAP7_75t_SL g627 ( .A(n_571), .B(n_529), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_582), .B(n_535), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_584), .B(n_528), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_584), .B(n_530), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_564), .B(n_537), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_575), .B(n_530), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_576), .B(n_530), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_587), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_551), .B(n_530), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_567), .Y(n_636) );
OR2x6_ASAP7_75t_L g637 ( .A(n_595), .B(n_529), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_587), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_575), .B(n_537), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_551), .B(n_553), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_568), .B(n_545), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_577), .B(n_544), .Y(n_642) );
AND2x4_ASAP7_75t_L g643 ( .A(n_560), .B(n_597), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_567), .Y(n_644) );
OR2x2_ASAP7_75t_L g645 ( .A(n_572), .B(n_553), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_565), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_544), .B(n_593), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_565), .B(n_566), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_593), .B(n_581), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_566), .Y(n_650) );
OR2x2_ASAP7_75t_L g651 ( .A(n_570), .B(n_585), .Y(n_651) );
INVx2_ASAP7_75t_SL g652 ( .A(n_543), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_580), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_585), .B(n_579), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_642), .B(n_579), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_645), .Y(n_656) );
OAI21xp5_ASAP7_75t_L g657 ( .A1(n_641), .A2(n_547), .B(n_562), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_640), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_641), .A2(n_581), .B1(n_558), .B2(n_554), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_646), .Y(n_660) );
NAND2xp5_ASAP7_75t_SL g661 ( .A(n_611), .B(n_549), .Y(n_661) );
INVx2_ASAP7_75t_SL g662 ( .A(n_652), .Y(n_662) );
NAND2x1p5_ASAP7_75t_L g663 ( .A(n_623), .B(n_571), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_605), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_620), .B(n_573), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_614), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_620), .B(n_573), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_650), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_642), .B(n_554), .Y(n_669) );
OAI21xp5_ASAP7_75t_L g670 ( .A1(n_615), .A2(n_549), .B(n_546), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_636), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_600), .A2(n_552), .B1(n_550), .B2(n_570), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_616), .Y(n_673) );
AND2x4_ASAP7_75t_SL g674 ( .A(n_632), .B(n_550), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_618), .Y(n_675) );
INVx1_ASAP7_75t_SL g676 ( .A(n_603), .Y(n_676) );
OR2x2_ASAP7_75t_L g677 ( .A(n_631), .B(n_591), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_647), .B(n_591), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_647), .B(n_555), .Y(n_679) );
AOI221xp5_ASAP7_75t_L g680 ( .A1(n_644), .A2(n_586), .B1(n_580), .B2(n_597), .C(n_560), .Y(n_680) );
INVx2_ASAP7_75t_L g681 ( .A(n_653), .Y(n_681) );
OR2x2_ASAP7_75t_L g682 ( .A(n_651), .B(n_592), .Y(n_682) );
AOI21xp33_ASAP7_75t_SL g683 ( .A1(n_615), .A2(n_597), .B(n_559), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_612), .B(n_586), .Y(n_684) );
NOR4xp25_ASAP7_75t_L g685 ( .A(n_648), .B(n_558), .C(n_555), .D(n_556), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_612), .B(n_556), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_613), .B(n_590), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_613), .B(n_590), .Y(n_688) );
NAND4xp25_ASAP7_75t_SL g689 ( .A(n_602), .B(n_552), .C(n_588), .D(n_589), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_621), .B(n_649), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_639), .Y(n_691) );
OAI222xp33_ASAP7_75t_L g692 ( .A1(n_637), .A2(n_559), .B1(n_589), .B2(n_592), .C1(n_598), .C2(n_594), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_639), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_634), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_655), .B(n_649), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_660), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_672), .A2(n_633), .B1(n_632), .B2(n_654), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_685), .B(n_621), .Y(n_698) );
AOI222xp33_ASAP7_75t_L g699 ( .A1(n_680), .A2(n_609), .B1(n_629), .B2(n_627), .C1(n_622), .C2(n_625), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_659), .A2(n_652), .B1(n_637), .B2(n_601), .Y(n_700) );
A2O1A1Ixp33_ASAP7_75t_L g701 ( .A1(n_683), .A2(n_627), .B(n_608), .C(n_607), .Y(n_701) );
OAI31xp33_ASAP7_75t_L g702 ( .A1(n_692), .A2(n_607), .A3(n_617), .B(n_643), .Y(n_702) );
INVx2_ASAP7_75t_L g703 ( .A(n_682), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g704 ( .A1(n_689), .A2(n_626), .B1(n_630), .B2(n_629), .Y(n_704) );
AOI211x1_ASAP7_75t_L g705 ( .A1(n_657), .A2(n_610), .B(n_606), .C(n_604), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_658), .B(n_610), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_668), .Y(n_707) );
O2A1O1Ixp33_ASAP7_75t_L g708 ( .A1(n_661), .A2(n_637), .B(n_635), .C(n_607), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_682), .Y(n_709) );
XNOR2x1_ASAP7_75t_L g710 ( .A(n_676), .B(n_630), .Y(n_710) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_694), .Y(n_711) );
INVx2_ASAP7_75t_SL g712 ( .A(n_674), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_655), .B(n_628), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_664), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_664), .Y(n_715) );
INVxp33_ASAP7_75t_L g716 ( .A(n_661), .Y(n_716) );
OR2x2_ASAP7_75t_L g717 ( .A(n_677), .B(n_619), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_673), .Y(n_718) );
INVx1_ASAP7_75t_SL g719 ( .A(n_674), .Y(n_719) );
NAND2x1p5_ASAP7_75t_L g720 ( .A(n_719), .B(n_662), .Y(n_720) );
AOI211xp5_ASAP7_75t_L g721 ( .A1(n_701), .A2(n_670), .B(n_662), .C(n_665), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_699), .A2(n_656), .B1(n_667), .B2(n_671), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_714), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_715), .Y(n_724) );
AOI221xp5_ASAP7_75t_L g725 ( .A1(n_705), .A2(n_684), .B1(n_669), .B2(n_679), .C(n_686), .Y(n_725) );
INVx4_ASAP7_75t_L g726 ( .A(n_712), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_698), .B(n_669), .Y(n_727) );
NOR2x1_ASAP7_75t_L g728 ( .A(n_701), .B(n_637), .Y(n_728) );
AOI21xp33_ASAP7_75t_L g729 ( .A1(n_716), .A2(n_675), .B(n_673), .Y(n_729) );
O2A1O1Ixp33_ASAP7_75t_L g730 ( .A1(n_708), .A2(n_663), .B(n_690), .C(n_675), .Y(n_730) );
AOI21xp33_ASAP7_75t_L g731 ( .A1(n_708), .A2(n_624), .B(n_681), .Y(n_731) );
AOI211xp5_ASAP7_75t_SL g732 ( .A1(n_700), .A2(n_643), .B(n_617), .C(n_559), .Y(n_732) );
AOI21xp33_ASAP7_75t_L g733 ( .A1(n_702), .A2(n_681), .B(n_666), .Y(n_733) );
AOI221xp5_ASAP7_75t_L g734 ( .A1(n_706), .A2(n_679), .B1(n_686), .B2(n_691), .C(n_693), .Y(n_734) );
AOI222xp33_ASAP7_75t_L g735 ( .A1(n_727), .A2(n_709), .B1(n_696), .B2(n_707), .C1(n_706), .C2(n_718), .Y(n_735) );
INVx1_ASAP7_75t_SL g736 ( .A(n_726), .Y(n_736) );
OAI221xp5_ASAP7_75t_L g737 ( .A1(n_721), .A2(n_697), .B1(n_710), .B2(n_704), .C(n_663), .Y(n_737) );
AOI31xp33_ASAP7_75t_L g738 ( .A1(n_728), .A2(n_663), .A3(n_711), .B(n_695), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_723), .Y(n_739) );
O2A1O1Ixp5_ASAP7_75t_SL g740 ( .A1(n_733), .A2(n_711), .B(n_713), .C(n_678), .Y(n_740) );
AOI211xp5_ASAP7_75t_L g741 ( .A1(n_730), .A2(n_643), .B(n_617), .C(n_703), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_722), .B(n_717), .Y(n_742) );
AO21x1_ASAP7_75t_L g743 ( .A1(n_726), .A2(n_666), .B(n_559), .Y(n_743) );
NOR2x1_ASAP7_75t_L g744 ( .A(n_736), .B(n_724), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_739), .Y(n_745) );
NAND2xp5_ASAP7_75t_SL g746 ( .A(n_743), .B(n_720), .Y(n_746) );
NAND4xp25_ASAP7_75t_L g747 ( .A(n_737), .B(n_732), .C(n_734), .D(n_725), .Y(n_747) );
AOI211xp5_ASAP7_75t_L g748 ( .A1(n_741), .A2(n_731), .B(n_729), .C(n_601), .Y(n_748) );
NOR3xp33_ASAP7_75t_L g749 ( .A(n_747), .B(n_738), .C(n_742), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_744), .B(n_735), .Y(n_750) );
NAND2x1p5_ASAP7_75t_L g751 ( .A(n_746), .B(n_677), .Y(n_751) );
XNOR2xp5_ASAP7_75t_L g752 ( .A(n_749), .B(n_748), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_751), .Y(n_753) );
INVx3_ASAP7_75t_L g754 ( .A(n_753), .Y(n_754) );
NOR4xp25_ASAP7_75t_L g755 ( .A(n_752), .B(n_750), .C(n_745), .D(n_740), .Y(n_755) );
OAI31xp33_ASAP7_75t_L g756 ( .A1(n_754), .A2(n_693), .A3(n_691), .B(n_606), .Y(n_756) );
AOI222xp33_ASAP7_75t_L g757 ( .A1(n_756), .A2(n_754), .B1(n_755), .B2(n_694), .C1(n_604), .C2(n_687), .Y(n_757) );
AO221x1_ASAP7_75t_L g758 ( .A1(n_757), .A2(n_638), .B1(n_634), .B2(n_598), .C(n_594), .Y(n_758) );
AO21x2_ASAP7_75t_L g759 ( .A1(n_758), .A2(n_688), .B(n_638), .Y(n_759) );
AOI22xp5_ASAP7_75t_L g760 ( .A1(n_759), .A2(n_628), .B1(n_625), .B2(n_599), .Y(n_760) );
endmodule