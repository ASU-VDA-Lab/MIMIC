module fake_jpeg_30103_n_51 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_51);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_51;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_43;
wire n_50;
wire n_37;
wire n_32;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx11_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_19),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_23),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_0),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_18),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_25),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_1),
.Y(n_25)
);

INVx4_ASAP7_75t_SL g26 ( 
.A(n_20),
.Y(n_26)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_22),
.B(n_1),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_22),
.B(n_2),
.Y(n_28)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_21),
.B(n_17),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_SL g35 ( 
.A(n_31),
.B(n_16),
.Y(n_35)
);

AO22x1_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_16),
.B1(n_17),
.B2(n_10),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_38),
.B(n_4),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_34),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_32),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_33),
.C(n_30),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_29),
.A2(n_9),
.B1(n_12),
.B2(n_11),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_43),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_44),
.Y(n_46)
);

NOR2x1_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_3),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_42),
.B(n_4),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_7),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_45),
.A2(n_5),
.B(n_6),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_48),
.A2(n_47),
.B(n_46),
.Y(n_49)
);

BUFx24_ASAP7_75t_SL g50 ( 
.A(n_49),
.Y(n_50)
);

AOI32xp33_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_42),
.A3(n_46),
.B1(n_37),
.B2(n_14),
.Y(n_51)
);


endmodule