module fake_ariane_644_n_2171 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2171);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2171;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_899;
wire n_352;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2116;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_2168;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_2129;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1769;
wire n_1632;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2143;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_223;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_44),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_74),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_134),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_88),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_32),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_37),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_162),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_176),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_195),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_53),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_68),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_51),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_74),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_150),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_30),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_148),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_92),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_91),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_87),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_153),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_193),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_216),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_75),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_109),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_80),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_42),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_32),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_58),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_166),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_24),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_155),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_28),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_63),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_46),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_169),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_198),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_26),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_189),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_41),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_217),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_0),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_158),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_29),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_2),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_1),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_165),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_185),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_105),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_111),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_178),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_90),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_119),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_24),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_188),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_108),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_180),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_58),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_130),
.Y(n_276)
);

BUFx8_ASAP7_75t_SL g277 ( 
.A(n_55),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_206),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_142),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_37),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_204),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_200),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_13),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_182),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_201),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_126),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_186),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_41),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_135),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_159),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_139),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_213),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_207),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_172),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_101),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_190),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_209),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_51),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_57),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_218),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_6),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_202),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_1),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_7),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_125),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_16),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_13),
.Y(n_307)
);

BUFx5_ASAP7_75t_L g308 ( 
.A(n_100),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_113),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_133),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_97),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_114),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_71),
.Y(n_313)
);

BUFx10_ASAP7_75t_L g314 ( 
.A(n_20),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_129),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_157),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_2),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_140),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_28),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_147),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_6),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_146),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_76),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_141),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_127),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_66),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_167),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_99),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_168),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_21),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_117),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_59),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_81),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_116),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_104),
.Y(n_335)
);

INVxp33_ASAP7_75t_SL g336 ( 
.A(n_19),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_120),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_42),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_170),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_54),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_179),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_83),
.Y(n_342)
);

BUFx2_ASAP7_75t_SL g343 ( 
.A(n_26),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_106),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_191),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_138),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_103),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_79),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_31),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_66),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_5),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_123),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_214),
.Y(n_353)
);

INVxp67_ASAP7_75t_SL g354 ( 
.A(n_69),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_34),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_163),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_215),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_22),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_85),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_72),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_144),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_84),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_36),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_47),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_210),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_39),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_124),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_56),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_78),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_33),
.Y(n_370)
);

BUFx2_ASAP7_75t_SL g371 ( 
.A(n_36),
.Y(n_371)
);

BUFx5_ASAP7_75t_L g372 ( 
.A(n_212),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_112),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_154),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_38),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_3),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_44),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_54),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_16),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_10),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_96),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_77),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_205),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_110),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_35),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_23),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g387 ( 
.A(n_145),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_12),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_38),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_194),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_10),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_60),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_98),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_94),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_177),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_115),
.Y(n_396)
);

INVxp67_ASAP7_75t_SL g397 ( 
.A(n_149),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_22),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_67),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_48),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_173),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_61),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_199),
.Y(n_403)
);

BUFx10_ASAP7_75t_L g404 ( 
.A(n_187),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_69),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_102),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_72),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_174),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_208),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_11),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_70),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_95),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_121),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_45),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_93),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_86),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_197),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_107),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_175),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_17),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_11),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_156),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_183),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_59),
.Y(n_424)
);

CKINVDCx14_ASAP7_75t_R g425 ( 
.A(n_57),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_43),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_18),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_70),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_122),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_68),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_23),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_277),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_307),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_414),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_336),
.B(n_309),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_424),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_225),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_227),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_261),
.Y(n_439)
);

INVxp67_ASAP7_75t_SL g440 ( 
.A(n_231),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_261),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_425),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_236),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_261),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_333),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_242),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_247),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_261),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_261),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_256),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_389),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_389),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_335),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_381),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_224),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_219),
.Y(n_456)
);

OR2x2_ASAP7_75t_L g457 ( 
.A(n_245),
.B(n_0),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_262),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_220),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_389),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_389),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_389),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_336),
.B(n_3),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_263),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_343),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_398),
.Y(n_466)
);

INVx1_ASAP7_75t_SL g467 ( 
.A(n_230),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_398),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_398),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_398),
.Y(n_470)
);

NAND2xp33_ASAP7_75t_R g471 ( 
.A(n_328),
.B(n_82),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_398),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_338),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_246),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_338),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_379),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_255),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_271),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_379),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_220),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_426),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_426),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_235),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_280),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_288),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_301),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_237),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_237),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_253),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_253),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_315),
.Y(n_491)
);

INVxp67_ASAP7_75t_SL g492 ( 
.A(n_231),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_315),
.Y(n_493)
);

INVxp33_ASAP7_75t_SL g494 ( 
.A(n_223),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_314),
.B(n_4),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_235),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_304),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_373),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_286),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_286),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_275),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_373),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_371),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_306),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_364),
.Y(n_505)
);

INVxp67_ASAP7_75t_SL g506 ( 
.A(n_340),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_313),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_413),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_413),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_317),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_228),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_248),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_321),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_375),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_377),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_251),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_259),
.Y(n_517)
);

INVxp67_ASAP7_75t_SL g518 ( 
.A(n_340),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_283),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_391),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_332),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_298),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_327),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_374),
.B(n_4),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_299),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_385),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_410),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_349),
.Y(n_528)
);

INVxp33_ASAP7_75t_L g529 ( 
.A(n_303),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_319),
.Y(n_530)
);

INVxp67_ASAP7_75t_SL g531 ( 
.A(n_391),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_327),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_355),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_360),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_326),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_387),
.B(n_305),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_330),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_363),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_350),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_411),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_366),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_368),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_370),
.Y(n_543)
);

BUFx6f_ASAP7_75t_SL g544 ( 
.A(n_404),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_359),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_427),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_452),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_452),
.Y(n_548)
);

OAI21x1_ASAP7_75t_L g549 ( 
.A1(n_439),
.A2(n_232),
.B(n_226),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_439),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_441),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_496),
.B(n_418),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_441),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_520),
.B(n_404),
.Y(n_554)
);

OA21x2_ASAP7_75t_L g555 ( 
.A1(n_444),
.A2(n_241),
.B(n_238),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_444),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_448),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_448),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_496),
.B(n_243),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_499),
.B(n_249),
.Y(n_560)
);

NAND3xp33_ASAP7_75t_L g561 ( 
.A(n_471),
.B(n_358),
.C(n_351),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_449),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_449),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_451),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_433),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_451),
.Y(n_566)
);

AND2x2_ASAP7_75t_SL g567 ( 
.A(n_495),
.B(n_287),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_456),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_460),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_460),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_434),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_520),
.B(n_404),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_520),
.B(n_386),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_499),
.B(n_500),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_436),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_529),
.B(n_440),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_461),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_461),
.Y(n_578)
);

INVxp67_ASAP7_75t_L g579 ( 
.A(n_459),
.Y(n_579)
);

AND2x6_ASAP7_75t_L g580 ( 
.A(n_487),
.B(n_359),
.Y(n_580)
);

NAND2xp33_ASAP7_75t_R g581 ( 
.A(n_494),
.B(n_223),
.Y(n_581)
);

AND2x2_ASAP7_75t_R g582 ( 
.A(n_544),
.B(n_399),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_462),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_462),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_483),
.B(n_402),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_466),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_492),
.B(n_314),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_466),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_SL g589 ( 
.A(n_544),
.B(n_314),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_483),
.B(n_267),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_468),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_468),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_469),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_536),
.B(n_268),
.Y(n_594)
);

HB1xp67_ASAP7_75t_L g595 ( 
.A(n_480),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_469),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_506),
.B(n_221),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_470),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_545),
.B(n_270),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_470),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_472),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_472),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_500),
.B(n_272),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_487),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_488),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_488),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_518),
.B(n_221),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_523),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_531),
.B(n_222),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_489),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_489),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_490),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_458),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_490),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_435),
.B(n_545),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_491),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_491),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_523),
.B(n_279),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_442),
.B(n_222),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_493),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_532),
.B(n_511),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_493),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_464),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_498),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g625 ( 
.A(n_478),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_498),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_502),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_502),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_508),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_532),
.B(n_234),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_495),
.B(n_281),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_508),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_509),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_524),
.B(n_234),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_455),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_509),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_473),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_473),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_588),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_567),
.A2(n_463),
.B1(n_457),
.B2(n_544),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_556),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_556),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_588),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_556),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_554),
.B(n_445),
.Y(n_645)
);

INVx5_ASAP7_75t_L g646 ( 
.A(n_580),
.Y(n_646)
);

AND2x6_ASAP7_75t_L g647 ( 
.A(n_554),
.B(n_287),
.Y(n_647)
);

INVx4_ASAP7_75t_L g648 ( 
.A(n_567),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_597),
.B(n_484),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_588),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_634),
.B(n_485),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_558),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_567),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_567),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_631),
.B(n_457),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_588),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_588),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_588),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_597),
.B(n_486),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_596),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_611),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_597),
.B(n_497),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_558),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_631),
.B(n_511),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_596),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_634),
.B(n_507),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_607),
.B(n_510),
.Y(n_667)
);

XNOR2xp5_ASAP7_75t_L g668 ( 
.A(n_635),
.B(n_474),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_596),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_611),
.Y(n_670)
);

BUFx2_ASAP7_75t_L g671 ( 
.A(n_565),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_596),
.Y(n_672)
);

BUFx8_ASAP7_75t_SL g673 ( 
.A(n_635),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_611),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_596),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_631),
.B(n_512),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_596),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_607),
.B(n_513),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_576),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_554),
.B(n_521),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_550),
.Y(n_681)
);

INVx4_ASAP7_75t_L g682 ( 
.A(n_580),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_558),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_550),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_576),
.B(n_512),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_615),
.B(n_528),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_562),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_562),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_550),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_576),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_611),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_621),
.B(n_516),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_562),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_563),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_550),
.Y(n_695)
);

AND3x2_ASAP7_75t_L g696 ( 
.A(n_589),
.B(n_503),
.C(n_465),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_563),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_551),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_563),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_608),
.Y(n_700)
);

INVx4_ASAP7_75t_L g701 ( 
.A(n_580),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_566),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_566),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_571),
.B(n_575),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_551),
.Y(n_705)
);

INVx2_ASAP7_75t_SL g706 ( 
.A(n_607),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_611),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_611),
.Y(n_708)
);

BUFx10_ASAP7_75t_L g709 ( 
.A(n_615),
.Y(n_709)
);

INVxp67_ASAP7_75t_SL g710 ( 
.A(n_574),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_551),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_561),
.A2(n_594),
.B1(n_631),
.B2(n_630),
.Y(n_712)
);

INVx1_ASAP7_75t_SL g713 ( 
.A(n_565),
.Y(n_713)
);

INVx4_ASAP7_75t_L g714 ( 
.A(n_580),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_611),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_566),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_551),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_608),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_572),
.B(n_533),
.Y(n_719)
);

INVxp67_ASAP7_75t_L g720 ( 
.A(n_581),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_578),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_609),
.B(n_534),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_557),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_572),
.B(n_538),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_578),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_611),
.Y(n_726)
);

AND2x6_ASAP7_75t_L g727 ( 
.A(n_572),
.B(n_287),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_609),
.B(n_541),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_578),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_630),
.B(n_542),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_608),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_568),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_583),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_557),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_557),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_608),
.Y(n_736)
);

OR2x2_ASAP7_75t_L g737 ( 
.A(n_571),
.B(n_467),
.Y(n_737)
);

OR2x6_ASAP7_75t_L g738 ( 
.A(n_568),
.B(n_516),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_594),
.B(n_543),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_630),
.B(n_609),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_557),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_564),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_609),
.B(n_517),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_583),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_631),
.B(n_517),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_611),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_583),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_631),
.B(n_519),
.Y(n_748)
);

BUFx2_ASAP7_75t_L g749 ( 
.A(n_568),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_587),
.B(n_519),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_585),
.A2(n_580),
.B1(n_587),
.B2(n_555),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_604),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_584),
.Y(n_753)
);

INVx2_ASAP7_75t_SL g754 ( 
.A(n_587),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_621),
.B(n_522),
.Y(n_755)
);

AND2x2_ASAP7_75t_SL g756 ( 
.A(n_589),
.B(n_287),
.Y(n_756)
);

AND2x4_ASAP7_75t_L g757 ( 
.A(n_590),
.B(n_522),
.Y(n_757)
);

OR2x6_ASAP7_75t_L g758 ( 
.A(n_625),
.B(n_525),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_625),
.B(n_437),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_584),
.Y(n_760)
);

NAND2x1p5_ASAP7_75t_L g761 ( 
.A(n_555),
.B(n_289),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_584),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_625),
.B(n_438),
.Y(n_763)
);

NAND3xp33_ASAP7_75t_L g764 ( 
.A(n_612),
.B(n_293),
.C(n_292),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_590),
.B(n_525),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_604),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_604),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_621),
.Y(n_768)
);

OR2x6_ASAP7_75t_L g769 ( 
.A(n_574),
.B(n_530),
.Y(n_769)
);

NAND2xp33_ASAP7_75t_L g770 ( 
.A(n_613),
.B(n_239),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_604),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_619),
.Y(n_772)
);

INVx2_ASAP7_75t_SL g773 ( 
.A(n_619),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_573),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_579),
.B(n_443),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_619),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_605),
.Y(n_777)
);

INVx5_ASAP7_75t_L g778 ( 
.A(n_580),
.Y(n_778)
);

INVx2_ASAP7_75t_SL g779 ( 
.A(n_590),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_590),
.Y(n_780)
);

NAND2xp33_ASAP7_75t_L g781 ( 
.A(n_613),
.B(n_239),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_605),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_605),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_612),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_564),
.Y(n_785)
);

AND2x2_ASAP7_75t_SL g786 ( 
.A(n_555),
.B(n_287),
.Y(n_786)
);

OR2x6_ASAP7_75t_L g787 ( 
.A(n_623),
.B(n_530),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_605),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_606),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_623),
.B(n_447),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_564),
.Y(n_791)
);

INVx3_ASAP7_75t_L g792 ( 
.A(n_606),
.Y(n_792)
);

OAI22xp33_ASAP7_75t_L g793 ( 
.A1(n_579),
.A2(n_428),
.B1(n_229),
.B2(n_407),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_648),
.B(n_590),
.Y(n_794)
);

NAND2xp33_ASAP7_75t_L g795 ( 
.A(n_680),
.B(n_719),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_752),
.Y(n_796)
);

INVx2_ASAP7_75t_SL g797 ( 
.A(n_737),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_784),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_784),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_739),
.B(n_595),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_641),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_648),
.B(n_756),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_641),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_686),
.B(n_590),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_756),
.A2(n_580),
.B1(n_555),
.B2(n_599),
.Y(n_805)
);

INVxp67_ASAP7_75t_L g806 ( 
.A(n_737),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_712),
.B(n_599),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_710),
.B(n_599),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_642),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_706),
.B(n_599),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_706),
.B(n_679),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_679),
.B(n_599),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_648),
.A2(n_599),
.B1(n_573),
.B2(n_580),
.Y(n_813)
);

NOR3xp33_ASAP7_75t_L g814 ( 
.A(n_713),
.B(n_454),
.C(n_354),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_752),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_690),
.B(n_573),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_709),
.B(n_552),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_740),
.B(n_552),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_749),
.B(n_575),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_648),
.B(n_756),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_754),
.B(n_585),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_754),
.B(n_585),
.Y(n_822)
);

NOR3xp33_ASAP7_75t_L g823 ( 
.A(n_775),
.B(n_432),
.C(n_233),
.Y(n_823)
);

OAI21xp5_ASAP7_75t_L g824 ( 
.A1(n_786),
.A2(n_549),
.B(n_555),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_709),
.B(n_240),
.Y(n_825)
);

NOR2xp67_ASAP7_75t_SL g826 ( 
.A(n_774),
.B(n_244),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_709),
.B(n_240),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_642),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_787),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_709),
.B(n_254),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_752),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_720),
.B(n_254),
.Y(n_832)
);

NOR2xp67_ASAP7_75t_L g833 ( 
.A(n_645),
.B(n_612),
.Y(n_833)
);

HB1xp67_ASAP7_75t_L g834 ( 
.A(n_738),
.Y(n_834)
);

NAND2x1_ASAP7_75t_L g835 ( 
.A(n_682),
.B(n_580),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_749),
.B(n_585),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_774),
.B(n_585),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_644),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_653),
.A2(n_580),
.B1(n_585),
.B2(n_397),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_783),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_653),
.B(n_258),
.Y(n_841)
);

NAND2xp33_ASAP7_75t_SL g842 ( 
.A(n_724),
.B(n_244),
.Y(n_842)
);

BUFx6f_ASAP7_75t_SL g843 ( 
.A(n_738),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_654),
.A2(n_651),
.B1(n_666),
.B2(n_640),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_644),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_673),
.Y(n_846)
);

INVx4_ASAP7_75t_L g847 ( 
.A(n_787),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_652),
.Y(n_848)
);

NAND2xp33_ASAP7_75t_L g849 ( 
.A(n_670),
.B(n_580),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_654),
.B(n_258),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_774),
.B(n_559),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_685),
.B(n_559),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_682),
.B(n_260),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_783),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_682),
.B(n_260),
.Y(n_855)
);

NAND3xp33_ASAP7_75t_SL g856 ( 
.A(n_732),
.B(n_450),
.C(n_446),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_682),
.B(n_382),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_652),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_685),
.B(n_560),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_783),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_743),
.B(n_560),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_671),
.B(n_453),
.Y(n_862)
);

AOI221xp5_ASAP7_75t_L g863 ( 
.A1(n_793),
.A2(n_407),
.B1(n_405),
.B2(n_400),
.C(n_392),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_730),
.B(n_603),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_792),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_664),
.B(n_603),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_769),
.A2(n_580),
.B1(n_555),
.B2(n_618),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_701),
.B(n_382),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_664),
.B(n_618),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_L g870 ( 
.A1(n_772),
.A2(n_620),
.B1(n_622),
.B2(n_617),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_671),
.B(n_477),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_792),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_SL g873 ( 
.A(n_738),
.B(n_501),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_664),
.B(n_617),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_792),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_663),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_681),
.Y(n_877)
);

OAI221xp5_ASAP7_75t_L g878 ( 
.A1(n_772),
.A2(n_421),
.B1(n_257),
.B2(n_252),
.C(n_250),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_664),
.B(n_617),
.Y(n_879)
);

INVx4_ASAP7_75t_L g880 ( 
.A(n_787),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_676),
.B(n_637),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_773),
.B(n_384),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_676),
.B(n_620),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_681),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_684),
.Y(n_885)
);

AND2x6_ASAP7_75t_SL g886 ( 
.A(n_738),
.B(n_758),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_684),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_676),
.B(n_622),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_676),
.B(n_627),
.Y(n_889)
);

AND2x4_ASAP7_75t_L g890 ( 
.A(n_787),
.B(n_637),
.Y(n_890)
);

NAND2xp33_ASAP7_75t_SL g891 ( 
.A(n_776),
.B(n_250),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_655),
.B(n_627),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_738),
.B(n_504),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_701),
.B(n_714),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_722),
.B(n_628),
.Y(n_895)
);

AOI22xp5_ASAP7_75t_L g896 ( 
.A1(n_776),
.A2(n_633),
.B1(n_628),
.B2(n_390),
.Y(n_896)
);

NOR2x1p5_ASAP7_75t_L g897 ( 
.A(n_704),
.B(n_252),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_728),
.B(n_628),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_701),
.B(n_384),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_649),
.B(n_633),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_718),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_663),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_689),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_683),
.Y(n_904)
);

OAI221xp5_ASAP7_75t_L g905 ( 
.A1(n_750),
.A2(n_420),
.B1(n_257),
.B2(n_430),
.C(n_378),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_655),
.B(n_633),
.Y(n_906)
);

NOR3xp33_ASAP7_75t_L g907 ( 
.A(n_770),
.B(n_380),
.C(n_378),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_659),
.B(n_637),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_655),
.B(n_638),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_655),
.B(n_638),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_689),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_692),
.B(n_638),
.Y(n_912)
);

INVxp67_ASAP7_75t_L g913 ( 
.A(n_668),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_758),
.B(n_505),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_692),
.B(n_606),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_683),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_755),
.B(n_606),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_687),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_662),
.B(n_636),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_667),
.B(n_636),
.Y(n_920)
);

INVx4_ASAP7_75t_L g921 ( 
.A(n_787),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_700),
.Y(n_922)
);

OR2x6_ASAP7_75t_L g923 ( 
.A(n_758),
.B(n_582),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_687),
.Y(n_924)
);

A2O1A1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_745),
.A2(n_549),
.B(n_632),
.C(n_629),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_695),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_695),
.Y(n_927)
);

AOI22xp33_ASAP7_75t_L g928 ( 
.A1(n_769),
.A2(n_624),
.B1(n_632),
.B2(n_629),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_701),
.B(n_390),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_755),
.B(n_610),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_768),
.B(n_610),
.Y(n_931)
);

NAND2xp33_ASAP7_75t_L g932 ( 
.A(n_670),
.B(n_393),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_688),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_698),
.Y(n_934)
);

NOR2xp67_ASAP7_75t_L g935 ( 
.A(n_704),
.B(n_764),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_688),
.Y(n_936)
);

BUFx8_ASAP7_75t_L g937 ( 
.A(n_757),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_768),
.B(n_610),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_698),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_714),
.B(n_393),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_678),
.B(n_610),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_758),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_693),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_705),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_768),
.B(n_636),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_748),
.B(n_614),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_693),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_769),
.B(n_614),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_718),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_769),
.B(n_614),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_705),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_769),
.B(n_636),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_757),
.B(n_614),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_696),
.B(n_632),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_668),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_759),
.B(n_514),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_694),
.Y(n_957)
);

AOI22xp33_ASAP7_75t_L g958 ( 
.A1(n_751),
.A2(n_632),
.B1(n_629),
.B2(n_626),
.Y(n_958)
);

AO221x1_ASAP7_75t_L g959 ( 
.A1(n_781),
.A2(n_582),
.B1(n_394),
.B2(n_294),
.C(n_416),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_779),
.B(n_616),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_763),
.B(n_515),
.Y(n_961)
);

OAI21xp5_ASAP7_75t_L g962 ( 
.A1(n_925),
.A2(n_786),
.B(n_697),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_824),
.A2(n_864),
.B(n_952),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_861),
.A2(n_643),
.B(n_639),
.Y(n_964)
);

NAND2x1p5_ASAP7_75t_L g965 ( 
.A(n_847),
.B(n_880),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_864),
.B(n_757),
.Y(n_966)
);

AOI22xp33_ASAP7_75t_L g967 ( 
.A1(n_802),
.A2(n_786),
.B1(n_764),
.B2(n_727),
.Y(n_967)
);

O2A1O1Ixp5_ASAP7_75t_L g968 ( 
.A1(n_804),
.A2(n_697),
.B(n_699),
.C(n_694),
.Y(n_968)
);

OAI21xp5_ASAP7_75t_L g969 ( 
.A1(n_952),
.A2(n_702),
.B(n_699),
.Y(n_969)
);

A2O1A1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_800),
.A2(n_780),
.B(n_779),
.C(n_639),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_800),
.B(n_790),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_796),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_795),
.A2(n_650),
.B(n_643),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_817),
.B(n_757),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_901),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_815),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_881),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_817),
.B(n_780),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_901),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_818),
.B(n_852),
.Y(n_980)
);

AOI22x1_ASAP7_75t_L g981 ( 
.A1(n_801),
.A2(n_703),
.B1(n_716),
.B2(n_702),
.Y(n_981)
);

AO21x1_ASAP7_75t_L g982 ( 
.A1(n_844),
.A2(n_761),
.B(n_716),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_859),
.B(n_647),
.Y(n_983)
);

NOR2xp67_ASAP7_75t_L g984 ( 
.A(n_806),
.B(n_765),
.Y(n_984)
);

NOR2x1p5_ASAP7_75t_SL g985 ( 
.A(n_815),
.B(n_650),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_866),
.B(n_647),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_847),
.B(n_700),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_869),
.B(n_647),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_881),
.Y(n_989)
);

NOR3xp33_ASAP7_75t_L g990 ( 
.A(n_905),
.B(n_537),
.C(n_535),
.Y(n_990)
);

AOI22xp5_ASAP7_75t_L g991 ( 
.A1(n_942),
.A2(n_727),
.B1(n_647),
.B2(n_718),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_946),
.A2(n_657),
.B(n_656),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_881),
.B(n_647),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_803),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_853),
.A2(n_657),
.B(n_656),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_SL g996 ( 
.A1(n_893),
.A2(n_527),
.B1(n_540),
.B2(n_526),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_890),
.A2(n_828),
.B1(n_838),
.B2(n_809),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_880),
.B(n_731),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_921),
.B(n_731),
.Y(n_999)
);

OAI21xp33_ASAP7_75t_L g1000 ( 
.A1(n_863),
.A2(n_388),
.B(n_380),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_921),
.B(n_731),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_853),
.A2(n_660),
.B(n_658),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_829),
.B(n_714),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_855),
.A2(n_660),
.B(n_658),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_890),
.B(n_714),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_855),
.A2(n_669),
.B(n_665),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_895),
.A2(n_669),
.B(n_672),
.C(n_665),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_811),
.B(n_647),
.Y(n_1008)
);

OAI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_948),
.A2(n_721),
.B(n_703),
.Y(n_1009)
);

AOI33xp33_ASAP7_75t_L g1010 ( 
.A1(n_819),
.A2(n_539),
.A3(n_537),
.B1(n_535),
.B2(n_729),
.B3(n_753),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_851),
.B(n_647),
.Y(n_1011)
);

NOR3xp33_ASAP7_75t_L g1012 ( 
.A(n_878),
.B(n_539),
.C(n_431),
.Y(n_1012)
);

BUFx8_ASAP7_75t_L g1013 ( 
.A(n_843),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_797),
.B(n_546),
.Y(n_1014)
);

AOI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_843),
.A2(n_727),
.B1(n_736),
.B2(n_725),
.Y(n_1015)
);

INVx4_ASAP7_75t_L g1016 ( 
.A(n_886),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_845),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_857),
.A2(n_675),
.B(n_672),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_834),
.B(n_736),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_833),
.B(n_727),
.Y(n_1020)
);

OAI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_950),
.A2(n_725),
.B(n_721),
.Y(n_1021)
);

OR2x2_ASAP7_75t_L g1022 ( 
.A(n_871),
.B(n_766),
.Y(n_1022)
);

OAI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_945),
.A2(n_733),
.B(n_729),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_857),
.A2(n_677),
.B(n_675),
.Y(n_1024)
);

NOR3xp33_ASAP7_75t_SL g1025 ( 
.A(n_825),
.B(n_392),
.C(n_388),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_848),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_890),
.B(n_727),
.Y(n_1027)
);

NOR2xp67_ASAP7_75t_L g1028 ( 
.A(n_856),
.B(n_616),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_895),
.B(n_727),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_935),
.B(n_937),
.Y(n_1030)
);

INVx1_ASAP7_75t_SL g1031 ( 
.A(n_862),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_868),
.A2(n_677),
.B(n_674),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_868),
.A2(n_674),
.B(n_661),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_899),
.A2(n_674),
.B(n_661),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_858),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_876),
.A2(n_744),
.B1(n_747),
.B2(n_733),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_898),
.B(n_727),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_831),
.Y(n_1038)
);

AOI33xp33_ASAP7_75t_L g1039 ( 
.A1(n_836),
.A2(n_744),
.A3(n_760),
.B1(n_762),
.B2(n_747),
.B3(n_753),
.Y(n_1039)
);

OAI321xp33_ASAP7_75t_L g1040 ( 
.A1(n_825),
.A2(n_482),
.A3(n_476),
.B1(n_475),
.B2(n_481),
.C(n_479),
.Y(n_1040)
);

NOR3xp33_ASAP7_75t_L g1041 ( 
.A(n_842),
.B(n_376),
.C(n_400),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_937),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_832),
.B(n_736),
.Y(n_1043)
);

AOI21xp33_ASAP7_75t_L g1044 ( 
.A1(n_954),
.A2(n_762),
.B(n_760),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_902),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_899),
.A2(n_691),
.B(n_661),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_904),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_916),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_827),
.A2(n_771),
.B1(n_789),
.B2(n_788),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_901),
.B(n_646),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_918),
.Y(n_1051)
);

NAND2x1p5_ASAP7_75t_L g1052 ( 
.A(n_802),
.B(n_646),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_898),
.A2(n_766),
.B(n_789),
.C(n_788),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_929),
.A2(n_707),
.B(n_691),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_831),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_929),
.A2(n_707),
.B(n_691),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_914),
.B(n_475),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_840),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_949),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_940),
.A2(n_708),
.B(n_707),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_940),
.A2(n_715),
.B(n_708),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_840),
.A2(n_715),
.B(n_708),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_949),
.Y(n_1063)
);

CKINVDCx8_ASAP7_75t_R g1064 ( 
.A(n_846),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_854),
.Y(n_1065)
);

AOI21x1_ASAP7_75t_L g1066 ( 
.A1(n_820),
.A2(n_771),
.B(n_767),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_949),
.B(n_873),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_854),
.A2(n_726),
.B(n_715),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_860),
.A2(n_746),
.B(n_726),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_860),
.A2(n_746),
.B(n_726),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_832),
.B(n_767),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_827),
.B(n_777),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_900),
.B(n_777),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_900),
.B(n_782),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_865),
.A2(n_746),
.B(n_782),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_830),
.B(n_761),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_865),
.A2(n_670),
.B(n_711),
.Y(n_1077)
);

OAI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_945),
.A2(n_761),
.B(n_791),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_908),
.B(n_711),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_872),
.A2(n_670),
.B(n_717),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_872),
.A2(n_670),
.B(n_717),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_875),
.A2(n_734),
.B(n_723),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_875),
.A2(n_734),
.B(n_723),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_908),
.B(n_735),
.Y(n_1084)
);

AOI21x1_ASAP7_75t_L g1085 ( 
.A1(n_820),
.A2(n_741),
.B(n_735),
.Y(n_1085)
);

OAI321xp33_ASAP7_75t_L g1086 ( 
.A1(n_830),
.A2(n_481),
.A3(n_479),
.B1(n_482),
.B2(n_616),
.C(n_629),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_894),
.A2(n_742),
.B(n_741),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_892),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_956),
.B(n_624),
.Y(n_1089)
);

OAI321xp33_ASAP7_75t_L g1090 ( 
.A1(n_896),
.A2(n_624),
.A3(n_626),
.B1(n_297),
.B2(n_383),
.C(n_323),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_894),
.A2(n_785),
.B(n_742),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_SL g1092 ( 
.A1(n_924),
.A2(n_791),
.B(n_785),
.C(n_422),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_919),
.A2(n_549),
.B(n_624),
.C(n_626),
.Y(n_1093)
);

O2A1O1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_915),
.A2(n_626),
.B(n_300),
.C(n_324),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_816),
.B(n_405),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_919),
.B(n_420),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_933),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_931),
.A2(n_778),
.B(n_646),
.Y(n_1098)
);

O2A1O1Ixp5_ASAP7_75t_L g1099 ( 
.A1(n_960),
.A2(n_602),
.B(n_569),
.C(n_564),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_920),
.A2(n_941),
.B(n_960),
.C(n_943),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_906),
.B(n_430),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_909),
.B(n_646),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_936),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_910),
.B(n_646),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_SL g1105 ( 
.A(n_923),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_938),
.A2(n_778),
.B(n_646),
.Y(n_1106)
);

NOR3xp33_ASAP7_75t_L g1107 ( 
.A(n_907),
.B(n_348),
.C(n_346),
.Y(n_1107)
);

AOI21x1_ASAP7_75t_L g1108 ( 
.A1(n_947),
.A2(n_549),
.B(n_569),
.Y(n_1108)
);

NOR2xp67_ASAP7_75t_L g1109 ( 
.A(n_913),
.B(n_547),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_912),
.B(n_778),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_957),
.A2(n_778),
.B1(n_352),
.B2(n_353),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_920),
.A2(n_417),
.B(n_401),
.C(n_357),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_917),
.A2(n_778),
.B(n_396),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_874),
.A2(n_879),
.B1(n_883),
.B2(n_888),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_930),
.A2(n_808),
.B(n_953),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_835),
.A2(n_778),
.B(n_396),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_949),
.Y(n_1117)
);

INVx2_ASAP7_75t_SL g1118 ( 
.A(n_955),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_889),
.B(n_395),
.Y(n_1119)
);

O2A1O1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_837),
.A2(n_602),
.B(n_593),
.C(n_586),
.Y(n_1120)
);

CKINVDCx8_ASAP7_75t_R g1121 ( 
.A(n_923),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_870),
.B(n_395),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_R g1123 ( 
.A(n_891),
.B(n_403),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_877),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_821),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_841),
.A2(n_412),
.B1(n_429),
.B2(n_423),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_884),
.A2(n_406),
.B(n_403),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_884),
.A2(n_408),
.B(n_406),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_885),
.A2(n_409),
.B(n_408),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_885),
.A2(n_412),
.B(n_409),
.Y(n_1130)
);

BUFx4f_ASAP7_75t_L g1131 ( 
.A(n_961),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_887),
.A2(n_911),
.B(n_903),
.Y(n_1132)
);

OAI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_941),
.A2(n_602),
.B(n_593),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_887),
.A2(n_415),
.B(n_429),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_903),
.A2(n_419),
.B(n_423),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_810),
.B(n_419),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_911),
.A2(n_334),
.B(n_265),
.Y(n_1137)
);

AO21x1_ASAP7_75t_L g1138 ( 
.A1(n_841),
.A2(n_602),
.B(n_586),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_798),
.B(n_264),
.Y(n_1139)
);

INVx3_ASAP7_75t_L g1140 ( 
.A(n_922),
.Y(n_1140)
);

HB1xp67_ASAP7_75t_L g1141 ( 
.A(n_794),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_926),
.A2(n_337),
.B(n_269),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_822),
.B(n_812),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_897),
.B(n_547),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_926),
.A2(n_570),
.B(n_586),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_927),
.A2(n_339),
.B(n_273),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_966),
.A2(n_799),
.B1(n_813),
.B2(n_794),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_994),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_963),
.B(n_922),
.Y(n_1149)
);

INVx4_ASAP7_75t_L g1150 ( 
.A(n_965),
.Y(n_1150)
);

AND2x4_ASAP7_75t_L g1151 ( 
.A(n_977),
.B(n_954),
.Y(n_1151)
);

A2O1A1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_971),
.A2(n_850),
.B(n_823),
.C(n_807),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_971),
.B(n_980),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_974),
.B(n_882),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1017),
.Y(n_1155)
);

AOI21xp33_ASAP7_75t_L g1156 ( 
.A1(n_1096),
.A2(n_850),
.B(n_805),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1100),
.A2(n_932),
.B(n_849),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1115),
.A2(n_939),
.B(n_927),
.Y(n_1158)
);

AOI22x1_ASAP7_75t_L g1159 ( 
.A1(n_973),
.A2(n_934),
.B1(n_951),
.B2(n_944),
.Y(n_1159)
);

AO21x1_ASAP7_75t_L g1160 ( 
.A1(n_1076),
.A2(n_934),
.B(n_951),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_1064),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1088),
.B(n_814),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_1076),
.B(n_939),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1023),
.A2(n_944),
.B(n_867),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_978),
.B(n_928),
.Y(n_1165)
);

OAI221xp5_ASAP7_75t_L g1166 ( 
.A1(n_1000),
.A2(n_826),
.B1(n_839),
.B2(n_958),
.C(n_302),
.Y(n_1166)
);

A2O1A1Ixp33_ASAP7_75t_SL g1167 ( 
.A1(n_978),
.A2(n_593),
.B(n_586),
.C(n_570),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_997),
.B(n_553),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1026),
.Y(n_1169)
);

INVx1_ASAP7_75t_SL g1170 ( 
.A(n_1014),
.Y(n_1170)
);

O2A1O1Ixp5_ASAP7_75t_L g1171 ( 
.A1(n_1138),
.A2(n_569),
.B(n_593),
.C(n_570),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_975),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1035),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_1031),
.B(n_266),
.Y(n_1174)
);

NAND3xp33_ASAP7_75t_SL g1175 ( 
.A(n_1012),
.B(n_325),
.C(n_274),
.Y(n_1175)
);

AOI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1096),
.A2(n_959),
.B1(n_344),
.B2(n_342),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1045),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1073),
.A2(n_345),
.B(n_278),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1088),
.B(n_569),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1131),
.B(n_276),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_1013),
.Y(n_1181)
);

OR2x2_ASAP7_75t_L g1182 ( 
.A(n_1118),
.B(n_547),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_1042),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_989),
.B(n_282),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_984),
.B(n_284),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1124),
.Y(n_1186)
);

O2A1O1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1012),
.A2(n_570),
.B(n_547),
.C(n_548),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1089),
.B(n_547),
.Y(n_1188)
);

A2O1A1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_1072),
.A2(n_547),
.B(n_548),
.C(n_598),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1072),
.A2(n_548),
.B(n_600),
.C(n_598),
.Y(n_1190)
);

O2A1O1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_990),
.A2(n_548),
.B(n_7),
.C(n_8),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_968),
.A2(n_341),
.B(n_290),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1047),
.Y(n_1193)
);

NAND3xp33_ASAP7_75t_L g1194 ( 
.A(n_1107),
.B(n_990),
.C(n_1112),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1085),
.A2(n_981),
.B(n_1066),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_SL g1196 ( 
.A(n_1016),
.B(n_285),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_975),
.Y(n_1197)
);

HB1xp67_ASAP7_75t_L g1198 ( 
.A(n_1141),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1141),
.B(n_8),
.Y(n_1199)
);

O2A1O1Ixp33_ASAP7_75t_SL g1200 ( 
.A1(n_970),
.A2(n_9),
.B(n_12),
.C(n_14),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1048),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_R g1202 ( 
.A(n_1121),
.B(n_291),
.Y(n_1202)
);

AOI21x1_ASAP7_75t_L g1203 ( 
.A1(n_982),
.A2(n_601),
.B(n_600),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1051),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1114),
.A2(n_356),
.B1(n_312),
.B2(n_316),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1057),
.B(n_9),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1074),
.A2(n_362),
.B(n_295),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1125),
.B(n_14),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_972),
.Y(n_1209)
);

INVxp67_ASAP7_75t_L g1210 ( 
.A(n_1019),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_962),
.A2(n_365),
.B(n_296),
.Y(n_1211)
);

CKINVDCx14_ASAP7_75t_R g1212 ( 
.A(n_1123),
.Y(n_1212)
);

NOR3xp33_ASAP7_75t_SL g1213 ( 
.A(n_1095),
.B(n_310),
.C(n_311),
.Y(n_1213)
);

A2O1A1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1071),
.A2(n_601),
.B(n_600),
.C(n_598),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_975),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_1030),
.B(n_1016),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_969),
.A2(n_369),
.B(n_320),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_1022),
.B(n_15),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1143),
.A2(n_322),
.B(n_329),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_976),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_SL g1221 ( 
.A(n_1019),
.B(n_331),
.Y(n_1221)
);

AND2x4_ASAP7_75t_L g1222 ( 
.A(n_1067),
.B(n_553),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1038),
.Y(n_1223)
);

INVx2_ASAP7_75t_SL g1224 ( 
.A(n_996),
.Y(n_1224)
);

NAND3xp33_ASAP7_75t_L g1225 ( 
.A(n_1107),
.B(n_601),
.C(n_600),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1078),
.A2(n_347),
.B(n_361),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1101),
.B(n_1010),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_964),
.A2(n_367),
.B(n_318),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1055),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_SL g1230 ( 
.A(n_1009),
.B(n_1021),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_SL g1231 ( 
.A(n_1044),
.B(n_553),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1097),
.B(n_17),
.Y(n_1232)
);

A2O1A1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1071),
.A2(n_601),
.B(n_600),
.C(n_598),
.Y(n_1233)
);

AOI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_998),
.A2(n_601),
.B1(n_600),
.B2(n_598),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1103),
.A2(n_601),
.B1(n_600),
.B2(n_598),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_SL g1236 ( 
.A(n_998),
.B(n_553),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_968),
.A2(n_294),
.B(n_318),
.Y(n_1237)
);

AO21x1_ASAP7_75t_L g1238 ( 
.A1(n_1043),
.A2(n_308),
.B(n_372),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1039),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1144),
.Y(n_1240)
);

CKINVDCx14_ASAP7_75t_R g1241 ( 
.A(n_975),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1036),
.A2(n_294),
.B(n_318),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_992),
.A2(n_1084),
.B(n_1079),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1058),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_999),
.B(n_553),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_1025),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1110),
.A2(n_294),
.B(n_318),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1087),
.A2(n_294),
.B(n_318),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1025),
.B(n_19),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1091),
.A2(n_394),
.B(n_416),
.Y(n_1250)
);

A2O1A1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1043),
.A2(n_601),
.B(n_600),
.C(n_598),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1065),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1028),
.A2(n_601),
.B1(n_600),
.B2(n_598),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1029),
.A2(n_553),
.B(n_598),
.C(n_592),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_1105),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_999),
.B(n_601),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1062),
.A2(n_416),
.B(n_394),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_SL g1258 ( 
.A(n_1105),
.B(n_592),
.Y(n_1258)
);

AOI21x1_ASAP7_75t_L g1259 ( 
.A1(n_995),
.A2(n_592),
.B(n_591),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1068),
.A2(n_416),
.B(n_394),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1109),
.B(n_20),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1069),
.A2(n_416),
.B(n_394),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_1139),
.Y(n_1263)
);

NAND2xp33_ASAP7_75t_L g1264 ( 
.A(n_979),
.B(n_372),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1070),
.A2(n_592),
.B(n_591),
.Y(n_1265)
);

NAND3xp33_ASAP7_75t_SL g1266 ( 
.A(n_1041),
.B(n_21),
.C(n_25),
.Y(n_1266)
);

OAI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1119),
.A2(n_591),
.B1(n_577),
.B2(n_553),
.Y(n_1267)
);

OAI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1136),
.A2(n_591),
.B1(n_577),
.B2(n_553),
.Y(n_1268)
);

INVx3_ASAP7_75t_L g1269 ( 
.A(n_965),
.Y(n_1269)
);

INVx1_ASAP7_75t_SL g1270 ( 
.A(n_1027),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_987),
.B(n_25),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_987),
.B(n_27),
.Y(n_1272)
);

INVx2_ASAP7_75t_SL g1273 ( 
.A(n_979),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1049),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_979),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1145),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1140),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1140),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1001),
.A2(n_592),
.B1(n_591),
.B2(n_577),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1001),
.B(n_27),
.Y(n_1280)
);

AO22x1_ASAP7_75t_L g1281 ( 
.A1(n_1041),
.A2(n_592),
.B1(n_591),
.B2(n_577),
.Y(n_1281)
);

O2A1O1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_1122),
.A2(n_29),
.B(n_30),
.C(n_33),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1075),
.A2(n_592),
.B(n_591),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1007),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1032),
.A2(n_592),
.B(n_591),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1063),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1033),
.A2(n_592),
.B(n_591),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_SL g1288 ( 
.A(n_993),
.B(n_577),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1034),
.A2(n_577),
.B(n_553),
.Y(n_1289)
);

NAND2xp33_ASAP7_75t_L g1290 ( 
.A(n_979),
.B(n_372),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1005),
.B(n_34),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_SL g1292 ( 
.A(n_1059),
.B(n_577),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1126),
.B(n_39),
.Y(n_1293)
);

INVx3_ASAP7_75t_L g1294 ( 
.A(n_1059),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1063),
.B(n_40),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_SL g1296 ( 
.A(n_1059),
.B(n_577),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_SL g1297 ( 
.A(n_1037),
.B(n_577),
.Y(n_1297)
);

BUFx6f_ASAP7_75t_L g1298 ( 
.A(n_1059),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1053),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1120),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1117),
.Y(n_1301)
);

AO21x2_ASAP7_75t_L g1302 ( 
.A1(n_1160),
.A2(n_1093),
.B(n_1133),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1148),
.Y(n_1303)
);

AO31x2_ASAP7_75t_L g1304 ( 
.A1(n_1238),
.A2(n_1164),
.A3(n_1243),
.B(n_1254),
.Y(n_1304)
);

NAND2x1p5_ASAP7_75t_L g1305 ( 
.A(n_1161),
.B(n_1117),
.Y(n_1305)
);

BUFx4_ASAP7_75t_SL g1306 ( 
.A(n_1181),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1195),
.A2(n_1132),
.B(n_1004),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1153),
.B(n_983),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1155),
.Y(n_1309)
);

AO31x2_ASAP7_75t_L g1310 ( 
.A1(n_1251),
.A2(n_1018),
.A3(n_1002),
.B(n_1006),
.Y(n_1310)
);

BUFx12f_ASAP7_75t_L g1311 ( 
.A(n_1255),
.Y(n_1311)
);

AOI31xp67_ASAP7_75t_L g1312 ( 
.A1(n_1230),
.A2(n_1149),
.A3(n_1168),
.B(n_1231),
.Y(n_1312)
);

AND2x4_ASAP7_75t_L g1313 ( 
.A(n_1151),
.B(n_1015),
.Y(n_1313)
);

A2O1A1Ixp33_ASAP7_75t_L g1314 ( 
.A1(n_1152),
.A2(n_1194),
.B(n_1156),
.C(n_1154),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1210),
.B(n_967),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1230),
.A2(n_1056),
.B(n_1046),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1206),
.B(n_40),
.Y(n_1317)
);

NOR2xp33_ASAP7_75t_L g1318 ( 
.A(n_1240),
.B(n_1040),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_1212),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1183),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_1216),
.Y(n_1321)
);

O2A1O1Ixp33_ASAP7_75t_SL g1322 ( 
.A1(n_1165),
.A2(n_1008),
.B(n_988),
.C(n_986),
.Y(n_1322)
);

A2O1A1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1154),
.A2(n_1090),
.B(n_1094),
.C(n_1086),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1210),
.B(n_967),
.Y(n_1324)
);

NOR2xp67_ASAP7_75t_L g1325 ( 
.A(n_1150),
.B(n_991),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1259),
.A2(n_1024),
.B(n_1108),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1157),
.A2(n_1054),
.B(n_1061),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_1216),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1165),
.A2(n_1060),
.B(n_1081),
.Y(n_1329)
);

OA21x2_ASAP7_75t_L g1330 ( 
.A1(n_1171),
.A2(n_1099),
.B(n_1080),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_1198),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1147),
.A2(n_1077),
.B(n_1011),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1158),
.A2(n_1092),
.B(n_1099),
.Y(n_1333)
);

AND2x4_ASAP7_75t_L g1334 ( 
.A(n_1151),
.B(n_985),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1170),
.B(n_1127),
.Y(n_1335)
);

BUFx2_ASAP7_75t_L g1336 ( 
.A(n_1241),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1169),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1218),
.B(n_1128),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1246),
.B(n_1129),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1173),
.Y(n_1340)
);

AO31x2_ASAP7_75t_L g1341 ( 
.A1(n_1237),
.A2(n_1247),
.A3(n_1214),
.B(n_1233),
.Y(n_1341)
);

AO31x2_ASAP7_75t_L g1342 ( 
.A1(n_1190),
.A2(n_1113),
.A3(n_1082),
.B(n_1083),
.Y(n_1342)
);

OR2x2_ASAP7_75t_L g1343 ( 
.A(n_1162),
.B(n_1134),
.Y(n_1343)
);

O2A1O1Ixp33_ASAP7_75t_SL g1344 ( 
.A1(n_1280),
.A2(n_1020),
.B(n_1102),
.C(n_1104),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1297),
.A2(n_1098),
.B(n_1106),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1186),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1276),
.A2(n_1116),
.B(n_1050),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1177),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1299),
.A2(n_1146),
.B(n_1142),
.Y(n_1349)
);

INVx5_ASAP7_75t_L g1350 ( 
.A(n_1172),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1171),
.A2(n_1135),
.B(n_1130),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1263),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1159),
.A2(n_1203),
.B(n_1248),
.Y(n_1353)
);

A2O1A1Ixp33_ASAP7_75t_L g1354 ( 
.A1(n_1208),
.A2(n_1111),
.B(n_1137),
.C(n_1003),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1209),
.Y(n_1355)
);

AOI221xp5_ASAP7_75t_L g1356 ( 
.A1(n_1218),
.A2(n_1052),
.B1(n_45),
.B2(n_46),
.C(n_47),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1274),
.A2(n_1052),
.B(n_372),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1193),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1167),
.A2(n_131),
.B(n_211),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1250),
.A2(n_372),
.B(n_308),
.Y(n_1360)
);

BUFx3_ASAP7_75t_L g1361 ( 
.A(n_1224),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1167),
.A2(n_128),
.B(n_203),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1285),
.A2(n_372),
.B(n_308),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1174),
.B(n_1198),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1201),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1257),
.A2(n_372),
.B(n_308),
.Y(n_1366)
);

AO31x2_ASAP7_75t_L g1367 ( 
.A1(n_1284),
.A2(n_372),
.A3(n_308),
.B(n_118),
.Y(n_1367)
);

INVxp33_ASAP7_75t_L g1368 ( 
.A(n_1202),
.Y(n_1368)
);

AOI221x1_ASAP7_75t_L g1369 ( 
.A1(n_1266),
.A2(n_308),
.B1(n_49),
.B2(n_50),
.C(n_52),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1204),
.Y(n_1370)
);

INVx3_ASAP7_75t_SL g1371 ( 
.A(n_1182),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1189),
.A2(n_308),
.B(n_49),
.Y(n_1372)
);

O2A1O1Ixp33_ASAP7_75t_L g1373 ( 
.A1(n_1266),
.A2(n_48),
.B(n_50),
.C(n_52),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1236),
.A2(n_136),
.B(n_196),
.Y(n_1374)
);

O2A1O1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1175),
.A2(n_53),
.B(n_55),
.C(n_56),
.Y(n_1375)
);

AOI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1208),
.A2(n_1199),
.B1(n_1293),
.B2(n_1291),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1252),
.Y(n_1377)
);

A2O1A1Ixp33_ASAP7_75t_L g1378 ( 
.A1(n_1191),
.A2(n_61),
.B(n_62),
.C(n_63),
.Y(n_1378)
);

INVx1_ASAP7_75t_SL g1379 ( 
.A(n_1270),
.Y(n_1379)
);

AND3x4_ASAP7_75t_L g1380 ( 
.A(n_1213),
.B(n_1301),
.C(n_1286),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1260),
.A2(n_308),
.B(n_151),
.Y(n_1381)
);

AO32x2_ASAP7_75t_L g1382 ( 
.A1(n_1267),
.A2(n_62),
.A3(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1245),
.A2(n_152),
.B(n_192),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1174),
.B(n_64),
.Y(n_1384)
);

AOI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1199),
.A2(n_65),
.B1(n_71),
.B2(n_73),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1239),
.B(n_73),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1271),
.B(n_89),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1220),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1202),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1223),
.Y(n_1390)
);

OAI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1300),
.A2(n_132),
.B(n_137),
.Y(n_1391)
);

BUFx2_ASAP7_75t_L g1392 ( 
.A(n_1172),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_1213),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1229),
.Y(n_1394)
);

AND2x6_ASAP7_75t_SL g1395 ( 
.A(n_1249),
.B(n_143),
.Y(n_1395)
);

BUFx5_ASAP7_75t_L g1396 ( 
.A(n_1277),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1262),
.A2(n_160),
.B(n_161),
.Y(n_1397)
);

OR2x6_ASAP7_75t_L g1398 ( 
.A(n_1150),
.B(n_164),
.Y(n_1398)
);

O2A1O1Ixp5_ASAP7_75t_SL g1399 ( 
.A1(n_1163),
.A2(n_171),
.B(n_181),
.C(n_184),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1244),
.Y(n_1400)
);

BUFx6f_ASAP7_75t_L g1401 ( 
.A(n_1172),
.Y(n_1401)
);

INVx3_ASAP7_75t_L g1402 ( 
.A(n_1172),
.Y(n_1402)
);

NOR2x1_ASAP7_75t_SL g1403 ( 
.A(n_1197),
.B(n_1298),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1256),
.A2(n_1192),
.B(n_1242),
.Y(n_1404)
);

OA21x2_ASAP7_75t_L g1405 ( 
.A1(n_1163),
.A2(n_1228),
.B(n_1287),
.Y(n_1405)
);

BUFx2_ASAP7_75t_L g1406 ( 
.A(n_1197),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1227),
.B(n_1291),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1232),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1269),
.B(n_1273),
.Y(n_1409)
);

AO31x2_ASAP7_75t_L g1410 ( 
.A1(n_1268),
.A2(n_1235),
.A3(n_1211),
.B(n_1289),
.Y(n_1410)
);

BUFx3_ASAP7_75t_L g1411 ( 
.A(n_1294),
.Y(n_1411)
);

OAI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1187),
.A2(n_1272),
.B(n_1225),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1292),
.A2(n_1296),
.B(n_1226),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1166),
.A2(n_1205),
.B1(n_1217),
.B2(n_1221),
.Y(n_1414)
);

AO31x2_ASAP7_75t_L g1415 ( 
.A1(n_1279),
.A2(n_1265),
.A3(n_1283),
.B(n_1179),
.Y(n_1415)
);

O2A1O1Ixp5_ASAP7_75t_L g1416 ( 
.A1(n_1281),
.A2(n_1185),
.B(n_1288),
.C(n_1295),
.Y(n_1416)
);

INVxp33_ASAP7_75t_L g1417 ( 
.A(n_1196),
.Y(n_1417)
);

NOR4xp25_ASAP7_75t_L g1418 ( 
.A(n_1175),
.B(n_1282),
.C(n_1200),
.D(n_1261),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1278),
.A2(n_1180),
.B1(n_1219),
.B2(n_1178),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1264),
.A2(n_1290),
.B(n_1234),
.Y(n_1420)
);

AOI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1207),
.A2(n_1188),
.B(n_1215),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1294),
.A2(n_1269),
.B(n_1253),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1253),
.A2(n_1176),
.B(n_1184),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1197),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1197),
.A2(n_1215),
.B1(n_1275),
.B2(n_1298),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1215),
.A2(n_1275),
.B(n_1298),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1215),
.A2(n_1275),
.B(n_1298),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1222),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1275),
.Y(n_1429)
);

BUFx2_ASAP7_75t_L g1430 ( 
.A(n_1222),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1258),
.A2(n_963),
.B(n_1243),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1243),
.A2(n_963),
.B(n_1230),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1148),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1210),
.A2(n_971),
.B1(n_800),
.B2(n_966),
.Y(n_1434)
);

INVx2_ASAP7_75t_SL g1435 ( 
.A(n_1161),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1151),
.B(n_977),
.Y(n_1436)
);

AND2x4_ASAP7_75t_L g1437 ( 
.A(n_1151),
.B(n_977),
.Y(n_1437)
);

NAND3xp33_ASAP7_75t_L g1438 ( 
.A(n_1194),
.B(n_971),
.C(n_800),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1148),
.Y(n_1439)
);

NOR2xp67_ASAP7_75t_SL g1440 ( 
.A(n_1161),
.B(n_1064),
.Y(n_1440)
);

AO31x2_ASAP7_75t_L g1441 ( 
.A1(n_1160),
.A2(n_1238),
.A3(n_982),
.B(n_1138),
.Y(n_1441)
);

OAI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1195),
.A2(n_1259),
.B(n_1158),
.Y(n_1442)
);

OAI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1164),
.A2(n_963),
.B(n_1100),
.Y(n_1443)
);

AO31x2_ASAP7_75t_L g1444 ( 
.A1(n_1160),
.A2(n_1238),
.A3(n_982),
.B(n_1138),
.Y(n_1444)
);

OA21x2_ASAP7_75t_L g1445 ( 
.A1(n_1195),
.A2(n_1171),
.B(n_1160),
.Y(n_1445)
);

AND2x6_ASAP7_75t_L g1446 ( 
.A(n_1269),
.B(n_890),
.Y(n_1446)
);

AOI31xp67_ASAP7_75t_L g1447 ( 
.A1(n_1230),
.A2(n_1149),
.A3(n_1168),
.B(n_1231),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1195),
.A2(n_1259),
.B(n_1158),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_SL g1449 ( 
.A1(n_1280),
.A2(n_963),
.B(n_1009),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_SL g1450 ( 
.A1(n_1280),
.A2(n_963),
.B(n_1009),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1148),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1243),
.A2(n_963),
.B(n_1230),
.Y(n_1452)
);

NOR4xp25_ASAP7_75t_L g1453 ( 
.A(n_1266),
.B(n_1194),
.C(n_1152),
.D(n_1191),
.Y(n_1453)
);

INVx2_ASAP7_75t_SL g1454 ( 
.A(n_1161),
.Y(n_1454)
);

AOI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1243),
.A2(n_963),
.B(n_1230),
.Y(n_1455)
);

NOR2xp33_ASAP7_75t_L g1456 ( 
.A(n_1153),
.B(n_800),
.Y(n_1456)
);

OAI21xp5_ASAP7_75t_L g1457 ( 
.A1(n_1164),
.A2(n_963),
.B(n_1100),
.Y(n_1457)
);

AOI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1243),
.A2(n_963),
.B(n_1230),
.Y(n_1458)
);

CKINVDCx11_ASAP7_75t_R g1459 ( 
.A(n_1161),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1195),
.A2(n_1259),
.B(n_1158),
.Y(n_1460)
);

AOI21xp33_ASAP7_75t_L g1461 ( 
.A1(n_1194),
.A2(n_800),
.B(n_1096),
.Y(n_1461)
);

A2O1A1Ixp33_ASAP7_75t_L g1462 ( 
.A1(n_1152),
.A2(n_971),
.B(n_1194),
.C(n_844),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1170),
.B(n_806),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1243),
.A2(n_963),
.B(n_1230),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_SL g1465 ( 
.A(n_1194),
.B(n_756),
.Y(n_1465)
);

O2A1O1Ixp33_ASAP7_75t_L g1466 ( 
.A1(n_1152),
.A2(n_800),
.B(n_739),
.C(n_971),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1243),
.A2(n_963),
.B(n_1230),
.Y(n_1467)
);

OA21x2_ASAP7_75t_L g1468 ( 
.A1(n_1195),
.A2(n_1171),
.B(n_1160),
.Y(n_1468)
);

OAI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1376),
.A2(n_1385),
.B1(n_1465),
.B2(n_1438),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1303),
.Y(n_1470)
);

BUFx12f_ASAP7_75t_L g1471 ( 
.A(n_1459),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1384),
.B(n_1317),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1376),
.A2(n_1461),
.B1(n_1438),
.B2(n_1465),
.Y(n_1473)
);

BUFx6f_ASAP7_75t_L g1474 ( 
.A(n_1350),
.Y(n_1474)
);

INVx6_ASAP7_75t_L g1475 ( 
.A(n_1350),
.Y(n_1475)
);

OAI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1385),
.A2(n_1434),
.B1(n_1369),
.B2(n_1417),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_SL g1477 ( 
.A1(n_1414),
.A2(n_1391),
.B1(n_1318),
.B2(n_1456),
.Y(n_1477)
);

INVx6_ASAP7_75t_L g1478 ( 
.A(n_1311),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1361),
.A2(n_1313),
.B1(n_1380),
.B2(n_1408),
.Y(n_1479)
);

BUFx6f_ASAP7_75t_L g1480 ( 
.A(n_1350),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1309),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_SL g1482 ( 
.A1(n_1391),
.A2(n_1372),
.B1(n_1407),
.B2(n_1338),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1356),
.A2(n_1352),
.B1(n_1379),
.B2(n_1355),
.Y(n_1483)
);

OAI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1371),
.A2(n_1364),
.B1(n_1315),
.B2(n_1324),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1379),
.A2(n_1346),
.B1(n_1463),
.B2(n_1334),
.Y(n_1485)
);

INVx6_ASAP7_75t_L g1486 ( 
.A(n_1320),
.Y(n_1486)
);

INVx1_ASAP7_75t_SL g1487 ( 
.A(n_1392),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1331),
.B(n_1336),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1337),
.Y(n_1489)
);

CKINVDCx11_ASAP7_75t_R g1490 ( 
.A(n_1389),
.Y(n_1490)
);

INVx2_ASAP7_75t_SL g1491 ( 
.A(n_1319),
.Y(n_1491)
);

CKINVDCx20_ASAP7_75t_R g1492 ( 
.A(n_1435),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1340),
.Y(n_1493)
);

OAI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1393),
.A2(n_1368),
.B1(n_1386),
.B2(n_1343),
.Y(n_1494)
);

OAI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1466),
.A2(n_1462),
.B1(n_1314),
.B2(n_1443),
.Y(n_1495)
);

OAI21xp5_ASAP7_75t_SL g1496 ( 
.A1(n_1373),
.A2(n_1378),
.B(n_1375),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1348),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1358),
.Y(n_1498)
);

OAI22x1_ASAP7_75t_L g1499 ( 
.A1(n_1339),
.A2(n_1433),
.B1(n_1365),
.B2(n_1370),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1334),
.A2(n_1400),
.B1(n_1388),
.B2(n_1390),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1443),
.A2(n_1457),
.B1(n_1323),
.B2(n_1431),
.Y(n_1501)
);

INVx6_ASAP7_75t_L g1502 ( 
.A(n_1436),
.Y(n_1502)
);

INVx3_ASAP7_75t_L g1503 ( 
.A(n_1401),
.Y(n_1503)
);

CKINVDCx20_ASAP7_75t_R g1504 ( 
.A(n_1454),
.Y(n_1504)
);

OAI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1398),
.A2(n_1335),
.B1(n_1328),
.B2(n_1321),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1439),
.Y(n_1506)
);

OAI21xp5_ASAP7_75t_SL g1507 ( 
.A1(n_1457),
.A2(n_1412),
.B(n_1354),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1394),
.A2(n_1437),
.B1(n_1428),
.B2(n_1377),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1451),
.Y(n_1509)
);

OAI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1398),
.A2(n_1308),
.B1(n_1412),
.B2(n_1432),
.Y(n_1510)
);

OAI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1430),
.A2(n_1305),
.B1(n_1325),
.B2(n_1395),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1437),
.A2(n_1449),
.B1(n_1450),
.B2(n_1446),
.Y(n_1512)
);

INVx6_ASAP7_75t_L g1513 ( 
.A(n_1446),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1406),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_SL g1515 ( 
.A1(n_1423),
.A2(n_1446),
.B1(n_1395),
.B2(n_1357),
.Y(n_1515)
);

BUFx2_ASAP7_75t_L g1516 ( 
.A(n_1429),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1382),
.Y(n_1517)
);

BUFx4_ASAP7_75t_R g1518 ( 
.A(n_1403),
.Y(n_1518)
);

BUFx10_ASAP7_75t_L g1519 ( 
.A(n_1306),
.Y(n_1519)
);

INVx1_ASAP7_75t_SL g1520 ( 
.A(n_1401),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1453),
.B(n_1452),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1325),
.A2(n_1419),
.B1(n_1357),
.B2(n_1387),
.Y(n_1522)
);

INVx3_ASAP7_75t_L g1523 ( 
.A(n_1424),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1455),
.A2(n_1467),
.B1(n_1464),
.B2(n_1458),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1349),
.A2(n_1351),
.B1(n_1409),
.B2(n_1404),
.Y(n_1525)
);

OAI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1453),
.A2(n_1420),
.B1(n_1411),
.B2(n_1382),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1351),
.A2(n_1302),
.B1(n_1421),
.B2(n_1396),
.Y(n_1527)
);

AOI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1440),
.A2(n_1418),
.B1(n_1396),
.B2(n_1422),
.Y(n_1528)
);

INVx6_ASAP7_75t_L g1529 ( 
.A(n_1424),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1382),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1332),
.A2(n_1333),
.B1(n_1413),
.B2(n_1402),
.Y(n_1531)
);

INVx1_ASAP7_75t_SL g1532 ( 
.A(n_1424),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_1402),
.Y(n_1533)
);

AOI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1418),
.A2(n_1396),
.B1(n_1322),
.B2(n_1425),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_SL g1535 ( 
.A1(n_1302),
.A2(n_1397),
.B1(n_1381),
.B2(n_1396),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1396),
.A2(n_1347),
.B1(n_1405),
.B2(n_1329),
.Y(n_1536)
);

INVx2_ASAP7_75t_SL g1537 ( 
.A(n_1426),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_SL g1538 ( 
.A(n_1416),
.B(n_1383),
.Y(n_1538)
);

INVx6_ASAP7_75t_L g1539 ( 
.A(n_1427),
.Y(n_1539)
);

BUFx12f_ASAP7_75t_L g1540 ( 
.A(n_1367),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1312),
.Y(n_1541)
);

INVx2_ASAP7_75t_SL g1542 ( 
.A(n_1441),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1447),
.Y(n_1543)
);

CKINVDCx20_ASAP7_75t_R g1544 ( 
.A(n_1374),
.Y(n_1544)
);

BUFx8_ASAP7_75t_L g1545 ( 
.A(n_1344),
.Y(n_1545)
);

OAI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1359),
.A2(n_1362),
.B1(n_1405),
.B2(n_1345),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1445),
.A2(n_1468),
.B1(n_1330),
.B2(n_1316),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1445),
.A2(n_1468),
.B1(n_1330),
.B2(n_1327),
.Y(n_1548)
);

AOI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1360),
.A2(n_1366),
.B1(n_1353),
.B2(n_1307),
.Y(n_1549)
);

INVx8_ASAP7_75t_L g1550 ( 
.A(n_1399),
.Y(n_1550)
);

AOI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1442),
.A2(n_1460),
.B(n_1448),
.Y(n_1551)
);

BUFx10_ASAP7_75t_L g1552 ( 
.A(n_1441),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1441),
.B(n_1444),
.Y(n_1553)
);

INVx6_ASAP7_75t_L g1554 ( 
.A(n_1444),
.Y(n_1554)
);

OAI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1304),
.A2(n_1341),
.B1(n_1410),
.B2(n_1444),
.Y(n_1555)
);

INVx1_ASAP7_75t_SL g1556 ( 
.A(n_1363),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1304),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1326),
.A2(n_1410),
.B1(n_1304),
.B2(n_1341),
.Y(n_1558)
);

BUFx2_ASAP7_75t_SL g1559 ( 
.A(n_1415),
.Y(n_1559)
);

BUFx6f_ASAP7_75t_L g1560 ( 
.A(n_1310),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1410),
.A2(n_1341),
.B1(n_1342),
.B2(n_1415),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_SL g1562 ( 
.A1(n_1342),
.A2(n_873),
.B1(n_1465),
.B2(n_450),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1310),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1310),
.Y(n_1564)
);

OAI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1466),
.A2(n_1438),
.B(n_1461),
.Y(n_1565)
);

AOI21xp5_ASAP7_75t_L g1566 ( 
.A1(n_1466),
.A2(n_1431),
.B(n_1443),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1376),
.A2(n_1224),
.B1(n_873),
.B2(n_756),
.Y(n_1567)
);

BUFx12f_ASAP7_75t_L g1568 ( 
.A(n_1459),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1376),
.A2(n_1224),
.B1(n_873),
.B2(n_756),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1438),
.A2(n_1376),
.B1(n_1434),
.B2(n_1466),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_SL g1571 ( 
.A1(n_1465),
.A2(n_873),
.B1(n_450),
.B2(n_453),
.Y(n_1571)
);

BUFx10_ASAP7_75t_L g1572 ( 
.A(n_1319),
.Y(n_1572)
);

INVx2_ASAP7_75t_SL g1573 ( 
.A(n_1336),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1303),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1303),
.Y(n_1575)
);

AOI22xp33_ASAP7_75t_SL g1576 ( 
.A1(n_1465),
.A2(n_873),
.B1(n_450),
.B2(n_453),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1376),
.A2(n_1224),
.B1(n_873),
.B2(n_756),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_SL g1578 ( 
.A1(n_1465),
.A2(n_873),
.B1(n_450),
.B2(n_453),
.Y(n_1578)
);

CKINVDCx11_ASAP7_75t_R g1579 ( 
.A(n_1459),
.Y(n_1579)
);

INVx2_ASAP7_75t_SL g1580 ( 
.A(n_1336),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_SL g1581 ( 
.A1(n_1465),
.A2(n_873),
.B1(n_450),
.B2(n_453),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_L g1582 ( 
.A1(n_1376),
.A2(n_1224),
.B1(n_873),
.B2(n_756),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1303),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1303),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1303),
.Y(n_1585)
);

CKINVDCx11_ASAP7_75t_R g1586 ( 
.A(n_1459),
.Y(n_1586)
);

CKINVDCx11_ASAP7_75t_R g1587 ( 
.A(n_1459),
.Y(n_1587)
);

CKINVDCx20_ASAP7_75t_R g1588 ( 
.A(n_1459),
.Y(n_1588)
);

BUFx4f_ASAP7_75t_SL g1589 ( 
.A(n_1311),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1303),
.Y(n_1590)
);

BUFx12f_ASAP7_75t_L g1591 ( 
.A(n_1459),
.Y(n_1591)
);

BUFx2_ASAP7_75t_L g1592 ( 
.A(n_1429),
.Y(n_1592)
);

OAI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1438),
.A2(n_1376),
.B1(n_1434),
.B2(n_1466),
.Y(n_1593)
);

AOI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1376),
.A2(n_800),
.B1(n_971),
.B2(n_873),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1303),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1376),
.A2(n_1224),
.B1(n_873),
.B2(n_756),
.Y(n_1596)
);

OAI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1376),
.A2(n_873),
.B1(n_1385),
.B2(n_1465),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1376),
.A2(n_1224),
.B1(n_873),
.B2(n_756),
.Y(n_1598)
);

INVx3_ASAP7_75t_L g1599 ( 
.A(n_1350),
.Y(n_1599)
);

INVx4_ASAP7_75t_SL g1600 ( 
.A(n_1446),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1376),
.A2(n_1224),
.B1(n_873),
.B2(n_756),
.Y(n_1601)
);

INVx2_ASAP7_75t_SL g1602 ( 
.A(n_1336),
.Y(n_1602)
);

BUFx4f_ASAP7_75t_SL g1603 ( 
.A(n_1311),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1303),
.Y(n_1604)
);

OAI21xp5_ASAP7_75t_SL g1605 ( 
.A1(n_1466),
.A2(n_1438),
.B(n_1376),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_SL g1606 ( 
.A1(n_1465),
.A2(n_873),
.B1(n_450),
.B2(n_453),
.Y(n_1606)
);

OAI21xp33_ASAP7_75t_SL g1607 ( 
.A1(n_1461),
.A2(n_1385),
.B(n_1376),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1303),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_SL g1609 ( 
.A1(n_1465),
.A2(n_873),
.B1(n_450),
.B2(n_453),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1376),
.A2(n_1224),
.B1(n_873),
.B2(n_756),
.Y(n_1610)
);

BUFx10_ASAP7_75t_L g1611 ( 
.A(n_1319),
.Y(n_1611)
);

BUFx2_ASAP7_75t_SL g1612 ( 
.A(n_1352),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_SL g1613 ( 
.A1(n_1465),
.A2(n_873),
.B1(n_450),
.B2(n_453),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1376),
.A2(n_1224),
.B1(n_873),
.B2(n_756),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1376),
.A2(n_800),
.B1(n_971),
.B2(n_873),
.Y(n_1615)
);

CKINVDCx11_ASAP7_75t_R g1616 ( 
.A(n_1459),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_SL g1617 ( 
.A1(n_1465),
.A2(n_873),
.B1(n_450),
.B2(n_453),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1384),
.B(n_1057),
.Y(n_1618)
);

AOI22xp33_ASAP7_75t_SL g1619 ( 
.A1(n_1465),
.A2(n_873),
.B1(n_450),
.B2(n_453),
.Y(n_1619)
);

OAI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1376),
.A2(n_873),
.B1(n_1385),
.B2(n_1465),
.Y(n_1620)
);

BUFx3_ASAP7_75t_L g1621 ( 
.A(n_1320),
.Y(n_1621)
);

BUFx4f_ASAP7_75t_L g1622 ( 
.A(n_1311),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1434),
.B(n_1462),
.Y(n_1623)
);

CKINVDCx11_ASAP7_75t_R g1624 ( 
.A(n_1459),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1376),
.A2(n_1224),
.B1(n_873),
.B2(n_756),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1303),
.Y(n_1626)
);

CKINVDCx20_ASAP7_75t_R g1627 ( 
.A(n_1459),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1541),
.Y(n_1628)
);

INVxp33_ASAP7_75t_L g1629 ( 
.A(n_1490),
.Y(n_1629)
);

INVx3_ASAP7_75t_L g1630 ( 
.A(n_1539),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1553),
.Y(n_1631)
);

BUFx12f_ASAP7_75t_SL g1632 ( 
.A(n_1474),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1521),
.Y(n_1633)
);

AOI222xp33_ASAP7_75t_L g1634 ( 
.A1(n_1597),
.A2(n_1620),
.B1(n_1607),
.B2(n_1567),
.C1(n_1625),
.C2(n_1569),
.Y(n_1634)
);

BUFx2_ASAP7_75t_L g1635 ( 
.A(n_1539),
.Y(n_1635)
);

OR2x6_ASAP7_75t_L g1636 ( 
.A(n_1513),
.B(n_1554),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1509),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1470),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1481),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1521),
.Y(n_1640)
);

BUFx2_ASAP7_75t_L g1641 ( 
.A(n_1539),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1517),
.B(n_1530),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1489),
.Y(n_1643)
);

BUFx6f_ASAP7_75t_L g1644 ( 
.A(n_1513),
.Y(n_1644)
);

HB1xp67_ASAP7_75t_L g1645 ( 
.A(n_1514),
.Y(n_1645)
);

INVx1_ASAP7_75t_SL g1646 ( 
.A(n_1486),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1493),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1497),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1498),
.Y(n_1649)
);

AO31x2_ASAP7_75t_L g1650 ( 
.A1(n_1501),
.A2(n_1566),
.A3(n_1531),
.B(n_1563),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1506),
.Y(n_1651)
);

BUFx3_ASAP7_75t_L g1652 ( 
.A(n_1486),
.Y(n_1652)
);

BUFx3_ASAP7_75t_L g1653 ( 
.A(n_1516),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1623),
.B(n_1605),
.Y(n_1654)
);

AOI22xp33_ASAP7_75t_SL g1655 ( 
.A1(n_1570),
.A2(n_1593),
.B1(n_1495),
.B2(n_1540),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1574),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1501),
.B(n_1605),
.Y(n_1657)
);

INVx3_ASAP7_75t_L g1658 ( 
.A(n_1560),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_L g1659 ( 
.A(n_1621),
.B(n_1492),
.Y(n_1659)
);

INVx3_ASAP7_75t_L g1660 ( 
.A(n_1560),
.Y(n_1660)
);

BUFx2_ASAP7_75t_L g1661 ( 
.A(n_1564),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1575),
.Y(n_1662)
);

INVx3_ASAP7_75t_L g1663 ( 
.A(n_1545),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1570),
.B(n_1593),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1583),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1584),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1585),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1623),
.B(n_1488),
.Y(n_1668)
);

AOI211x1_ASAP7_75t_L g1669 ( 
.A1(n_1476),
.A2(n_1494),
.B(n_1469),
.C(n_1472),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1557),
.B(n_1507),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1590),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1595),
.Y(n_1672)
);

INVx3_ASAP7_75t_L g1673 ( 
.A(n_1545),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1604),
.B(n_1608),
.Y(n_1674)
);

BUFx2_ASAP7_75t_L g1675 ( 
.A(n_1537),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1507),
.B(n_1484),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1626),
.Y(n_1677)
);

AND2x4_ASAP7_75t_L g1678 ( 
.A(n_1600),
.B(n_1528),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1499),
.B(n_1487),
.Y(n_1679)
);

INVx1_ASAP7_75t_SL g1680 ( 
.A(n_1504),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1543),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1561),
.B(n_1473),
.Y(n_1682)
);

INVx2_ASAP7_75t_SL g1683 ( 
.A(n_1475),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1487),
.Y(n_1684)
);

BUFx3_ASAP7_75t_L g1685 ( 
.A(n_1592),
.Y(n_1685)
);

OAI21x1_ASAP7_75t_L g1686 ( 
.A1(n_1551),
.A2(n_1524),
.B(n_1531),
.Y(n_1686)
);

INVx2_ASAP7_75t_SL g1687 ( 
.A(n_1475),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1571),
.A2(n_1617),
.B1(n_1609),
.B2(n_1613),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1542),
.Y(n_1689)
);

INVx6_ASAP7_75t_L g1690 ( 
.A(n_1600),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1500),
.Y(n_1691)
);

BUFx6f_ASAP7_75t_L g1692 ( 
.A(n_1513),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1510),
.Y(n_1693)
);

AO21x2_ASAP7_75t_L g1694 ( 
.A1(n_1546),
.A2(n_1555),
.B(n_1566),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1552),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1559),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1618),
.B(n_1558),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1527),
.B(n_1477),
.Y(n_1698)
);

AO21x2_ASAP7_75t_L g1699 ( 
.A1(n_1551),
.A2(n_1549),
.B(n_1526),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1524),
.Y(n_1700)
);

INVx3_ASAP7_75t_L g1701 ( 
.A(n_1599),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1510),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1534),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1556),
.Y(n_1704)
);

OAI21x1_ASAP7_75t_SL g1705 ( 
.A1(n_1565),
.A2(n_1495),
.B(n_1615),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1594),
.B(n_1565),
.Y(n_1706)
);

INVx3_ASAP7_75t_L g1707 ( 
.A(n_1599),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1556),
.Y(n_1708)
);

BUFx2_ASAP7_75t_L g1709 ( 
.A(n_1533),
.Y(n_1709)
);

OA21x2_ASAP7_75t_L g1710 ( 
.A1(n_1548),
.A2(n_1547),
.B(n_1536),
.Y(n_1710)
);

INVxp67_ASAP7_75t_SL g1711 ( 
.A(n_1525),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1482),
.B(n_1479),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1505),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1550),
.Y(n_1714)
);

INVx5_ASAP7_75t_L g1715 ( 
.A(n_1475),
.Y(n_1715)
);

HB1xp67_ASAP7_75t_L g1716 ( 
.A(n_1520),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1503),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1485),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1508),
.Y(n_1719)
);

BUFx3_ASAP7_75t_L g1720 ( 
.A(n_1529),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1503),
.Y(n_1721)
);

AO21x2_ASAP7_75t_L g1722 ( 
.A1(n_1538),
.A2(n_1496),
.B(n_1511),
.Y(n_1722)
);

OAI21x1_ASAP7_75t_L g1723 ( 
.A1(n_1522),
.A2(n_1512),
.B(n_1523),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1535),
.Y(n_1724)
);

BUFx2_ASAP7_75t_R g1725 ( 
.A(n_1612),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1573),
.B(n_1602),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1515),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1532),
.Y(n_1728)
);

INVx3_ASAP7_75t_L g1729 ( 
.A(n_1529),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1532),
.Y(n_1730)
);

NOR2xp67_ASAP7_75t_L g1731 ( 
.A(n_1580),
.B(n_1491),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1562),
.Y(n_1732)
);

OA21x2_ASAP7_75t_L g1733 ( 
.A1(n_1496),
.A2(n_1601),
.B(n_1610),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1480),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_1579),
.Y(n_1735)
);

BUFx2_ASAP7_75t_L g1736 ( 
.A(n_1544),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1518),
.Y(n_1737)
);

AOI22xp33_ASAP7_75t_L g1738 ( 
.A1(n_1576),
.A2(n_1581),
.B1(n_1578),
.B2(n_1606),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1483),
.B(n_1502),
.Y(n_1739)
);

OA21x2_ASAP7_75t_L g1740 ( 
.A1(n_1577),
.A2(n_1582),
.B(n_1596),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1598),
.B(n_1614),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_1586),
.Y(n_1742)
);

INVx3_ASAP7_75t_L g1743 ( 
.A(n_1478),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1478),
.Y(n_1744)
);

INVx3_ASAP7_75t_L g1745 ( 
.A(n_1622),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1619),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1572),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1622),
.B(n_1519),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1572),
.Y(n_1749)
);

AOI22xp33_ASAP7_75t_L g1750 ( 
.A1(n_1471),
.A2(n_1591),
.B1(n_1568),
.B2(n_1587),
.Y(n_1750)
);

NOR2x1_ASAP7_75t_SL g1751 ( 
.A(n_1722),
.B(n_1624),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1633),
.B(n_1611),
.Y(n_1752)
);

OAI21xp33_ASAP7_75t_L g1753 ( 
.A1(n_1657),
.A2(n_1588),
.B(n_1627),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1678),
.B(n_1589),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1733),
.A2(n_1616),
.B1(n_1603),
.B2(n_1519),
.Y(n_1755)
);

OAI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1655),
.A2(n_1664),
.B1(n_1657),
.B2(n_1654),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1736),
.B(n_1697),
.Y(n_1757)
);

AOI221xp5_ASAP7_75t_L g1758 ( 
.A1(n_1669),
.A2(n_1712),
.B1(n_1698),
.B2(n_1640),
.C(n_1705),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1643),
.Y(n_1759)
);

AND2x4_ASAP7_75t_L g1760 ( 
.A(n_1678),
.B(n_1630),
.Y(n_1760)
);

NOR2x1_ASAP7_75t_SL g1761 ( 
.A(n_1722),
.B(n_1676),
.Y(n_1761)
);

OAI21xp5_ASAP7_75t_L g1762 ( 
.A1(n_1664),
.A2(n_1676),
.B(n_1706),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1670),
.B(n_1702),
.Y(n_1763)
);

OAI21xp5_ASAP7_75t_L g1764 ( 
.A1(n_1706),
.A2(n_1698),
.B(n_1711),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1670),
.B(n_1702),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1693),
.B(n_1674),
.Y(n_1766)
);

AND2x4_ASAP7_75t_L g1767 ( 
.A(n_1678),
.B(n_1630),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1674),
.B(n_1643),
.Y(n_1768)
);

CKINVDCx5p33_ASAP7_75t_R g1769 ( 
.A(n_1652),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1647),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1637),
.B(n_1668),
.Y(n_1771)
);

OAI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1703),
.A2(n_1724),
.B(n_1723),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1648),
.Y(n_1773)
);

OAI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1703),
.A2(n_1723),
.B(n_1727),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1645),
.B(n_1684),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1649),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1651),
.Y(n_1777)
);

OA21x2_ASAP7_75t_L g1778 ( 
.A1(n_1686),
.A2(n_1700),
.B(n_1714),
.Y(n_1778)
);

INVx3_ASAP7_75t_L g1779 ( 
.A(n_1701),
.Y(n_1779)
);

HB1xp67_ASAP7_75t_L g1780 ( 
.A(n_1716),
.Y(n_1780)
);

INVx3_ASAP7_75t_L g1781 ( 
.A(n_1701),
.Y(n_1781)
);

OR2x6_ASAP7_75t_L g1782 ( 
.A(n_1636),
.B(n_1690),
.Y(n_1782)
);

AOI22xp33_ASAP7_75t_L g1783 ( 
.A1(n_1733),
.A2(n_1634),
.B1(n_1740),
.B2(n_1732),
.Y(n_1783)
);

AOI211xp5_ASAP7_75t_L g1784 ( 
.A1(n_1727),
.A2(n_1682),
.B(n_1732),
.C(n_1737),
.Y(n_1784)
);

AO32x2_ASAP7_75t_L g1785 ( 
.A1(n_1683),
.A2(n_1687),
.A3(n_1642),
.B1(n_1631),
.B2(n_1679),
.Y(n_1785)
);

BUFx3_ASAP7_75t_L g1786 ( 
.A(n_1652),
.Y(n_1786)
);

HB1xp67_ASAP7_75t_L g1787 ( 
.A(n_1730),
.Y(n_1787)
);

AOI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1733),
.A2(n_1722),
.B1(n_1741),
.B2(n_1738),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1665),
.B(n_1667),
.Y(n_1789)
);

INVxp67_ASAP7_75t_L g1790 ( 
.A(n_1726),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1635),
.B(n_1641),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1733),
.A2(n_1688),
.B1(n_1737),
.B2(n_1673),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1665),
.Y(n_1793)
);

CKINVDCx5p33_ASAP7_75t_R g1794 ( 
.A(n_1735),
.Y(n_1794)
);

OAI22xp5_ASAP7_75t_L g1795 ( 
.A1(n_1663),
.A2(n_1673),
.B1(n_1725),
.B2(n_1731),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1667),
.Y(n_1796)
);

AOI221xp5_ASAP7_75t_L g1797 ( 
.A1(n_1705),
.A2(n_1746),
.B1(n_1639),
.B2(n_1638),
.C(n_1671),
.Y(n_1797)
);

AND2x4_ASAP7_75t_L g1798 ( 
.A(n_1635),
.B(n_1641),
.Y(n_1798)
);

BUFx2_ASAP7_75t_L g1799 ( 
.A(n_1653),
.Y(n_1799)
);

HB1xp67_ASAP7_75t_L g1800 ( 
.A(n_1730),
.Y(n_1800)
);

OAI221xp5_ASAP7_75t_SL g1801 ( 
.A1(n_1746),
.A2(n_1679),
.B1(n_1713),
.B2(n_1700),
.C(n_1750),
.Y(n_1801)
);

NOR2xp33_ASAP7_75t_L g1802 ( 
.A(n_1747),
.B(n_1749),
.Y(n_1802)
);

NAND4xp25_ASAP7_75t_L g1803 ( 
.A(n_1747),
.B(n_1749),
.C(n_1653),
.D(n_1685),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1685),
.B(n_1709),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1709),
.B(n_1646),
.Y(n_1805)
);

O2A1O1Ixp33_ASAP7_75t_SL g1806 ( 
.A1(n_1663),
.A2(n_1673),
.B(n_1745),
.C(n_1629),
.Y(n_1806)
);

AOI221xp5_ASAP7_75t_L g1807 ( 
.A1(n_1713),
.A2(n_1691),
.B1(n_1718),
.B2(n_1719),
.C(n_1677),
.Y(n_1807)
);

NOR2x1_ASAP7_75t_R g1808 ( 
.A(n_1735),
.B(n_1742),
.Y(n_1808)
);

AOI22xp5_ASAP7_75t_SL g1809 ( 
.A1(n_1742),
.A2(n_1663),
.B1(n_1748),
.B2(n_1743),
.Y(n_1809)
);

OAI22xp5_ASAP7_75t_SL g1810 ( 
.A1(n_1745),
.A2(n_1659),
.B1(n_1743),
.B2(n_1680),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1694),
.B(n_1650),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1656),
.B(n_1662),
.Y(n_1812)
);

OAI22xp5_ASAP7_75t_L g1813 ( 
.A1(n_1740),
.A2(n_1744),
.B1(n_1690),
.B2(n_1729),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1694),
.B(n_1650),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1694),
.B(n_1650),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1666),
.Y(n_1816)
);

OA21x2_ASAP7_75t_L g1817 ( 
.A1(n_1681),
.A2(n_1696),
.B(n_1704),
.Y(n_1817)
);

BUFx3_ASAP7_75t_L g1818 ( 
.A(n_1720),
.Y(n_1818)
);

OAI211xp5_ASAP7_75t_L g1819 ( 
.A1(n_1675),
.A2(n_1707),
.B(n_1710),
.C(n_1717),
.Y(n_1819)
);

OA21x2_ASAP7_75t_L g1820 ( 
.A1(n_1708),
.A2(n_1689),
.B(n_1628),
.Y(n_1820)
);

O2A1O1Ixp33_ASAP7_75t_L g1821 ( 
.A1(n_1699),
.A2(n_1734),
.B(n_1721),
.C(n_1729),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1766),
.B(n_1672),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1820),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1759),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1763),
.B(n_1650),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1763),
.B(n_1650),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1770),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1773),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1765),
.B(n_1699),
.Y(n_1829)
);

AOI22xp5_ASAP7_75t_L g1830 ( 
.A1(n_1756),
.A2(n_1740),
.B1(n_1739),
.B2(n_1690),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1776),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1777),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1765),
.B(n_1699),
.Y(n_1833)
);

HB1xp67_ASAP7_75t_L g1834 ( 
.A(n_1780),
.Y(n_1834)
);

OR2x2_ASAP7_75t_L g1835 ( 
.A(n_1771),
.B(n_1642),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1793),
.Y(n_1836)
);

BUFx3_ASAP7_75t_L g1837 ( 
.A(n_1786),
.Y(n_1837)
);

INVx8_ASAP7_75t_L g1838 ( 
.A(n_1754),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1796),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1768),
.B(n_1710),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1817),
.Y(n_1841)
);

OR2x2_ASAP7_75t_L g1842 ( 
.A(n_1775),
.B(n_1631),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1768),
.B(n_1710),
.Y(n_1843)
);

HB1xp67_ASAP7_75t_L g1844 ( 
.A(n_1787),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1757),
.B(n_1710),
.Y(n_1845)
);

INVx4_ASAP7_75t_L g1846 ( 
.A(n_1769),
.Y(n_1846)
);

CKINVDCx20_ASAP7_75t_R g1847 ( 
.A(n_1794),
.Y(n_1847)
);

INVxp67_ASAP7_75t_SL g1848 ( 
.A(n_1817),
.Y(n_1848)
);

AND2x4_ASAP7_75t_L g1849 ( 
.A(n_1760),
.B(n_1767),
.Y(n_1849)
);

INVxp67_ASAP7_75t_L g1850 ( 
.A(n_1802),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1800),
.B(n_1661),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1785),
.B(n_1661),
.Y(n_1852)
);

AOI22xp5_ASAP7_75t_L g1853 ( 
.A1(n_1788),
.A2(n_1740),
.B1(n_1644),
.B2(n_1692),
.Y(n_1853)
);

BUFx6f_ASAP7_75t_L g1854 ( 
.A(n_1818),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1762),
.B(n_1728),
.Y(n_1855)
);

BUFx3_ASAP7_75t_L g1856 ( 
.A(n_1786),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1785),
.B(n_1695),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1785),
.B(n_1695),
.Y(n_1858)
);

CKINVDCx20_ASAP7_75t_R g1859 ( 
.A(n_1794),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1785),
.B(n_1660),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1791),
.B(n_1798),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1791),
.B(n_1658),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1798),
.B(n_1789),
.Y(n_1863)
);

NOR2xp33_ASAP7_75t_L g1864 ( 
.A(n_1753),
.B(n_1632),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1824),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1863),
.B(n_1799),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1824),
.Y(n_1867)
);

OAI21xp5_ASAP7_75t_L g1868 ( 
.A1(n_1830),
.A2(n_1758),
.B(n_1764),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1827),
.Y(n_1869)
);

OR2x2_ASAP7_75t_L g1870 ( 
.A(n_1835),
.B(n_1790),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1827),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1840),
.B(n_1811),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1823),
.Y(n_1873)
);

BUFx3_ASAP7_75t_L g1874 ( 
.A(n_1854),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1828),
.Y(n_1875)
);

INVx5_ASAP7_75t_L g1876 ( 
.A(n_1852),
.Y(n_1876)
);

INVx1_ASAP7_75t_SL g1877 ( 
.A(n_1851),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1823),
.Y(n_1878)
);

OAI221xp5_ASAP7_75t_SL g1879 ( 
.A1(n_1830),
.A2(n_1783),
.B1(n_1755),
.B2(n_1797),
.C(n_1811),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1825),
.B(n_1814),
.Y(n_1880)
);

NOR2xp33_ASAP7_75t_L g1881 ( 
.A(n_1846),
.B(n_1808),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1840),
.B(n_1814),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1828),
.Y(n_1883)
);

HB1xp67_ASAP7_75t_L g1884 ( 
.A(n_1844),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1843),
.B(n_1815),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1831),
.Y(n_1886)
);

INVxp67_ASAP7_75t_L g1887 ( 
.A(n_1834),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1832),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1863),
.B(n_1804),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1832),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1861),
.B(n_1752),
.Y(n_1891)
);

NOR2x1_ASAP7_75t_L g1892 ( 
.A(n_1837),
.B(n_1803),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1843),
.B(n_1815),
.Y(n_1893)
);

HB1xp67_ASAP7_75t_L g1894 ( 
.A(n_1851),
.Y(n_1894)
);

AND2x2_ASAP7_75t_SL g1895 ( 
.A(n_1852),
.B(n_1754),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1836),
.Y(n_1896)
);

INVx4_ASAP7_75t_L g1897 ( 
.A(n_1838),
.Y(n_1897)
);

AOI21xp5_ASAP7_75t_SL g1898 ( 
.A1(n_1848),
.A2(n_1751),
.B(n_1761),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1861),
.B(n_1829),
.Y(n_1899)
);

INVxp67_ASAP7_75t_SL g1900 ( 
.A(n_1841),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1846),
.B(n_1769),
.Y(n_1901)
);

AOI22xp33_ASAP7_75t_SL g1902 ( 
.A1(n_1829),
.A2(n_1792),
.B1(n_1819),
.B2(n_1774),
.Y(n_1902)
);

AND2x4_ASAP7_75t_L g1903 ( 
.A(n_1849),
.B(n_1779),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1836),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1833),
.B(n_1778),
.Y(n_1905)
);

AND2x4_ASAP7_75t_L g1906 ( 
.A(n_1849),
.B(n_1779),
.Y(n_1906)
);

OAI221xp5_ASAP7_75t_L g1907 ( 
.A1(n_1853),
.A2(n_1801),
.B1(n_1783),
.B2(n_1784),
.C(n_1772),
.Y(n_1907)
);

OAI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1850),
.A2(n_1807),
.B1(n_1809),
.B2(n_1810),
.Y(n_1908)
);

HB1xp67_ASAP7_75t_L g1909 ( 
.A(n_1857),
.Y(n_1909)
);

AND2x4_ASAP7_75t_L g1910 ( 
.A(n_1849),
.B(n_1781),
.Y(n_1910)
);

OAI33xp33_ASAP7_75t_L g1911 ( 
.A1(n_1855),
.A2(n_1795),
.A3(n_1813),
.B1(n_1821),
.B2(n_1812),
.B3(n_1816),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1833),
.B(n_1778),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1845),
.B(n_1752),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1845),
.B(n_1825),
.Y(n_1914)
);

NAND4xp25_ASAP7_75t_L g1915 ( 
.A(n_1846),
.B(n_1802),
.C(n_1805),
.D(n_1853),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1865),
.Y(n_1916)
);

AND2x4_ASAP7_75t_L g1917 ( 
.A(n_1876),
.B(n_1860),
.Y(n_1917)
);

HB1xp67_ASAP7_75t_L g1918 ( 
.A(n_1884),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1895),
.B(n_1837),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1873),
.Y(n_1920)
);

OR2x6_ASAP7_75t_L g1921 ( 
.A(n_1898),
.B(n_1782),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1873),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1865),
.B(n_1826),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1895),
.B(n_1856),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1867),
.Y(n_1925)
);

OAI31xp33_ASAP7_75t_SL g1926 ( 
.A1(n_1892),
.A2(n_1864),
.A3(n_1826),
.B(n_1860),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1867),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1895),
.B(n_1899),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1869),
.Y(n_1929)
);

AND2x4_ASAP7_75t_L g1930 ( 
.A(n_1876),
.B(n_1857),
.Y(n_1930)
);

BUFx3_ASAP7_75t_L g1931 ( 
.A(n_1874),
.Y(n_1931)
);

OR2x2_ASAP7_75t_L g1932 ( 
.A(n_1877),
.B(n_1835),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1899),
.B(n_1856),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1914),
.B(n_1876),
.Y(n_1934)
);

OR2x2_ASAP7_75t_L g1935 ( 
.A(n_1877),
.B(n_1842),
.Y(n_1935)
);

NAND2x1p5_ASAP7_75t_L g1936 ( 
.A(n_1892),
.B(n_1715),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1869),
.B(n_1839),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1871),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1876),
.B(n_1913),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1875),
.Y(n_1940)
);

HB1xp67_ASAP7_75t_L g1941 ( 
.A(n_1884),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1875),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1883),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1883),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1886),
.Y(n_1945)
);

AND2x4_ASAP7_75t_L g1946 ( 
.A(n_1903),
.B(n_1858),
.Y(n_1946)
);

INVx3_ASAP7_75t_L g1947 ( 
.A(n_1903),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1888),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1888),
.B(n_1822),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1890),
.Y(n_1950)
);

OR2x2_ASAP7_75t_L g1951 ( 
.A(n_1894),
.B(n_1842),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1878),
.Y(n_1952)
);

AND2x4_ASAP7_75t_L g1953 ( 
.A(n_1903),
.B(n_1906),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1903),
.B(n_1862),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1906),
.B(n_1862),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1896),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1928),
.B(n_1909),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1918),
.B(n_1887),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1916),
.Y(n_1959)
);

INVx2_ASAP7_75t_SL g1960 ( 
.A(n_1919),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1916),
.Y(n_1961)
);

INVx1_ASAP7_75t_SL g1962 ( 
.A(n_1919),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1928),
.B(n_1909),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1924),
.B(n_1894),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1925),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1924),
.B(n_1906),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1918),
.B(n_1887),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1934),
.B(n_1910),
.Y(n_1968)
);

AOI21xp33_ASAP7_75t_L g1969 ( 
.A1(n_1926),
.A2(n_1908),
.B(n_1902),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1920),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1925),
.Y(n_1971)
);

OAI21xp33_ASAP7_75t_SL g1972 ( 
.A1(n_1926),
.A2(n_1915),
.B(n_1866),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1934),
.B(n_1910),
.Y(n_1973)
);

HB1xp67_ASAP7_75t_L g1974 ( 
.A(n_1941),
.Y(n_1974)
);

OR2x2_ASAP7_75t_L g1975 ( 
.A(n_1932),
.B(n_1880),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1927),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1954),
.B(n_1910),
.Y(n_1977)
);

AND2x4_ASAP7_75t_L g1978 ( 
.A(n_1953),
.B(n_1897),
.Y(n_1978)
);

OR2x2_ASAP7_75t_L g1979 ( 
.A(n_1932),
.B(n_1880),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1954),
.B(n_1910),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1955),
.B(n_1891),
.Y(n_1981)
);

OR2x6_ASAP7_75t_L g1982 ( 
.A(n_1936),
.B(n_1898),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1955),
.B(n_1891),
.Y(n_1983)
);

OR2x2_ASAP7_75t_L g1984 ( 
.A(n_1951),
.B(n_1915),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1953),
.B(n_1889),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1920),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1941),
.B(n_1872),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1953),
.B(n_1889),
.Y(n_1988)
);

AOI221xp5_ASAP7_75t_L g1989 ( 
.A1(n_1923),
.A2(n_1911),
.B1(n_1879),
.B2(n_1908),
.C(n_1905),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1920),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1927),
.Y(n_1991)
);

NOR2xp33_ASAP7_75t_L g1992 ( 
.A(n_1931),
.B(n_1847),
.Y(n_1992)
);

OR2x2_ASAP7_75t_L g1993 ( 
.A(n_1951),
.B(n_1870),
.Y(n_1993)
);

HB1xp67_ASAP7_75t_L g1994 ( 
.A(n_1937),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1929),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1929),
.Y(n_1996)
);

AOI33xp33_ASAP7_75t_L g1997 ( 
.A1(n_1938),
.A2(n_1902),
.A3(n_1912),
.B1(n_1905),
.B2(n_1885),
.B3(n_1893),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1938),
.Y(n_1998)
);

OR3x2_ASAP7_75t_L g1999 ( 
.A(n_1935),
.B(n_1879),
.C(n_1870),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1940),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1953),
.B(n_1866),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1940),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1942),
.Y(n_2003)
);

INVx1_ASAP7_75t_SL g2004 ( 
.A(n_1933),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1922),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1942),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1939),
.B(n_1874),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1949),
.B(n_1872),
.Y(n_2008)
);

OR2x2_ASAP7_75t_L g2009 ( 
.A(n_1935),
.B(n_1904),
.Y(n_2009)
);

NOR2xp67_ASAP7_75t_L g2010 ( 
.A(n_1947),
.B(n_1897),
.Y(n_2010)
);

CKINVDCx5p33_ASAP7_75t_R g2011 ( 
.A(n_1992),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1985),
.B(n_1931),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1999),
.Y(n_2013)
);

AND3x2_ASAP7_75t_L g2014 ( 
.A(n_1989),
.B(n_1868),
.C(n_1881),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1985),
.B(n_1931),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1959),
.Y(n_2016)
);

INVxp67_ASAP7_75t_L g2017 ( 
.A(n_1958),
.Y(n_2017)
);

INVx1_ASAP7_75t_SL g2018 ( 
.A(n_1974),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1969),
.B(n_1943),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1959),
.Y(n_2020)
);

OAI22xp5_ASAP7_75t_SL g2021 ( 
.A1(n_1982),
.A2(n_1936),
.B1(n_1859),
.B2(n_1921),
.Y(n_2021)
);

INVxp33_ASAP7_75t_L g2022 ( 
.A(n_1964),
.Y(n_2022)
);

INVx1_ASAP7_75t_SL g2023 ( 
.A(n_1967),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1994),
.B(n_1993),
.Y(n_2024)
);

INVx2_ASAP7_75t_SL g2025 ( 
.A(n_1978),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1961),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1961),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1993),
.B(n_1943),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1988),
.B(n_1939),
.Y(n_2029)
);

NOR2xp33_ASAP7_75t_L g2030 ( 
.A(n_2004),
.B(n_1911),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1997),
.B(n_1944),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1965),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1988),
.B(n_1946),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1981),
.B(n_1983),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1975),
.B(n_1944),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1975),
.B(n_1945),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1981),
.B(n_1946),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_SL g2038 ( 
.A(n_1972),
.B(n_1936),
.Y(n_2038)
);

OR2x2_ASAP7_75t_L g2039 ( 
.A(n_1979),
.B(n_1923),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1964),
.B(n_1872),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1999),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1965),
.Y(n_2042)
);

INVx2_ASAP7_75t_SL g2043 ( 
.A(n_1978),
.Y(n_2043)
);

OR2x2_ASAP7_75t_L g2044 ( 
.A(n_1979),
.B(n_1949),
.Y(n_2044)
);

INVx2_ASAP7_75t_SL g2045 ( 
.A(n_1978),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_1983),
.B(n_2001),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_2001),
.B(n_1946),
.Y(n_2047)
);

INVx1_ASAP7_75t_SL g2048 ( 
.A(n_1962),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_1970),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_1966),
.B(n_1977),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_2034),
.B(n_1978),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_2014),
.B(n_1984),
.Y(n_2052)
);

A2O1A1Ixp33_ASAP7_75t_L g2053 ( 
.A1(n_2013),
.A2(n_2041),
.B(n_2030),
.C(n_2031),
.Y(n_2053)
);

OAI221xp5_ASAP7_75t_L g2054 ( 
.A1(n_2013),
.A2(n_1984),
.B1(n_1868),
.B2(n_1936),
.C(n_1982),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_2048),
.B(n_1957),
.Y(n_2055)
);

AOI22xp5_ASAP7_75t_L g2056 ( 
.A1(n_2013),
.A2(n_1907),
.B1(n_1960),
.B2(n_1957),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_2046),
.B(n_2050),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_2016),
.Y(n_2058)
);

NAND3xp33_ASAP7_75t_L g2059 ( 
.A(n_2041),
.B(n_1960),
.C(n_1971),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2016),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2020),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_2034),
.B(n_1966),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_2046),
.B(n_1977),
.Y(n_2063)
);

INVx1_ASAP7_75t_SL g2064 ( 
.A(n_2011),
.Y(n_2064)
);

OAI21xp5_ASAP7_75t_L g2065 ( 
.A1(n_2041),
.A2(n_1982),
.B(n_1963),
.Y(n_2065)
);

AOI22xp5_ASAP7_75t_L g2066 ( 
.A1(n_2031),
.A2(n_1907),
.B1(n_1963),
.B2(n_1921),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2020),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_2048),
.B(n_2008),
.Y(n_2068)
);

NOR3xp33_ASAP7_75t_L g2069 ( 
.A(n_2019),
.B(n_2023),
.C(n_2018),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2026),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2026),
.Y(n_2071)
);

OR2x2_ASAP7_75t_L g2072 ( 
.A(n_2019),
.B(n_2009),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2027),
.Y(n_2073)
);

AOI21xp5_ASAP7_75t_L g2074 ( 
.A1(n_2038),
.A2(n_1982),
.B(n_2010),
.Y(n_2074)
);

INVx2_ASAP7_75t_SL g2075 ( 
.A(n_2012),
.Y(n_2075)
);

AOI22xp5_ASAP7_75t_L g2076 ( 
.A1(n_2021),
.A2(n_1921),
.B1(n_1912),
.B2(n_1905),
.Y(n_2076)
);

AOI211xp5_ASAP7_75t_L g2077 ( 
.A1(n_2021),
.A2(n_2010),
.B(n_1806),
.C(n_1987),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_2027),
.Y(n_2078)
);

AOI322xp5_ASAP7_75t_L g2079 ( 
.A1(n_2023),
.A2(n_1885),
.A3(n_1893),
.B1(n_1882),
.B2(n_1912),
.C1(n_1930),
.C2(n_1917),
.Y(n_2079)
);

INVxp67_ASAP7_75t_SL g2080 ( 
.A(n_2069),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2058),
.Y(n_2081)
);

NAND2x2_ASAP7_75t_L g2082 ( 
.A(n_2075),
.B(n_2025),
.Y(n_2082)
);

INVx2_ASAP7_75t_L g2083 ( 
.A(n_2062),
.Y(n_2083)
);

OAI21xp5_ASAP7_75t_L g2084 ( 
.A1(n_2053),
.A2(n_2017),
.B(n_2022),
.Y(n_2084)
);

AOI32xp33_ASAP7_75t_L g2085 ( 
.A1(n_2069),
.A2(n_2018),
.A3(n_2024),
.B1(n_2028),
.B2(n_2015),
.Y(n_2085)
);

NOR2xp33_ASAP7_75t_L g2086 ( 
.A(n_2064),
.B(n_2025),
.Y(n_2086)
);

OAI22xp5_ASAP7_75t_L g2087 ( 
.A1(n_2056),
.A2(n_2066),
.B1(n_2053),
.B2(n_2076),
.Y(n_2087)
);

AOI21xp5_ASAP7_75t_L g2088 ( 
.A1(n_2052),
.A2(n_2059),
.B(n_2054),
.Y(n_2088)
);

AOI22xp5_ASAP7_75t_L g2089 ( 
.A1(n_2055),
.A2(n_2049),
.B1(n_2012),
.B2(n_2015),
.Y(n_2089)
);

AOI22xp33_ASAP7_75t_L g2090 ( 
.A1(n_2072),
.A2(n_2049),
.B1(n_2065),
.B2(n_2068),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_2057),
.B(n_2050),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_2062),
.B(n_2033),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_2075),
.B(n_2024),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_2060),
.Y(n_2094)
);

OR2x2_ASAP7_75t_L g2095 ( 
.A(n_2063),
.B(n_2044),
.Y(n_2095)
);

OAI221xp5_ASAP7_75t_SL g2096 ( 
.A1(n_2079),
.A2(n_1982),
.B1(n_2039),
.B2(n_2044),
.C(n_2032),
.Y(n_2096)
);

OAI22xp33_ASAP7_75t_L g2097 ( 
.A1(n_2074),
.A2(n_1921),
.B1(n_2039),
.B2(n_2028),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_2061),
.Y(n_2098)
);

NAND4xp75_ASAP7_75t_L g2099 ( 
.A(n_2051),
.B(n_2043),
.C(n_2045),
.D(n_2049),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_2051),
.B(n_2043),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2067),
.Y(n_2101)
);

OAI221xp5_ASAP7_75t_L g2102 ( 
.A1(n_2077),
.A2(n_2035),
.B1(n_2036),
.B2(n_2045),
.C(n_2040),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2095),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_2091),
.B(n_2070),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_2083),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_2092),
.B(n_2033),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2080),
.Y(n_2107)
);

OAI21xp5_ASAP7_75t_L g2108 ( 
.A1(n_2080),
.A2(n_2073),
.B(n_2071),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_2085),
.B(n_2078),
.Y(n_2109)
);

INVxp67_ASAP7_75t_L g2110 ( 
.A(n_2086),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2093),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_2081),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2094),
.Y(n_2113)
);

OAI221xp5_ASAP7_75t_L g2114 ( 
.A1(n_2087),
.A2(n_2035),
.B1(n_2036),
.B2(n_2032),
.C(n_2042),
.Y(n_2114)
);

XOR2x2_ASAP7_75t_L g2115 ( 
.A(n_2084),
.B(n_2047),
.Y(n_2115)
);

INVxp67_ASAP7_75t_L g2116 ( 
.A(n_2088),
.Y(n_2116)
);

AOI22xp33_ASAP7_75t_L g2117 ( 
.A1(n_2088),
.A2(n_1986),
.B1(n_1990),
.B2(n_1970),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2103),
.Y(n_2118)
);

NOR3xp33_ASAP7_75t_L g2119 ( 
.A(n_2116),
.B(n_2099),
.C(n_2096),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_2106),
.Y(n_2120)
);

AND2x4_ASAP7_75t_L g2121 ( 
.A(n_2105),
.B(n_2100),
.Y(n_2121)
);

NOR2x1_ASAP7_75t_L g2122 ( 
.A(n_2107),
.B(n_2108),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_2115),
.Y(n_2123)
);

NOR4xp25_ASAP7_75t_L g2124 ( 
.A(n_2116),
.B(n_2096),
.C(n_2101),
.D(n_2098),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2104),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_2112),
.Y(n_2126)
);

OR2x2_ASAP7_75t_L g2127 ( 
.A(n_2109),
.B(n_2089),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_2110),
.B(n_2090),
.Y(n_2128)
);

AOI221xp5_ASAP7_75t_L g2129 ( 
.A1(n_2117),
.A2(n_2102),
.B1(n_2097),
.B2(n_2042),
.C(n_1990),
.Y(n_2129)
);

NAND2xp33_ASAP7_75t_L g2130 ( 
.A(n_2111),
.B(n_2047),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_2110),
.B(n_2037),
.Y(n_2131)
);

AOI322xp5_ASAP7_75t_L g2132 ( 
.A1(n_2119),
.A2(n_2113),
.A3(n_2097),
.B1(n_2114),
.B2(n_1885),
.C1(n_1893),
.C2(n_1882),
.Y(n_2132)
);

O2A1O1Ixp33_ASAP7_75t_SL g2133 ( 
.A1(n_2131),
.A2(n_2082),
.B(n_1901),
.C(n_2003),
.Y(n_2133)
);

OAI22xp33_ASAP7_75t_L g2134 ( 
.A1(n_2128),
.A2(n_1921),
.B1(n_1986),
.B2(n_2005),
.Y(n_2134)
);

OAI22xp5_ASAP7_75t_L g2135 ( 
.A1(n_2122),
.A2(n_2009),
.B1(n_2037),
.B2(n_1930),
.Y(n_2135)
);

AOI211xp5_ASAP7_75t_L g2136 ( 
.A1(n_2124),
.A2(n_2029),
.B(n_1806),
.C(n_1930),
.Y(n_2136)
);

NOR2x1_ASAP7_75t_L g2137 ( 
.A(n_2123),
.B(n_1971),
.Y(n_2137)
);

OAI211xp5_ASAP7_75t_SL g2138 ( 
.A1(n_2127),
.A2(n_2000),
.B(n_2006),
.C(n_1991),
.Y(n_2138)
);

NOR2x1_ASAP7_75t_L g2139 ( 
.A(n_2118),
.B(n_2126),
.Y(n_2139)
);

INVx1_ASAP7_75t_SL g2140 ( 
.A(n_2137),
.Y(n_2140)
);

NOR3xp33_ASAP7_75t_SL g2141 ( 
.A(n_2138),
.B(n_2125),
.C(n_2129),
.Y(n_2141)
);

NOR2x1_ASAP7_75t_L g2142 ( 
.A(n_2139),
.B(n_2121),
.Y(n_2142)
);

AOI211xp5_ASAP7_75t_L g2143 ( 
.A1(n_2136),
.A2(n_2124),
.B(n_2121),
.C(n_2130),
.Y(n_2143)
);

AOI222xp33_ASAP7_75t_L g2144 ( 
.A1(n_2135),
.A2(n_2134),
.B1(n_2120),
.B2(n_2132),
.C1(n_2005),
.C2(n_1900),
.Y(n_2144)
);

AOI21xp5_ASAP7_75t_L g2145 ( 
.A1(n_2133),
.A2(n_1991),
.B(n_1976),
.Y(n_2145)
);

NAND3xp33_ASAP7_75t_SL g2146 ( 
.A(n_2136),
.B(n_2029),
.C(n_2007),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2139),
.Y(n_2147)
);

NAND4xp75_ASAP7_75t_L g2148 ( 
.A(n_2142),
.B(n_2007),
.C(n_1976),
.D(n_2006),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_2147),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_2140),
.Y(n_2150)
);

OR2x2_ASAP7_75t_L g2151 ( 
.A(n_2146),
.B(n_1995),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2141),
.Y(n_2152)
);

INVx1_ASAP7_75t_SL g2153 ( 
.A(n_2145),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_2153),
.B(n_2143),
.Y(n_2154)
);

OAI31xp33_ASAP7_75t_L g2155 ( 
.A1(n_2152),
.A2(n_2144),
.A3(n_1930),
.B(n_1917),
.Y(n_2155)
);

OR3x2_ASAP7_75t_L g2156 ( 
.A(n_2152),
.B(n_1996),
.C(n_1995),
.Y(n_2156)
);

A2O1A1Ixp33_ASAP7_75t_L g2157 ( 
.A1(n_2150),
.A2(n_2003),
.B(n_2002),
.C(n_2000),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_2154),
.B(n_2149),
.Y(n_2158)
);

NOR2x1_ASAP7_75t_L g2159 ( 
.A(n_2157),
.B(n_2148),
.Y(n_2159)
);

AO22x1_ASAP7_75t_L g2160 ( 
.A1(n_2158),
.A2(n_2159),
.B1(n_2156),
.B2(n_2155),
.Y(n_2160)
);

OA21x2_ASAP7_75t_L g2161 ( 
.A1(n_2160),
.A2(n_2151),
.B(n_1998),
.Y(n_2161)
);

BUFx3_ASAP7_75t_L g2162 ( 
.A(n_2160),
.Y(n_2162)
);

AOI22xp5_ASAP7_75t_L g2163 ( 
.A1(n_2162),
.A2(n_2002),
.B1(n_1998),
.B2(n_1996),
.Y(n_2163)
);

HB1xp67_ASAP7_75t_L g2164 ( 
.A(n_2162),
.Y(n_2164)
);

AOI22xp33_ASAP7_75t_L g2165 ( 
.A1(n_2164),
.A2(n_2161),
.B1(n_1922),
.B2(n_1952),
.Y(n_2165)
);

OAI21xp5_ASAP7_75t_L g2166 ( 
.A1(n_2163),
.A2(n_2161),
.B(n_1946),
.Y(n_2166)
);

AOI21xp33_ASAP7_75t_SL g2167 ( 
.A1(n_2166),
.A2(n_1921),
.B(n_1922),
.Y(n_2167)
);

AO21x2_ASAP7_75t_L g2168 ( 
.A1(n_2167),
.A2(n_2165),
.B(n_1980),
.Y(n_2168)
);

XNOR2xp5_ASAP7_75t_L g2169 ( 
.A(n_2168),
.B(n_1968),
.Y(n_2169)
);

AOI221xp5_ASAP7_75t_L g2170 ( 
.A1(n_2169),
.A2(n_1948),
.B1(n_1950),
.B2(n_1945),
.C(n_1956),
.Y(n_2170)
);

AOI211xp5_ASAP7_75t_L g2171 ( 
.A1(n_2170),
.A2(n_1973),
.B(n_1968),
.C(n_1980),
.Y(n_2171)
);


endmodule