module fake_aes_58_n_18 (n_1, n_2, n_0, n_18);
input n_1;
input n_2;
input n_0;
output n_18;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_17;
wire n_5;
wire n_14;
wire n_8;
wire n_15;
wire n_10;
wire n_7;
CKINVDCx5p33_ASAP7_75t_R g3 ( .A(n_2), .Y(n_3) );
INVx1_ASAP7_75t_L g4 ( .A(n_0), .Y(n_4) );
INVx2_ASAP7_75t_L g5 ( .A(n_0), .Y(n_5) );
A2O1A1Ixp33_ASAP7_75t_L g6 ( .A1(n_4), .A2(n_0), .B(n_1), .C(n_2), .Y(n_6) );
OAI22x1_ASAP7_75t_L g7 ( .A1(n_3), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_7) );
AND2x4_ASAP7_75t_L g8 ( .A(n_4), .B(n_1), .Y(n_8) );
OR2x2_ASAP7_75t_L g9 ( .A(n_8), .B(n_5), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_8), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_9), .Y(n_11) );
NAND2xp5_ASAP7_75t_L g12 ( .A(n_10), .B(n_5), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_12), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_11), .B(n_6), .Y(n_14) );
NOR2x1_ASAP7_75t_L g15 ( .A(n_14), .B(n_11), .Y(n_15) );
AND2x2_ASAP7_75t_L g16 ( .A(n_13), .B(n_7), .Y(n_16) );
OAI21x1_ASAP7_75t_SL g17 ( .A1(n_15), .A2(n_13), .B(n_5), .Y(n_17) );
NAND2xp5_ASAP7_75t_SL g18 ( .A(n_17), .B(n_16), .Y(n_18) );
endmodule