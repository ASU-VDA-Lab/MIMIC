module fake_ariane_2754_n_823 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_823);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_823;

wire n_295;
wire n_356;
wire n_556;
wire n_190;
wire n_698;
wire n_695;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_423;
wire n_347;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_801;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_672;
wire n_487;
wire n_740;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_259;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_173;
wire n_242;
wire n_645;
wire n_320;
wire n_309;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_381;
wire n_344;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_821;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_780;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_181;
wire n_723;
wire n_617;
wire n_658;
wire n_616;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_747;
wire n_772;
wire n_741;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_742;
wire n_716;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_804;
wire n_280;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_793;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_428;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_317;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g172 ( 
.A(n_80),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_136),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_17),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_69),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_37),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_116),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_128),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_48),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_92),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_15),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_12),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_0),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_46),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_155),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_22),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

BUFx5_ASAP7_75t_L g188 ( 
.A(n_60),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_96),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_63),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_143),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_159),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_10),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_31),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_122),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_132),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_76),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_95),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_84),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_161),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_154),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_10),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_45),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_139),
.Y(n_204)
);

BUFx10_ASAP7_75t_L g205 ( 
.A(n_113),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_127),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_101),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_125),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_150),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_148),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_108),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_99),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_22),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_44),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_74),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_12),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_119),
.Y(n_217)
);

BUFx8_ASAP7_75t_SL g218 ( 
.A(n_8),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_137),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_64),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_152),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_88),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_41),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_67),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_55),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_146),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_141),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_157),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_26),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_151),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_153),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_166),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_193),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_218),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_188),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_181),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_208),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_228),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_186),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_183),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_183),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_194),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_202),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_190),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_229),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_190),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_204),
.Y(n_247)
);

INVxp67_ASAP7_75t_SL g248 ( 
.A(n_203),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_182),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_173),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_204),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_174),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_172),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_175),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_176),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_213),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_177),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_188),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_178),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_187),
.B(n_0),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_179),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_180),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_211),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_210),
.B(n_1),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_184),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_210),
.B(n_1),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_224),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_216),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_221),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_232),
.Y(n_270)
);

INVxp67_ASAP7_75t_SL g271 ( 
.A(n_203),
.Y(n_271)
);

NOR2xp67_ASAP7_75t_L g272 ( 
.A(n_185),
.B(n_2),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_222),
.Y(n_273)
);

INVxp33_ASAP7_75t_L g274 ( 
.A(n_227),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_189),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_205),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_205),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_221),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_205),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_244),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_252),
.Y(n_281)
);

NAND2xp33_ASAP7_75t_SL g282 ( 
.A(n_264),
.B(n_227),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_244),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_235),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_246),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_279),
.B(n_223),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_248),
.B(n_226),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_269),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_279),
.B(n_191),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_235),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_246),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_237),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_235),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_249),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_247),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_192),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_247),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_236),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_239),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_242),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_258),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_250),
.Y(n_302)
);

NAND2xp33_ASAP7_75t_R g303 ( 
.A(n_243),
.B(n_195),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_251),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_251),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_256),
.Y(n_306)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_264),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_254),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_238),
.Y(n_309)
);

INVx6_ASAP7_75t_L g310 ( 
.A(n_266),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_257),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_253),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_278),
.B(n_196),
.Y(n_313)
);

AND2x4_ASAP7_75t_L g314 ( 
.A(n_266),
.B(n_227),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_268),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_253),
.Y(n_316)
);

OR2x6_ASAP7_75t_L g317 ( 
.A(n_276),
.B(n_227),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_261),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_262),
.B(n_197),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_258),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_265),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_234),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_275),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_245),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_255),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_R g326 ( 
.A(n_277),
.B(n_231),
.Y(n_326)
);

NAND3xp33_ASAP7_75t_L g327 ( 
.A(n_276),
.B(n_199),
.C(n_198),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_277),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_255),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_259),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_307),
.B(n_259),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_281),
.Y(n_332)
);

OAI221xp5_ASAP7_75t_L g333 ( 
.A1(n_312),
.A2(n_233),
.B1(n_260),
.B2(n_263),
.C(n_270),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_316),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_328),
.A2(n_272),
.B1(n_263),
.B2(n_270),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_284),
.Y(n_336)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_320),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g338 ( 
.A(n_294),
.B(n_267),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_284),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_325),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_320),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_298),
.B(n_267),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_329),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_290),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_296),
.B(n_273),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_330),
.Y(n_346)
);

NAND2xp33_ASAP7_75t_SL g347 ( 
.A(n_302),
.B(n_200),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_307),
.B(n_273),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_290),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_299),
.B(n_274),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_320),
.Y(n_351)
);

NAND2x1p5_ASAP7_75t_L g352 ( 
.A(n_308),
.B(n_272),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_293),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_320),
.Y(n_354)
);

INVx4_ASAP7_75t_L g355 ( 
.A(n_314),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_311),
.B(n_201),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_307),
.B(n_319),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_280),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_314),
.B(n_206),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_293),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_281),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_324),
.B(n_240),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_288),
.B(n_207),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_300),
.B(n_240),
.Y(n_364)
);

OR2x2_ASAP7_75t_L g365 ( 
.A(n_302),
.B(n_318),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_287),
.B(n_258),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_301),
.Y(n_367)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_314),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_283),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_285),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_291),
.Y(n_371)
);

AND2x6_ASAP7_75t_L g372 ( 
.A(n_308),
.B(n_241),
.Y(n_372)
);

NAND2x1p5_ASAP7_75t_L g373 ( 
.A(n_286),
.B(n_289),
.Y(n_373)
);

OAI221xp5_ASAP7_75t_L g374 ( 
.A1(n_282),
.A2(n_241),
.B1(n_230),
.B2(n_225),
.C(n_220),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_301),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_292),
.Y(n_376)
);

OR2x6_ASAP7_75t_L g377 ( 
.A(n_317),
.B(n_2),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_318),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_295),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_297),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_321),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g382 ( 
.A(n_317),
.B(n_3),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_309),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_304),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_305),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_310),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_310),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_310),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_321),
.B(n_209),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_323),
.B(n_212),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_323),
.B(n_214),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_306),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_306),
.B(n_3),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_317),
.B(n_4),
.Y(n_394)
);

OR2x6_ASAP7_75t_L g395 ( 
.A(n_317),
.B(n_4),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_327),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_288),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_366),
.B(n_313),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_382),
.B(n_326),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_366),
.B(n_282),
.Y(n_400)
);

NOR2xp67_ASAP7_75t_L g401 ( 
.A(n_365),
.B(n_303),
.Y(n_401)
);

NAND2x1_ASAP7_75t_L g402 ( 
.A(n_372),
.B(n_188),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_357),
.B(n_215),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_382),
.B(n_188),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_360),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_334),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_345),
.B(n_217),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_345),
.B(n_348),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_340),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_350),
.B(n_322),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_355),
.B(n_368),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_355),
.B(n_5),
.Y(n_412)
);

INVx5_ASAP7_75t_L g413 ( 
.A(n_341),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_348),
.B(n_219),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_361),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_343),
.Y(n_416)
);

OR2x2_ASAP7_75t_L g417 ( 
.A(n_338),
.B(n_315),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_355),
.B(n_5),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_346),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_358),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_392),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_331),
.B(n_188),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g423 ( 
.A(n_342),
.B(n_378),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_L g424 ( 
.A1(n_382),
.A2(n_188),
.B1(n_315),
.B2(n_8),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_372),
.A2(n_188),
.B1(n_7),
.B2(n_9),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_332),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_376),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_372),
.A2(n_6),
.B1(n_11),
.B2(n_13),
.Y(n_428)
);

AO221x1_ASAP7_75t_L g429 ( 
.A1(n_377),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.C(n_15),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_368),
.B(n_14),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_368),
.B(n_16),
.Y(n_431)
);

INVxp67_ASAP7_75t_SL g432 ( 
.A(n_394),
.Y(n_432)
);

INVx8_ASAP7_75t_L g433 ( 
.A(n_372),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_397),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_362),
.B(n_16),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_372),
.B(n_17),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_364),
.B(n_18),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_360),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_369),
.B(n_18),
.Y(n_439)
);

INVx2_ASAP7_75t_SL g440 ( 
.A(n_397),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g441 ( 
.A(n_381),
.B(n_19),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_381),
.B(n_19),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_336),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_394),
.B(n_356),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_389),
.B(n_20),
.Y(n_445)
);

OR2x2_ASAP7_75t_SL g446 ( 
.A(n_393),
.B(n_20),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_370),
.B(n_21),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_337),
.A2(n_89),
.B(n_170),
.Y(n_448)
);

AND2x6_ASAP7_75t_SL g449 ( 
.A(n_390),
.B(n_21),
.Y(n_449)
);

AND2x6_ASAP7_75t_SL g450 ( 
.A(n_377),
.B(n_23),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_394),
.B(n_23),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_359),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_452)
);

AOI22xp33_ASAP7_75t_L g453 ( 
.A1(n_377),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_371),
.B(n_27),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_379),
.B(n_28),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_L g456 ( 
.A1(n_395),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_375),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_332),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_359),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_380),
.B(n_32),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_384),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_375),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_336),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_389),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_385),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_L g466 ( 
.A1(n_395),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_L g467 ( 
.A1(n_395),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_467)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_458),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_R g469 ( 
.A(n_433),
.B(n_376),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_434),
.B(n_386),
.Y(n_470)
);

BUFx4f_ASAP7_75t_L g471 ( 
.A(n_440),
.Y(n_471)
);

NAND2x1_ASAP7_75t_L g472 ( 
.A(n_457),
.B(n_337),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g473 ( 
.A(n_421),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_408),
.B(n_396),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_398),
.B(n_352),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_443),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_433),
.Y(n_477)
);

OR2x6_ASAP7_75t_L g478 ( 
.A(n_433),
.B(n_352),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_423),
.B(n_383),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_427),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_R g481 ( 
.A(n_434),
.B(n_383),
.Y(n_481)
);

A2O1A1Ixp33_ASAP7_75t_L g482 ( 
.A1(n_445),
.A2(n_333),
.B(n_335),
.C(n_396),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_406),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_410),
.B(n_363),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_401),
.B(n_337),
.Y(n_485)
);

BUFx2_ASAP7_75t_L g486 ( 
.A(n_415),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_413),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_417),
.B(n_391),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_432),
.B(n_407),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_409),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_443),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_442),
.Y(n_492)
);

CKINVDCx6p67_ASAP7_75t_R g493 ( 
.A(n_442),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_413),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_416),
.Y(n_495)
);

AO22x1_ASAP7_75t_L g496 ( 
.A1(n_445),
.A2(n_388),
.B1(n_387),
.B2(n_347),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g497 ( 
.A(n_441),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_411),
.B(n_391),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_449),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_411),
.B(n_373),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_451),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_414),
.B(n_373),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_463),
.Y(n_503)
);

INVx5_ASAP7_75t_L g504 ( 
.A(n_413),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_444),
.B(n_341),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_419),
.B(n_420),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_451),
.Y(n_507)
);

BUFx8_ASAP7_75t_L g508 ( 
.A(n_461),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_465),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_413),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_463),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_444),
.B(n_374),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_399),
.B(n_341),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_405),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_R g515 ( 
.A(n_400),
.B(n_347),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_412),
.B(n_339),
.Y(n_516)
);

NOR2xp67_ASAP7_75t_L g517 ( 
.A(n_399),
.B(n_339),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_412),
.B(n_344),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_462),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_450),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_438),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_422),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_475),
.B(n_424),
.Y(n_523)
);

AOI21x1_ASAP7_75t_L g524 ( 
.A1(n_496),
.A2(n_402),
.B(n_430),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_506),
.B(n_424),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_522),
.A2(n_448),
.B(n_436),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_498),
.B(n_500),
.Y(n_527)
);

INVx4_ASAP7_75t_L g528 ( 
.A(n_504),
.Y(n_528)
);

BUFx2_ASAP7_75t_L g529 ( 
.A(n_481),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_489),
.B(n_435),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_482),
.B(n_437),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_479),
.B(n_453),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_483),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_484),
.A2(n_426),
.B1(n_453),
.B2(n_456),
.Y(n_534)
);

AOI221xp5_ASAP7_75t_L g535 ( 
.A1(n_488),
.A2(n_456),
.B1(n_459),
.B2(n_452),
.C(n_466),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_482),
.B(n_418),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_501),
.B(n_418),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_490),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_476),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_495),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_509),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g542 ( 
.A1(n_474),
.A2(n_431),
.B(n_403),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_473),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_511),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_474),
.A2(n_431),
.B(n_439),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_516),
.A2(n_404),
.B(n_460),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_L g547 ( 
.A1(n_502),
.A2(n_455),
.B(n_454),
.Y(n_547)
);

OAI21x1_ASAP7_75t_L g548 ( 
.A1(n_522),
.A2(n_447),
.B(n_404),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_518),
.A2(n_467),
.B(n_466),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_501),
.B(n_507),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_504),
.Y(n_551)
);

OAI21xp33_ASAP7_75t_L g552 ( 
.A1(n_481),
.A2(n_428),
.B(n_425),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_485),
.A2(n_467),
.B(n_354),
.Y(n_553)
);

AO31x2_ASAP7_75t_L g554 ( 
.A1(n_512),
.A2(n_344),
.A3(n_367),
.B(n_349),
.Y(n_554)
);

NOR2xp67_ASAP7_75t_L g555 ( 
.A(n_504),
.B(n_464),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_485),
.A2(n_341),
.B(n_351),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_L g557 ( 
.A1(n_512),
.A2(n_367),
.B(n_353),
.Y(n_557)
);

OAI21x1_ASAP7_75t_L g558 ( 
.A1(n_476),
.A2(n_353),
.B(n_349),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_507),
.B(n_429),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_514),
.Y(n_560)
);

OAI21x1_ASAP7_75t_L g561 ( 
.A1(n_491),
.A2(n_375),
.B(n_354),
.Y(n_561)
);

AO31x2_ASAP7_75t_L g562 ( 
.A1(n_491),
.A2(n_375),
.A3(n_354),
.B(n_351),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_515),
.B(n_351),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_515),
.B(n_351),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_L g565 ( 
.A1(n_521),
.A2(n_354),
.B(n_43),
.Y(n_565)
);

OAI21x1_ASAP7_75t_L g566 ( 
.A1(n_503),
.A2(n_42),
.B(n_47),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_472),
.A2(n_49),
.B(n_50),
.Y(n_567)
);

OR2x2_ASAP7_75t_L g568 ( 
.A(n_523),
.B(n_492),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_539),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_L g570 ( 
.A1(n_549),
.A2(n_471),
.B(n_517),
.Y(n_570)
);

A2O1A1Ixp33_ASAP7_75t_L g571 ( 
.A1(n_535),
.A2(n_513),
.B(n_505),
.C(n_497),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_536),
.B(n_532),
.Y(n_572)
);

OAI21x1_ASAP7_75t_L g573 ( 
.A1(n_526),
.A2(n_503),
.B(n_519),
.Y(n_573)
);

OA21x2_ASAP7_75t_L g574 ( 
.A1(n_545),
.A2(n_505),
.B(n_513),
.Y(n_574)
);

AOI221x1_ASAP7_75t_L g575 ( 
.A1(n_536),
.A2(n_505),
.B1(n_513),
.B2(n_519),
.C(n_470),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g576 ( 
.A1(n_534),
.A2(n_493),
.B1(n_471),
.B2(n_480),
.Y(n_576)
);

OR2x2_ASAP7_75t_SL g577 ( 
.A(n_525),
.B(n_469),
.Y(n_577)
);

OAI21xp5_ASAP7_75t_L g578 ( 
.A1(n_527),
.A2(n_470),
.B(n_504),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_L g579 ( 
.A1(n_537),
.A2(n_532),
.B1(n_530),
.B2(n_531),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_533),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_543),
.B(n_480),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_552),
.A2(n_508),
.B1(n_559),
.B2(n_468),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_543),
.Y(n_583)
);

OAI21x1_ASAP7_75t_L g584 ( 
.A1(n_526),
.A2(n_519),
.B(n_510),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_528),
.B(n_478),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_544),
.B(n_470),
.Y(n_586)
);

OAI21x1_ASAP7_75t_L g587 ( 
.A1(n_561),
.A2(n_519),
.B(n_510),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_529),
.B(n_486),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_538),
.Y(n_589)
);

OAI21x1_ASAP7_75t_L g590 ( 
.A1(n_561),
.A2(n_510),
.B(n_494),
.Y(n_590)
);

AOI21xp5_ASAP7_75t_L g591 ( 
.A1(n_542),
.A2(n_478),
.B(n_510),
.Y(n_591)
);

OAI21x1_ASAP7_75t_SL g592 ( 
.A1(n_547),
.A2(n_469),
.B(n_520),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_540),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_560),
.A2(n_508),
.B1(n_478),
.B2(n_520),
.Y(n_594)
);

O2A1O1Ixp33_ASAP7_75t_L g595 ( 
.A1(n_550),
.A2(n_487),
.B(n_446),
.C(n_499),
.Y(n_595)
);

INVx6_ASAP7_75t_L g596 ( 
.A(n_551),
.Y(n_596)
);

OAI21x1_ASAP7_75t_L g597 ( 
.A1(n_566),
.A2(n_494),
.B(n_487),
.Y(n_597)
);

OAI21x1_ASAP7_75t_L g598 ( 
.A1(n_566),
.A2(n_494),
.B(n_477),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_541),
.Y(n_599)
);

OA21x2_ASAP7_75t_L g600 ( 
.A1(n_546),
.A2(n_494),
.B(n_52),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_539),
.B(n_477),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_528),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_551),
.Y(n_603)
);

INVx6_ASAP7_75t_L g604 ( 
.A(n_551),
.Y(n_604)
);

OR2x6_ASAP7_75t_L g605 ( 
.A(n_528),
.B(n_477),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_562),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_557),
.B(n_477),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_551),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_524),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_554),
.Y(n_610)
);

OAI221xp5_ASAP7_75t_L g611 ( 
.A1(n_582),
.A2(n_555),
.B1(n_565),
.B2(n_564),
.C(n_563),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_579),
.A2(n_548),
.B1(n_553),
.B2(n_558),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_SL g613 ( 
.A1(n_589),
.A2(n_548),
.B1(n_558),
.B2(n_567),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_572),
.B(n_562),
.Y(n_614)
);

INVx1_ASAP7_75t_SL g615 ( 
.A(n_583),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_589),
.A2(n_556),
.B1(n_562),
.B2(n_554),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_583),
.B(n_562),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_608),
.B(n_554),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_596),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_608),
.B(n_51),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_581),
.B(n_53),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_586),
.B(n_54),
.Y(n_622)
);

OR2x6_ASAP7_75t_L g623 ( 
.A(n_578),
.B(n_56),
.Y(n_623)
);

NAND2xp33_ASAP7_75t_SL g624 ( 
.A(n_602),
.B(n_57),
.Y(n_624)
);

AO21x1_ASAP7_75t_SL g625 ( 
.A1(n_570),
.A2(n_58),
.B(n_59),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_576),
.A2(n_61),
.B1(n_62),
.B2(n_65),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_568),
.A2(n_171),
.B1(n_68),
.B2(n_70),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_585),
.B(n_66),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_L g629 ( 
.A1(n_577),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_596),
.Y(n_630)
);

NOR2x1_ASAP7_75t_SL g631 ( 
.A(n_605),
.B(n_75),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_580),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_593),
.Y(n_633)
);

A2O1A1Ixp33_ASAP7_75t_L g634 ( 
.A1(n_571),
.A2(n_77),
.B(n_78),
.C(n_79),
.Y(n_634)
);

INVx3_ASAP7_75t_SL g635 ( 
.A(n_577),
.Y(n_635)
);

AOI21x1_ASAP7_75t_L g636 ( 
.A1(n_597),
.A2(n_81),
.B(n_82),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_599),
.Y(n_637)
);

NAND2xp33_ASAP7_75t_R g638 ( 
.A(n_600),
.B(n_574),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_596),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_L g640 ( 
.A1(n_588),
.A2(n_83),
.B1(n_85),
.B2(n_86),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_596),
.Y(n_641)
);

OAI221xp5_ASAP7_75t_L g642 ( 
.A1(n_568),
.A2(n_87),
.B1(n_90),
.B2(n_91),
.C(n_93),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_569),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_586),
.B(n_94),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_569),
.Y(n_645)
);

BUFx2_ASAP7_75t_L g646 ( 
.A(n_604),
.Y(n_646)
);

AOI21xp33_ASAP7_75t_L g647 ( 
.A1(n_610),
.A2(n_97),
.B(n_98),
.Y(n_647)
);

NAND2xp33_ASAP7_75t_L g648 ( 
.A(n_602),
.B(n_100),
.Y(n_648)
);

NAND3xp33_ASAP7_75t_SL g649 ( 
.A(n_595),
.B(n_102),
.C(n_103),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_604),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_L g651 ( 
.A1(n_594),
.A2(n_591),
.B1(n_602),
.B2(n_574),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_574),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_585),
.B(n_601),
.Y(n_653)
);

OAI22xp33_ASAP7_75t_L g654 ( 
.A1(n_575),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_585),
.B(n_107),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_603),
.B(n_109),
.Y(n_656)
);

OR2x6_ASAP7_75t_L g657 ( 
.A(n_607),
.B(n_110),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_604),
.B(n_603),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_604),
.Y(n_659)
);

INVx3_ASAP7_75t_SL g660 ( 
.A(n_605),
.Y(n_660)
);

OR2x2_ASAP7_75t_L g661 ( 
.A(n_606),
.B(n_111),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_654),
.A2(n_606),
.B1(n_592),
.B2(n_607),
.Y(n_662)
);

OAI22xp5_ASAP7_75t_L g663 ( 
.A1(n_627),
.A2(n_605),
.B1(n_609),
.B2(n_600),
.Y(n_663)
);

AOI221xp5_ASAP7_75t_L g664 ( 
.A1(n_654),
.A2(n_592),
.B1(n_609),
.B2(n_600),
.C(n_575),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_615),
.B(n_590),
.Y(n_665)
);

NOR4xp25_ASAP7_75t_L g666 ( 
.A(n_642),
.B(n_609),
.C(n_573),
.D(n_584),
.Y(n_666)
);

OA21x2_ASAP7_75t_L g667 ( 
.A1(n_612),
.A2(n_597),
.B(n_598),
.Y(n_667)
);

OR2x6_ASAP7_75t_L g668 ( 
.A(n_623),
.B(n_573),
.Y(n_668)
);

OAI221xp5_ASAP7_75t_L g669 ( 
.A1(n_626),
.A2(n_605),
.B1(n_598),
.B2(n_584),
.C(n_590),
.Y(n_669)
);

CKINVDCx16_ASAP7_75t_R g670 ( 
.A(n_620),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_627),
.A2(n_587),
.B1(n_114),
.B2(n_115),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_617),
.B(n_587),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_632),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_633),
.Y(n_674)
);

AOI221xp5_ASAP7_75t_L g675 ( 
.A1(n_649),
.A2(n_112),
.B1(n_117),
.B2(n_118),
.C(n_120),
.Y(n_675)
);

OAI22xp33_ASAP7_75t_L g676 ( 
.A1(n_642),
.A2(n_121),
.B1(n_123),
.B2(n_124),
.Y(n_676)
);

OAI21x1_ASAP7_75t_L g677 ( 
.A1(n_636),
.A2(n_612),
.B(n_651),
.Y(n_677)
);

INVx4_ASAP7_75t_L g678 ( 
.A(n_641),
.Y(n_678)
);

OAI22xp33_ASAP7_75t_L g679 ( 
.A1(n_623),
.A2(n_126),
.B1(n_129),
.B2(n_130),
.Y(n_679)
);

INVx2_ASAP7_75t_SL g680 ( 
.A(n_650),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_649),
.A2(n_131),
.B1(n_133),
.B2(n_134),
.Y(n_681)
);

BUFx2_ASAP7_75t_L g682 ( 
.A(n_635),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_618),
.A2(n_135),
.B1(n_138),
.B2(n_140),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_637),
.B(n_142),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_623),
.A2(n_144),
.B1(n_145),
.B2(n_147),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g686 ( 
.A1(n_620),
.A2(n_624),
.B1(n_657),
.B2(n_621),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_643),
.Y(n_687)
);

AOI221xp5_ASAP7_75t_L g688 ( 
.A1(n_634),
.A2(n_149),
.B1(n_158),
.B2(n_160),
.C(n_162),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_618),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_645),
.Y(n_690)
);

OR2x2_ASAP7_75t_L g691 ( 
.A(n_614),
.B(n_167),
.Y(n_691)
);

HB1xp67_ASAP7_75t_L g692 ( 
.A(n_652),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_SL g693 ( 
.A1(n_648),
.A2(n_168),
.B1(n_169),
.B2(n_611),
.Y(n_693)
);

AO221x2_ASAP7_75t_L g694 ( 
.A1(n_629),
.A2(n_640),
.B1(n_635),
.B2(n_653),
.C(n_624),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_646),
.B(n_658),
.Y(n_695)
);

OAI221xp5_ASAP7_75t_L g696 ( 
.A1(n_634),
.A2(n_616),
.B1(n_613),
.B2(n_611),
.C(n_657),
.Y(n_696)
);

AOI221xp5_ASAP7_75t_SL g697 ( 
.A1(n_658),
.A2(n_659),
.B1(n_630),
.B2(n_644),
.C(n_622),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_630),
.B(n_659),
.Y(n_698)
);

OAI22xp5_ASAP7_75t_L g699 ( 
.A1(n_657),
.A2(n_628),
.B1(n_661),
.B2(n_613),
.Y(n_699)
);

OAI22xp33_ASAP7_75t_L g700 ( 
.A1(n_638),
.A2(n_660),
.B1(n_628),
.B2(n_619),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_687),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_696),
.A2(n_625),
.B1(n_647),
.B2(n_655),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_672),
.B(n_639),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_690),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_692),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_665),
.B(n_631),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_692),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_673),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_674),
.Y(n_709)
);

BUFx2_ASAP7_75t_L g710 ( 
.A(n_682),
.Y(n_710)
);

INVx4_ASAP7_75t_R g711 ( 
.A(n_680),
.Y(n_711)
);

HB1xp67_ASAP7_75t_L g712 ( 
.A(n_695),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_668),
.Y(n_713)
);

OR2x2_ASAP7_75t_L g714 ( 
.A(n_670),
.B(n_660),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_668),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_668),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_667),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_667),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_677),
.B(n_656),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_697),
.B(n_638),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_694),
.A2(n_699),
.B1(n_676),
.B2(n_693),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_698),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_666),
.B(n_662),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_662),
.B(n_664),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_691),
.B(n_700),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_669),
.Y(n_726)
);

AND2x4_ASAP7_75t_L g727 ( 
.A(n_678),
.B(n_686),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_700),
.Y(n_728)
);

OR2x2_ASAP7_75t_L g729 ( 
.A(n_694),
.B(n_678),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_703),
.B(n_663),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_703),
.B(n_693),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_707),
.Y(n_732)
);

AO21x2_ASAP7_75t_L g733 ( 
.A1(n_723),
.A2(n_676),
.B(n_679),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_707),
.Y(n_734)
);

HB1xp67_ASAP7_75t_L g735 ( 
.A(n_705),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_705),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_705),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_717),
.Y(n_738)
);

OAI22xp33_ASAP7_75t_L g739 ( 
.A1(n_726),
.A2(n_679),
.B1(n_671),
.B2(n_688),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_704),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_717),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_710),
.Y(n_742)
);

NOR4xp25_ASAP7_75t_SL g743 ( 
.A(n_710),
.B(n_675),
.C(n_685),
.D(n_681),
.Y(n_743)
);

OAI211xp5_ASAP7_75t_SL g744 ( 
.A1(n_721),
.A2(n_681),
.B(n_685),
.C(n_684),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_704),
.Y(n_745)
);

AND4x1_ASAP7_75t_L g746 ( 
.A(n_723),
.B(n_683),
.C(n_689),
.D(n_724),
.Y(n_746)
);

OAI21x1_ASAP7_75t_L g747 ( 
.A1(n_718),
.A2(n_726),
.B(n_720),
.Y(n_747)
);

OAI22xp5_ASAP7_75t_L g748 ( 
.A1(n_702),
.A2(n_729),
.B1(n_724),
.B2(n_726),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_740),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_732),
.B(n_708),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_732),
.B(n_734),
.Y(n_751)
);

OAI21x1_ASAP7_75t_L g752 ( 
.A1(n_747),
.A2(n_718),
.B(n_728),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_742),
.B(n_712),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_740),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_742),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_730),
.B(n_729),
.Y(n_756)
);

AND3x2_ASAP7_75t_L g757 ( 
.A(n_731),
.B(n_727),
.C(n_728),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_730),
.B(n_727),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_735),
.B(n_727),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_734),
.B(n_708),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_736),
.B(n_727),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_733),
.B(n_713),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_761),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_761),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_758),
.B(n_731),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_762),
.A2(n_733),
.B1(n_744),
.B2(n_748),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_758),
.B(n_733),
.Y(n_767)
);

OR2x2_ASAP7_75t_L g768 ( 
.A(n_753),
.B(n_733),
.Y(n_768)
);

OAI322xp33_ASAP7_75t_L g769 ( 
.A1(n_766),
.A2(n_756),
.A3(n_739),
.B1(n_760),
.B2(n_750),
.C1(n_751),
.C2(n_754),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_765),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_763),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_764),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_767),
.B(n_753),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_770),
.B(n_766),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_770),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_773),
.Y(n_776)
);

INVx3_ASAP7_75t_SL g777 ( 
.A(n_773),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_777),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_776),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_778),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_779),
.B(n_775),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_778),
.Y(n_782)
);

O2A1O1Ixp33_ASAP7_75t_L g783 ( 
.A1(n_780),
.A2(n_774),
.B(n_769),
.C(n_768),
.Y(n_783)
);

NOR2x1_ASAP7_75t_L g784 ( 
.A(n_782),
.B(n_774),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_781),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_781),
.B(n_772),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_781),
.B(n_771),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_785),
.B(n_755),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_784),
.A2(n_743),
.B(n_751),
.Y(n_789)
);

AND4x1_ASAP7_75t_L g790 ( 
.A(n_786),
.B(n_711),
.C(n_759),
.D(n_743),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_787),
.B(n_760),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_783),
.A2(n_762),
.B1(n_747),
.B2(n_757),
.Y(n_792)
);

O2A1O1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_784),
.A2(n_762),
.B(n_746),
.C(n_750),
.Y(n_793)
);

OAI211xp5_ASAP7_75t_SL g794 ( 
.A1(n_793),
.A2(n_711),
.B(n_714),
.C(n_746),
.Y(n_794)
);

AOI311xp33_ASAP7_75t_L g795 ( 
.A1(n_791),
.A2(n_754),
.A3(n_749),
.B(n_736),
.C(n_737),
.Y(n_795)
);

NOR3xp33_ASAP7_75t_L g796 ( 
.A(n_789),
.B(n_752),
.C(n_762),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_788),
.Y(n_797)
);

NAND4xp25_ASAP7_75t_L g798 ( 
.A(n_792),
.B(n_714),
.C(n_759),
.D(n_706),
.Y(n_798)
);

OAI211xp5_ASAP7_75t_L g799 ( 
.A1(n_797),
.A2(n_790),
.B(n_749),
.C(n_737),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_796),
.B(n_706),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_794),
.A2(n_719),
.B1(n_752),
.B2(n_725),
.Y(n_801)
);

BUFx2_ASAP7_75t_L g802 ( 
.A(n_798),
.Y(n_802)
);

NOR2xp67_ASAP7_75t_L g803 ( 
.A(n_795),
.B(n_701),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_797),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_804),
.B(n_701),
.Y(n_805)
);

OAI221xp5_ASAP7_75t_L g806 ( 
.A1(n_799),
.A2(n_725),
.B1(n_741),
.B2(n_738),
.C(n_709),
.Y(n_806)
);

NAND4xp75_ASAP7_75t_L g807 ( 
.A(n_803),
.B(n_801),
.C(n_802),
.D(n_800),
.Y(n_807)
);

OA22x2_ASAP7_75t_L g808 ( 
.A1(n_804),
.A2(n_719),
.B1(n_716),
.B2(n_715),
.Y(n_808)
);

INVxp67_ASAP7_75t_L g809 ( 
.A(n_804),
.Y(n_809)
);

XNOR2xp5_ASAP7_75t_L g810 ( 
.A(n_807),
.B(n_719),
.Y(n_810)
);

NOR2x1_ASAP7_75t_L g811 ( 
.A(n_805),
.B(n_719),
.Y(n_811)
);

CKINVDCx20_ASAP7_75t_R g812 ( 
.A(n_809),
.Y(n_812)
);

AND2x4_ASAP7_75t_L g813 ( 
.A(n_808),
.B(n_722),
.Y(n_813)
);

NAND3xp33_ASAP7_75t_SL g814 ( 
.A(n_806),
.B(n_715),
.C(n_716),
.Y(n_814)
);

INVxp67_ASAP7_75t_SL g815 ( 
.A(n_809),
.Y(n_815)
);

XNOR2xp5_ASAP7_75t_L g816 ( 
.A(n_812),
.B(n_713),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_816),
.B(n_815),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_817),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_818),
.Y(n_819)
);

INVxp67_ASAP7_75t_L g820 ( 
.A(n_819),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_820),
.A2(n_818),
.B1(n_811),
.B2(n_810),
.Y(n_821)
);

OAI221xp5_ASAP7_75t_R g822 ( 
.A1(n_821),
.A2(n_814),
.B1(n_813),
.B2(n_745),
.C(n_738),
.Y(n_822)
);

AOI211xp5_ASAP7_75t_L g823 ( 
.A1(n_822),
.A2(n_745),
.B(n_741),
.C(n_738),
.Y(n_823)
);


endmodule