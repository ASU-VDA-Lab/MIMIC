module real_jpeg_28630_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_202;
wire n_128;
wire n_216;
wire n_179;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_206;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_0),
.A2(n_36),
.B1(n_41),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_0),
.A2(n_46),
.B1(n_54),
.B2(n_55),
.Y(n_126)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_1),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_61),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_2),
.A2(n_36),
.B1(n_41),
.B2(n_61),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_2),
.A2(n_54),
.B1(n_55),
.B2(n_61),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_3),
.A2(n_36),
.B1(n_41),
.B2(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_3),
.Y(n_124)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_5),
.A2(n_36),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_5),
.A2(n_42),
.B1(n_54),
.B2(n_55),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_6),
.A2(n_36),
.B1(n_41),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_6),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_8),
.A2(n_54),
.B1(n_55),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_8),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_85),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_8),
.A2(n_36),
.B1(n_41),
.B2(n_85),
.Y(n_143)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

O2A1O1Ixp33_ASAP7_75t_SL g23 ( 
.A1(n_10),
.A2(n_24),
.B(n_25),
.C(n_30),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_10),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_10),
.B(n_72),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_10),
.B(n_55),
.Y(n_155)
);

A2O1A1O1Ixp25_ASAP7_75t_L g157 ( 
.A1(n_10),
.A2(n_55),
.B(n_87),
.C(n_155),
.D(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_10),
.B(n_52),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_10),
.A2(n_35),
.B(n_168),
.Y(n_187)
);

A2O1A1O1Ixp25_ASAP7_75t_L g199 ( 
.A1(n_10),
.A2(n_28),
.B(n_51),
.C(n_63),
.D(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_10),
.B(n_28),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_65),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_11),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_65),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_11),
.A2(n_54),
.B1(n_55),
.B2(n_65),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_11),
.A2(n_36),
.B1(n_41),
.B2(n_65),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_12),
.A2(n_30),
.B1(n_31),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_12),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_70),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_12),
.A2(n_54),
.B1(n_55),
.B2(n_70),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_12),
.A2(n_36),
.B1(n_41),
.B2(n_70),
.Y(n_175)
);

O2A1O1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_13),
.A2(n_55),
.B(n_88),
.C(n_91),
.Y(n_87)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_13),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_13),
.B(n_36),
.Y(n_156)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_15),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

INVx11_ASAP7_75t_SL g37 ( 
.A(n_16),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_132),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_130),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_107),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_20),
.B(n_107),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_78),
.C(n_94),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_21),
.B(n_147),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_47),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_22),
.B(n_48),
.C(n_77),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_32),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_23),
.A2(n_32),
.B1(n_33),
.B2(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_23),
.Y(n_139)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_24),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_24),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B(n_28),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_26),
.B(n_93),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_26),
.B(n_190),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_28),
.A2(n_29),
.B1(n_53),
.B2(n_57),
.Y(n_56)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI32xp33_ASAP7_75t_L g207 ( 
.A1(n_29),
.A2(n_55),
.A3(n_200),
.B1(n_208),
.B2(n_210),
.Y(n_207)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_39),
.B1(n_43),
.B2(n_45),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_34),
.A2(n_174),
.B1(n_176),
.B2(n_177),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_35),
.A2(n_44),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_35),
.A2(n_81),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_35),
.A2(n_40),
.B1(n_44),
.B2(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_35),
.A2(n_167),
.B(n_168),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_35),
.B(n_170),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_36),
.A2(n_41),
.B1(n_89),
.B2(n_90),
.Y(n_91)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI32xp33_ASAP7_75t_L g154 ( 
.A1(n_41),
.A2(n_54),
.A3(n_90),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_41),
.B(n_189),
.Y(n_188)
);

INVx5_ASAP7_75t_SL g122 ( 
.A(n_43),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_43),
.B(n_169),
.Y(n_168)
);

INVx11_ASAP7_75t_L g178 ( 
.A(n_43),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_43),
.A2(n_185),
.B(n_206),
.Y(n_205)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_45),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_67),
.B2(n_77),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_59),
.B(n_62),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_51),
.A2(n_52),
.B1(n_60),
.B2(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_51),
.B(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_56),
.Y(n_51)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_53),
.Y(n_209)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

NAND2xp33_ASAP7_75t_SL g210 ( 
.A(n_54),
.B(n_209),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_55),
.B(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_64),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_66),
.A2(n_117),
.B(n_118),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_66),
.A2(n_106),
.B(n_118),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_67),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_71),
.B(n_73),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_69),
.A2(n_72),
.B1(n_74),
.B2(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_72),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_72),
.B(n_76),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_76),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_74),
.A2(n_101),
.B(n_102),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_78),
.B(n_94),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_83),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_83),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_86),
.B1(n_92),
.B2(n_93),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_84),
.A2(n_93),
.B(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_86),
.A2(n_92),
.B1(n_93),
.B2(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_86),
.A2(n_221),
.B(n_222),
.Y(n_220)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_87),
.B(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_87),
.A2(n_91),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_93),
.B(n_99),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_93),
.A2(n_97),
.B(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_100),
.C(n_104),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_95),
.A2(n_96),
.B1(n_104),
.B2(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_100),
.B(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_107)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_120),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_115),
.B2(n_116),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.Y(n_120)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_127),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_148),
.B(n_229),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_146),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_134),
.B(n_146),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_138),
.C(n_140),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_135),
.B(n_227),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_138),
.B(n_140),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.C(n_144),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_141),
.B(n_216),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_142),
.A2(n_144),
.B1(n_145),
.B2(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_142),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_143),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_224),
.B(n_228),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_212),
.B(n_223),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_195),
.B(n_211),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_171),
.B(n_194),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_159),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_153),
.B(n_159),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_157),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_158),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_166),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_164),
.C(n_166),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_165),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_167),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_180),
.B(n_193),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_179),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_173),
.B(n_179),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_175),
.A2(n_178),
.B(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_186),
.B(n_192),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_182),
.B(n_183),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_196),
.B(n_197),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_204),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_201),
.C(n_204),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_203),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_207),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_207),
.Y(n_219)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_213),
.B(n_214),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_218),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_219),
.C(n_220),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_225),
.B(n_226),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);


endmodule