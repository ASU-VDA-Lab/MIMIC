module fake_jpeg_28586_n_353 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_353);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_353;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_37),
.Y(n_81)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_47),
.Y(n_60)
);

BUFx2_ASAP7_75t_R g45 ( 
.A(n_19),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_50),
.Y(n_78)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_19),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

CKINVDCx6p67_ASAP7_75t_R g53 ( 
.A(n_49),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_34),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_49),
.A2(n_23),
.B1(n_28),
.B2(n_32),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_54),
.A2(n_59),
.B1(n_67),
.B2(n_75),
.Y(n_95)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_30),
.B1(n_33),
.B2(n_32),
.Y(n_59)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_45),
.A2(n_30),
.B1(n_34),
.B2(n_35),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_68),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_48),
.A2(n_34),
.B1(n_35),
.B2(n_28),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_48),
.A2(n_34),
.B1(n_28),
.B2(n_27),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_16),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_66),
.B(n_80),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_38),
.A2(n_36),
.B1(n_33),
.B2(n_32),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_40),
.A2(n_28),
.B1(n_19),
.B2(n_18),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_42),
.A2(n_47),
.B(n_19),
.C(n_18),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_70),
.A2(n_77),
.B(n_73),
.C(n_60),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_40),
.A2(n_28),
.B1(n_19),
.B2(n_18),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_71),
.A2(n_79),
.B1(n_37),
.B2(n_41),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_44),
.A2(n_24),
.B1(n_17),
.B2(n_29),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_17),
.C(n_25),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_16),
.B1(n_24),
.B2(n_29),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_26),
.B1(n_25),
.B2(n_22),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_28),
.B1(n_33),
.B2(n_36),
.Y(n_75)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_38),
.B(n_26),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_21),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_40),
.A2(n_36),
.B1(n_22),
.B2(n_21),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_46),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_66),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_82),
.B(n_88),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_86),
.A2(n_89),
.B1(n_114),
.B2(n_81),
.Y(n_145)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

OR2x2_ASAP7_75t_SL g89 ( 
.A(n_73),
.B(n_46),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_52),
.A2(n_37),
.B1(n_41),
.B2(n_22),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_91),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_92),
.A2(n_104),
.B1(n_111),
.B2(n_119),
.Y(n_128)
);

BUFx4f_ASAP7_75t_SL g93 ( 
.A(n_53),
.Y(n_93)
);

INVx4_ASAP7_75t_SL g139 ( 
.A(n_93),
.Y(n_139)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_96),
.B(n_105),
.Y(n_123)
);

AO22x1_ASAP7_75t_SL g97 ( 
.A1(n_70),
.A2(n_43),
.B1(n_50),
.B2(n_51),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_53),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_60),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_100),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_70),
.B(n_69),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_109),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_56),
.B(n_15),
.Y(n_100)
);

INVxp33_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_102),
.Y(n_141)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_54),
.A2(n_51),
.B1(n_50),
.B2(n_43),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_108),
.Y(n_142)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_21),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_74),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_115),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_59),
.A2(n_51),
.B1(n_43),
.B2(n_14),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_56),
.B(n_13),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_113),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_56),
.B(n_78),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_81),
.A2(n_13),
.B1(n_1),
.B2(n_2),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_76),
.A2(n_62),
.B1(n_65),
.B2(n_63),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_116),
.A2(n_2),
.B(n_3),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_78),
.B(n_0),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_120),
.Y(n_140)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_121),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_67),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_80),
.B(n_76),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_76),
.B(n_61),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_122),
.A2(n_145),
.B(n_113),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_107),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_147),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_115),
.A2(n_79),
.B1(n_71),
.B2(n_68),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_126),
.A2(n_130),
.B1(n_135),
.B2(n_137),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_96),
.A2(n_56),
.B(n_53),
.C(n_75),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_129),
.A2(n_148),
.B(n_112),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_110),
.A2(n_57),
.B1(n_64),
.B2(n_53),
.Y(n_130)
);

AO21x1_ASAP7_75t_L g154 ( 
.A1(n_133),
.A2(n_120),
.B(n_85),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_57),
.B1(n_53),
.B2(n_58),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_84),
.A2(n_57),
.B1(n_53),
.B2(n_58),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_58),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_146),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_83),
.B(n_1),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_83),
.B(n_12),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_97),
.B(n_2),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_152),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_82),
.B(n_3),
.Y(n_152)
);

AO22x1_ASAP7_75t_L g205 ( 
.A1(n_154),
.A2(n_122),
.B1(n_125),
.B2(n_133),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_97),
.B1(n_85),
.B2(n_98),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_156),
.A2(n_160),
.B1(n_162),
.B2(n_186),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_157),
.A2(n_139),
.B(n_5),
.Y(n_217)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_158),
.Y(n_193)
);

AO22x1_ASAP7_75t_SL g159 ( 
.A1(n_149),
.A2(n_97),
.B1(n_89),
.B2(n_95),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_175),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_128),
.A2(n_95),
.B1(n_107),
.B2(n_109),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_119),
.B(n_117),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_165),
.B(n_170),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_128),
.A2(n_88),
.B1(n_111),
.B2(n_87),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_127),
.Y(n_164)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_164),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_144),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_166),
.B(n_168),
.Y(n_199)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_167),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_124),
.B(n_94),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_169),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_129),
.A2(n_92),
.B(n_106),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_134),
.Y(n_171)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_171),
.Y(n_203)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_172),
.Y(n_214)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_174),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_103),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_103),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_178),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_129),
.A2(n_102),
.B(n_103),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_145),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_90),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_139),
.A2(n_118),
.B1(n_108),
.B2(n_121),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_SL g204 ( 
.A1(n_179),
.A2(n_137),
.B(n_139),
.C(n_93),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_136),
.B(n_93),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_185),
.Y(n_208)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_142),
.Y(n_181)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_134),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_182),
.Y(n_194)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_183),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_144),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_184),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_143),
.B(n_93),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_149),
.A2(n_133),
.B1(n_123),
.B2(n_145),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_123),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_188),
.B(n_201),
.C(n_216),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_156),
.A2(n_126),
.B1(n_135),
.B2(n_148),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_192),
.A2(n_212),
.B1(n_173),
.B2(n_184),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_161),
.A2(n_148),
.B(n_122),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_196),
.A2(n_204),
.B(n_185),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_197),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_125),
.C(n_140),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_180),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_213),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_205),
.B(n_159),
.Y(n_234)
);

OA21x2_ASAP7_75t_L g207 ( 
.A1(n_177),
.A2(n_141),
.B(n_131),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_207),
.A2(n_217),
.B(n_155),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_153),
.B(n_132),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_211),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_163),
.B(n_140),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_210),
.B(n_205),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_169),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_162),
.A2(n_130),
.B1(n_104),
.B2(n_132),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_169),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_173),
.A2(n_131),
.B1(n_152),
.B2(n_141),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_215),
.A2(n_160),
.B1(n_153),
.B2(n_155),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_163),
.B(n_151),
.Y(n_216)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_221),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_222),
.A2(n_233),
.B1(n_190),
.B2(n_159),
.Y(n_255)
);

BUFx5_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_224),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_168),
.Y(n_226)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_226),
.Y(n_260)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_198),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_228),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_178),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_230),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_231),
.A2(n_187),
.B1(n_206),
.B2(n_189),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_192),
.A2(n_173),
.B1(n_212),
.B2(n_187),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_235),
.Y(n_253)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_214),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_193),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_236),
.B(n_237),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_219),
.B(n_166),
.Y(n_237)
);

AOI32xp33_ASAP7_75t_L g238 ( 
.A1(n_190),
.A2(n_197),
.A3(n_196),
.B1(n_217),
.B2(n_205),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_238),
.B(n_242),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_188),
.B(n_165),
.C(n_183),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_241),
.Y(n_261)
);

AOI21x1_ASAP7_75t_L g264 ( 
.A1(n_240),
.A2(n_245),
.B(n_246),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_201),
.B(n_181),
.C(n_174),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_218),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_176),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_243),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_154),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_244),
.B(n_248),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_245),
.A2(n_203),
.B(n_200),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_220),
.B(n_175),
.Y(n_246)
);

OAI322xp33_ASAP7_75t_L g265 ( 
.A1(n_246),
.A2(n_208),
.A3(n_206),
.B1(n_154),
.B2(n_204),
.C1(n_167),
.C2(n_158),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_220),
.B(n_170),
.Y(n_247)
);

INVxp67_ASAP7_75t_SL g256 ( 
.A(n_247),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_249),
.A2(n_257),
.B1(n_272),
.B2(n_225),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_224),
.Y(n_251)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_251),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_255),
.A2(n_263),
.B1(n_266),
.B2(n_179),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_234),
.A2(n_189),
.B1(n_207),
.B2(n_208),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_239),
.B(n_210),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_259),
.B(n_242),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_236),
.Y(n_262)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_262),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_222),
.A2(n_207),
.B1(n_159),
.B2(n_204),
.Y(n_263)
);

HB1xp67_ASAP7_75t_SL g278 ( 
.A(n_264),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_265),
.A2(n_237),
.B1(n_240),
.B2(n_231),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_233),
.A2(n_204),
.B1(n_164),
.B2(n_172),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_229),
.B(n_203),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_171),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_272),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_264),
.Y(n_299)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_269),
.Y(n_275)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_275),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_229),
.C(n_241),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_277),
.C(n_279),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_232),
.C(n_244),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_232),
.C(n_248),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_260),
.A2(n_225),
.B1(n_223),
.B2(n_235),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_280),
.A2(n_287),
.B1(n_291),
.B2(n_267),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_283),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_271),
.A2(n_238),
.B1(n_221),
.B2(n_230),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_289),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_257),
.A2(n_227),
.B1(n_200),
.B2(n_194),
.Y(n_285)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_285),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_182),
.C(n_171),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_258),
.C(n_263),
.Y(n_301)
);

INVxp33_ASAP7_75t_L g288 ( 
.A(n_269),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_288),
.Y(n_310)
);

A2O1A1O1Ixp25_ASAP7_75t_L g290 ( 
.A1(n_253),
.A2(n_139),
.B(n_169),
.C(n_7),
.D(n_8),
.Y(n_290)
);

NAND4xp25_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_266),
.C(n_256),
.D(n_250),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_255),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_268),
.B(n_4),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_293),
.B(n_252),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_294),
.B(n_297),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_281),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_307),
.C(n_295),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_258),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_303),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_276),
.B(n_253),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_305),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_254),
.C(n_7),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_278),
.A2(n_6),
.B(n_7),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_306),
.A2(n_291),
.B(n_8),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_279),
.B(n_277),
.C(n_284),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_309),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_283),
.B(n_6),
.C(n_8),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_311),
.B(n_312),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_287),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_313),
.B(n_315),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_285),
.Y(n_315)
);

INVx5_ASAP7_75t_L g316 ( 
.A(n_299),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_317),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_292),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_295),
.B(n_275),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_318),
.B(n_324),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_320),
.A2(n_273),
.B1(n_8),
.B2(n_9),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_298),
.B(n_282),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_298),
.C(n_296),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_305),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_325),
.B(n_331),
.C(n_312),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_310),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_326),
.B(n_330),
.Y(n_338)
);

A2O1A1Ixp33_ASAP7_75t_SL g327 ( 
.A1(n_311),
.A2(n_288),
.B(n_300),
.C(n_308),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_327),
.A2(n_316),
.B1(n_324),
.B2(n_315),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_323),
.B(n_273),
.Y(n_330)
);

FAx1_ASAP7_75t_SL g331 ( 
.A(n_321),
.B(n_309),
.CI(n_290),
.CON(n_331),
.SN(n_331)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_332),
.B(n_11),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_319),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_333),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_340)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_336),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_334),
.B(n_314),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_337),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_339),
.B(n_343),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_340),
.B(n_342),
.Y(n_344)
);

AOI221x1_ASAP7_75t_L g341 ( 
.A1(n_327),
.A2(n_326),
.B1(n_331),
.B2(n_329),
.C(n_325),
.Y(n_341)
);

AOI322xp5_ASAP7_75t_L g345 ( 
.A1(n_341),
.A2(n_12),
.A3(n_327),
.B1(n_328),
.B2(n_338),
.C1(n_336),
.C2(n_337),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_335),
.B(n_11),
.Y(n_343)
);

OAI21x1_ASAP7_75t_SL g350 ( 
.A1(n_345),
.A2(n_344),
.B(n_348),
.Y(n_350)
);

OAI21xp33_ASAP7_75t_L g349 ( 
.A1(n_347),
.A2(n_327),
.B(n_328),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_349),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_351),
.A2(n_350),
.B(n_348),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_352),
.B(n_346),
.Y(n_353)
);


endmodule