module fake_ibex_1690_n_2003 (n_151, n_85, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_108, n_350, n_165, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_357, n_88, n_412, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_421, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_417, n_265, n_158, n_259, n_276, n_339, n_210, n_348, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_384, n_373, n_244, n_73, n_343, n_310, n_426, n_323, n_143, n_106, n_386, n_8, n_224, n_183, n_67, n_333, n_110, n_306, n_400, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_434, n_296, n_120, n_168, n_155, n_315, n_13, n_122, n_116, n_370, n_431, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_22, n_136, n_261, n_30, n_367, n_221, n_437, n_355, n_407, n_102, n_52, n_99, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_420, n_141, n_222, n_186, n_349, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_427, n_157, n_219, n_246, n_31, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_139, n_429, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_347, n_335, n_413, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_257, n_77, n_44, n_401, n_66, n_305, n_307, n_192, n_140, n_416, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_26, n_188, n_200, n_199, n_410, n_308, n_411, n_135, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_225, n_360, n_272, n_23, n_223, n_381, n_382, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_378, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_303, n_362, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_345, n_408, n_119, n_361, n_419, n_72, n_319, n_195, n_212, n_311, n_406, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_344, n_393, n_436, n_428, n_297, n_435, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_399, n_254, n_213, n_424, n_271, n_241, n_68, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_380, n_281, n_425, n_2003);

input n_151;
input n_85;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_108;
input n_350;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_417;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_210;
input n_348;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_67;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_434;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_13;
input n_122;
input n_116;
input n_370;
input n_431;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_367;
input n_221;
input n_437;
input n_355;
input n_407;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_141;
input n_222;
input n_186;
input n_349;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_427;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_139;
input n_429;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_347;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_257;
input n_77;
input n_44;
input n_401;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_416;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_26;
input n_188;
input n_200;
input n_199;
input n_410;
input n_308;
input n_411;
input n_135;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_225;
input n_360;
input n_272;
input n_23;
input n_223;
input n_381;
input n_382;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_378;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_345;
input n_408;
input n_119;
input n_361;
input n_419;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_344;
input n_393;
input n_436;
input n_428;
input n_297;
input n_435;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_399;
input n_254;
input n_213;
input n_424;
input n_271;
input n_241;
input n_68;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_380;
input n_281;
input n_425;

output n_2003;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_1983;
wire n_992;
wire n_1582;
wire n_766;
wire n_1110;
wire n_1382;
wire n_1998;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_1930;
wire n_452;
wire n_1234;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_1954;
wire n_1883;
wire n_1125;
wire n_733;
wire n_622;
wire n_1226;
wire n_1034;
wire n_1765;
wire n_872;
wire n_1873;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_1722;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_1391;
wire n_884;
wire n_667;
wire n_850;
wire n_1971;
wire n_879;
wire n_1957;
wire n_723;
wire n_1144;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_1766;
wire n_550;
wire n_1922;
wire n_557;
wire n_641;
wire n_1937;
wire n_893;
wire n_527;
wire n_1654;
wire n_496;
wire n_1258;
wire n_1344;
wire n_1929;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_824;
wire n_1945;
wire n_441;
wire n_694;
wire n_787;
wire n_523;
wire n_614;
wire n_1130;
wire n_1228;
wire n_1081;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_1926;
wire n_904;
wire n_1970;
wire n_1778;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_1910;
wire n_715;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_1606;
wire n_769;
wire n_1595;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_1886;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_777;
wire n_1955;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_558;
wire n_666;
wire n_1638;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_793;
wire n_937;
wire n_1645;
wire n_973;
wire n_1038;
wire n_618;
wire n_1943;
wire n_1863;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_1588;
wire n_1301;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_553;
wire n_554;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_745;
wire n_447;
wire n_1753;
wire n_562;
wire n_564;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_978;
wire n_579;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_1936;
wire n_1717;
wire n_1609;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_695;
wire n_1549;
wire n_639;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_1742;
wire n_1818;
wire n_870;
wire n_1709;
wire n_1610;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_455;
wire n_1701;
wire n_1243;
wire n_1121;
wire n_693;
wire n_606;
wire n_737;
wire n_1571;
wire n_1980;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_1543;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_1441;
wire n_1924;
wire n_1921;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_981;
wire n_1591;
wire n_583;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_974;
wire n_1036;
wire n_1831;
wire n_608;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1733;
wire n_1634;
wire n_1932;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1421;
wire n_1203;
wire n_561;
wire n_471;
wire n_846;
wire n_1793;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_1032;
wire n_936;
wire n_469;
wire n_1884;
wire n_1825;
wire n_1589;
wire n_1210;
wire n_591;
wire n_1933;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_623;
wire n_585;
wire n_1982;
wire n_1334;
wire n_1963;
wire n_483;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1977;
wire n_1200;
wire n_1120;
wire n_576;
wire n_1602;
wire n_1776;
wire n_1852;
wire n_1522;
wire n_1279;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1935;
wire n_1146;
wire n_488;
wire n_705;
wire n_1548;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_472;
wire n_1704;
wire n_847;
wire n_1436;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_1545;
wire n_456;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_814;
wire n_1864;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_1470;
wire n_444;
wire n_1761;
wire n_1836;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1875;
wire n_1615;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_650;
wire n_1575;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_951;
wire n_468;
wire n_1580;
wire n_1574;
wire n_780;
wire n_502;
wire n_1705;
wire n_633;
wire n_1746;
wire n_726;
wire n_532;
wire n_1439;
wire n_863;
wire n_597;
wire n_1832;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_1785;
wire n_486;
wire n_1870;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1967;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_1925;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_890;
wire n_628;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_1972;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1941;
wire n_1679;
wire n_1497;
wire n_2002;
wire n_1578;
wire n_1143;
wire n_1783;
wire n_510;
wire n_972;
wire n_1815;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_2000;
wire n_1857;
wire n_1920;
wire n_545;
wire n_887;
wire n_1162;
wire n_1997;
wire n_1894;
wire n_961;
wire n_991;
wire n_634;
wire n_1349;
wire n_1331;
wire n_1223;
wire n_1323;
wire n_578;
wire n_1739;
wire n_1777;
wire n_1353;
wire n_1429;
wire n_1546;
wire n_1432;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1874;
wire n_1834;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_1830;
wire n_1629;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_1340;
wire n_1626;
wire n_674;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_1612;
wire n_703;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_1517;
wire n_690;
wire n_1225;
wire n_1962;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_604;
wire n_1598;
wire n_977;
wire n_1895;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_1625;
wire n_933;
wire n_1774;
wire n_1797;
wire n_1037;
wire n_1899;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_742;
wire n_1191;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_636;
wire n_1259;
wire n_490;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_1538;
wire n_487;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_1889;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_922;
wire n_1790;
wire n_993;
wire n_851;
wire n_1725;
wire n_1135;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_1066;
wire n_648;
wire n_571;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_826;
wire n_1976;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_839;
wire n_768;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_722;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_804;
wire n_1455;
wire n_484;
wire n_1642;
wire n_1871;
wire n_480;
wire n_1057;
wire n_1473;
wire n_516;
wire n_1403;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_950;
wire n_512;
wire n_685;
wire n_1222;
wire n_1630;
wire n_1879;
wire n_1959;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_1779;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_1956;
wire n_681;
wire n_1718;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_1788;
wire n_786;
wire n_505;
wire n_1621;
wire n_1919;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_1893;
wire n_1570;
wire n_701;
wire n_995;
wire n_1000;
wire n_1931;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_812;
wire n_1961;
wire n_1050;
wire n_599;
wire n_1769;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_1632;
wire n_688;
wire n_1547;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1542;
wire n_1097;
wire n_1909;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_1872;
wire n_1940;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_1978;
wire n_1767;
wire n_1939;
wire n_1768;
wire n_1443;
wire n_478;
wire n_1585;
wire n_1861;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1584;
wire n_1481;
wire n_1928;
wire n_828;
wire n_1438;
wire n_1973;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_1693;
wire n_698;
wire n_1892;
wire n_1061;
wire n_682;
wire n_1373;
wire n_1686;
wire n_1302;
wire n_886;
wire n_1010;
wire n_883;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_854;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_914;
wire n_1986;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_1720;
wire n_880;
wire n_654;
wire n_1911;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1397;
wire n_1211;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1866;
wire n_1220;
wire n_467;
wire n_1398;
wire n_1262;
wire n_1904;
wire n_442;
wire n_1692;
wire n_1012;
wire n_1805;
wire n_960;
wire n_689;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1385;
wire n_1142;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_1868;
wire n_966;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_477;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_918;
wire n_1913;
wire n_672;
wire n_1039;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_566;
wire n_581;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_548;
wire n_1158;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_1404;
wire n_546;
wire n_788;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_888;
wire n_1325;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_955;
wire n_1333;
wire n_1916;
wire n_952;
wire n_1675;
wire n_1947;
wire n_1640;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1732;
wire n_1354;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_1934;
wire n_1900;
wire n_519;
wire n_1843;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_1902;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;

INVx1_ASAP7_75t_L g441 ( 
.A(n_89),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_387),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_115),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_91),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_124),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_339),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_208),
.Y(n_447)
);

CKINVDCx14_ASAP7_75t_R g448 ( 
.A(n_351),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_286),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_170),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_67),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_402),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_189),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_411),
.Y(n_454)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_51),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_231),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_398),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_33),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_108),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_1),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_366),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_381),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_373),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_12),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_316),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_257),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_317),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_261),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_143),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_307),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_169),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_424),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_146),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_256),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_87),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_377),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_102),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_33),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_235),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_99),
.Y(n_480)
);

CKINVDCx14_ASAP7_75t_R g481 ( 
.A(n_407),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_163),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_439),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_62),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_414),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_340),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_30),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_406),
.Y(n_488)
);

BUFx5_ASAP7_75t_L g489 ( 
.A(n_412),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_277),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_268),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_319),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_308),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_142),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_210),
.Y(n_495)
);

INVx1_ASAP7_75t_SL g496 ( 
.A(n_65),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_278),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_222),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_353),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_282),
.Y(n_500)
);

INVx2_ASAP7_75t_SL g501 ( 
.A(n_4),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_259),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_253),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_132),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_203),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_69),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_75),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_88),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_386),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_72),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_15),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_161),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_101),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_117),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_225),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_295),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_63),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_389),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_410),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_280),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_226),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_153),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_378),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_73),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_315),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_399),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_273),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_144),
.Y(n_528)
);

CKINVDCx16_ASAP7_75t_R g529 ( 
.A(n_195),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_26),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_112),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_155),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_28),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_194),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_285),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_220),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_165),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_248),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_270),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_11),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_27),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_374),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_97),
.Y(n_543)
);

BUFx10_ASAP7_75t_L g544 ( 
.A(n_385),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_364),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_209),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_156),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_131),
.Y(n_548)
);

INVxp67_ASAP7_75t_SL g549 ( 
.A(n_427),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_417),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_48),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_350),
.Y(n_552)
);

INVx1_ASAP7_75t_SL g553 ( 
.A(n_59),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_236),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_311),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_352),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_38),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_292),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_400),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_420),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_423),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_116),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_13),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_395),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_1),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_43),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_376),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_260),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_48),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_393),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_81),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_233),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_279),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_118),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_11),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_181),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_30),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_314),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_435),
.Y(n_579)
);

CKINVDCx16_ASAP7_75t_R g580 ( 
.A(n_196),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_240),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_358),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_135),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_408),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_75),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_425),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_28),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_43),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_405),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_148),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_383),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_382),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_52),
.Y(n_593)
);

INVxp67_ASAP7_75t_SL g594 ( 
.A(n_432),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_375),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_172),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_45),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_102),
.Y(n_598)
);

CKINVDCx16_ASAP7_75t_R g599 ( 
.A(n_5),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_368),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_87),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_66),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_324),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_205),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_422),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_372),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_16),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_394),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_68),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_42),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_437),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_388),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_404),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_430),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_365),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_80),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_188),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_313),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_409),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_362),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_349),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_171),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_401),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_283),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_294),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_298),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_321),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_440),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_413),
.Y(n_629)
);

CKINVDCx16_ASAP7_75t_R g630 ( 
.A(n_238),
.Y(n_630)
);

BUFx10_ASAP7_75t_L g631 ( 
.A(n_200),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_379),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_241),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_162),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_137),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_151),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_182),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_396),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_355),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_149),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_176),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_22),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_103),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_334),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_112),
.Y(n_645)
);

BUFx2_ASAP7_75t_L g646 ( 
.A(n_369),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_341),
.Y(n_647)
);

BUFx10_ASAP7_75t_L g648 ( 
.A(n_27),
.Y(n_648)
);

INVx1_ASAP7_75t_SL g649 ( 
.A(n_35),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_23),
.Y(n_650)
);

BUFx2_ASAP7_75t_L g651 ( 
.A(n_73),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_55),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_419),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_403),
.Y(n_654)
);

CKINVDCx11_ASAP7_75t_R g655 ( 
.A(n_12),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_213),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_245),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_60),
.Y(n_658)
);

BUFx10_ASAP7_75t_L g659 ( 
.A(n_290),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_343),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_113),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_18),
.Y(n_662)
);

BUFx10_ASAP7_75t_L g663 ( 
.A(n_348),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_363),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_66),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_59),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_223),
.Y(n_667)
);

CKINVDCx20_ASAP7_75t_R g668 ( 
.A(n_384),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_434),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_354),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_202),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_31),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_342),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_118),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_25),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_416),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_415),
.Y(n_677)
);

BUFx10_ASAP7_75t_L g678 ( 
.A(n_360),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_359),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_109),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_310),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_126),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_21),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_335),
.Y(n_684)
);

INVx1_ASAP7_75t_SL g685 ( 
.A(n_92),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_121),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_199),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_356),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_214),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g690 ( 
.A(n_347),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_421),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_85),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_54),
.Y(n_693)
);

CKINVDCx20_ASAP7_75t_R g694 ( 
.A(n_436),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_370),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_119),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_429),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_84),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_104),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_428),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_179),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_186),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_367),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_216),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_41),
.Y(n_705)
);

CKINVDCx14_ASAP7_75t_R g706 ( 
.A(n_139),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_31),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_397),
.Y(n_708)
);

CKINVDCx14_ASAP7_75t_R g709 ( 
.A(n_107),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_361),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_380),
.Y(n_711)
);

CKINVDCx20_ASAP7_75t_R g712 ( 
.A(n_76),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_40),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_390),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_392),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_56),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_154),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_371),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_57),
.Y(n_719)
);

CKINVDCx14_ASAP7_75t_R g720 ( 
.A(n_24),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_391),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_433),
.Y(n_722)
);

INVx1_ASAP7_75t_SL g723 ( 
.A(n_300),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_84),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_357),
.Y(n_725)
);

CKINVDCx20_ASAP7_75t_R g726 ( 
.A(n_288),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_60),
.Y(n_727)
);

BUFx8_ASAP7_75t_SL g728 ( 
.A(n_431),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_418),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_9),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_42),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_47),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_333),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_72),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_53),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_323),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_168),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_426),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_728),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_442),
.Y(n_740)
);

INVxp67_ASAP7_75t_SL g741 ( 
.A(n_517),
.Y(n_741)
);

INVxp67_ASAP7_75t_SL g742 ( 
.A(n_517),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_447),
.Y(n_743)
);

CKINVDCx20_ASAP7_75t_R g744 ( 
.A(n_709),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_709),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_608),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_646),
.Y(n_747)
);

INVxp67_ASAP7_75t_SL g748 ( 
.A(n_610),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_452),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_720),
.Y(n_750)
);

CKINVDCx20_ASAP7_75t_R g751 ( 
.A(n_720),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_610),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_457),
.Y(n_753)
);

HB1xp67_ASAP7_75t_L g754 ( 
.A(n_651),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_492),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_692),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_692),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_480),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_503),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_480),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_455),
.Y(n_761)
);

INVxp33_ASAP7_75t_L g762 ( 
.A(n_655),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_686),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_686),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_501),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_645),
.Y(n_766)
);

CKINVDCx14_ASAP7_75t_R g767 ( 
.A(n_448),
.Y(n_767)
);

INVxp67_ASAP7_75t_L g768 ( 
.A(n_441),
.Y(n_768)
);

CKINVDCx16_ASAP7_75t_R g769 ( 
.A(n_599),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_444),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_451),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_458),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_460),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_506),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_508),
.Y(n_775)
);

CKINVDCx16_ASAP7_75t_R g776 ( 
.A(n_529),
.Y(n_776)
);

CKINVDCx16_ASAP7_75t_R g777 ( 
.A(n_580),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_510),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_533),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_509),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_515),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_556),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_551),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_586),
.Y(n_784)
);

INVxp67_ASAP7_75t_SL g785 ( 
.A(n_565),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_489),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_566),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_595),
.Y(n_788)
);

CKINVDCx20_ASAP7_75t_R g789 ( 
.A(n_477),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_575),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_600),
.Y(n_791)
);

CKINVDCx16_ASAP7_75t_R g792 ( 
.A(n_630),
.Y(n_792)
);

BUFx6f_ASAP7_75t_L g793 ( 
.A(n_482),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_443),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_611),
.Y(n_795)
);

HB1xp67_ASAP7_75t_L g796 ( 
.A(n_459),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_577),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_587),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_601),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_653),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_602),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_657),
.Y(n_802)
);

INVxp67_ASAP7_75t_SL g803 ( 
.A(n_607),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_668),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_643),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_489),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_696),
.Y(n_807)
);

INVxp67_ASAP7_75t_L g808 ( 
.A(n_707),
.Y(n_808)
);

INVxp33_ASAP7_75t_SL g809 ( 
.A(n_464),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_730),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_731),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_734),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_544),
.Y(n_813)
);

INVxp67_ASAP7_75t_L g814 ( 
.A(n_648),
.Y(n_814)
);

HB1xp67_ASAP7_75t_L g815 ( 
.A(n_475),
.Y(n_815)
);

INVxp33_ASAP7_75t_SL g816 ( 
.A(n_478),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_544),
.Y(n_817)
);

CKINVDCx20_ASAP7_75t_R g818 ( 
.A(n_530),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_489),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_631),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_631),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_671),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_659),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_659),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_676),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_663),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_663),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_678),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_678),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_453),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_690),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_694),
.Y(n_832)
);

CKINVDCx20_ASAP7_75t_R g833 ( 
.A(n_574),
.Y(n_833)
);

INVxp67_ASAP7_75t_L g834 ( 
.A(n_648),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_726),
.Y(n_835)
);

INVxp33_ASAP7_75t_L g836 ( 
.A(n_650),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_465),
.Y(n_837)
);

CKINVDCx16_ASAP7_75t_R g838 ( 
.A(n_609),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_466),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_472),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_479),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_484),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_786),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_744),
.A2(n_750),
.B1(n_751),
.B2(n_745),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_765),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_749),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_753),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_766),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_793),
.Y(n_849)
);

INVx3_ASAP7_75t_L g850 ( 
.A(n_786),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_740),
.B(n_650),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_813),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_793),
.Y(n_853)
);

INVx3_ASAP7_75t_L g854 ( 
.A(n_806),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_752),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_806),
.Y(n_856)
);

BUFx2_ASAP7_75t_L g857 ( 
.A(n_767),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_756),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_757),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_819),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_743),
.B(n_700),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_819),
.Y(n_862)
);

BUFx12f_ASAP7_75t_L g863 ( 
.A(n_739),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_758),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_741),
.Y(n_865)
);

OA21x2_ASAP7_75t_L g866 ( 
.A1(n_830),
.A2(n_500),
.B(n_499),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_742),
.B(n_721),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_794),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_796),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_R g870 ( 
.A(n_767),
.B(n_448),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_748),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_793),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_760),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_755),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_759),
.Y(n_875)
);

BUFx8_ASAP7_75t_L g876 ( 
.A(n_762),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_770),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_771),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_772),
.Y(n_879)
);

AND2x6_ASAP7_75t_L g880 ( 
.A(n_837),
.B(n_476),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_817),
.Y(n_881)
);

NAND2xp33_ASAP7_75t_SL g882 ( 
.A(n_762),
.B(n_487),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_773),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_774),
.Y(n_884)
);

HB1xp67_ASAP7_75t_SL g885 ( 
.A(n_780),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_793),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_775),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_763),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_764),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_746),
.B(n_481),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_820),
.B(n_445),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_778),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_839),
.B(n_499),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_779),
.Y(n_894)
);

NOR2x1_ASAP7_75t_L g895 ( 
.A(n_821),
.B(n_476),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_754),
.B(n_481),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_783),
.Y(n_897)
);

AND2x2_ASAP7_75t_SL g898 ( 
.A(n_776),
.B(n_650),
.Y(n_898)
);

OAI22xp5_ASAP7_75t_SL g899 ( 
.A1(n_789),
.A2(n_724),
.B1(n_732),
.B2(n_712),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_787),
.Y(n_900)
);

OR2x6_ASAP7_75t_L g901 ( 
.A(n_814),
.B(n_650),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_790),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_797),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_798),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_799),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_777),
.B(n_706),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_823),
.B(n_446),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_840),
.B(n_500),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_815),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_SL g910 ( 
.A1(n_789),
.A2(n_507),
.B1(n_513),
.B2(n_511),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_801),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_805),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_841),
.B(n_537),
.Y(n_913)
);

CKINVDCx6p67_ASAP7_75t_R g914 ( 
.A(n_792),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_842),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_807),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_810),
.Y(n_917)
);

CKINVDCx20_ASAP7_75t_R g918 ( 
.A(n_818),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_781),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_811),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_812),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_768),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_769),
.B(n_706),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_824),
.B(n_449),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_782),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_808),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_785),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_747),
.B(n_514),
.Y(n_928)
);

INVxp67_ASAP7_75t_L g929 ( 
.A(n_834),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_803),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_836),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_826),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_827),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_828),
.B(n_483),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_784),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_829),
.B(n_537),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_788),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_836),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_744),
.Y(n_939)
);

NOR2x1_ASAP7_75t_L g940 ( 
.A(n_745),
.B(n_573),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_809),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_816),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_750),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_791),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_751),
.B(n_524),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_795),
.Y(n_946)
);

AND2x2_ASAP7_75t_SL g947 ( 
.A(n_838),
.B(n_490),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_800),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_761),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_802),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_761),
.B(n_573),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_804),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_822),
.Y(n_953)
);

BUFx2_ASAP7_75t_L g954 ( 
.A(n_818),
.Y(n_954)
);

INVx4_ASAP7_75t_L g955 ( 
.A(n_825),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_831),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_832),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_835),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_833),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_833),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_794),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_765),
.Y(n_962)
);

INVx3_ASAP7_75t_L g963 ( 
.A(n_765),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_749),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_754),
.B(n_531),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_793),
.Y(n_966)
);

AOI22xp5_ASAP7_75t_SL g967 ( 
.A1(n_789),
.A2(n_540),
.B1(n_543),
.B2(n_541),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_765),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_754),
.B(n_557),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_741),
.B(n_545),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_749),
.Y(n_971)
);

BUFx3_ASAP7_75t_L g972 ( 
.A(n_765),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_793),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_741),
.B(n_545),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_765),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_765),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_765),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_786),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_786),
.Y(n_979)
);

INVx4_ASAP7_75t_L g980 ( 
.A(n_786),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_765),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_765),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_765),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_749),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_765),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_741),
.B(n_589),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_765),
.Y(n_987)
);

CKINVDCx20_ASAP7_75t_R g988 ( 
.A(n_789),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_765),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_765),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_813),
.B(n_450),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_793),
.Y(n_992)
);

INVx3_ASAP7_75t_L g993 ( 
.A(n_765),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_749),
.Y(n_994)
);

NOR2xp67_ASAP7_75t_L g995 ( 
.A(n_752),
.B(n_738),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_786),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_765),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_754),
.B(n_562),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_765),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_754),
.B(n_563),
.Y(n_1000)
);

AND2x4_ASAP7_75t_L g1001 ( 
.A(n_740),
.B(n_620),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_741),
.B(n_589),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_765),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_765),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_740),
.B(n_620),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_741),
.B(n_606),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_765),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_786),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_922),
.B(n_454),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_926),
.B(n_456),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_889),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_866),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_889),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_921),
.B(n_461),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_932),
.B(n_462),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_889),
.Y(n_1016)
);

AND2x2_ASAP7_75t_SL g1017 ( 
.A(n_947),
.B(n_498),
.Y(n_1017)
);

INVxp67_ASAP7_75t_L g1018 ( 
.A(n_868),
.Y(n_1018)
);

NAND2xp33_ASAP7_75t_L g1019 ( 
.A(n_880),
.B(n_489),
.Y(n_1019)
);

NAND3xp33_ASAP7_75t_L g1020 ( 
.A(n_896),
.B(n_571),
.C(n_569),
.Y(n_1020)
);

INVx4_ASAP7_75t_L g1021 ( 
.A(n_901),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_900),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_866),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_900),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_931),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_932),
.B(n_463),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_921),
.B(n_467),
.Y(n_1027)
);

OAI21xp33_ASAP7_75t_SL g1028 ( 
.A1(n_867),
.A2(n_519),
.B(n_504),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_938),
.Y(n_1029)
);

OR2x2_ASAP7_75t_L g1030 ( 
.A(n_909),
.B(n_496),
.Y(n_1030)
);

BUFx2_ASAP7_75t_L g1031 ( 
.A(n_915),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_900),
.Y(n_1032)
);

INVxp33_ASAP7_75t_SL g1033 ( 
.A(n_870),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_845),
.Y(n_1034)
);

NAND3xp33_ASAP7_75t_L g1035 ( 
.A(n_928),
.B(n_588),
.C(n_585),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_917),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_845),
.Y(n_1037)
);

BUFx2_ASAP7_75t_L g1038 ( 
.A(n_961),
.Y(n_1038)
);

OR2x6_ASAP7_75t_L g1039 ( 
.A(n_863),
.B(n_522),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_963),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_963),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_975),
.Y(n_1042)
);

INVx1_ASAP7_75t_SL g1043 ( 
.A(n_941),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_930),
.B(n_468),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_965),
.B(n_553),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_917),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_917),
.Y(n_1047)
);

AND3x2_ASAP7_75t_L g1048 ( 
.A(n_954),
.B(n_594),
.C(n_549),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_890),
.B(n_623),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_865),
.B(n_469),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_920),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_940),
.A2(n_597),
.B1(n_598),
.B2(n_593),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_975),
.Y(n_1053)
);

BUFx2_ASAP7_75t_L g1054 ( 
.A(n_876),
.Y(n_1054)
);

OR2x6_ASAP7_75t_L g1055 ( 
.A(n_955),
.B(n_535),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_920),
.Y(n_1056)
);

BUFx2_ASAP7_75t_L g1057 ( 
.A(n_876),
.Y(n_1057)
);

AOI22xp33_ASAP7_75t_L g1058 ( 
.A1(n_871),
.A2(n_536),
.B1(n_542),
.B2(n_539),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_920),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_981),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_929),
.B(n_702),
.Y(n_1061)
);

INVx2_ASAP7_75t_SL g1062 ( 
.A(n_901),
.Y(n_1062)
);

INVx8_ASAP7_75t_L g1063 ( 
.A(n_901),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_927),
.A2(n_642),
.B1(n_652),
.B2(n_616),
.Y(n_1064)
);

INVx3_ASAP7_75t_L g1065 ( 
.A(n_981),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_864),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_989),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_932),
.B(n_470),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_877),
.B(n_471),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_989),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_933),
.B(n_473),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_855),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_891),
.B(n_723),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_873),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_888),
.Y(n_1075)
);

AOI22x1_ASAP7_75t_L g1076 ( 
.A1(n_993),
.A2(n_621),
.B1(n_637),
.B2(n_606),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_869),
.B(n_474),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_907),
.B(n_485),
.Y(n_1078)
);

BUFx10_ASAP7_75t_L g1079 ( 
.A(n_898),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_993),
.Y(n_1080)
);

NAND3xp33_ASAP7_75t_L g1081 ( 
.A(n_940),
.B(n_661),
.C(n_658),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_850),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_852),
.B(n_881),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_924),
.B(n_486),
.Y(n_1084)
);

INVx3_ASAP7_75t_L g1085 ( 
.A(n_851),
.Y(n_1085)
);

INVx1_ASAP7_75t_SL g1086 ( 
.A(n_969),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_851),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_848),
.Y(n_1088)
);

INVx2_ASAP7_75t_SL g1089 ( 
.A(n_998),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_878),
.B(n_879),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_962),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_968),
.Y(n_1092)
);

AO22x2_ASAP7_75t_L g1093 ( 
.A1(n_844),
.A2(n_685),
.B1(n_649),
.B2(n_550),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_850),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_1000),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_976),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_880),
.Y(n_1097)
);

INVx6_ASAP7_75t_L g1098 ( 
.A(n_955),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_854),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_977),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_854),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_1001),
.B(n_488),
.Y(n_1102)
);

OAI22xp33_ASAP7_75t_L g1103 ( 
.A1(n_914),
.A2(n_665),
.B1(n_666),
.B2(n_662),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_858),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_972),
.Y(n_1105)
);

INVx4_ASAP7_75t_L g1106 ( 
.A(n_880),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_883),
.B(n_491),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_884),
.B(n_493),
.Y(n_1108)
);

BUFx3_ASAP7_75t_L g1109 ( 
.A(n_857),
.Y(n_1109)
);

INVx2_ASAP7_75t_SL g1110 ( 
.A(n_923),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_880),
.Y(n_1111)
);

INVx2_ASAP7_75t_SL g1112 ( 
.A(n_906),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_856),
.Y(n_1113)
);

INVxp33_ASAP7_75t_SL g1114 ( 
.A(n_846),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_982),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_856),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_951),
.B(n_672),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_859),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_1001),
.B(n_494),
.Y(n_1119)
);

OAI22xp33_ASAP7_75t_L g1120 ( 
.A1(n_942),
.A2(n_675),
.B1(n_680),
.B2(n_674),
.Y(n_1120)
);

AOI21x1_ASAP7_75t_L g1121 ( 
.A1(n_843),
.A2(n_554),
.B(n_548),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_860),
.Y(n_1122)
);

OAI22xp33_ASAP7_75t_L g1123 ( 
.A1(n_948),
.A2(n_693),
.B1(n_698),
.B2(n_683),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_1005),
.B(n_497),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_980),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_862),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_978),
.Y(n_1127)
);

NAND2xp33_ASAP7_75t_L g1128 ( 
.A(n_887),
.B(n_892),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_980),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_894),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_916),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_L g1132 ( 
.A1(n_897),
.A2(n_568),
.B1(n_578),
.B2(n_559),
.Y(n_1132)
);

AOI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_1005),
.A2(n_705),
.B1(n_713),
.B2(n_699),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_983),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_985),
.Y(n_1135)
);

INVx3_ASAP7_75t_L g1136 ( 
.A(n_987),
.Y(n_1136)
);

INVx2_ASAP7_75t_SL g1137 ( 
.A(n_895),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_990),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_979),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_997),
.Y(n_1140)
);

AND3x2_ASAP7_75t_L g1141 ( 
.A(n_949),
.B(n_583),
.C(n_579),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_991),
.B(n_502),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_999),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1003),
.Y(n_1144)
);

BUFx3_ASAP7_75t_L g1145 ( 
.A(n_950),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_995),
.B(n_505),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_861),
.B(n_512),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_996),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1008),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_1004),
.B(n_716),
.Y(n_1150)
);

BUFx4f_ASAP7_75t_L g1151 ( 
.A(n_950),
.Y(n_1151)
);

AOI22xp33_ASAP7_75t_L g1152 ( 
.A1(n_902),
.A2(n_903),
.B1(n_905),
.B2(n_904),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1007),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_911),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_849),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_867),
.B(n_516),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_936),
.B(n_518),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_912),
.Y(n_1158)
);

BUFx10_ASAP7_75t_L g1159 ( 
.A(n_951),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_849),
.Y(n_1160)
);

INVx8_ASAP7_75t_L g1161 ( 
.A(n_950),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_970),
.Y(n_1162)
);

BUFx3_ASAP7_75t_L g1163 ( 
.A(n_958),
.Y(n_1163)
);

AND2x6_ASAP7_75t_L g1164 ( 
.A(n_895),
.B(n_654),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_970),
.Y(n_1165)
);

BUFx3_ASAP7_75t_L g1166 ( 
.A(n_958),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_893),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_936),
.B(n_520),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_893),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_974),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_967),
.B(n_719),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_974),
.B(n_986),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_995),
.B(n_521),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_986),
.Y(n_1174)
);

OAI22x1_ASAP7_75t_L g1175 ( 
.A1(n_960),
.A2(n_735),
.B1(n_727),
.B2(n_592),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1002),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_967),
.B(n_654),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_908),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_934),
.B(n_1006),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1002),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_908),
.Y(n_1181)
);

AND2x2_ASAP7_75t_SL g1182 ( 
.A(n_945),
.B(n_584),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_913),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1006),
.B(n_523),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_953),
.A2(n_737),
.B1(n_617),
.B2(n_618),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_913),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_956),
.A2(n_667),
.B1(n_670),
.B2(n_603),
.Y(n_1187)
);

INVxp67_ASAP7_75t_SL g1188 ( 
.A(n_952),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_882),
.B(n_525),
.Y(n_1189)
);

INVxp67_ASAP7_75t_SL g1190 ( 
.A(n_952),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_946),
.B(n_679),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_849),
.Y(n_1192)
);

INVx4_ASAP7_75t_L g1193 ( 
.A(n_958),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_957),
.Y(n_1194)
);

BUFx10_ASAP7_75t_L g1195 ( 
.A(n_847),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_939),
.B(n_526),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_853),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_910),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_853),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_853),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_910),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_SL g1202 ( 
.A(n_874),
.B(n_527),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_872),
.Y(n_1203)
);

INVxp67_ASAP7_75t_L g1204 ( 
.A(n_885),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_872),
.Y(n_1205)
);

INVxp33_ASAP7_75t_SL g1206 ( 
.A(n_875),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_872),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_886),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_886),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_886),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_966),
.Y(n_1211)
);

AND2x4_ASAP7_75t_L g1212 ( 
.A(n_943),
.B(n_679),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_966),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_966),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_973),
.Y(n_1215)
);

NOR3xp33_ASAP7_75t_L g1216 ( 
.A(n_844),
.B(n_684),
.C(n_681),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_919),
.B(n_528),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_973),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_973),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_L g1220 ( 
.A(n_992),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_992),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_SL g1222 ( 
.A(n_959),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_992),
.Y(n_1223)
);

BUFx2_ASAP7_75t_L g1224 ( 
.A(n_925),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_935),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_937),
.B(n_532),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_959),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_959),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_944),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_964),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_971),
.B(n_534),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_984),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_994),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_899),
.Y(n_1234)
);

INVx2_ASAP7_75t_SL g1235 ( 
.A(n_918),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_899),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_SL g1237 ( 
.A(n_988),
.B(n_538),
.Y(n_1237)
);

INVx3_ASAP7_75t_L g1238 ( 
.A(n_889),
.Y(n_1238)
);

BUFx10_ASAP7_75t_L g1239 ( 
.A(n_898),
.Y(n_1239)
);

INVx4_ASAP7_75t_L g1240 ( 
.A(n_901),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_SL g1241 ( 
.A(n_932),
.B(n_546),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1018),
.B(n_547),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1162),
.B(n_552),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1125),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1162),
.Y(n_1245)
);

NAND2x1_ASAP7_75t_L g1246 ( 
.A(n_1021),
.B(n_1240),
.Y(n_1246)
);

OAI221xp5_ASAP7_75t_L g1247 ( 
.A1(n_1086),
.A2(n_691),
.B1(n_701),
.B2(n_688),
.C(n_687),
.Y(n_1247)
);

OR2x6_ASAP7_75t_L g1248 ( 
.A(n_1054),
.B(n_703),
.Y(n_1248)
);

NOR2xp67_ASAP7_75t_L g1249 ( 
.A(n_1204),
.B(n_0),
.Y(n_1249)
);

INVxp67_ASAP7_75t_L g1250 ( 
.A(n_1031),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1165),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_SL g1252 ( 
.A1(n_1236),
.A2(n_558),
.B1(n_560),
.B2(n_555),
.Y(n_1252)
);

BUFx12f_ASAP7_75t_L g1253 ( 
.A(n_1057),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1165),
.Y(n_1254)
);

AOI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1017),
.A2(n_708),
.B1(n_710),
.B2(n_704),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1170),
.B(n_561),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1174),
.B(n_1176),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1167),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1188),
.B(n_715),
.Y(n_1259)
);

OR2x6_ASAP7_75t_L g1260 ( 
.A(n_1063),
.B(n_718),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_1125),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1169),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1125),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1129),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1198),
.A2(n_736),
.B1(n_722),
.B2(n_637),
.Y(n_1265)
);

OR2x2_ASAP7_75t_L g1266 ( 
.A(n_1038),
.B(n_0),
.Y(n_1266)
);

AOI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1216),
.A2(n_567),
.B1(n_570),
.B2(n_564),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1021),
.B(n_733),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1110),
.B(n_572),
.Y(n_1269)
);

AOI22x1_ASAP7_75t_L g1270 ( 
.A1(n_1012),
.A2(n_639),
.B1(n_640),
.B2(n_621),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1178),
.Y(n_1271)
);

INVxp33_ASAP7_75t_L g1272 ( 
.A(n_1030),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1181),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1180),
.B(n_576),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1043),
.B(n_2),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1171),
.B(n_2),
.Y(n_1276)
);

NAND2x1_ASAP7_75t_L g1277 ( 
.A(n_1240),
.B(n_639),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1172),
.B(n_581),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_SL g1279 ( 
.A(n_1062),
.B(n_582),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1112),
.B(n_590),
.Y(n_1280)
);

OR2x2_ASAP7_75t_L g1281 ( 
.A(n_1045),
.B(n_3),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1136),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1183),
.Y(n_1283)
);

INVx2_ASAP7_75t_SL g1284 ( 
.A(n_1063),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1136),
.Y(n_1285)
);

INVx4_ASAP7_75t_L g1286 ( 
.A(n_1098),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1186),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1034),
.B(n_591),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1072),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_SL g1290 ( 
.A(n_1106),
.B(n_729),
.Y(n_1290)
);

OAI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1236),
.A2(n_604),
.B1(n_605),
.B2(n_596),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_SL g1292 ( 
.A(n_1195),
.Y(n_1292)
);

AOI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1150),
.A2(n_613),
.B1(n_614),
.B2(n_612),
.Y(n_1293)
);

OAI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1201),
.A2(n_619),
.B1(n_622),
.B2(n_615),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_1089),
.B(n_624),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1034),
.B(n_625),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1095),
.B(n_627),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1065),
.B(n_628),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1065),
.B(n_629),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1156),
.B(n_632),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_1150),
.B(n_633),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1037),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1072),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1040),
.Y(n_1304)
);

BUFx6f_ASAP7_75t_SL g1305 ( 
.A(n_1195),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1090),
.B(n_634),
.Y(n_1306)
);

INVx2_ASAP7_75t_SL g1307 ( 
.A(n_1098),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1088),
.B(n_635),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1091),
.B(n_636),
.Y(n_1309)
);

AOI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1182),
.A2(n_641),
.B1(n_644),
.B2(n_638),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1104),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1092),
.B(n_647),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1096),
.B(n_656),
.Y(n_1313)
);

AND2x4_ASAP7_75t_L g1314 ( 
.A(n_1190),
.B(n_3),
.Y(n_1314)
);

NOR2xp67_ASAP7_75t_L g1315 ( 
.A(n_1106),
.B(n_122),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1100),
.B(n_660),
.Y(n_1316)
);

CKINVDCx14_ASAP7_75t_R g1317 ( 
.A(n_1224),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1194),
.A2(n_640),
.B1(n_489),
.B2(n_664),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_L g1319 ( 
.A(n_1020),
.B(n_669),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_L g1320 ( 
.A(n_1117),
.B(n_673),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1104),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1115),
.B(n_677),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_SL g1323 ( 
.A(n_1097),
.B(n_682),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_SL g1324 ( 
.A(n_1097),
.B(n_725),
.Y(n_1324)
);

INVxp67_ASAP7_75t_L g1325 ( 
.A(n_1109),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1134),
.B(n_689),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1093),
.B(n_1159),
.Y(n_1327)
);

NAND2xp33_ASAP7_75t_L g1328 ( 
.A(n_1097),
.B(n_489),
.Y(n_1328)
);

NOR2xp67_ASAP7_75t_L g1329 ( 
.A(n_1081),
.B(n_123),
.Y(n_1329)
);

O2A1O1Ixp33_ASAP7_75t_L g1330 ( 
.A1(n_1179),
.A2(n_6),
.B(n_4),
.C(n_5),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_SL g1331 ( 
.A(n_1111),
.B(n_717),
.Y(n_1331)
);

INVxp67_ASAP7_75t_L g1332 ( 
.A(n_1225),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1041),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1042),
.Y(n_1334)
);

BUFx3_ASAP7_75t_L g1335 ( 
.A(n_1161),
.Y(n_1335)
);

INVx8_ASAP7_75t_L g1336 ( 
.A(n_1161),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1105),
.B(n_6),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_SL g1338 ( 
.A(n_1111),
.B(n_714),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1118),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_SL g1340 ( 
.A(n_1111),
.B(n_697),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1118),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1053),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1135),
.B(n_1138),
.Y(n_1343)
);

NAND2xp33_ASAP7_75t_L g1344 ( 
.A(n_1012),
.B(n_711),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1140),
.B(n_7),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1143),
.B(n_7),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_SL g1347 ( 
.A(n_1105),
.B(n_482),
.Y(n_1347)
);

BUFx3_ASAP7_75t_L g1348 ( 
.A(n_1145),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1060),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_SL g1350 ( 
.A(n_1123),
.B(n_482),
.Y(n_1350)
);

NOR3xp33_ASAP7_75t_L g1351 ( 
.A(n_1103),
.B(n_8),
.C(n_9),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1144),
.B(n_8),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1153),
.B(n_10),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1067),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1154),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_SL g1356 ( 
.A(n_1184),
.B(n_482),
.Y(n_1356)
);

OAI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1152),
.A2(n_626),
.B1(n_695),
.B2(n_495),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1055),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1158),
.B(n_10),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1102),
.B(n_13),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1114),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1093),
.B(n_14),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1157),
.B(n_14),
.Y(n_1363)
);

NAND3xp33_ASAP7_75t_SL g1364 ( 
.A(n_1229),
.B(n_15),
.C(n_16),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1168),
.B(n_17),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1131),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1055),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1177),
.A2(n_626),
.B1(n_495),
.B2(n_695),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1085),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_SL g1370 ( 
.A(n_1028),
.B(n_495),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1070),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_SL g1372 ( 
.A(n_1014),
.B(n_495),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1025),
.B(n_17),
.Y(n_1373)
);

INVx3_ASAP7_75t_L g1374 ( 
.A(n_1131),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_SL g1375 ( 
.A(n_1027),
.B(n_626),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1085),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1087),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1029),
.Y(n_1378)
);

AND2x6_ASAP7_75t_L g1379 ( 
.A(n_1023),
.B(n_695),
.Y(n_1379)
);

INVx2_ASAP7_75t_SL g1380 ( 
.A(n_1159),
.Y(n_1380)
);

AOI22x1_ASAP7_75t_SL g1381 ( 
.A1(n_1206),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_1381)
);

NOR2xp33_ASAP7_75t_L g1382 ( 
.A(n_1119),
.B(n_19),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_SL g1383 ( 
.A(n_1151),
.B(n_626),
.Y(n_1383)
);

NOR2x1p5_ASAP7_75t_L g1384 ( 
.A(n_1234),
.B(n_695),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1083),
.B(n_20),
.Y(n_1385)
);

OAI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1023),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_1386)
);

INVxp67_ASAP7_75t_L g1387 ( 
.A(n_1225),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_SL g1388 ( 
.A(n_1033),
.B(n_24),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_1124),
.B(n_1133),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_SL g1390 ( 
.A(n_1151),
.B(n_25),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1049),
.B(n_26),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1128),
.B(n_29),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_SL g1393 ( 
.A(n_1069),
.B(n_29),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_1235),
.B(n_32),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_SL g1395 ( 
.A(n_1107),
.B(n_32),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1080),
.A2(n_127),
.B(n_125),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1130),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1052),
.B(n_1061),
.Y(n_1398)
);

AOI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1064),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1066),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1058),
.B(n_34),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1122),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1074),
.Y(n_1403)
);

AOI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1035),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_1404)
);

INVx2_ASAP7_75t_SL g1405 ( 
.A(n_1163),
.Y(n_1405)
);

AOI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1229),
.A2(n_40),
.B1(n_37),
.B2(n_39),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1075),
.B(n_39),
.Y(n_1407)
);

INVxp67_ASAP7_75t_SL g1408 ( 
.A(n_1225),
.Y(n_1408)
);

INVxp67_ASAP7_75t_L g1409 ( 
.A(n_1044),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1108),
.B(n_1050),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1120),
.B(n_41),
.Y(n_1411)
);

OAI221xp5_ASAP7_75t_L g1412 ( 
.A1(n_1132),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.C(n_47),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1082),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1094),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1122),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1079),
.B(n_44),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1126),
.Y(n_1417)
);

NAND2x1_ASAP7_75t_L g1418 ( 
.A(n_1238),
.B(n_1126),
.Y(n_1418)
);

NAND3xp33_ASAP7_75t_L g1419 ( 
.A(n_1231),
.B(n_46),
.C(n_49),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1099),
.Y(n_1420)
);

NAND2xp33_ASAP7_75t_L g1421 ( 
.A(n_1024),
.B(n_128),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1232),
.B(n_49),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1222),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1137),
.B(n_50),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1191),
.B(n_50),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1191),
.B(n_51),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1147),
.B(n_52),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1232),
.B(n_53),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1234),
.B(n_54),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1077),
.B(n_55),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1127),
.Y(n_1431)
);

BUFx6f_ASAP7_75t_L g1432 ( 
.A(n_1024),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_SL g1433 ( 
.A(n_1230),
.B(n_56),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1127),
.A2(n_61),
.B1(n_57),
.B2(n_58),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1233),
.A2(n_62),
.B1(n_58),
.B2(n_61),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1101),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1164),
.A2(n_1076),
.B1(n_1148),
.B2(n_1139),
.Y(n_1437)
);

BUFx6f_ASAP7_75t_L g1438 ( 
.A(n_1024),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_1432),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1272),
.B(n_1237),
.Y(n_1440)
);

INVx3_ASAP7_75t_L g1441 ( 
.A(n_1261),
.Y(n_1441)
);

AO22x1_ASAP7_75t_L g1442 ( 
.A1(n_1361),
.A2(n_1234),
.B1(n_1166),
.B2(n_1193),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1336),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1257),
.Y(n_1444)
);

NOR3xp33_ASAP7_75t_SL g1445 ( 
.A(n_1247),
.B(n_1189),
.C(n_1202),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1327),
.A2(n_1212),
.B1(n_1228),
.B2(n_1227),
.Y(n_1446)
);

AOI21xp33_ASAP7_75t_L g1447 ( 
.A1(n_1242),
.A2(n_1226),
.B(n_1217),
.Y(n_1447)
);

BUFx3_ASAP7_75t_L g1448 ( 
.A(n_1336),
.Y(n_1448)
);

BUFx2_ASAP7_75t_L g1449 ( 
.A(n_1250),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_SL g1450 ( 
.A(n_1325),
.B(n_1079),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_SL g1451 ( 
.A(n_1261),
.B(n_1239),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1258),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1262),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_SL g1454 ( 
.A(n_1292),
.B(n_1039),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1271),
.B(n_1141),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1273),
.B(n_1212),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1317),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1358),
.B(n_1239),
.Y(n_1458)
);

AND2x6_ASAP7_75t_SL g1459 ( 
.A(n_1248),
.B(n_1039),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1283),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1287),
.B(n_1073),
.Y(n_1461)
);

NAND2xp33_ASAP7_75t_SL g1462 ( 
.A(n_1292),
.B(n_1222),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1355),
.Y(n_1463)
);

AND2x4_ASAP7_75t_L g1464 ( 
.A(n_1378),
.B(n_1409),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1343),
.B(n_1185),
.Y(n_1465)
);

INVx2_ASAP7_75t_SL g1466 ( 
.A(n_1335),
.Y(n_1466)
);

AOI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1398),
.A2(n_1187),
.B1(n_1164),
.B2(n_1175),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1261),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1289),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1303),
.Y(n_1470)
);

BUFx6f_ASAP7_75t_L g1471 ( 
.A(n_1432),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1311),
.Y(n_1472)
);

BUFx2_ASAP7_75t_L g1473 ( 
.A(n_1253),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1321),
.B(n_1009),
.Y(n_1474)
);

INVx5_ASAP7_75t_L g1475 ( 
.A(n_1260),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1345),
.Y(n_1476)
);

NOR2x1_ASAP7_75t_L g1477 ( 
.A(n_1384),
.B(n_1019),
.Y(n_1477)
);

INVxp67_ASAP7_75t_SL g1478 ( 
.A(n_1337),
.Y(n_1478)
);

INVx3_ASAP7_75t_L g1479 ( 
.A(n_1246),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1346),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1352),
.Y(n_1481)
);

INVx4_ASAP7_75t_L g1482 ( 
.A(n_1305),
.Y(n_1482)
);

INVx4_ASAP7_75t_L g1483 ( 
.A(n_1305),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1339),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1276),
.A2(n_1389),
.B1(n_1314),
.B2(n_1385),
.Y(n_1485)
);

INVx4_ASAP7_75t_L g1486 ( 
.A(n_1260),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1341),
.B(n_1010),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1245),
.Y(n_1488)
);

AOI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1410),
.A2(n_1173),
.B(n_1146),
.Y(n_1489)
);

CKINVDCx16_ASAP7_75t_R g1490 ( 
.A(n_1248),
.Y(n_1490)
);

INVx2_ASAP7_75t_SL g1491 ( 
.A(n_1423),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1278),
.B(n_1193),
.Y(n_1492)
);

INVx3_ASAP7_75t_L g1493 ( 
.A(n_1402),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1255),
.B(n_1078),
.Y(n_1494)
);

INVx3_ASAP7_75t_L g1495 ( 
.A(n_1415),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1353),
.Y(n_1496)
);

CKINVDCx20_ASAP7_75t_R g1497 ( 
.A(n_1367),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1377),
.Y(n_1498)
);

AND3x1_ASAP7_75t_L g1499 ( 
.A(n_1388),
.B(n_1142),
.C(n_1084),
.Y(n_1499)
);

INVx1_ASAP7_75t_SL g1500 ( 
.A(n_1337),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1251),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1254),
.B(n_1048),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_L g1503 ( 
.A(n_1301),
.B(n_1320),
.Y(n_1503)
);

NAND3xp33_ASAP7_75t_SL g1504 ( 
.A(n_1351),
.B(n_1196),
.C(n_1026),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1397),
.Y(n_1505)
);

INVx2_ASAP7_75t_SL g1506 ( 
.A(n_1284),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_SL g1507 ( 
.A(n_1266),
.B(n_1380),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1400),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1281),
.B(n_1164),
.Y(n_1509)
);

AND2x2_ASAP7_75t_SL g1510 ( 
.A(n_1362),
.B(n_1113),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1259),
.B(n_1164),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1403),
.Y(n_1512)
);

INVxp67_ASAP7_75t_L g1513 ( 
.A(n_1314),
.Y(n_1513)
);

AND2x4_ASAP7_75t_L g1514 ( 
.A(n_1332),
.B(n_1015),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1373),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1428),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_SL g1517 ( 
.A(n_1286),
.B(n_1293),
.Y(n_1517)
);

INVx4_ASAP7_75t_L g1518 ( 
.A(n_1286),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1417),
.Y(n_1519)
);

BUFx6f_ASAP7_75t_L g1520 ( 
.A(n_1432),
.Y(n_1520)
);

OAI21xp33_ASAP7_75t_SL g1521 ( 
.A1(n_1437),
.A2(n_1241),
.B(n_1068),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1359),
.Y(n_1522)
);

AO21x1_ASAP7_75t_L g1523 ( 
.A1(n_1357),
.A2(n_1121),
.B(n_1032),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1385),
.A2(n_1411),
.B1(n_1259),
.B2(n_1401),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1306),
.B(n_1071),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1302),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1387),
.B(n_1269),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1304),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1280),
.B(n_1116),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1408),
.B(n_1238),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1275),
.B(n_1149),
.Y(n_1531)
);

AOI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1360),
.A2(n_1013),
.B1(n_1016),
.B2(n_1011),
.Y(n_1532)
);

NOR2xp67_ASAP7_75t_L g1533 ( 
.A(n_1419),
.B(n_129),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1295),
.B(n_1022),
.Y(n_1534)
);

INVxp67_ASAP7_75t_SL g1535 ( 
.A(n_1438),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1310),
.B(n_63),
.Y(n_1536)
);

CKINVDCx20_ASAP7_75t_R g1537 ( 
.A(n_1348),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1394),
.A2(n_1076),
.B1(n_1046),
.B2(n_1047),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1265),
.B(n_1431),
.Y(n_1539)
);

AOI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1412),
.A2(n_1051),
.B1(n_1056),
.B2(n_1036),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_SL g1541 ( 
.A(n_1294),
.B(n_1059),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1264),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1333),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1382),
.B(n_64),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1334),
.Y(n_1545)
);

BUFx6f_ASAP7_75t_L g1546 ( 
.A(n_1438),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1342),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_1381),
.Y(n_1548)
);

INVx5_ASAP7_75t_L g1549 ( 
.A(n_1379),
.Y(n_1549)
);

HB1xp67_ASAP7_75t_L g1550 ( 
.A(n_1405),
.Y(n_1550)
);

AOI22xp5_ASAP7_75t_SL g1551 ( 
.A1(n_1416),
.A2(n_67),
.B1(n_64),
.B2(n_65),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_SL g1552 ( 
.A(n_1291),
.B(n_1155),
.Y(n_1552)
);

INVx2_ASAP7_75t_SL g1553 ( 
.A(n_1307),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_1252),
.Y(n_1554)
);

BUFx3_ASAP7_75t_L g1555 ( 
.A(n_1277),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1297),
.B(n_68),
.Y(n_1556)
);

INVx1_ASAP7_75t_SL g1557 ( 
.A(n_1429),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1430),
.A2(n_1211),
.B1(n_1219),
.B2(n_1218),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1349),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1256),
.B(n_69),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1243),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1274),
.B(n_70),
.Y(n_1562)
);

INVx3_ASAP7_75t_L g1563 ( 
.A(n_1282),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1350),
.A2(n_1211),
.B1(n_1219),
.B2(n_1218),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_1399),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1425),
.B(n_70),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1267),
.B(n_71),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_SL g1568 ( 
.A(n_1438),
.B(n_1155),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1354),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_SL g1570 ( 
.A(n_1285),
.B(n_1155),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1426),
.B(n_71),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1391),
.B(n_74),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1371),
.Y(n_1573)
);

INVxp67_ASAP7_75t_L g1574 ( 
.A(n_1422),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1268),
.B(n_74),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1369),
.Y(n_1576)
);

BUFx2_ASAP7_75t_L g1577 ( 
.A(n_1244),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1370),
.A2(n_1221),
.B1(n_1207),
.B2(n_1209),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_SL g1579 ( 
.A(n_1249),
.B(n_1160),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1308),
.B(n_76),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1407),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_1263),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1309),
.B(n_77),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_1406),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1413),
.Y(n_1585)
);

NOR2x1_ASAP7_75t_R g1586 ( 
.A(n_1390),
.B(n_1160),
.Y(n_1586)
);

AND2x4_ASAP7_75t_SL g1587 ( 
.A(n_1366),
.B(n_1160),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_1565),
.B(n_1279),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_L g1589 ( 
.A(n_1584),
.B(n_1319),
.Y(n_1589)
);

AO21x1_ASAP7_75t_L g1590 ( 
.A1(n_1552),
.A2(n_1386),
.B(n_1330),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1444),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1503),
.B(n_1312),
.Y(n_1592)
);

A2O1A1Ixp33_ASAP7_75t_SL g1593 ( 
.A1(n_1527),
.A2(n_1368),
.B(n_1427),
.C(n_1365),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1524),
.B(n_1464),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1464),
.B(n_1313),
.Y(n_1595)
);

OAI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1485),
.A2(n_1392),
.B1(n_1363),
.B2(n_1270),
.Y(n_1596)
);

INVx3_ASAP7_75t_L g1597 ( 
.A(n_1518),
.Y(n_1597)
);

AOI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1490),
.A2(n_1433),
.B1(n_1393),
.B2(n_1395),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1465),
.B(n_1316),
.Y(n_1599)
);

OAI22x1_ASAP7_75t_L g1600 ( 
.A1(n_1475),
.A2(n_1404),
.B1(n_1364),
.B2(n_1424),
.Y(n_1600)
);

AOI21xp5_ASAP7_75t_L g1601 ( 
.A1(n_1521),
.A2(n_1356),
.B(n_1344),
.Y(n_1601)
);

INVx1_ASAP7_75t_SL g1602 ( 
.A(n_1537),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_L g1603 ( 
.A(n_1486),
.B(n_1322),
.Y(n_1603)
);

NOR2xp67_ASAP7_75t_L g1604 ( 
.A(n_1475),
.B(n_1434),
.Y(n_1604)
);

INVx1_ASAP7_75t_SL g1605 ( 
.A(n_1443),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1469),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1516),
.B(n_1326),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_SL g1608 ( 
.A(n_1475),
.B(n_1315),
.Y(n_1608)
);

INVxp67_ASAP7_75t_L g1609 ( 
.A(n_1449),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1470),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1472),
.Y(n_1611)
);

O2A1O1Ixp33_ASAP7_75t_L g1612 ( 
.A1(n_1494),
.A2(n_1435),
.B(n_1300),
.C(n_1288),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_SL g1613 ( 
.A(n_1486),
.B(n_1315),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_SL g1614 ( 
.A(n_1454),
.B(n_1329),
.Y(n_1614)
);

O2A1O1Ixp33_ASAP7_75t_L g1615 ( 
.A1(n_1447),
.A2(n_1298),
.B(n_1299),
.C(n_1296),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1457),
.B(n_1414),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1463),
.B(n_1376),
.Y(n_1617)
);

BUFx6f_ASAP7_75t_L g1618 ( 
.A(n_1439),
.Y(n_1618)
);

CKINVDCx8_ASAP7_75t_R g1619 ( 
.A(n_1459),
.Y(n_1619)
);

A2O1A1Ixp33_ASAP7_75t_L g1620 ( 
.A1(n_1521),
.A2(n_1329),
.B(n_1374),
.C(n_1366),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1498),
.B(n_1420),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1557),
.B(n_1374),
.Y(n_1622)
);

NOR2xp67_ASAP7_75t_L g1623 ( 
.A(n_1448),
.B(n_1323),
.Y(n_1623)
);

AOI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1581),
.A2(n_1375),
.B(n_1372),
.Y(n_1624)
);

BUFx3_ASAP7_75t_L g1625 ( 
.A(n_1473),
.Y(n_1625)
);

BUFx6f_ASAP7_75t_L g1626 ( 
.A(n_1439),
.Y(n_1626)
);

BUFx3_ASAP7_75t_L g1627 ( 
.A(n_1497),
.Y(n_1627)
);

CKINVDCx20_ASAP7_75t_R g1628 ( 
.A(n_1462),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1484),
.B(n_1318),
.Y(n_1629)
);

AOI21xp5_ASAP7_75t_L g1630 ( 
.A1(n_1522),
.A2(n_1328),
.B(n_1347),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1478),
.B(n_1436),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1452),
.Y(n_1632)
);

BUFx8_ASAP7_75t_L g1633 ( 
.A(n_1466),
.Y(n_1633)
);

BUFx2_ASAP7_75t_L g1634 ( 
.A(n_1491),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_SL g1635 ( 
.A(n_1510),
.B(n_1396),
.Y(n_1635)
);

AO21x1_ASAP7_75t_L g1636 ( 
.A1(n_1572),
.A2(n_1421),
.B(n_1383),
.Y(n_1636)
);

O2A1O1Ixp33_ASAP7_75t_L g1637 ( 
.A1(n_1544),
.A2(n_1290),
.B(n_1331),
.C(n_1324),
.Y(n_1637)
);

OAI21x1_ASAP7_75t_L g1638 ( 
.A1(n_1568),
.A2(n_1418),
.B(n_1221),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1499),
.B(n_1338),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1513),
.B(n_1440),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1460),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1561),
.B(n_1340),
.Y(n_1642)
);

NAND2xp33_ASAP7_75t_SL g1643 ( 
.A(n_1445),
.B(n_1379),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1507),
.B(n_77),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1505),
.Y(n_1645)
);

AOI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1476),
.A2(n_1214),
.B(n_1205),
.Y(n_1646)
);

OAI21x1_ASAP7_75t_L g1647 ( 
.A1(n_1523),
.A2(n_1570),
.B(n_1441),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1508),
.Y(n_1648)
);

O2A1O1Ixp33_ASAP7_75t_L g1649 ( 
.A1(n_1560),
.A2(n_1199),
.B(n_1200),
.C(n_1197),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1500),
.A2(n_1379),
.B1(n_1210),
.B2(n_1220),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1502),
.B(n_78),
.Y(n_1651)
);

NAND3xp33_ASAP7_75t_SL g1652 ( 
.A(n_1548),
.B(n_1208),
.C(n_1203),
.Y(n_1652)
);

BUFx5_ASAP7_75t_L g1653 ( 
.A(n_1526),
.Y(n_1653)
);

O2A1O1Ixp33_ASAP7_75t_L g1654 ( 
.A1(n_1562),
.A2(n_1215),
.B(n_1223),
.C(n_1213),
.Y(n_1654)
);

NAND2x1p5_ASAP7_75t_L g1655 ( 
.A(n_1482),
.B(n_1192),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1474),
.B(n_1379),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1512),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1453),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1480),
.A2(n_1210),
.B(n_1192),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1519),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1487),
.B(n_78),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1458),
.B(n_79),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1554),
.B(n_79),
.Y(n_1663)
);

AOI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1536),
.A2(n_1210),
.B1(n_1220),
.B2(n_1192),
.Y(n_1664)
);

AOI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1481),
.A2(n_1220),
.B(n_133),
.Y(n_1665)
);

AOI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1496),
.A2(n_134),
.B(n_130),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1493),
.Y(n_1667)
);

AOI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1515),
.A2(n_138),
.B(n_136),
.Y(n_1668)
);

AND2x4_ASAP7_75t_L g1669 ( 
.A(n_1528),
.B(n_80),
.Y(n_1669)
);

BUFx2_ASAP7_75t_L g1670 ( 
.A(n_1482),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1543),
.B(n_81),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_SL g1672 ( 
.A(n_1575),
.B(n_82),
.Y(n_1672)
);

O2A1O1Ixp33_ASAP7_75t_L g1673 ( 
.A1(n_1580),
.A2(n_85),
.B(n_82),
.C(n_83),
.Y(n_1673)
);

BUFx3_ASAP7_75t_L g1674 ( 
.A(n_1483),
.Y(n_1674)
);

INVx2_ASAP7_75t_SL g1675 ( 
.A(n_1483),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1585),
.Y(n_1676)
);

OAI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1467),
.A2(n_88),
.B1(n_83),
.B2(n_86),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1461),
.B(n_86),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1467),
.B(n_89),
.Y(n_1679)
);

INVx1_ASAP7_75t_SL g1680 ( 
.A(n_1605),
.Y(n_1680)
);

AO31x2_ASAP7_75t_L g1681 ( 
.A1(n_1620),
.A2(n_1566),
.A3(n_1571),
.B(n_1468),
.Y(n_1681)
);

AOI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1593),
.A2(n_1471),
.B(n_1439),
.Y(n_1682)
);

OAI22x1_ASAP7_75t_L g1683 ( 
.A1(n_1663),
.A2(n_1575),
.B1(n_1551),
.B2(n_1567),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1591),
.Y(n_1684)
);

BUFx10_ASAP7_75t_L g1685 ( 
.A(n_1669),
.Y(n_1685)
);

AOI21xp5_ASAP7_75t_L g1686 ( 
.A1(n_1601),
.A2(n_1520),
.B(n_1471),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_SL g1687 ( 
.A(n_1619),
.B(n_1518),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1606),
.Y(n_1688)
);

AOI21xp5_ASAP7_75t_L g1689 ( 
.A1(n_1596),
.A2(n_1520),
.B(n_1471),
.Y(n_1689)
);

AO21x2_ASAP7_75t_L g1690 ( 
.A1(n_1647),
.A2(n_1533),
.B(n_1579),
.Y(n_1690)
);

AOI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1635),
.A2(n_1546),
.B(n_1520),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1662),
.B(n_1545),
.Y(n_1692)
);

AOI21xp5_ASAP7_75t_L g1693 ( 
.A1(n_1659),
.A2(n_1546),
.B(n_1533),
.Y(n_1693)
);

AND2x4_ASAP7_75t_L g1694 ( 
.A(n_1597),
.B(n_1549),
.Y(n_1694)
);

OAI21x1_ASAP7_75t_L g1695 ( 
.A1(n_1650),
.A2(n_1441),
.B(n_1477),
.Y(n_1695)
);

OAI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1669),
.A2(n_1446),
.B1(n_1583),
.B2(n_1456),
.Y(n_1696)
);

AO21x2_ASAP7_75t_L g1697 ( 
.A1(n_1604),
.A2(n_1509),
.B(n_1504),
.Y(n_1697)
);

OAI21x1_ASAP7_75t_L g1698 ( 
.A1(n_1638),
.A2(n_1665),
.B(n_1636),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1632),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1592),
.B(n_1547),
.Y(n_1700)
);

INVx1_ASAP7_75t_SL g1701 ( 
.A(n_1602),
.Y(n_1701)
);

A2O1A1Ixp33_ASAP7_75t_L g1702 ( 
.A1(n_1612),
.A2(n_1529),
.B(n_1534),
.C(n_1574),
.Y(n_1702)
);

AND2x4_ASAP7_75t_L g1703 ( 
.A(n_1597),
.B(n_1549),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1653),
.Y(n_1704)
);

OAI21xp5_ASAP7_75t_L g1705 ( 
.A1(n_1615),
.A2(n_1489),
.B(n_1556),
.Y(n_1705)
);

BUFx6f_ASAP7_75t_L g1706 ( 
.A(n_1618),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1594),
.B(n_1559),
.Y(n_1707)
);

OAI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1672),
.A2(n_1455),
.B1(n_1539),
.B2(n_1538),
.Y(n_1708)
);

INVx1_ASAP7_75t_SL g1709 ( 
.A(n_1625),
.Y(n_1709)
);

INVx3_ASAP7_75t_L g1710 ( 
.A(n_1653),
.Y(n_1710)
);

OAI21x1_ASAP7_75t_L g1711 ( 
.A1(n_1649),
.A2(n_1477),
.B(n_1535),
.Y(n_1711)
);

OAI21x1_ASAP7_75t_L g1712 ( 
.A1(n_1654),
.A2(n_1495),
.B(n_1493),
.Y(n_1712)
);

OAI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1599),
.A2(n_1540),
.B(n_1525),
.Y(n_1713)
);

BUFx3_ASAP7_75t_L g1714 ( 
.A(n_1633),
.Y(n_1714)
);

O2A1O1Ixp33_ASAP7_75t_SL g1715 ( 
.A1(n_1613),
.A2(n_1517),
.B(n_1511),
.C(n_1451),
.Y(n_1715)
);

OAI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1678),
.A2(n_1661),
.B(n_1679),
.Y(n_1716)
);

OAI22x1_ASAP7_75t_L g1717 ( 
.A1(n_1670),
.A2(n_1609),
.B1(n_1634),
.B2(n_1675),
.Y(n_1717)
);

AOI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1643),
.A2(n_1546),
.B(n_1586),
.Y(n_1718)
);

A2O1A1Ixp33_ASAP7_75t_L g1719 ( 
.A1(n_1673),
.A2(n_1492),
.B(n_1495),
.C(n_1569),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1589),
.B(n_1506),
.Y(n_1720)
);

OAI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1656),
.A2(n_1540),
.B(n_1541),
.Y(n_1721)
);

AO31x2_ASAP7_75t_L g1722 ( 
.A1(n_1590),
.A2(n_1576),
.A3(n_1501),
.B(n_1488),
.Y(n_1722)
);

A2O1A1Ixp33_ASAP7_75t_L g1723 ( 
.A1(n_1644),
.A2(n_1573),
.B(n_1531),
.C(n_1514),
.Y(n_1723)
);

OAI21xp5_ASAP7_75t_L g1724 ( 
.A1(n_1598),
.A2(n_1564),
.B(n_1558),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1607),
.B(n_1641),
.Y(n_1725)
);

AOI21xp5_ASAP7_75t_L g1726 ( 
.A1(n_1608),
.A2(n_1586),
.B(n_1549),
.Y(n_1726)
);

AO21x2_ASAP7_75t_L g1727 ( 
.A1(n_1639),
.A2(n_1532),
.B(n_1514),
.Y(n_1727)
);

AOI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1640),
.A2(n_1553),
.B1(n_1450),
.B2(n_1442),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1653),
.Y(n_1729)
);

NAND3x1_ASAP7_75t_L g1730 ( 
.A(n_1588),
.B(n_1479),
.C(n_1563),
.Y(n_1730)
);

CKINVDCx14_ASAP7_75t_R g1731 ( 
.A(n_1714),
.Y(n_1731)
);

CKINVDCx20_ASAP7_75t_R g1732 ( 
.A(n_1709),
.Y(n_1732)
);

CKINVDCx6p67_ASAP7_75t_R g1733 ( 
.A(n_1680),
.Y(n_1733)
);

OA21x2_ASAP7_75t_L g1734 ( 
.A1(n_1698),
.A2(n_1664),
.B(n_1624),
.Y(n_1734)
);

OAI21x1_ASAP7_75t_L g1735 ( 
.A1(n_1689),
.A2(n_1630),
.B(n_1666),
.Y(n_1735)
);

NOR2xp67_ASAP7_75t_L g1736 ( 
.A(n_1717),
.B(n_1674),
.Y(n_1736)
);

OAI21x1_ASAP7_75t_L g1737 ( 
.A1(n_1682),
.A2(n_1668),
.B(n_1614),
.Y(n_1737)
);

AOI22xp33_ASAP7_75t_L g1738 ( 
.A1(n_1683),
.A2(n_1677),
.B1(n_1600),
.B2(n_1651),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_SL g1739 ( 
.A1(n_1685),
.A2(n_1628),
.B1(n_1653),
.B2(n_1627),
.Y(n_1739)
);

OAI21x1_ASAP7_75t_L g1740 ( 
.A1(n_1686),
.A2(n_1655),
.B(n_1646),
.Y(n_1740)
);

OAI21x1_ASAP7_75t_L g1741 ( 
.A1(n_1693),
.A2(n_1578),
.B(n_1610),
.Y(n_1741)
);

OAI21x1_ASAP7_75t_SL g1742 ( 
.A1(n_1718),
.A2(n_1595),
.B(n_1631),
.Y(n_1742)
);

OAI221xp5_ASAP7_75t_L g1743 ( 
.A1(n_1716),
.A2(n_1603),
.B1(n_1642),
.B2(n_1616),
.C(n_1622),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1684),
.B(n_1611),
.Y(n_1744)
);

INVxp67_ASAP7_75t_L g1745 ( 
.A(n_1704),
.Y(n_1745)
);

INVx4_ASAP7_75t_L g1746 ( 
.A(n_1694),
.Y(n_1746)
);

OAI21x1_ASAP7_75t_L g1747 ( 
.A1(n_1712),
.A2(n_1637),
.B(n_1479),
.Y(n_1747)
);

O2A1O1Ixp33_ASAP7_75t_L g1748 ( 
.A1(n_1702),
.A2(n_1723),
.B(n_1696),
.C(n_1719),
.Y(n_1748)
);

AOI22xp33_ASAP7_75t_L g1749 ( 
.A1(n_1713),
.A2(n_1652),
.B1(n_1671),
.B2(n_1667),
.Y(n_1749)
);

OAI21x1_ASAP7_75t_L g1750 ( 
.A1(n_1691),
.A2(n_1660),
.B(n_1648),
.Y(n_1750)
);

OA21x2_ASAP7_75t_L g1751 ( 
.A1(n_1705),
.A2(n_1629),
.B(n_1645),
.Y(n_1751)
);

OA21x2_ASAP7_75t_L g1752 ( 
.A1(n_1721),
.A2(n_1676),
.B(n_1657),
.Y(n_1752)
);

AND2x4_ASAP7_75t_L g1753 ( 
.A(n_1704),
.B(n_1618),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1699),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1688),
.Y(n_1755)
);

BUFx6f_ASAP7_75t_L g1756 ( 
.A(n_1706),
.Y(n_1756)
);

OAI22xp33_ASAP7_75t_L g1757 ( 
.A1(n_1725),
.A2(n_1658),
.B1(n_1621),
.B2(n_1617),
.Y(n_1757)
);

BUFx4f_ASAP7_75t_SL g1758 ( 
.A(n_1701),
.Y(n_1758)
);

INVx3_ASAP7_75t_L g1759 ( 
.A(n_1694),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1692),
.Y(n_1760)
);

OAI21x1_ASAP7_75t_L g1761 ( 
.A1(n_1695),
.A2(n_1563),
.B(n_1542),
.Y(n_1761)
);

OAI21xp5_ASAP7_75t_L g1762 ( 
.A1(n_1708),
.A2(n_1623),
.B(n_1550),
.Y(n_1762)
);

OAI22xp33_ASAP7_75t_L g1763 ( 
.A1(n_1687),
.A2(n_1555),
.B1(n_1577),
.B2(n_1618),
.Y(n_1763)
);

AOI221xp5_ASAP7_75t_L g1764 ( 
.A1(n_1700),
.A2(n_1582),
.B1(n_1530),
.B2(n_1626),
.C(n_1587),
.Y(n_1764)
);

NOR2xp33_ASAP7_75t_L g1765 ( 
.A(n_1720),
.B(n_1633),
.Y(n_1765)
);

OAI21x1_ASAP7_75t_L g1766 ( 
.A1(n_1711),
.A2(n_1653),
.B(n_1626),
.Y(n_1766)
);

AO21x2_ASAP7_75t_L g1767 ( 
.A1(n_1690),
.A2(n_1530),
.B(n_1626),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1760),
.B(n_1707),
.Y(n_1768)
);

A2O1A1Ixp33_ASAP7_75t_L g1769 ( 
.A1(n_1736),
.A2(n_1748),
.B(n_1762),
.C(n_1739),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1754),
.B(n_1722),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1755),
.Y(n_1771)
);

OAI22xp5_ASAP7_75t_L g1772 ( 
.A1(n_1739),
.A2(n_1730),
.B1(n_1728),
.B2(n_1729),
.Y(n_1772)
);

HB1xp67_ASAP7_75t_L g1773 ( 
.A(n_1745),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1745),
.B(n_1722),
.Y(n_1774)
);

CKINVDCx9p33_ASAP7_75t_R g1775 ( 
.A(n_1765),
.Y(n_1775)
);

AOI21xp5_ASAP7_75t_SL g1776 ( 
.A1(n_1757),
.A2(n_1748),
.B(n_1746),
.Y(n_1776)
);

O2A1O1Ixp33_ASAP7_75t_L g1777 ( 
.A1(n_1743),
.A2(n_1715),
.B(n_1724),
.C(n_1727),
.Y(n_1777)
);

AOI21x1_ASAP7_75t_SL g1778 ( 
.A1(n_1731),
.A2(n_1703),
.B(n_1685),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1751),
.B(n_1722),
.Y(n_1779)
);

CKINVDCx20_ASAP7_75t_R g1780 ( 
.A(n_1732),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1751),
.B(n_1729),
.Y(n_1781)
);

O2A1O1Ixp5_ASAP7_75t_L g1782 ( 
.A1(n_1757),
.A2(n_1703),
.B(n_1710),
.C(n_1726),
.Y(n_1782)
);

OAI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1738),
.A2(n_1710),
.B1(n_1706),
.B2(n_1697),
.Y(n_1783)
);

OAI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1743),
.A2(n_1706),
.B1(n_1681),
.B2(n_92),
.Y(n_1784)
);

AOI21xp5_ASAP7_75t_SL g1785 ( 
.A1(n_1746),
.A2(n_1681),
.B(n_90),
.Y(n_1785)
);

AOI21x1_ASAP7_75t_SL g1786 ( 
.A1(n_1753),
.A2(n_90),
.B(n_91),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1744),
.B(n_1681),
.Y(n_1787)
);

BUFx3_ASAP7_75t_L g1788 ( 
.A(n_1759),
.Y(n_1788)
);

NOR2xp67_ASAP7_75t_L g1789 ( 
.A(n_1759),
.B(n_93),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1750),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1733),
.B(n_93),
.Y(n_1791)
);

AOI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1763),
.A2(n_94),
.B(n_95),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1752),
.Y(n_1793)
);

HB1xp67_ASAP7_75t_L g1794 ( 
.A(n_1753),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1752),
.B(n_94),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1767),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1762),
.B(n_95),
.Y(n_1797)
);

BUFx3_ASAP7_75t_L g1798 ( 
.A(n_1788),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1793),
.Y(n_1799)
);

AO21x2_ASAP7_75t_L g1800 ( 
.A1(n_1785),
.A2(n_1742),
.B(n_1767),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1771),
.Y(n_1801)
);

OR2x6_ASAP7_75t_L g1802 ( 
.A(n_1776),
.B(n_1766),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1773),
.Y(n_1803)
);

AND2x4_ASAP7_75t_L g1804 ( 
.A(n_1781),
.B(n_1756),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1770),
.Y(n_1805)
);

INVx4_ASAP7_75t_SL g1806 ( 
.A(n_1788),
.Y(n_1806)
);

INVx3_ASAP7_75t_L g1807 ( 
.A(n_1793),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1768),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1774),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1774),
.Y(n_1810)
);

OA21x2_ASAP7_75t_L g1811 ( 
.A1(n_1796),
.A2(n_1747),
.B(n_1735),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1781),
.Y(n_1812)
);

HB1xp67_ASAP7_75t_L g1813 ( 
.A(n_1794),
.Y(n_1813)
);

CKINVDCx8_ASAP7_75t_R g1814 ( 
.A(n_1775),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1787),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1787),
.B(n_1749),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1779),
.B(n_1734),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1795),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1779),
.Y(n_1819)
);

OAI21xp5_ASAP7_75t_L g1820 ( 
.A1(n_1769),
.A2(n_1764),
.B(n_1737),
.Y(n_1820)
);

HB1xp67_ASAP7_75t_L g1821 ( 
.A(n_1795),
.Y(n_1821)
);

NOR4xp25_ASAP7_75t_SL g1822 ( 
.A(n_1814),
.B(n_1778),
.C(n_1764),
.D(n_1785),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1819),
.B(n_1796),
.Y(n_1823)
);

HB1xp67_ASAP7_75t_L g1824 ( 
.A(n_1803),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1799),
.Y(n_1825)
);

BUFx3_ASAP7_75t_L g1826 ( 
.A(n_1798),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1799),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1808),
.B(n_1809),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1801),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1801),
.Y(n_1830)
);

HB1xp67_ASAP7_75t_L g1831 ( 
.A(n_1813),
.Y(n_1831)
);

INVx2_ASAP7_75t_SL g1832 ( 
.A(n_1798),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1809),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1819),
.B(n_1790),
.Y(n_1834)
);

HB1xp67_ASAP7_75t_L g1835 ( 
.A(n_1812),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1807),
.Y(n_1836)
);

INVx4_ASAP7_75t_R g1837 ( 
.A(n_1814),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1810),
.Y(n_1838)
);

OR2x2_ASAP7_75t_L g1839 ( 
.A(n_1810),
.B(n_1783),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1821),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1812),
.B(n_1790),
.Y(n_1841)
);

AOI22xp33_ASAP7_75t_SL g1842 ( 
.A1(n_1826),
.A2(n_1832),
.B1(n_1772),
.B2(n_1824),
.Y(n_1842)
);

AO21x2_ASAP7_75t_L g1843 ( 
.A1(n_1840),
.A2(n_1820),
.B(n_1791),
.Y(n_1843)
);

AOI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1831),
.A2(n_1816),
.B1(n_1818),
.B2(n_1758),
.Y(n_1844)
);

CKINVDCx20_ASAP7_75t_R g1845 ( 
.A(n_1826),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1835),
.Y(n_1846)
);

OR2x2_ASAP7_75t_L g1847 ( 
.A(n_1828),
.B(n_1833),
.Y(n_1847)
);

BUFx2_ASAP7_75t_L g1848 ( 
.A(n_1832),
.Y(n_1848)
);

AOI22xp33_ASAP7_75t_SL g1849 ( 
.A1(n_1839),
.A2(n_1802),
.B1(n_1780),
.B2(n_1800),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_SL g1850 ( 
.A(n_1839),
.B(n_1806),
.Y(n_1850)
);

OAI22xp33_ASAP7_75t_L g1851 ( 
.A1(n_1837),
.A2(n_1802),
.B1(n_1818),
.B2(n_1789),
.Y(n_1851)
);

AOI22xp33_ASAP7_75t_L g1852 ( 
.A1(n_1833),
.A2(n_1797),
.B1(n_1817),
.B2(n_1802),
.Y(n_1852)
);

AOI222xp33_ASAP7_75t_SL g1853 ( 
.A1(n_1838),
.A2(n_1784),
.B1(n_1780),
.B2(n_1805),
.C1(n_1815),
.C2(n_1807),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1825),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1838),
.B(n_1805),
.Y(n_1855)
);

OR2x2_ASAP7_75t_L g1856 ( 
.A(n_1825),
.B(n_1815),
.Y(n_1856)
);

INVx1_ASAP7_75t_SL g1857 ( 
.A(n_1823),
.Y(n_1857)
);

OAI22xp33_ASAP7_75t_L g1858 ( 
.A1(n_1836),
.A2(n_1802),
.B1(n_1792),
.B2(n_1807),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1829),
.B(n_1817),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1829),
.B(n_1804),
.Y(n_1860)
);

AOI22xp33_ASAP7_75t_L g1861 ( 
.A1(n_1830),
.A2(n_1800),
.B1(n_1804),
.B2(n_1806),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1823),
.B(n_1804),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1855),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1847),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1846),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1843),
.B(n_1830),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1859),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1848),
.B(n_1841),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1860),
.Y(n_1869)
);

INVx3_ASAP7_75t_L g1870 ( 
.A(n_1854),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1868),
.B(n_1842),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1865),
.B(n_1856),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1864),
.B(n_1862),
.Y(n_1873)
);

INVx2_ASAP7_75t_SL g1874 ( 
.A(n_1865),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1871),
.B(n_1867),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1873),
.B(n_1869),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1875),
.B(n_1876),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1876),
.B(n_1874),
.Y(n_1878)
);

NAND2x1p5_ASAP7_75t_L g1879 ( 
.A(n_1876),
.B(n_1850),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1875),
.B(n_1874),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1880),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1878),
.Y(n_1882)
);

AOI21xp33_ASAP7_75t_SL g1883 ( 
.A1(n_1879),
.A2(n_1877),
.B(n_1851),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1880),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1878),
.B(n_1863),
.Y(n_1885)
);

O2A1O1Ixp5_ASAP7_75t_L g1886 ( 
.A1(n_1877),
.A2(n_1866),
.B(n_1851),
.C(n_1858),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1880),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1881),
.B(n_1866),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1884),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1887),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1882),
.B(n_1845),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1882),
.B(n_1872),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1885),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1886),
.Y(n_1894)
);

INVx3_ASAP7_75t_L g1895 ( 
.A(n_1883),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1886),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1881),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1894),
.B(n_1843),
.Y(n_1898)
);

NAND3xp33_ASAP7_75t_L g1899 ( 
.A(n_1896),
.B(n_1849),
.C(n_1853),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1895),
.B(n_1844),
.Y(n_1900)
);

AOI21xp33_ASAP7_75t_SL g1901 ( 
.A1(n_1889),
.A2(n_1858),
.B(n_96),
.Y(n_1901)
);

AOI22xp5_ASAP7_75t_L g1902 ( 
.A1(n_1891),
.A2(n_1844),
.B1(n_1852),
.B2(n_1870),
.Y(n_1902)
);

INVxp67_ASAP7_75t_SL g1903 ( 
.A(n_1890),
.Y(n_1903)
);

OAI221xp5_ASAP7_75t_L g1904 ( 
.A1(n_1895),
.A2(n_1861),
.B1(n_1852),
.B2(n_1777),
.C(n_1870),
.Y(n_1904)
);

OAI21xp5_ASAP7_75t_SL g1905 ( 
.A1(n_1897),
.A2(n_1822),
.B(n_1857),
.Y(n_1905)
);

OAI21xp33_ASAP7_75t_L g1906 ( 
.A1(n_1893),
.A2(n_1836),
.B(n_1834),
.Y(n_1906)
);

AND5x1_ASAP7_75t_L g1907 ( 
.A(n_1888),
.B(n_1786),
.C(n_97),
.D(n_98),
.E(n_99),
.Y(n_1907)
);

AOI221xp5_ASAP7_75t_L g1908 ( 
.A1(n_1888),
.A2(n_1782),
.B1(n_1800),
.B2(n_1827),
.C(n_1834),
.Y(n_1908)
);

AOI21xp5_ASAP7_75t_L g1909 ( 
.A1(n_1892),
.A2(n_1811),
.B(n_1827),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1894),
.B(n_1841),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1894),
.B(n_96),
.Y(n_1911)
);

OAI21xp5_ASAP7_75t_L g1912 ( 
.A1(n_1894),
.A2(n_1741),
.B(n_1740),
.Y(n_1912)
);

AOI211xp5_ASAP7_75t_L g1913 ( 
.A1(n_1894),
.A2(n_101),
.B(n_98),
.C(n_100),
.Y(n_1913)
);

O2A1O1Ixp5_ASAP7_75t_L g1914 ( 
.A1(n_1894),
.A2(n_104),
.B(n_100),
.C(n_103),
.Y(n_1914)
);

OAI221xp5_ASAP7_75t_L g1915 ( 
.A1(n_1905),
.A2(n_1756),
.B1(n_106),
.B2(n_107),
.C(n_108),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1911),
.Y(n_1916)
);

AOI221xp5_ASAP7_75t_L g1917 ( 
.A1(n_1914),
.A2(n_1756),
.B1(n_106),
.B2(n_109),
.C(n_110),
.Y(n_1917)
);

AOI22xp5_ASAP7_75t_L g1918 ( 
.A1(n_1899),
.A2(n_1806),
.B1(n_1811),
.B2(n_1734),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1910),
.Y(n_1919)
);

AOI22xp5_ASAP7_75t_L g1920 ( 
.A1(n_1900),
.A2(n_1806),
.B1(n_1811),
.B2(n_1761),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1898),
.Y(n_1921)
);

OAI21xp5_ASAP7_75t_L g1922 ( 
.A1(n_1913),
.A2(n_1903),
.B(n_1904),
.Y(n_1922)
);

AOI311xp33_ASAP7_75t_L g1923 ( 
.A1(n_1912),
.A2(n_105),
.A3(n_110),
.B(n_111),
.C(n_113),
.Y(n_1923)
);

OAI32xp33_ASAP7_75t_L g1924 ( 
.A1(n_1906),
.A2(n_105),
.A3(n_111),
.B1(n_114),
.B2(n_115),
.Y(n_1924)
);

A2O1A1Ixp33_ASAP7_75t_L g1925 ( 
.A1(n_1901),
.A2(n_114),
.B(n_116),
.C(n_117),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1902),
.B(n_1908),
.Y(n_1926)
);

NAND4xp25_ASAP7_75t_L g1927 ( 
.A(n_1909),
.B(n_119),
.C(n_120),
.D(n_121),
.Y(n_1927)
);

NAND5xp2_ASAP7_75t_L g1928 ( 
.A(n_1907),
.B(n_120),
.C(n_140),
.D(n_141),
.E(n_145),
.Y(n_1928)
);

OAI211xp5_ASAP7_75t_L g1929 ( 
.A1(n_1913),
.A2(n_1811),
.B(n_150),
.C(n_152),
.Y(n_1929)
);

AOI22xp5_ASAP7_75t_L g1930 ( 
.A1(n_1899),
.A2(n_147),
.B1(n_157),
.B2(n_158),
.Y(n_1930)
);

AOI22xp33_ASAP7_75t_L g1931 ( 
.A1(n_1899),
.A2(n_159),
.B1(n_160),
.B2(n_164),
.Y(n_1931)
);

NOR3xp33_ASAP7_75t_L g1932 ( 
.A(n_1915),
.B(n_166),
.C(n_167),
.Y(n_1932)
);

INVx2_ASAP7_75t_SL g1933 ( 
.A(n_1919),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1925),
.B(n_173),
.Y(n_1934)
);

INVx2_ASAP7_75t_SL g1935 ( 
.A(n_1921),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1924),
.Y(n_1936)
);

INVxp67_ASAP7_75t_L g1937 ( 
.A(n_1928),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1916),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1922),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1931),
.B(n_174),
.Y(n_1940)
);

BUFx12f_ASAP7_75t_L g1941 ( 
.A(n_1923),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1926),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1930),
.B(n_175),
.Y(n_1943)
);

OR2x2_ASAP7_75t_L g1944 ( 
.A(n_1927),
.B(n_1918),
.Y(n_1944)
);

NAND3xp33_ASAP7_75t_L g1945 ( 
.A(n_1917),
.B(n_177),
.C(n_178),
.Y(n_1945)
);

INVx1_ASAP7_75t_SL g1946 ( 
.A(n_1920),
.Y(n_1946)
);

AND3x1_ASAP7_75t_L g1947 ( 
.A(n_1929),
.B(n_180),
.C(n_183),
.Y(n_1947)
);

HB1xp67_ASAP7_75t_L g1948 ( 
.A(n_1921),
.Y(n_1948)
);

HB1xp67_ASAP7_75t_L g1949 ( 
.A(n_1948),
.Y(n_1949)
);

NAND3xp33_ASAP7_75t_L g1950 ( 
.A(n_1942),
.B(n_184),
.C(n_185),
.Y(n_1950)
);

OAI221xp5_ASAP7_75t_L g1951 ( 
.A1(n_1937),
.A2(n_187),
.B1(n_190),
.B2(n_191),
.C(n_192),
.Y(n_1951)
);

OAI21xp33_ASAP7_75t_L g1952 ( 
.A1(n_1939),
.A2(n_193),
.B(n_197),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1935),
.B(n_198),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1933),
.B(n_201),
.Y(n_1954)
);

OAI321xp33_ASAP7_75t_L g1955 ( 
.A1(n_1936),
.A2(n_204),
.A3(n_206),
.B1(n_207),
.B2(n_211),
.C(n_212),
.Y(n_1955)
);

AOI221xp5_ASAP7_75t_L g1956 ( 
.A1(n_1932),
.A2(n_215),
.B1(n_217),
.B2(n_218),
.C(n_219),
.Y(n_1956)
);

NAND3xp33_ASAP7_75t_L g1957 ( 
.A(n_1934),
.B(n_221),
.C(n_224),
.Y(n_1957)
);

OAI21xp5_ASAP7_75t_L g1958 ( 
.A1(n_1945),
.A2(n_227),
.B(n_228),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1944),
.Y(n_1959)
);

OAI211xp5_ASAP7_75t_SL g1960 ( 
.A1(n_1938),
.A2(n_229),
.B(n_230),
.C(n_232),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1941),
.Y(n_1961)
);

OR2x2_ASAP7_75t_L g1962 ( 
.A(n_1946),
.B(n_234),
.Y(n_1962)
);

OR2x2_ASAP7_75t_L g1963 ( 
.A(n_1961),
.B(n_1943),
.Y(n_1963)
);

OAI22xp5_ASAP7_75t_SL g1964 ( 
.A1(n_1959),
.A2(n_1947),
.B1(n_1940),
.B2(n_242),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1949),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1962),
.Y(n_1966)
);

NOR4xp75_ASAP7_75t_SL g1967 ( 
.A(n_1953),
.B(n_1947),
.C(n_239),
.D(n_243),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1954),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1956),
.B(n_1958),
.Y(n_1969)
);

NOR2x1p5_ASAP7_75t_L g1970 ( 
.A(n_1957),
.B(n_237),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1952),
.B(n_244),
.Y(n_1971)
);

AOI22xp5_ASAP7_75t_L g1972 ( 
.A1(n_1951),
.A2(n_246),
.B1(n_247),
.B2(n_249),
.Y(n_1972)
);

OAI221xp5_ASAP7_75t_L g1973 ( 
.A1(n_1950),
.A2(n_1960),
.B1(n_1955),
.B2(n_252),
.C(n_254),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1949),
.B(n_250),
.Y(n_1974)
);

XNOR2x1_ASAP7_75t_L g1975 ( 
.A(n_1970),
.B(n_251),
.Y(n_1975)
);

NOR2x1_ASAP7_75t_L g1976 ( 
.A(n_1965),
.B(n_255),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1966),
.Y(n_1977)
);

AND3x1_ASAP7_75t_L g1978 ( 
.A(n_1974),
.B(n_258),
.C(n_262),
.Y(n_1978)
);

OR3x1_ASAP7_75t_L g1979 ( 
.A(n_1968),
.B(n_263),
.C(n_264),
.Y(n_1979)
);

CKINVDCx5p33_ASAP7_75t_R g1980 ( 
.A(n_1964),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1972),
.B(n_265),
.Y(n_1981)
);

AOI22xp5_ASAP7_75t_L g1982 ( 
.A1(n_1980),
.A2(n_1973),
.B1(n_1969),
.B2(n_1963),
.Y(n_1982)
);

NAND3xp33_ASAP7_75t_SL g1983 ( 
.A(n_1977),
.B(n_1971),
.C(n_1967),
.Y(n_1983)
);

AOI322xp5_ASAP7_75t_L g1984 ( 
.A1(n_1981),
.A2(n_266),
.A3(n_267),
.B1(n_269),
.B2(n_271),
.C1(n_272),
.C2(n_274),
.Y(n_1984)
);

A2O1A1Ixp33_ASAP7_75t_L g1985 ( 
.A1(n_1976),
.A2(n_275),
.B(n_276),
.C(n_281),
.Y(n_1985)
);

AOI322xp5_ASAP7_75t_L g1986 ( 
.A1(n_1979),
.A2(n_284),
.A3(n_287),
.B1(n_289),
.B2(n_291),
.C1(n_293),
.C2(n_296),
.Y(n_1986)
);

AOI21x1_ASAP7_75t_L g1987 ( 
.A1(n_1982),
.A2(n_1975),
.B(n_1978),
.Y(n_1987)
);

OAI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1985),
.A2(n_297),
.B1(n_299),
.B2(n_301),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_SL g1989 ( 
.A(n_1986),
.B(n_302),
.Y(n_1989)
);

AND2x4_ASAP7_75t_L g1990 ( 
.A(n_1987),
.B(n_1983),
.Y(n_1990)
);

AOI21xp5_ASAP7_75t_L g1991 ( 
.A1(n_1989),
.A2(n_1984),
.B(n_304),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1988),
.B(n_303),
.Y(n_1992)
);

XNOR2xp5_ASAP7_75t_L g1993 ( 
.A(n_1987),
.B(n_305),
.Y(n_1993)
);

OAI22xp5_ASAP7_75t_L g1994 ( 
.A1(n_1993),
.A2(n_306),
.B1(n_309),
.B2(n_312),
.Y(n_1994)
);

AO22x2_ASAP7_75t_L g1995 ( 
.A1(n_1990),
.A2(n_438),
.B1(n_320),
.B2(n_322),
.Y(n_1995)
);

AOI22xp5_ASAP7_75t_L g1996 ( 
.A1(n_1991),
.A2(n_318),
.B1(n_325),
.B2(n_326),
.Y(n_1996)
);

INVxp67_ASAP7_75t_SL g1997 ( 
.A(n_1996),
.Y(n_1997)
);

CKINVDCx20_ASAP7_75t_R g1998 ( 
.A(n_1994),
.Y(n_1998)
);

AOI21xp5_ASAP7_75t_L g1999 ( 
.A1(n_1997),
.A2(n_1995),
.B(n_1992),
.Y(n_1999)
);

AOI22xp5_ASAP7_75t_L g2000 ( 
.A1(n_1999),
.A2(n_1998),
.B1(n_328),
.B2(n_329),
.Y(n_2000)
);

AOI22x1_ASAP7_75t_L g2001 ( 
.A1(n_2000),
.A2(n_327),
.B1(n_330),
.B2(n_331),
.Y(n_2001)
);

AOI221xp5_ASAP7_75t_L g2002 ( 
.A1(n_2001),
.A2(n_332),
.B1(n_336),
.B2(n_337),
.C(n_338),
.Y(n_2002)
);

AOI211xp5_ASAP7_75t_L g2003 ( 
.A1(n_2002),
.A2(n_344),
.B(n_345),
.C(n_346),
.Y(n_2003)
);


endmodule