module fake_jpeg_1694_n_190 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_190);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_190;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_30),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_14),
.B(n_1),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_20),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_22),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_8),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_33),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_1),
.Y(n_66)
);

NAND3xp33_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_67),
.C(n_68),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_21),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_65),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx6_ASAP7_75t_SL g70 ( 
.A(n_52),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_70),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_72),
.A2(n_64),
.B1(n_50),
.B2(n_53),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_50),
.B1(n_62),
.B2(n_49),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_78),
.A2(n_73),
.B1(n_61),
.B2(n_60),
.Y(n_99)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_62),
.B1(n_64),
.B2(n_57),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_64),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_84),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_70),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_71),
.Y(n_88)
);

NAND5xp2_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_83),
.C(n_48),
.D(n_46),
.E(n_59),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_54),
.C(n_3),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_98),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_57),
.B1(n_47),
.B2(n_60),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_46),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_94),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_59),
.B(n_51),
.C(n_63),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_91),
.B(n_93),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_77),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_51),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_53),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_101),
.Y(n_112)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_100),
.Y(n_104)
);

INVxp67_ASAP7_75t_SL g100 ( 
.A(n_75),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_84),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_102),
.B(n_6),
.Y(n_123)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_71),
.B(n_63),
.Y(n_105)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_61),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_111),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_120),
.B1(n_10),
.B2(n_11),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_2),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_115),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_86),
.Y(n_115)
);

INVx3_ASAP7_75t_SL g116 ( 
.A(n_95),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_103),
.A2(n_23),
.B1(n_44),
.B2(n_43),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_117),
.A2(n_118),
.B1(n_92),
.B2(n_99),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_89),
.A2(n_103),
.B1(n_99),
.B2(n_87),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_97),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_123),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_99),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_26),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_110),
.B(n_6),
.Y(n_126)
);

NAND3xp33_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_133),
.C(n_136),
.Y(n_159)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_135),
.Y(n_148)
);

FAx1_ASAP7_75t_SL g130 ( 
.A(n_111),
.B(n_120),
.CI(n_122),
.CON(n_130),
.SN(n_130)
);

AOI322xp5_ASAP7_75t_L g145 ( 
.A1(n_130),
.A2(n_105),
.A3(n_108),
.B1(n_117),
.B2(n_29),
.C1(n_45),
.C2(n_38),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_104),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_131),
.A2(n_142),
.B1(n_12),
.B2(n_14),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_107),
.B(n_9),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_119),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_139),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_27),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_15),
.C(n_16),
.Y(n_158)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_141),
.Y(n_154)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_104),
.A2(n_28),
.B1(n_42),
.B2(n_40),
.Y(n_142)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_144),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_145),
.B(n_146),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_128),
.B(n_121),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_143),
.B(n_37),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_155),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_150),
.A2(n_152),
.B1(n_135),
.B2(n_142),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_134),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_36),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_158),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_15),
.Y(n_157)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_157),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_125),
.Y(n_160)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_160),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_167),
.Y(n_176)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_154),
.Y(n_163)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_163),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_153),
.A2(n_130),
.B1(n_131),
.B2(n_127),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_166),
.Y(n_173)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_127),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_170),
.A2(n_153),
.B(n_163),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_171),
.B(n_155),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_174),
.C(n_178),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_171),
.B(n_147),
.C(n_156),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_177),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_151),
.C(n_158),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_179),
.B(n_181),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_176),
.A2(n_169),
.B(n_161),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_170),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_182),
.A2(n_165),
.B1(n_164),
.B2(n_168),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_183),
.A2(n_182),
.B1(n_180),
.B2(n_159),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_185),
.A2(n_184),
.B(n_183),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_152),
.Y(n_187)
);

AOI322xp5_ASAP7_75t_L g188 ( 
.A1(n_187),
.A2(n_144),
.A3(n_17),
.B1(n_18),
.B2(n_19),
.C1(n_20),
.C2(n_16),
.Y(n_188)
);

OAI221xp5_ASAP7_75t_SL g189 ( 
.A1(n_188),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.C(n_25),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_34),
.Y(n_190)
);


endmodule