module fake_jpeg_31684_n_448 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_448);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_448;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx8_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_12),
.B(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

BUFx24_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_30),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_52),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_50),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_51),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_15),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_15),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_58),
.Y(n_95)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_55),
.Y(n_142)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_18),
.B(n_1),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_18),
.B(n_32),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_59),
.B(n_60),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_22),
.B(n_2),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_61),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_22),
.B(n_2),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_62),
.B(n_63),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_19),
.B(n_2),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_30),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_70),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_19),
.B(n_3),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_66),
.B(n_72),
.Y(n_114)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_32),
.B(n_3),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_33),
.B(n_3),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_33),
.B(n_3),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_73),
.Y(n_113)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

BUFx10_ASAP7_75t_L g75 ( 
.A(n_16),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_75),
.Y(n_124)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_16),
.Y(n_76)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_76),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_40),
.B(n_4),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_79),
.Y(n_133)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_83),
.Y(n_129)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_88),
.A2(n_89),
.B1(n_55),
.B2(n_76),
.Y(n_94)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_16),
.Y(n_90)
);

NAND2x1_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_30),
.Y(n_125)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_89),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_46),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_92),
.A2(n_46),
.B1(n_24),
.B2(n_27),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_94),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_100),
.A2(n_9),
.B(n_10),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_74),
.A2(n_24),
.B1(n_44),
.B2(n_39),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_110),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_63),
.A2(n_24),
.B1(n_44),
.B2(n_39),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_82),
.A2(n_23),
.B1(n_44),
.B2(n_39),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_66),
.A2(n_20),
.B1(n_38),
.B2(n_35),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_64),
.A2(n_20),
.B1(n_38),
.B2(n_35),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_119),
.B(n_121),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_61),
.A2(n_20),
.B1(n_38),
.B2(n_35),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_122),
.A2(n_128),
.B1(n_48),
.B2(n_55),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_125),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_67),
.A2(n_17),
.B1(n_34),
.B2(n_28),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_80),
.B(n_17),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_137),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_83),
.A2(n_17),
.B1(n_34),
.B2(n_28),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_71),
.A2(n_45),
.B1(n_27),
.B2(n_34),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_138),
.A2(n_140),
.B1(n_144),
.B2(n_29),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_81),
.B(n_45),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_75),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_87),
.A2(n_88),
.B1(n_85),
.B2(n_68),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_69),
.A2(n_45),
.B1(n_28),
.B2(n_27),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_145),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_107),
.B(n_23),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_147),
.B(n_160),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_148),
.A2(n_169),
.B1(n_172),
.B2(n_179),
.Y(n_212)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_111),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_149),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_98),
.B(n_53),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_150),
.B(n_173),
.Y(n_230)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_97),
.Y(n_151)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_151),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_152),
.B(n_165),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_98),
.B(n_56),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_153),
.B(n_170),
.Y(n_203)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_97),
.Y(n_154)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_154),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_23),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_155),
.B(n_159),
.Y(n_198)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_105),
.Y(n_156)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_156),
.Y(n_227)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_105),
.Y(n_158)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_158),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_114),
.B(n_75),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_121),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_161),
.Y(n_200)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_164),
.Y(n_210)
);

OA22x2_ASAP7_75t_L g165 ( 
.A1(n_125),
.A2(n_48),
.B1(n_75),
.B2(n_90),
.Y(n_165)
);

INVx11_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_166),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_109),
.Y(n_167)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_167),
.Y(n_213)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_120),
.Y(n_168)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_168),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_113),
.A2(n_47),
.B1(n_57),
.B2(n_50),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_29),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_171),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_103),
.A2(n_51),
.B1(n_50),
.B2(n_78),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_130),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_136),
.B(n_30),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_174),
.B(n_180),
.Y(n_209)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_131),
.Y(n_176)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_176),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_106),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_177),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_104),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_178),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_134),
.A2(n_51),
.B1(n_77),
.B2(n_30),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_130),
.Y(n_180)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_111),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_181),
.B(n_184),
.Y(n_229)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_129),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_182),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_109),
.A2(n_30),
.B1(n_42),
.B2(n_29),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_183),
.A2(n_186),
.B1(n_188),
.B2(n_190),
.Y(n_195)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_127),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_139),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_185),
.Y(n_196)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_129),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_187),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_123),
.A2(n_29),
.B1(n_6),
.B2(n_8),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_136),
.B(n_5),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_191),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_123),
.A2(n_101),
.B1(n_115),
.B2(n_96),
.Y(n_190)
);

O2A1O1Ixp33_ASAP7_75t_L g191 ( 
.A1(n_116),
.A2(n_29),
.B(n_6),
.C(n_8),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_136),
.B(n_5),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_9),
.Y(n_214)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_115),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_193),
.B(n_141),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_194),
.A2(n_118),
.B1(n_95),
.B2(n_93),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_197),
.A2(n_146),
.B1(n_152),
.B2(n_147),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_159),
.B(n_101),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_207),
.B(n_217),
.C(n_220),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_161),
.A2(n_135),
.B1(n_112),
.B2(n_106),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_211),
.A2(n_234),
.B1(n_173),
.B2(n_180),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_214),
.B(n_11),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_135),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_191),
.Y(n_246)
);

MAJx2_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_104),
.C(n_96),
.Y(n_217)
);

FAx1_ASAP7_75t_SL g219 ( 
.A(n_155),
.B(n_126),
.CI(n_142),
.CON(n_219),
.SN(n_219)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_219),
.B(n_163),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_108),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_175),
.B(n_108),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_221),
.B(n_231),
.C(n_99),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_145),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_224),
.B(n_225),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_150),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_175),
.B(n_126),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_164),
.A2(n_102),
.B1(n_112),
.B2(n_132),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_233),
.A2(n_162),
.B1(n_193),
.B2(n_177),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_146),
.A2(n_102),
.B1(n_143),
.B2(n_141),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_165),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_175),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_157),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_236),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_239),
.B(n_245),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_160),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_240),
.B(n_256),
.Y(n_293)
);

BUFx5_ASAP7_75t_L g241 ( 
.A(n_232),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_241),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_242),
.B(n_251),
.Y(n_305)
);

A2O1A1O1Ixp25_ASAP7_75t_L g243 ( 
.A1(n_198),
.A2(n_199),
.B(n_216),
.C(n_209),
.D(n_235),
.Y(n_243)
);

A2O1A1Ixp33_ASAP7_75t_L g304 ( 
.A1(n_243),
.A2(n_211),
.B(n_226),
.C(n_204),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_244),
.A2(n_263),
.B1(n_269),
.B2(n_275),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_236),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_246),
.B(n_255),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_247),
.B(n_250),
.Y(n_302)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_200),
.Y(n_248)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_248),
.Y(n_285)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_200),
.Y(n_249)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_249),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_203),
.B(n_157),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_252),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_229),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_253),
.B(n_254),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_197),
.B(n_184),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_198),
.B(n_194),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_207),
.B(n_151),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_258),
.A2(n_237),
.B1(n_227),
.B2(n_206),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_223),
.A2(n_199),
.B(n_210),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_259),
.A2(n_271),
.B(n_204),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_215),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_260),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_230),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_261),
.B(n_267),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_196),
.B(n_154),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_262),
.B(n_274),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_210),
.A2(n_162),
.B1(n_158),
.B2(n_156),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_223),
.B(n_165),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_264),
.Y(n_290)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_205),
.Y(n_266)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_266),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_230),
.B(n_165),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_223),
.B(n_187),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_268),
.A2(n_270),
.B(n_195),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_235),
.A2(n_182),
.B1(n_168),
.B2(n_171),
.Y(n_269)
);

AO21x1_ASAP7_75t_L g270 ( 
.A1(n_212),
.A2(n_142),
.B(n_143),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_219),
.A2(n_142),
.B(n_149),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_218),
.B(n_99),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_272),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_195),
.A2(n_166),
.B1(n_181),
.B2(n_127),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_273),
.A2(n_208),
.B1(n_13),
.B2(n_14),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_231),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_220),
.B(n_221),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_217),
.C(n_214),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_257),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_265),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_279),
.B(n_295),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_282),
.A2(n_304),
.B(n_307),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_283),
.B(n_289),
.C(n_292),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_284),
.B(n_297),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g341 ( 
.A1(n_287),
.A2(n_311),
.B1(n_241),
.B2(n_263),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_257),
.B(n_234),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_213),
.C(n_202),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_202),
.C(n_201),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_294),
.B(n_301),
.Y(n_326)
);

BUFx24_ASAP7_75t_SL g295 ( 
.A(n_250),
.Y(n_295)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_256),
.B(n_228),
.C(n_222),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_262),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_298),
.B(n_253),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_240),
.B(n_232),
.C(n_227),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_271),
.A2(n_204),
.B(n_226),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_308),
.A2(n_267),
.B(n_252),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_243),
.B(n_206),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_309),
.B(n_268),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_264),
.A2(n_205),
.B1(n_208),
.B2(n_13),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_310),
.Y(n_322)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_285),
.Y(n_314)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_314),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_312),
.A2(n_260),
.B1(n_240),
.B2(n_259),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_315),
.A2(n_340),
.B1(n_296),
.B2(n_305),
.Y(n_344)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_285),
.Y(n_316)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_316),
.Y(n_349)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_286),
.Y(n_317)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_317),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_282),
.A2(n_270),
.B(n_264),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_319),
.B(n_323),
.Y(n_356)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_286),
.Y(n_320)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_320),
.Y(n_357)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_299),
.Y(n_321)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_321),
.Y(n_360)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_299),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_298),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_324),
.A2(n_329),
.B1(n_331),
.B2(n_333),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_278),
.B(n_255),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_325),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_330),
.B(n_334),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_278),
.B(n_293),
.Y(n_331)
);

BUFx24_ASAP7_75t_L g332 ( 
.A(n_300),
.Y(n_332)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_332),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_293),
.B(n_246),
.Y(n_333)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_301),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_335),
.A2(n_336),
.B1(n_338),
.B2(n_283),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_306),
.B(n_244),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_307),
.A2(n_247),
.B(n_268),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_337),
.B(n_306),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_291),
.B(n_239),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_288),
.B(n_277),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_339),
.B(n_284),
.C(n_292),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_308),
.A2(n_270),
.B(n_252),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_341),
.A2(n_242),
.B1(n_310),
.B2(n_273),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_343),
.B(n_346),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_344),
.A2(n_351),
.B1(n_353),
.B2(n_355),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_313),
.B(n_288),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_315),
.A2(n_305),
.B1(n_289),
.B2(n_309),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_340),
.A2(n_305),
.B1(n_302),
.B2(n_290),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_354),
.A2(n_280),
.B1(n_320),
.B2(n_317),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_335),
.A2(n_290),
.B1(n_296),
.B2(n_303),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_322),
.A2(n_304),
.B1(n_311),
.B2(n_258),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_358),
.B(n_362),
.Y(n_368)
);

BUFx24_ASAP7_75t_SL g359 ( 
.A(n_318),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_359),
.B(n_280),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_361),
.B(n_364),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_322),
.A2(n_312),
.B1(n_336),
.B2(n_325),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_363),
.B(n_339),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_313),
.B(n_294),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_327),
.B(n_297),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_365),
.B(n_366),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_326),
.B(n_281),
.C(n_279),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_367),
.B(n_372),
.Y(n_398)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_347),
.Y(n_369)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_369),
.Y(n_392)
);

OAI31xp33_ASAP7_75t_L g370 ( 
.A1(n_356),
.A2(n_331),
.A3(n_333),
.B(n_319),
.Y(n_370)
);

A2O1A1Ixp33_ASAP7_75t_L g393 ( 
.A1(n_370),
.A2(n_351),
.B(n_248),
.C(n_357),
.Y(n_393)
);

FAx1_ASAP7_75t_SL g371 ( 
.A(n_361),
.B(n_334),
.CI(n_327),
.CON(n_371),
.SN(n_371)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_371),
.B(n_373),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_352),
.B(n_338),
.Y(n_372)
);

FAx1_ASAP7_75t_SL g373 ( 
.A(n_342),
.B(n_337),
.CI(n_326),
.CON(n_373),
.SN(n_373)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_355),
.B(n_324),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_374),
.B(n_375),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_360),
.B(n_316),
.Y(n_376)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_376),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_377),
.B(n_378),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_342),
.A2(n_328),
.B1(n_314),
.B2(n_330),
.Y(n_378)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_345),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_381),
.B(n_384),
.Y(n_388)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_349),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_350),
.B(n_323),
.Y(n_385)
);

INVx13_ASAP7_75t_L g396 ( 
.A(n_385),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_358),
.A2(n_328),
.B1(n_321),
.B2(n_249),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_386),
.A2(n_332),
.B(n_348),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_382),
.B(n_364),
.C(n_346),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_389),
.B(n_390),
.C(n_394),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_382),
.B(n_343),
.C(n_366),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_383),
.A2(n_344),
.B(n_353),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_391),
.A2(n_401),
.B(n_373),
.Y(n_412)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_393),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_379),
.B(n_365),
.C(n_348),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_399),
.B(n_376),
.Y(n_408)
);

INVxp33_ASAP7_75t_SL g400 ( 
.A(n_370),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_400),
.B(n_386),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_383),
.A2(n_332),
.B(n_275),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_391),
.A2(n_374),
.B1(n_369),
.B2(n_368),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_403),
.A2(n_412),
.B1(n_405),
.B2(n_407),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_398),
.B(n_377),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_404),
.B(n_406),
.Y(n_422)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_405),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_399),
.A2(n_378),
.B(n_368),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_408),
.B(n_409),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_388),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_397),
.B(n_375),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_410),
.B(n_394),
.C(n_390),
.Y(n_420)
);

OR2x2_ASAP7_75t_L g411 ( 
.A(n_396),
.B(n_385),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_411),
.A2(n_414),
.B1(n_388),
.B2(n_332),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_402),
.A2(n_395),
.B1(n_397),
.B2(n_393),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_413),
.A2(n_401),
.B1(n_388),
.B2(n_392),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_402),
.A2(n_384),
.B(n_381),
.Y(n_414)
);

AOI21x1_ASAP7_75t_SL g416 ( 
.A1(n_411),
.A2(n_396),
.B(n_395),
.Y(n_416)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_416),
.Y(n_432)
);

BUFx24_ASAP7_75t_SL g417 ( 
.A(n_410),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_417),
.B(n_419),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_418),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_420),
.B(n_415),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_421),
.B(n_414),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_403),
.A2(n_387),
.B1(n_380),
.B2(n_373),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_423),
.A2(n_413),
.B1(n_406),
.B2(n_408),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_415),
.B(n_389),
.C(n_379),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_424),
.A2(n_412),
.B(n_387),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_429),
.B(n_430),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_431),
.B(n_434),
.Y(n_437)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_433),
.Y(n_436)
);

A2O1A1Ixp33_ASAP7_75t_L g434 ( 
.A1(n_416),
.A2(n_371),
.B(n_269),
.C(n_266),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_427),
.B(n_422),
.Y(n_438)
);

OAI21x1_ASAP7_75t_L g440 ( 
.A1(n_438),
.A2(n_439),
.B(n_426),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_432),
.B(n_418),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_440),
.B(n_441),
.C(n_437),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_436),
.A2(n_428),
.B1(n_425),
.B2(n_419),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_435),
.B(n_424),
.C(n_420),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_442),
.A2(n_428),
.B(n_437),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_443),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_445),
.B(n_444),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_446),
.A2(n_434),
.B(n_371),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_447),
.B(n_13),
.Y(n_448)
);


endmodule