module fake_jpeg_10448_n_247 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_247);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_247;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_45;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_31),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_8),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_16),
.C(n_28),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_35),
.C(n_29),
.Y(n_61)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_29),
.B(n_22),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_55),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_66),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_74),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVxp33_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_39),
.A2(n_27),
.B1(n_15),
.B2(n_24),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_64),
.A2(n_72),
.B1(n_73),
.B2(n_24),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_44),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_36),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_17),
.B1(n_27),
.B2(n_25),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_25),
.B1(n_27),
.B2(n_17),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_28),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_18),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_18),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_68),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_83),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_79),
.B(n_81),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_64),
.A2(n_17),
.B1(n_51),
.B2(n_15),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_89),
.B1(n_91),
.B2(n_65),
.Y(n_99)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_65),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_87),
.Y(n_100)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_47),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

OAI32xp33_ASAP7_75t_L g91 ( 
.A1(n_66),
.A2(n_61),
.A3(n_73),
.B1(n_60),
.B2(n_28),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_92),
.A2(n_70),
.B(n_69),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_30),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_38),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_62),
.Y(n_94)
);

INVxp33_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

BUFx12_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_85),
.B(n_57),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_103),
.B(n_81),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_99),
.B(n_107),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_76),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_109),
.Y(n_117)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_0),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_70),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_65),
.B1(n_59),
.B2(n_51),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_63),
.B1(n_19),
.B2(n_28),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_69),
.B1(n_36),
.B2(n_40),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_108),
.A2(n_112),
.B1(n_82),
.B2(n_94),
.Y(n_125)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_36),
.B1(n_40),
.B2(n_47),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_93),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_79),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_88),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_118),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_34),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_91),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_90),
.B1(n_86),
.B2(n_84),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_119),
.A2(n_133),
.B1(n_104),
.B2(n_97),
.Y(n_144)
);

NAND3xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_57),
.C(n_83),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_122),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_23),
.B(n_14),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_121),
.A2(n_125),
.B(n_106),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_100),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_124),
.B(n_128),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_30),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_129),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_68),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_109),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_108),
.A2(n_63),
.B1(n_62),
.B2(n_19),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_131),
.A2(n_112),
.B1(n_114),
.B2(n_101),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_14),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_23),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_145),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_96),
.Y(n_140)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_142),
.A2(n_150),
.B1(n_154),
.B2(n_32),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_103),
.Y(n_143)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_144),
.Y(n_170)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_121),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_148),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_96),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_123),
.A2(n_104),
.B1(n_97),
.B2(n_107),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_151),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_123),
.A2(n_129),
.B(n_125),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_32),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_133),
.A2(n_95),
.B1(n_96),
.B2(n_56),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_153),
.A2(n_26),
.B1(n_21),
.B2(n_34),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_118),
.A2(n_95),
.B1(n_32),
.B2(n_45),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_127),
.C(n_116),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_157),
.C(n_161),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_155),
.B(n_115),
.C(n_131),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_138),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_167),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_126),
.C(n_32),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_135),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_160),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_147),
.Y(n_167)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_144),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_169),
.B(n_151),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_32),
.C(n_45),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_174),
.C(n_154),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_135),
.B(n_32),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_190),
.Y(n_201)
);

FAx1_ASAP7_75t_SL g176 ( 
.A(n_164),
.B(n_143),
.CI(n_136),
.CON(n_176),
.SN(n_176)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_10),
.Y(n_200)
);

NAND3xp33_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_137),
.C(n_146),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_182),
.Y(n_196)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_179),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_180),
.B(n_161),
.C(n_172),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_158),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_160),
.A2(n_152),
.B1(n_145),
.B2(n_150),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_183),
.A2(n_187),
.B1(n_170),
.B2(n_165),
.Y(n_191)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_162),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_185),
.Y(n_198)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_166),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_173),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_188),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_142),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_141),
.C(n_153),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_174),
.B(n_141),
.Y(n_190)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_193),
.C(n_197),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_157),
.C(n_163),
.Y(n_193)
);

MAJx2_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_175),
.C(n_189),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_194),
.B(n_26),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_186),
.A2(n_171),
.B1(n_168),
.B2(n_26),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_199),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_200),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_180),
.C(n_190),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_181),
.C(n_45),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_10),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_203),
.B(n_176),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_206),
.B(n_210),
.Y(n_221)
);

NOR2xp67_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_188),
.Y(n_207)
);

NOR2xp67_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_194),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_216),
.C(n_205),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_9),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_198),
.B(n_195),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_201),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_9),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_214),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_21),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_38),
.C(n_26),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_195),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_217),
.B(n_220),
.Y(n_232)
);

NOR2xp67_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_216),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_201),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_222),
.B(n_223),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_208),
.A2(n_8),
.B(n_13),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_225),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_38),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_6),
.C(n_12),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_4),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_219),
.A2(n_209),
.B1(n_21),
.B2(n_6),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_228),
.B(n_230),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_217),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_223),
.C(n_225),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_232),
.B(n_221),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_235),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_230),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_231),
.C(n_233),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_237),
.A2(n_4),
.B1(n_5),
.B2(n_11),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_13),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_241),
.B(n_238),
.Y(n_242)
);

OAI321xp33_ASAP7_75t_L g244 ( 
.A1(n_242),
.A2(n_243),
.A3(n_240),
.B1(n_4),
.B2(n_5),
.C(n_11),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_244),
.B(n_12),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_245),
.B(n_1),
.C(n_2),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_246),
.A2(n_1),
.B(n_2),
.Y(n_247)
);


endmodule