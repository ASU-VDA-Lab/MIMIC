module fake_jpeg_12408_n_564 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_564);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_564;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_18),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_12),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_55),
.Y(n_129)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_56),
.Y(n_127)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_57),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_58),
.Y(n_124)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_59),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_61),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_21),
.B(n_7),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_62),
.B(n_93),
.Y(n_117)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_21),
.B(n_7),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_64),
.B(n_89),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_27),
.B(n_8),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_65),
.B(n_87),
.Y(n_142)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_67),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_34),
.Y(n_68)
);

INVxp67_ASAP7_75t_SL g115 ( 
.A(n_68),
.Y(n_115)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_69),
.Y(n_141)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_71),
.Y(n_145)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_72),
.Y(n_143)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_74),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_76),
.Y(n_148)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_77),
.Y(n_144)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_79),
.Y(n_160)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_81),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_82),
.Y(n_163)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_38),
.Y(n_86)
);

INVx13_ASAP7_75t_L g171 ( 
.A(n_86),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_27),
.B(n_8),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_8),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx6_ASAP7_75t_SL g120 ( 
.A(n_92),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_42),
.B(n_8),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_94),
.Y(n_140)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_95),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_96),
.Y(n_167)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_42),
.B(n_6),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_99),
.B(n_108),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_40),
.Y(n_100)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_100),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_40),
.Y(n_102)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_45),
.Y(n_104)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_104),
.Y(n_150)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_105),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_106),
.Y(n_166)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_26),
.Y(n_107)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_107),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_52),
.B(n_6),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_78),
.A2(n_49),
.B1(n_41),
.B2(n_26),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_116),
.A2(n_125),
.B1(n_134),
.B2(n_136),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_68),
.A2(n_49),
.B1(n_41),
.B2(n_26),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_57),
.A2(n_49),
.B1(n_43),
.B2(n_41),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_63),
.A2(n_43),
.B1(n_41),
.B2(n_47),
.Y(n_136)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_72),
.Y(n_149)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_95),
.A2(n_43),
.B1(n_50),
.B2(n_47),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_151),
.A2(n_172),
.B1(n_45),
.B2(n_50),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_89),
.B(n_52),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_155),
.B(n_159),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_84),
.B(n_35),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_156),
.B(n_162),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_54),
.B(n_35),
.Y(n_159)
);

HAxp5_ASAP7_75t_SL g161 ( 
.A(n_59),
.B(n_24),
.CON(n_161),
.SN(n_161)
);

AOI21xp33_ASAP7_75t_L g215 ( 
.A1(n_161),
.A2(n_44),
.B(n_53),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_107),
.B(n_35),
.Y(n_162)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_102),
.Y(n_165)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

AOI21xp33_ASAP7_75t_L g170 ( 
.A1(n_92),
.A2(n_28),
.B(n_24),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_170),
.B(n_36),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_61),
.A2(n_43),
.B1(n_50),
.B2(n_47),
.Y(n_172)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_74),
.Y(n_174)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_174),
.Y(n_214)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_79),
.Y(n_175)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_175),
.Y(n_205)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_176),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_122),
.B(n_86),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_177),
.B(n_202),
.C(n_212),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_120),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_178),
.B(n_198),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_142),
.B(n_24),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_179),
.B(n_187),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_171),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_180),
.B(n_203),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_121),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_181),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_182),
.Y(n_245)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_184),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_137),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_185),
.Y(n_292)
);

BUFx12f_ASAP7_75t_L g186 ( 
.A(n_114),
.Y(n_186)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_186),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_131),
.B(n_28),
.Y(n_187)
);

AOI32xp33_ASAP7_75t_L g188 ( 
.A1(n_117),
.A2(n_54),
.A3(n_60),
.B1(n_103),
.B2(n_91),
.Y(n_188)
);

FAx1_ASAP7_75t_SL g251 ( 
.A(n_188),
.B(n_172),
.CI(n_151),
.CON(n_251),
.SN(n_251)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_139),
.Y(n_189)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_189),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_132),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_190),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_115),
.A2(n_37),
.B1(n_53),
.B2(n_19),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_191),
.Y(n_293)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_133),
.Y(n_192)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_192),
.Y(n_266)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_135),
.Y(n_193)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_193),
.Y(n_271)
);

NAND2xp33_ASAP7_75t_SL g195 ( 
.A(n_145),
.B(n_36),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_195),
.A2(n_215),
.B(n_19),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_129),
.Y(n_196)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_196),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_115),
.A2(n_37),
.B1(n_53),
.B2(n_19),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_197),
.A2(n_125),
.B1(n_116),
.B2(n_130),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_154),
.B(n_28),
.Y(n_198)
);

BUFx2_ASAP7_75t_SL g199 ( 
.A(n_171),
.Y(n_199)
);

INVx4_ASAP7_75t_SL g278 ( 
.A(n_199),
.Y(n_278)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_152),
.Y(n_200)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_200),
.Y(n_268)
);

AO22x1_ASAP7_75t_L g295 ( 
.A1(n_201),
.A2(n_227),
.B1(n_1),
.B2(n_2),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_148),
.B(n_36),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_126),
.B(n_44),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_168),
.Y(n_206)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_206),
.Y(n_250)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_207),
.Y(n_265)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_113),
.Y(n_209)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_209),
.Y(n_269)
);

AND2x2_ASAP7_75t_SL g210 ( 
.A(n_109),
.B(n_0),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_210),
.B(n_211),
.Y(n_263)
);

AND2x2_ASAP7_75t_SL g211 ( 
.A(n_112),
.B(n_0),
.Y(n_211)
);

AND2x2_ASAP7_75t_SL g212 ( 
.A(n_118),
.B(n_0),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_134),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_216),
.B(n_220),
.Y(n_255)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_166),
.Y(n_217)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_217),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_119),
.B(n_0),
.Y(n_218)
);

OAI21xp33_ASAP7_75t_L g257 ( 
.A1(n_218),
.A2(n_225),
.B(n_23),
.Y(n_257)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_153),
.Y(n_219)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_219),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_141),
.B(n_44),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_158),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_221),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_127),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_222),
.B(n_232),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_113),
.Y(n_223)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_223),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_144),
.B(n_37),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_224),
.B(n_230),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_111),
.B(n_143),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_164),
.Y(n_226)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_226),
.Y(n_260)
);

A2O1A1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_161),
.A2(n_29),
.B(n_23),
.C(n_22),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_157),
.Y(n_228)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_228),
.Y(n_288)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_138),
.Y(n_229)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_229),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_157),
.B(n_29),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_147),
.Y(n_231)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_231),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_127),
.B(n_29),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_124),
.Y(n_233)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_233),
.Y(n_272)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_147),
.Y(n_234)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_234),
.Y(n_277)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_110),
.Y(n_235)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_235),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_236),
.A2(n_123),
.B1(n_167),
.B2(n_140),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_173),
.B(n_23),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_22),
.Y(n_262)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_158),
.Y(n_238)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_238),
.Y(n_282)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_110),
.Y(n_239)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_239),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_202),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_243),
.B(n_284),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_208),
.B(n_123),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_246),
.B(n_212),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_R g335 ( 
.A(n_247),
.B(n_2),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_249),
.A2(n_259),
.B1(n_238),
.B2(n_200),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_251),
.B(n_257),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_252),
.A2(n_264),
.B1(n_283),
.B2(n_163),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_213),
.A2(n_167),
.B1(n_140),
.B2(n_128),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_262),
.B(n_276),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_227),
.A2(n_136),
.B1(n_82),
.B2(n_98),
.Y(n_264)
);

FAx1_ASAP7_75t_SL g274 ( 
.A(n_195),
.B(n_1),
.CI(n_2),
.CON(n_274),
.SN(n_274)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_274),
.B(n_1),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_194),
.B(n_183),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_210),
.A2(n_100),
.B1(n_88),
.B2(n_90),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_202),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_177),
.A2(n_225),
.B1(n_128),
.B2(n_160),
.Y(n_285)
);

AO21x2_ASAP7_75t_L g310 ( 
.A1(n_285),
.A2(n_290),
.B(n_205),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_177),
.A2(n_163),
.B1(n_160),
.B2(n_106),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_204),
.B(n_22),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_291),
.B(n_46),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_295),
.A2(n_218),
.B(n_189),
.Y(n_308)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_270),
.Y(n_296)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_296),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_293),
.A2(n_225),
.B(n_233),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_297),
.A2(n_326),
.B(n_329),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_275),
.Y(n_298)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_298),
.Y(n_380)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_277),
.Y(n_300)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_300),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_211),
.C(n_212),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_301),
.B(n_320),
.C(n_336),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_303),
.B(n_313),
.Y(n_351)
);

O2A1O1Ixp33_ASAP7_75t_L g304 ( 
.A1(n_293),
.A2(n_210),
.B(n_211),
.C(n_218),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_304),
.A2(n_311),
.B(n_337),
.Y(n_356)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_288),
.Y(n_305)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_305),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_255),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_306),
.B(n_308),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_245),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_307),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_309),
.B(n_319),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_L g373 ( 
.A1(n_310),
.A2(n_318),
.B1(n_334),
.B2(n_287),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_247),
.A2(n_181),
.B(n_196),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_245),
.Y(n_312)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_312),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_267),
.B(n_176),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_288),
.Y(n_314)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_314),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_316),
.A2(n_323),
.B1(n_328),
.B2(n_332),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_317),
.A2(n_269),
.B1(n_286),
.B2(n_265),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_L g318 ( 
.A1(n_264),
.A2(n_223),
.B1(n_229),
.B2(n_207),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_246),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_281),
.B(n_219),
.C(n_192),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_294),
.Y(n_321)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_321),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_263),
.B(n_217),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_322),
.B(n_324),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_259),
.A2(n_228),
.B1(n_234),
.B2(n_231),
.Y(n_323)
);

OAI32xp33_ASAP7_75t_L g324 ( 
.A1(n_295),
.A2(n_214),
.A3(n_185),
.B1(n_104),
.B2(n_101),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_263),
.B(n_184),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_325),
.B(n_331),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_263),
.A2(n_222),
.B(n_193),
.Y(n_326)
);

AOI21xp33_ASAP7_75t_L g327 ( 
.A1(n_254),
.A2(n_186),
.B(n_209),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_327),
.A2(n_335),
.B(n_278),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_249),
.A2(n_96),
.B1(n_94),
.B2(n_85),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_261),
.A2(n_239),
.B(n_186),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_278),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_330),
.B(n_341),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_274),
.B(n_221),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_251),
.A2(n_182),
.B1(n_50),
.B2(n_47),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_271),
.Y(n_333)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_333),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_251),
.A2(n_46),
.B1(n_3),
.B2(n_4),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_257),
.B(n_244),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_274),
.A2(n_3),
.B(n_4),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_283),
.A2(n_46),
.B1(n_5),
.B2(n_9),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_338),
.A2(n_266),
.B1(n_275),
.B2(n_292),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_280),
.B(n_4),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_339),
.B(n_342),
.Y(n_379)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_253),
.Y(n_340)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_340),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_248),
.B(n_46),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_260),
.B(n_5),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_343),
.B(n_266),
.Y(n_370)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_253),
.Y(n_344)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_344),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_317),
.A2(n_282),
.B1(n_268),
.B2(n_242),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_346),
.A2(n_347),
.B1(n_348),
.B2(n_358),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_319),
.A2(n_268),
.B1(n_269),
.B2(n_271),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_336),
.B(n_250),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_349),
.B(n_352),
.C(n_330),
.Y(n_408)
);

MAJx2_ASAP7_75t_L g352 ( 
.A(n_301),
.B(n_272),
.C(n_265),
.Y(n_352)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_315),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_353),
.B(n_382),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_310),
.A2(n_258),
.B1(n_286),
.B2(n_240),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_339),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_360),
.B(n_367),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_362),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_335),
.A2(n_241),
.B(n_289),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_363),
.A2(n_368),
.B(n_326),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_310),
.A2(n_258),
.B1(n_240),
.B2(n_289),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_366),
.A2(n_385),
.B1(n_316),
.B2(n_323),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_329),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_299),
.A2(n_279),
.B(n_273),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_370),
.B(n_371),
.Y(n_418)
);

BUFx5_ASAP7_75t_L g371 ( 
.A(n_321),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_372),
.A2(n_373),
.B1(n_310),
.B2(n_311),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_313),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_375),
.B(n_305),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_306),
.B(n_273),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_310),
.A2(n_279),
.B1(n_287),
.B2(n_292),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_386),
.B(n_320),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_387),
.B(n_403),
.C(n_405),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_354),
.A2(n_299),
.B(n_297),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_388),
.A2(n_398),
.B(n_400),
.Y(n_429)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_376),
.Y(n_390)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_390),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_L g437 ( 
.A1(n_391),
.A2(n_419),
.B1(n_374),
.B2(n_383),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_382),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_392),
.B(n_415),
.Y(n_451)
);

AO22x1_ASAP7_75t_L g393 ( 
.A1(n_356),
.A2(n_361),
.B1(n_365),
.B2(n_355),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_393),
.A2(n_394),
.B(n_395),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_367),
.A2(n_299),
.B1(n_334),
.B2(n_332),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_354),
.A2(n_308),
.B(n_331),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_396),
.B(n_420),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_361),
.A2(n_310),
.B1(n_303),
.B2(n_322),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_397),
.A2(n_366),
.B1(n_350),
.B2(n_368),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_378),
.B(n_325),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_376),
.Y(n_399)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_399),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_355),
.A2(n_337),
.B(n_304),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_345),
.Y(n_401)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_401),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_386),
.B(n_342),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_360),
.B(n_375),
.Y(n_404)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_404),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_349),
.B(n_351),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_352),
.B(n_302),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_406),
.B(n_423),
.C(n_374),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_407),
.A2(n_409),
.B1(n_417),
.B2(n_359),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_408),
.B(n_357),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_346),
.A2(n_328),
.B1(n_338),
.B2(n_324),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_351),
.B(n_296),
.Y(n_411)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_411),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_378),
.B(n_379),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_412),
.B(n_413),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_379),
.B(n_300),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_365),
.B(n_314),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_414),
.B(n_416),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_347),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_345),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_348),
.A2(n_309),
.B1(n_312),
.B2(n_307),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_353),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_377),
.B(n_333),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_421),
.B(n_371),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_352),
.B(n_340),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_409),
.A2(n_359),
.B1(n_356),
.B2(n_372),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_426),
.A2(n_431),
.B1(n_434),
.B2(n_393),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_422),
.A2(n_362),
.B1(n_385),
.B2(n_358),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_428),
.A2(n_430),
.B1(n_437),
.B2(n_439),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_387),
.B(n_406),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_433),
.B(n_435),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_394),
.A2(n_377),
.B1(n_370),
.B2(n_350),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_408),
.B(n_363),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_436),
.B(n_393),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_403),
.B(n_383),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_438),
.B(n_448),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_391),
.A2(n_357),
.B1(n_364),
.B2(n_381),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_397),
.A2(n_422),
.B1(n_404),
.B2(n_414),
.Y(n_440)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_440),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_398),
.A2(n_369),
.B1(n_380),
.B2(n_381),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_445),
.A2(n_396),
.B(n_410),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_446),
.B(n_453),
.C(n_454),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_405),
.B(n_384),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_449),
.B(n_452),
.Y(n_474)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_418),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_423),
.B(n_384),
.C(n_344),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_412),
.B(n_364),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_407),
.A2(n_380),
.B1(n_312),
.B2(n_307),
.Y(n_455)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_455),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_442),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_456),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_458),
.B(n_477),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_461),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_432),
.B(n_398),
.C(n_411),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_462),
.B(n_463),
.C(n_467),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_432),
.B(n_395),
.C(n_400),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_434),
.B(n_438),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_465),
.B(n_475),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_429),
.A2(n_388),
.B(n_402),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_466),
.A2(n_445),
.B(n_439),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_433),
.B(n_413),
.C(n_402),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_442),
.Y(n_468)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_468),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_469),
.A2(n_479),
.B1(n_481),
.B2(n_425),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_441),
.B(n_416),
.Y(n_470)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_470),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_446),
.B(n_453),
.C(n_448),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_473),
.B(n_457),
.C(n_471),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_443),
.B(n_401),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_441),
.B(n_390),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_476),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_424),
.B(n_417),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_424),
.B(n_389),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_478),
.B(n_482),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_426),
.A2(n_389),
.B1(n_298),
.B2(n_256),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_435),
.B(n_256),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_480),
.B(n_9),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_444),
.A2(n_5),
.B1(n_9),
.B2(n_10),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_451),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_SL g483 ( 
.A(n_458),
.B(n_436),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_SL g512 ( 
.A(n_483),
.B(n_488),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_460),
.A2(n_444),
.B1(n_454),
.B2(n_440),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_484),
.B(n_501),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_463),
.A2(n_447),
.B1(n_429),
.B2(n_428),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_485),
.B(n_461),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_487),
.A2(n_490),
.B(n_464),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_SL g488 ( 
.A(n_471),
.B(n_447),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_466),
.A2(n_430),
.B(n_450),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_491),
.A2(n_502),
.B1(n_468),
.B2(n_464),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_462),
.B(n_427),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_497),
.B(n_486),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_499),
.B(n_481),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_500),
.B(n_504),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_473),
.B(n_10),
.C(n_11),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_469),
.A2(n_10),
.B1(n_15),
.B2(n_16),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_457),
.B(n_10),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_SL g522 ( 
.A(n_504),
.B(n_470),
.Y(n_522)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_505),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_494),
.B(n_480),
.C(n_472),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_507),
.B(n_509),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_508),
.B(n_519),
.Y(n_532)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_493),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_492),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_510),
.B(n_515),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_511),
.B(n_514),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_486),
.A2(n_459),
.B1(n_478),
.B2(n_477),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_513),
.B(n_521),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_488),
.B(n_472),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_492),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_498),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_516),
.B(n_517),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_494),
.B(n_467),
.C(n_459),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_518),
.B(n_522),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_500),
.B(n_479),
.C(n_456),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_520),
.B(n_496),
.C(n_484),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_520),
.A2(n_485),
.B(n_503),
.Y(n_523)
);

OAI21x1_ASAP7_75t_L g541 ( 
.A1(n_523),
.A2(n_529),
.B(n_512),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_524),
.B(n_531),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_517),
.B(n_496),
.Y(n_526)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_526),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_506),
.Y(n_528)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_528),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_518),
.A2(n_474),
.B(n_490),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_507),
.B(n_483),
.C(n_487),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_514),
.B(n_491),
.C(n_498),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_535),
.B(n_511),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_530),
.B(n_505),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_538),
.B(n_539),
.Y(n_552)
);

NAND3xp33_ASAP7_75t_L g539 ( 
.A(n_536),
.B(n_476),
.C(n_489),
.Y(n_539)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_541),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_527),
.A2(n_513),
.B1(n_495),
.B2(n_522),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_542),
.B(n_546),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_544),
.B(n_532),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_526),
.B(n_512),
.C(n_499),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_535),
.A2(n_534),
.B1(n_502),
.B2(n_524),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_547),
.A2(n_537),
.B1(n_534),
.B2(n_533),
.Y(n_553)
);

NOR2x1_ASAP7_75t_L g550 ( 
.A(n_540),
.B(n_531),
.Y(n_550)
);

AOI21xp5_ASAP7_75t_SL g554 ( 
.A1(n_550),
.A2(n_543),
.B(n_537),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_551),
.B(n_553),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_L g558 ( 
.A1(n_554),
.A2(n_556),
.B(n_557),
.Y(n_558)
);

INVxp33_ASAP7_75t_L g556 ( 
.A(n_551),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_549),
.B(n_545),
.Y(n_557)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_555),
.A2(n_552),
.B(n_548),
.Y(n_559)
);

AOI321xp33_ASAP7_75t_L g560 ( 
.A1(n_559),
.A2(n_548),
.A3(n_547),
.B1(n_539),
.B2(n_546),
.C(n_525),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_L g561 ( 
.A1(n_560),
.A2(n_558),
.B(n_501),
.Y(n_561)
);

AO21x2_ASAP7_75t_L g562 ( 
.A1(n_561),
.A2(n_15),
.B(n_16),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_562),
.A2(n_16),
.B1(n_18),
.B2(n_489),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_563),
.B(n_18),
.Y(n_564)
);


endmodule