module real_aes_7162_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g167 ( .A1(n_0), .A2(n_168), .B(n_171), .C(n_175), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_1), .B(n_159), .Y(n_178) );
INVx1_ASAP7_75t_L g110 ( .A(n_2), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_3), .B(n_169), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_4), .A2(n_128), .B(n_471), .Y(n_470) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_5), .A2(n_133), .B(n_136), .C(n_498), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_6), .A2(n_128), .B(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_7), .B(n_159), .Y(n_477) );
AO21x2_ASAP7_75t_L g235 ( .A1(n_8), .A2(n_161), .B(n_236), .Y(n_235) );
AND2x6_ASAP7_75t_L g133 ( .A(n_9), .B(n_134), .Y(n_133) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_10), .A2(n_133), .B(n_136), .C(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g511 ( .A(n_11), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g111 ( .A(n_12), .B(n_41), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_13), .B(n_174), .Y(n_500) );
INVx1_ASAP7_75t_L g154 ( .A(n_14), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_15), .B(n_169), .Y(n_242) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_16), .A2(n_170), .B(n_531), .C(n_533), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_17), .B(n_159), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_18), .B(n_148), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_L g135 ( .A1(n_19), .A2(n_136), .B(n_139), .C(n_147), .Y(n_135) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_20), .A2(n_173), .B(n_229), .C(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_21), .B(n_174), .Y(n_449) );
AOI222xp33_ASAP7_75t_L g113 ( .A1(n_22), .A2(n_23), .B1(n_114), .B2(n_695), .C1(n_700), .C2(n_701), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_22), .Y(n_700) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_24), .B(n_174), .Y(n_485) );
CKINVDCx16_ASAP7_75t_R g445 ( .A(n_25), .Y(n_445) );
INVx1_ASAP7_75t_L g484 ( .A(n_26), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_27), .A2(n_136), .B(n_147), .C(n_239), .Y(n_238) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_28), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_29), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_30), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g462 ( .A(n_31), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_32), .A2(n_128), .B(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g131 ( .A(n_33), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_L g186 ( .A1(n_34), .A2(n_187), .B(n_188), .C(n_192), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_35), .Y(n_502) );
A2O1A1Ixp33_ASAP7_75t_L g473 ( .A1(n_36), .A2(n_173), .B(n_474), .C(n_476), .Y(n_473) );
INVxp67_ASAP7_75t_L g463 ( .A(n_37), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_38), .B(n_241), .Y(n_240) );
CKINVDCx14_ASAP7_75t_R g472 ( .A(n_39), .Y(n_472) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_40), .A2(n_136), .B(n_147), .C(n_483), .Y(n_482) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_42), .A2(n_175), .B(n_509), .C(n_510), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_43), .B(n_127), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g232 ( .A(n_44), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_45), .B(n_169), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_46), .B(n_128), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_47), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_48), .Y(n_459) );
A2O1A1Ixp33_ASAP7_75t_L g213 ( .A1(n_49), .A2(n_187), .B(n_192), .C(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g172 ( .A(n_50), .Y(n_172) );
INVx1_ASAP7_75t_L g215 ( .A(n_51), .Y(n_215) );
INVx1_ASAP7_75t_L g517 ( .A(n_52), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_53), .B(n_128), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_54), .Y(n_156) );
CKINVDCx14_ASAP7_75t_R g507 ( .A(n_55), .Y(n_507) );
INVx1_ASAP7_75t_L g134 ( .A(n_56), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_57), .B(n_128), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_58), .B(n_159), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_59), .A2(n_146), .B(n_202), .C(n_204), .Y(n_201) );
INVx1_ASAP7_75t_L g153 ( .A(n_60), .Y(n_153) );
INVx1_ASAP7_75t_SL g475 ( .A(n_61), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_62), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_63), .B(n_169), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_64), .B(n_159), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_65), .B(n_170), .Y(n_226) );
INVx1_ASAP7_75t_L g448 ( .A(n_66), .Y(n_448) );
CKINVDCx16_ASAP7_75t_R g165 ( .A(n_67), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_68), .B(n_141), .Y(n_140) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_69), .A2(n_136), .B(n_192), .C(n_255), .Y(n_254) );
CKINVDCx16_ASAP7_75t_R g200 ( .A(n_70), .Y(n_200) );
INVx1_ASAP7_75t_L g103 ( .A(n_71), .Y(n_103) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_72), .A2(n_128), .B(n_506), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_73), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_74), .A2(n_128), .B(n_528), .Y(n_527) );
AOI222xp33_ASAP7_75t_SL g98 ( .A1(n_75), .A2(n_99), .B1(n_112), .B2(n_704), .C1(n_709), .C2(n_716), .Y(n_98) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_75), .A2(n_118), .B1(n_711), .B2(n_712), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_75), .Y(n_712) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_76), .A2(n_127), .B(n_458), .Y(n_457) );
CKINVDCx16_ASAP7_75t_R g481 ( .A(n_77), .Y(n_481) );
INVx1_ASAP7_75t_L g529 ( .A(n_78), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g143 ( .A(n_79), .B(n_144), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_80), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_81), .A2(n_128), .B(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g532 ( .A(n_82), .Y(n_532) );
INVx2_ASAP7_75t_L g151 ( .A(n_83), .Y(n_151) );
INVx1_ASAP7_75t_L g499 ( .A(n_84), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g262 ( .A(n_85), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_86), .B(n_174), .Y(n_227) );
OR2x2_ASAP7_75t_L g107 ( .A(n_87), .B(n_108), .Y(n_107) );
OR2x2_ASAP7_75t_L g117 ( .A(n_87), .B(n_109), .Y(n_117) );
INVx2_ASAP7_75t_L g433 ( .A(n_87), .Y(n_433) );
A2O1A1Ixp33_ASAP7_75t_L g446 ( .A1(n_88), .A2(n_136), .B(n_192), .C(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_89), .B(n_128), .Y(n_185) );
INVx1_ASAP7_75t_L g189 ( .A(n_90), .Y(n_189) );
INVxp67_ASAP7_75t_L g205 ( .A(n_91), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_92), .B(n_161), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_93), .B(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g222 ( .A(n_94), .Y(n_222) );
INVx1_ASAP7_75t_L g256 ( .A(n_95), .Y(n_256) );
INVx2_ASAP7_75t_L g520 ( .A(n_96), .Y(n_520) );
AND2x2_ASAP7_75t_L g217 ( .A(n_97), .B(n_150), .Y(n_217) );
INVx1_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
NAND2xp33_ASAP7_75t_L g100 ( .A(n_101), .B(n_105), .Y(n_100) );
NOR2xp33_ASAP7_75t_SL g101 ( .A(n_102), .B(n_104), .Y(n_101) );
INVx1_ASAP7_75t_SL g708 ( .A(n_102), .Y(n_708) );
INVx1_ASAP7_75t_L g707 ( .A(n_104), .Y(n_707) );
OA21x2_ASAP7_75t_L g717 ( .A1(n_104), .A2(n_708), .B(n_718), .Y(n_717) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
OAI21xp5_ASAP7_75t_L g709 ( .A1(n_106), .A2(n_710), .B(n_713), .Y(n_709) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
HB1xp67_ASAP7_75t_L g715 ( .A(n_107), .Y(n_715) );
BUFx2_ASAP7_75t_L g718 ( .A(n_107), .Y(n_718) );
NOR2x2_ASAP7_75t_L g703 ( .A(n_108), .B(n_433), .Y(n_703) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g432 ( .A(n_109), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
INVxp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
OAI22xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_118), .B1(n_432), .B2(n_434), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g696 ( .A(n_116), .Y(n_696) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g711 ( .A(n_118), .Y(n_711) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI22xp5_ASAP7_75t_SL g695 ( .A1(n_119), .A2(n_696), .B1(n_697), .B2(n_698), .Y(n_695) );
AND2x2_ASAP7_75t_SL g119 ( .A(n_120), .B(n_368), .Y(n_119) );
NOR5xp2_ASAP7_75t_L g120 ( .A(n_121), .B(n_299), .C(n_328), .D(n_348), .E(n_355), .Y(n_120) );
OAI211xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_179), .B(n_243), .C(n_286), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_123), .A2(n_371), .B1(n_373), .B2(n_374), .Y(n_370) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_158), .Y(n_123) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_124), .Y(n_246) );
AND2x4_ASAP7_75t_L g279 ( .A(n_124), .B(n_280), .Y(n_279) );
INVx5_ASAP7_75t_L g297 ( .A(n_124), .Y(n_297) );
AND2x2_ASAP7_75t_L g306 ( .A(n_124), .B(n_298), .Y(n_306) );
AND2x2_ASAP7_75t_L g318 ( .A(n_124), .B(n_183), .Y(n_318) );
AND2x2_ASAP7_75t_L g414 ( .A(n_124), .B(n_282), .Y(n_414) );
OR2x6_ASAP7_75t_L g124 ( .A(n_125), .B(n_155), .Y(n_124) );
AOI21xp5_ASAP7_75t_SL g125 ( .A1(n_126), .A2(n_135), .B(n_148), .Y(n_125) );
BUFx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x4_ASAP7_75t_L g128 ( .A(n_129), .B(n_133), .Y(n_128) );
NAND2x1p5_ASAP7_75t_L g223 ( .A(n_129), .B(n_133), .Y(n_223) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_132), .Y(n_129) );
INVx1_ASAP7_75t_L g146 ( .A(n_130), .Y(n_146) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g137 ( .A(n_131), .Y(n_137) );
INVx1_ASAP7_75t_L g230 ( .A(n_131), .Y(n_230) );
INVx1_ASAP7_75t_L g138 ( .A(n_132), .Y(n_138) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_132), .Y(n_142) );
INVx3_ASAP7_75t_L g170 ( .A(n_132), .Y(n_170) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_132), .Y(n_174) );
INVx1_ASAP7_75t_L g241 ( .A(n_132), .Y(n_241) );
BUFx3_ASAP7_75t_L g147 ( .A(n_133), .Y(n_147) );
INVx4_ASAP7_75t_SL g177 ( .A(n_133), .Y(n_177) );
INVx5_ASAP7_75t_L g166 ( .A(n_136), .Y(n_166) );
AND2x6_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
BUFx3_ASAP7_75t_L g176 ( .A(n_137), .Y(n_176) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_137), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_143), .B(n_145), .Y(n_139) );
INVx2_ASAP7_75t_L g144 ( .A(n_141), .Y(n_144) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx4_ASAP7_75t_L g203 ( .A(n_142), .Y(n_203) );
O2A1O1Ixp33_ASAP7_75t_L g188 ( .A1(n_144), .A2(n_189), .B(n_190), .C(n_191), .Y(n_188) );
O2A1O1Ixp33_ASAP7_75t_L g214 ( .A1(n_144), .A2(n_191), .B(n_215), .C(n_216), .Y(n_214) );
O2A1O1Ixp33_ASAP7_75t_L g447 ( .A1(n_144), .A2(n_448), .B(n_449), .C(n_450), .Y(n_447) );
O2A1O1Ixp5_ASAP7_75t_L g498 ( .A1(n_144), .A2(n_450), .B(n_499), .C(n_500), .Y(n_498) );
O2A1O1Ixp33_ASAP7_75t_L g483 ( .A1(n_145), .A2(n_169), .B(n_484), .C(n_485), .Y(n_483) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_146), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_149), .B(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g157 ( .A(n_150), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_150), .A2(n_185), .B(n_186), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_150), .A2(n_212), .B(n_213), .Y(n_211) );
O2A1O1Ixp33_ASAP7_75t_L g480 ( .A1(n_150), .A2(n_223), .B(n_481), .C(n_482), .Y(n_480) );
OA21x2_ASAP7_75t_L g504 ( .A1(n_150), .A2(n_505), .B(n_512), .Y(n_504) );
AND2x2_ASAP7_75t_SL g150 ( .A(n_151), .B(n_152), .Y(n_150) );
AND2x2_ASAP7_75t_L g162 ( .A(n_151), .B(n_152), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
AO21x2_ASAP7_75t_L g494 ( .A1(n_157), .A2(n_495), .B(n_501), .Y(n_494) );
INVx2_ASAP7_75t_L g280 ( .A(n_158), .Y(n_280) );
AND2x2_ASAP7_75t_L g298 ( .A(n_158), .B(n_252), .Y(n_298) );
AND2x2_ASAP7_75t_L g317 ( .A(n_158), .B(n_251), .Y(n_317) );
AND2x2_ASAP7_75t_L g357 ( .A(n_158), .B(n_297), .Y(n_357) );
OA21x2_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_163), .B(n_178), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_160), .B(n_194), .Y(n_193) );
AO21x2_ASAP7_75t_L g220 ( .A1(n_160), .A2(n_221), .B(n_231), .Y(n_220) );
AO21x2_ASAP7_75t_L g252 ( .A1(n_160), .A2(n_253), .B(n_261), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_160), .B(n_262), .Y(n_261) );
AO21x2_ASAP7_75t_L g443 ( .A1(n_160), .A2(n_444), .B(n_451), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_160), .B(n_487), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_160), .B(n_502), .Y(n_501) );
INVx4_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_161), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_161), .A2(n_237), .B(n_238), .Y(n_236) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g233 ( .A(n_162), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_SL g164 ( .A1(n_165), .A2(n_166), .B(n_167), .C(n_177), .Y(n_164) );
INVx2_ASAP7_75t_L g187 ( .A(n_166), .Y(n_187) );
O2A1O1Ixp33_ASAP7_75t_L g199 ( .A1(n_166), .A2(n_177), .B(n_200), .C(n_201), .Y(n_199) );
O2A1O1Ixp33_ASAP7_75t_SL g458 ( .A1(n_166), .A2(n_177), .B(n_459), .C(n_460), .Y(n_458) );
O2A1O1Ixp33_ASAP7_75t_L g471 ( .A1(n_166), .A2(n_177), .B(n_472), .C(n_473), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_SL g506 ( .A1(n_166), .A2(n_177), .B(n_507), .C(n_508), .Y(n_506) );
O2A1O1Ixp33_ASAP7_75t_SL g516 ( .A1(n_166), .A2(n_177), .B(n_517), .C(n_518), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_SL g528 ( .A1(n_166), .A2(n_177), .B(n_529), .C(n_530), .Y(n_528) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_169), .B(n_205), .Y(n_204) );
OAI22xp33_ASAP7_75t_L g461 ( .A1(n_169), .A2(n_203), .B1(n_462), .B2(n_463), .Y(n_461) );
INVx5_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_170), .B(n_511), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_172), .B(n_173), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_173), .B(n_475), .Y(n_474) );
INVx4_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g509 ( .A(n_174), .Y(n_509) );
INVx2_ASAP7_75t_L g450 ( .A(n_175), .Y(n_450) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_176), .Y(n_191) );
INVx1_ASAP7_75t_L g533 ( .A(n_176), .Y(n_533) );
INVx1_ASAP7_75t_L g192 ( .A(n_177), .Y(n_192) );
INVxp67_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_181), .B(n_207), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AOI322xp5_ASAP7_75t_L g416 ( .A1(n_182), .A2(n_218), .A3(n_271), .B1(n_279), .B2(n_333), .C1(n_417), .C2(n_420), .Y(n_416) );
AND2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_195), .Y(n_182) );
INVx5_ASAP7_75t_L g248 ( .A(n_183), .Y(n_248) );
AND2x2_ASAP7_75t_L g265 ( .A(n_183), .B(n_250), .Y(n_265) );
BUFx2_ASAP7_75t_L g343 ( .A(n_183), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_183), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g420 ( .A(n_183), .B(n_327), .Y(n_420) );
OR2x6_ASAP7_75t_L g183 ( .A(n_184), .B(n_193), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_195), .B(n_209), .Y(n_274) );
INVx1_ASAP7_75t_L g301 ( .A(n_195), .Y(n_301) );
AND2x2_ASAP7_75t_L g314 ( .A(n_195), .B(n_234), .Y(n_314) );
AND2x2_ASAP7_75t_L g415 ( .A(n_195), .B(n_333), .Y(n_415) );
INVx3_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
OR2x2_ASAP7_75t_L g269 ( .A(n_196), .B(n_209), .Y(n_269) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_196), .Y(n_277) );
OR2x2_ASAP7_75t_L g284 ( .A(n_196), .B(n_234), .Y(n_284) );
AND2x2_ASAP7_75t_L g294 ( .A(n_196), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_196), .B(n_220), .Y(n_323) );
INVxp67_ASAP7_75t_L g347 ( .A(n_196), .Y(n_347) );
AND2x2_ASAP7_75t_L g354 ( .A(n_196), .B(n_218), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_196), .B(n_234), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_196), .B(n_219), .Y(n_380) );
OA21x2_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B(n_206), .Y(n_196) );
OA21x2_ASAP7_75t_L g469 ( .A1(n_197), .A2(n_470), .B(n_477), .Y(n_469) );
OA21x2_ASAP7_75t_L g514 ( .A1(n_197), .A2(n_515), .B(n_521), .Y(n_514) );
OA21x2_ASAP7_75t_L g526 ( .A1(n_197), .A2(n_527), .B(n_534), .Y(n_526) );
O2A1O1Ixp33_ASAP7_75t_L g255 ( .A1(n_202), .A2(n_256), .B(n_257), .C(n_258), .Y(n_255) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_203), .B(n_520), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_203), .B(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_218), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_209), .B(n_235), .Y(n_324) );
OR2x2_ASAP7_75t_L g346 ( .A(n_209), .B(n_219), .Y(n_346) );
AND2x2_ASAP7_75t_L g359 ( .A(n_209), .B(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_209), .B(n_314), .Y(n_365) );
OAI211xp5_ASAP7_75t_SL g369 ( .A1(n_209), .A2(n_370), .B(n_375), .C(n_384), .Y(n_369) );
AND2x2_ASAP7_75t_L g430 ( .A(n_209), .B(n_234), .Y(n_430) );
INVx5_ASAP7_75t_SL g209 ( .A(n_210), .Y(n_209) );
OR2x2_ASAP7_75t_L g283 ( .A(n_210), .B(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_210), .B(n_289), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_210), .B(n_278), .Y(n_290) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_210), .Y(n_292) );
OR2x2_ASAP7_75t_L g303 ( .A(n_210), .B(n_219), .Y(n_303) );
AND2x2_ASAP7_75t_SL g308 ( .A(n_210), .B(n_294), .Y(n_308) );
AND2x2_ASAP7_75t_L g333 ( .A(n_210), .B(n_219), .Y(n_333) );
AND2x2_ASAP7_75t_L g353 ( .A(n_210), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g391 ( .A(n_210), .B(n_218), .Y(n_391) );
OR2x2_ASAP7_75t_L g394 ( .A(n_210), .B(n_380), .Y(n_394) );
OR2x6_ASAP7_75t_L g210 ( .A(n_211), .B(n_217), .Y(n_210) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_234), .Y(n_218) );
A2O1A1Ixp33_ASAP7_75t_L g337 ( .A1(n_219), .A2(n_338), .B(n_341), .C(n_347), .Y(n_337) );
INVx5_ASAP7_75t_SL g219 ( .A(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_220), .B(n_234), .Y(n_268) );
AND2x2_ASAP7_75t_L g272 ( .A(n_220), .B(n_235), .Y(n_272) );
OR2x2_ASAP7_75t_L g278 ( .A(n_220), .B(n_234), .Y(n_278) );
OAI21xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_224), .Y(n_221) );
OAI21xp5_ASAP7_75t_L g444 ( .A1(n_223), .A2(n_445), .B(n_446), .Y(n_444) );
OAI21xp5_ASAP7_75t_L g495 ( .A1(n_223), .A2(n_496), .B(n_497), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_228), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_228), .A2(n_240), .B(n_242), .Y(n_239) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx3_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_232), .B(n_233), .Y(n_231) );
INVx2_ASAP7_75t_L g455 ( .A(n_233), .Y(n_455) );
INVx1_ASAP7_75t_SL g295 ( .A(n_234), .Y(n_295) );
OR2x2_ASAP7_75t_L g423 ( .A(n_234), .B(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_263), .B(n_266), .C(n_275), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AOI31xp33_ASAP7_75t_L g348 ( .A1(n_245), .A2(n_349), .A3(n_351), .B(n_352), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_246), .B(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_247), .B(n_279), .Y(n_285) );
AND2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_248), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g305 ( .A(n_248), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g310 ( .A(n_248), .B(n_280), .Y(n_310) );
AND2x2_ASAP7_75t_L g320 ( .A(n_248), .B(n_279), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_248), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g340 ( .A(n_248), .B(n_297), .Y(n_340) );
AND2x2_ASAP7_75t_L g345 ( .A(n_248), .B(n_317), .Y(n_345) );
OR2x2_ASAP7_75t_L g364 ( .A(n_248), .B(n_250), .Y(n_364) );
OR2x2_ASAP7_75t_L g366 ( .A(n_248), .B(n_367), .Y(n_366) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_248), .Y(n_413) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g313 ( .A(n_250), .B(n_280), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_250), .B(n_297), .Y(n_336) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
BUFx2_ASAP7_75t_L g282 ( .A(n_252), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_254), .B(n_260), .Y(n_253) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx3_ASAP7_75t_L g476 ( .A(n_259), .Y(n_476) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g373 ( .A(n_265), .B(n_297), .Y(n_373) );
AOI322xp5_ASAP7_75t_L g375 ( .A1(n_265), .A2(n_279), .A3(n_317), .B1(n_376), .B2(n_377), .C1(n_378), .C2(n_381), .Y(n_375) );
INVx1_ASAP7_75t_L g383 ( .A(n_265), .Y(n_383) );
NAND2xp33_ASAP7_75t_L g266 ( .A(n_267), .B(n_270), .Y(n_266) );
INVx1_ASAP7_75t_SL g377 ( .A(n_267), .Y(n_377) );
OR2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
OR2x2_ASAP7_75t_L g329 ( .A(n_268), .B(n_274), .Y(n_329) );
INVx1_ASAP7_75t_L g360 ( .A(n_268), .Y(n_360) );
INVx2_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
AND2x4_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OAI32xp33_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_279), .A3(n_281), .B1(n_283), .B2(n_285), .Y(n_275) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
AOI21xp33_ASAP7_75t_SL g315 ( .A1(n_278), .A2(n_293), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_SL g330 ( .A(n_279), .Y(n_330) );
AND2x4_ASAP7_75t_L g327 ( .A(n_280), .B(n_297), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_280), .B(n_363), .Y(n_362) );
AOI322xp5_ASAP7_75t_L g392 ( .A1(n_281), .A2(n_308), .A3(n_327), .B1(n_360), .B2(n_393), .C1(n_395), .C2(n_396), .Y(n_392) );
OAI221xp5_ASAP7_75t_L g421 ( .A1(n_281), .A2(n_358), .B1(n_422), .B2(n_423), .C(n_425), .Y(n_421) );
AND2x2_ASAP7_75t_L g309 ( .A(n_282), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_SL g289 ( .A(n_284), .Y(n_289) );
OR2x2_ASAP7_75t_L g361 ( .A(n_284), .B(n_346), .Y(n_361) );
OAI31xp33_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_290), .A3(n_291), .B(n_296), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_287), .A2(n_320), .B1(n_321), .B2(n_325), .Y(n_319) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g332 ( .A(n_289), .B(n_333), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_291), .A2(n_332), .B1(n_385), .B2(n_388), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g374 ( .A(n_294), .B(n_343), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_294), .B(n_333), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_295), .B(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g408 ( .A(n_295), .B(n_346), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_296), .A2(n_391), .B1(n_404), .B2(n_407), .Y(n_403) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
INVx2_ASAP7_75t_L g312 ( .A(n_297), .Y(n_312) );
AND2x2_ASAP7_75t_L g395 ( .A(n_297), .B(n_317), .Y(n_395) );
OR2x2_ASAP7_75t_L g397 ( .A(n_297), .B(n_364), .Y(n_397) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_297), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_298), .B(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_298), .B(n_343), .Y(n_351) );
OAI211xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_304), .B(n_307), .C(n_319), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AOI221xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_309), .B1(n_311), .B2(n_314), .C(n_315), .Y(n_307) );
INVxp67_ASAP7_75t_L g419 ( .A(n_310), .Y(n_419) );
INVx1_ASAP7_75t_L g386 ( .A(n_311), .Y(n_386) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
AND2x2_ASAP7_75t_L g350 ( .A(n_312), .B(n_317), .Y(n_350) );
INVx1_ASAP7_75t_L g367 ( .A(n_313), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_313), .B(n_340), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx1_ASAP7_75t_L g382 ( .A(n_317), .Y(n_382) );
AND2x2_ASAP7_75t_L g388 ( .A(n_317), .B(n_343), .Y(n_388) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
OR2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx1_ASAP7_75t_SL g376 ( .A(n_324), .Y(n_376) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_327), .B(n_363), .Y(n_387) );
OAI221xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_330), .B1(n_331), .B2(n_334), .C(n_337), .Y(n_328) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g424 ( .A(n_333), .Y(n_424) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g342 ( .A(n_336), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_340), .B(n_399), .Y(n_398) );
AOI21xp33_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_344), .B(n_346), .Y(n_341) );
OAI211xp5_ASAP7_75t_SL g389 ( .A1(n_344), .A2(n_390), .B(n_392), .C(n_398), .Y(n_389) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g401 ( .A(n_346), .Y(n_401) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OAI222xp33_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_358), .B1(n_361), .B2(n_362), .C1(n_365), .C2(n_366), .Y(n_355) );
INVx1_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g431 ( .A(n_362), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_363), .B(n_406), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_363), .A2(n_410), .B1(n_412), .B2(n_415), .Y(n_409) );
INVx2_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
NOR4xp25_ASAP7_75t_L g368 ( .A(n_369), .B(n_389), .C(n_402), .D(n_421), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_371), .B(n_401), .Y(n_411) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g378 ( .A(n_376), .B(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_379), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
NAND2xp5_ASAP7_75t_SL g385 ( .A(n_386), .B(n_387), .Y(n_385) );
INVx1_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NAND3xp33_ASAP7_75t_L g402 ( .A(n_403), .B(n_409), .C(n_416), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .Y(n_412) );
INVx2_ASAP7_75t_L g418 ( .A(n_414), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
OAI21xp5_ASAP7_75t_SL g425 ( .A1(n_426), .A2(n_428), .B(n_431), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g699 ( .A(n_432), .Y(n_699) );
INVx2_ASAP7_75t_L g697 ( .A(n_434), .Y(n_697) );
OR2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_629), .Y(n_434) );
NAND5xp2_ASAP7_75t_L g435 ( .A(n_436), .B(n_558), .C(n_588), .D(n_609), .E(n_615), .Y(n_435) );
AOI221xp5_ASAP7_75t_SL g436 ( .A1(n_437), .A2(n_491), .B1(n_522), .B2(n_524), .C(n_535), .Y(n_436) );
INVxp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_439), .B(n_488), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_440), .B(n_466), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
A2O1A1Ixp33_ASAP7_75t_SL g609 ( .A1(n_441), .A2(n_478), .B(n_610), .C(n_613), .Y(n_609) );
AND2x2_ASAP7_75t_L g679 ( .A(n_441), .B(n_479), .Y(n_679) );
AND2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_453), .Y(n_441) );
AND2x2_ASAP7_75t_L g537 ( .A(n_442), .B(n_538), .Y(n_537) );
OR2x2_ASAP7_75t_L g541 ( .A(n_442), .B(n_538), .Y(n_541) );
OR2x2_ASAP7_75t_L g567 ( .A(n_442), .B(n_479), .Y(n_567) );
AND2x2_ASAP7_75t_L g569 ( .A(n_442), .B(n_469), .Y(n_569) );
AND2x2_ASAP7_75t_L g587 ( .A(n_442), .B(n_468), .Y(n_587) );
INVx1_ASAP7_75t_L g620 ( .A(n_442), .Y(n_620) );
INVx2_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
BUFx2_ASAP7_75t_L g490 ( .A(n_443), .Y(n_490) );
AND2x2_ASAP7_75t_L g523 ( .A(n_443), .B(n_469), .Y(n_523) );
AND2x2_ASAP7_75t_L g676 ( .A(n_443), .B(n_479), .Y(n_676) );
AND2x2_ASAP7_75t_L g557 ( .A(n_453), .B(n_467), .Y(n_557) );
OR2x2_ASAP7_75t_L g561 ( .A(n_453), .B(n_479), .Y(n_561) );
AND2x2_ASAP7_75t_L g586 ( .A(n_453), .B(n_587), .Y(n_586) );
INVx1_ASAP7_75t_SL g633 ( .A(n_453), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_453), .B(n_595), .Y(n_681) );
AO21x2_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_456), .B(n_464), .Y(n_453) );
INVx1_ASAP7_75t_L g539 ( .A(n_454), .Y(n_539) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OA21x2_ASAP7_75t_L g538 ( .A1(n_457), .A2(n_465), .B(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
OAI322xp33_ASAP7_75t_L g682 ( .A1(n_466), .A2(n_618), .A3(n_641), .B1(n_662), .B2(n_683), .C1(n_685), .C2(n_686), .Y(n_682) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_467), .B(n_538), .Y(n_685) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_478), .Y(n_467) );
AND2x2_ASAP7_75t_L g489 ( .A(n_468), .B(n_490), .Y(n_489) );
AND2x4_ASAP7_75t_L g554 ( .A(n_468), .B(n_479), .Y(n_554) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g595 ( .A(n_469), .B(n_479), .Y(n_595) );
AND2x2_ASAP7_75t_L g639 ( .A(n_469), .B(n_478), .Y(n_639) );
AND2x2_ASAP7_75t_L g522 ( .A(n_478), .B(n_523), .Y(n_522) );
OR2x2_ASAP7_75t_L g540 ( .A(n_478), .B(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_478), .B(n_569), .Y(n_693) );
INVx3_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g488 ( .A(n_479), .B(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_479), .B(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g607 ( .A(n_479), .B(n_538), .Y(n_607) );
AND2x2_ASAP7_75t_L g634 ( .A(n_479), .B(n_569), .Y(n_634) );
OR2x2_ASAP7_75t_L g690 ( .A(n_479), .B(n_541), .Y(n_690) );
OR2x6_ASAP7_75t_L g479 ( .A(n_480), .B(n_486), .Y(n_479) );
INVx1_ASAP7_75t_SL g576 ( .A(n_488), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_489), .B(n_607), .Y(n_608) );
AND2x2_ASAP7_75t_L g642 ( .A(n_489), .B(n_632), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_489), .B(n_565), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_489), .B(n_687), .Y(n_686) );
OAI31xp33_ASAP7_75t_L g660 ( .A1(n_491), .A2(n_522), .A3(n_661), .B(n_663), .Y(n_660) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_503), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g627 ( .A(n_492), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g643 ( .A(n_492), .B(n_578), .Y(n_643) );
OR2x2_ASAP7_75t_L g650 ( .A(n_492), .B(n_651), .Y(n_650) );
OR2x2_ASAP7_75t_L g662 ( .A(n_492), .B(n_551), .Y(n_662) );
CKINVDCx16_ASAP7_75t_R g492 ( .A(n_493), .Y(n_492) );
OR2x2_ASAP7_75t_L g596 ( .A(n_493), .B(n_597), .Y(n_596) );
BUFx3_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g524 ( .A(n_494), .B(n_525), .Y(n_524) );
INVx4_ASAP7_75t_L g545 ( .A(n_494), .Y(n_545) );
AND2x2_ASAP7_75t_L g582 ( .A(n_494), .B(n_526), .Y(n_582) );
AND2x2_ASAP7_75t_L g581 ( .A(n_503), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_SL g651 ( .A(n_503), .Y(n_651) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_513), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_504), .B(n_545), .Y(n_544) );
OR2x2_ASAP7_75t_L g551 ( .A(n_504), .B(n_514), .Y(n_551) );
INVx2_ASAP7_75t_L g571 ( .A(n_504), .Y(n_571) );
AND2x2_ASAP7_75t_L g585 ( .A(n_504), .B(n_514), .Y(n_585) );
AND2x2_ASAP7_75t_L g592 ( .A(n_504), .B(n_548), .Y(n_592) );
BUFx3_ASAP7_75t_L g602 ( .A(n_504), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_504), .B(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g547 ( .A(n_513), .Y(n_547) );
AND2x2_ASAP7_75t_L g555 ( .A(n_513), .B(n_545), .Y(n_555) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g525 ( .A(n_514), .B(n_526), .Y(n_525) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_514), .Y(n_579) );
INVx2_ASAP7_75t_SL g562 ( .A(n_523), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_523), .B(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_523), .B(n_632), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g655 ( .A(n_524), .B(n_602), .Y(n_655) );
INVx1_ASAP7_75t_SL g689 ( .A(n_524), .Y(n_689) );
INVx1_ASAP7_75t_SL g597 ( .A(n_525), .Y(n_597) );
INVx1_ASAP7_75t_SL g548 ( .A(n_526), .Y(n_548) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_526), .Y(n_559) );
OR2x2_ASAP7_75t_L g570 ( .A(n_526), .B(n_545), .Y(n_570) );
AND2x2_ASAP7_75t_L g584 ( .A(n_526), .B(n_545), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_526), .B(n_574), .Y(n_636) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_540), .B(n_542), .C(n_553), .Y(n_535) );
AOI31xp33_ASAP7_75t_L g652 ( .A1(n_536), .A2(n_653), .A3(n_654), .B(n_655), .Y(n_652) );
AND2x2_ASAP7_75t_L g625 ( .A(n_537), .B(n_554), .Y(n_625) );
BUFx3_ASAP7_75t_L g565 ( .A(n_538), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_538), .B(n_569), .Y(n_568) );
OR2x2_ASAP7_75t_L g601 ( .A(n_538), .B(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_538), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_SL g556 ( .A(n_541), .Y(n_556) );
OAI222xp33_ASAP7_75t_L g665 ( .A1(n_541), .A2(n_666), .B1(n_669), .B2(n_670), .C1(n_671), .C2(n_672), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_543), .B(n_549), .Y(n_542) );
INVx1_ASAP7_75t_L g671 ( .A(n_543), .Y(n_671) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_546), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_545), .B(n_548), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_545), .B(n_571), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_545), .B(n_546), .Y(n_641) );
INVx1_ASAP7_75t_L g692 ( .A(n_545), .Y(n_692) );
NAND2xp5_ASAP7_75t_SL g622 ( .A(n_546), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g694 ( .A(n_546), .Y(n_694) );
AND2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
INVx2_ASAP7_75t_L g574 ( .A(n_547), .Y(n_574) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_548), .Y(n_617) );
AOI32xp33_ASAP7_75t_L g553 ( .A1(n_549), .A2(n_554), .A3(n_555), .B1(n_556), .B2(n_557), .Y(n_553) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_551), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g628 ( .A(n_551), .Y(n_628) );
OR2x2_ASAP7_75t_L g669 ( .A(n_551), .B(n_570), .Y(n_669) );
INVx1_ASAP7_75t_L g605 ( .A(n_552), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_554), .B(n_565), .Y(n_590) );
INVx3_ASAP7_75t_L g599 ( .A(n_554), .Y(n_599) );
AOI322xp5_ASAP7_75t_L g615 ( .A1(n_554), .A2(n_599), .A3(n_616), .B1(n_618), .B2(n_621), .C1(n_625), .C2(n_626), .Y(n_615) );
AND2x2_ASAP7_75t_L g591 ( .A(n_555), .B(n_592), .Y(n_591) );
INVxp67_ASAP7_75t_L g668 ( .A(n_555), .Y(n_668) );
A2O1A1O1Ixp25_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_560), .B(n_563), .C(n_571), .D(n_572), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_559), .B(n_602), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
OAI221xp5_ASAP7_75t_L g572 ( .A1(n_561), .A2(n_573), .B1(n_576), .B2(n_577), .C(n_580), .Y(n_572) );
INVx1_ASAP7_75t_SL g687 ( .A(n_561), .Y(n_687) );
AOI21xp33_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_568), .B(n_570), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g675 ( .A(n_565), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OAI221xp5_ASAP7_75t_SL g657 ( .A1(n_567), .A2(n_651), .B1(n_658), .B2(n_659), .C(n_660), .Y(n_657) );
OAI222xp33_ASAP7_75t_L g688 ( .A1(n_568), .A2(n_689), .B1(n_690), .B2(n_691), .C1(n_693), .C2(n_694), .Y(n_688) );
AND2x2_ASAP7_75t_L g646 ( .A(n_569), .B(n_632), .Y(n_646) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_569), .A2(n_584), .B(n_631), .Y(n_658) );
INVx1_ASAP7_75t_L g672 ( .A(n_569), .Y(n_672) );
INVx2_ASAP7_75t_SL g575 ( .A(n_570), .Y(n_575) );
AND2x2_ASAP7_75t_L g578 ( .A(n_571), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
INVx1_ASAP7_75t_SL g612 ( .A(n_574), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_574), .B(n_584), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_575), .B(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_575), .B(n_585), .Y(n_614) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OAI21xp5_ASAP7_75t_SL g580 ( .A1(n_581), .A2(n_583), .B(n_586), .Y(n_580) );
INVx1_ASAP7_75t_SL g598 ( .A(n_582), .Y(n_598) );
AND2x2_ASAP7_75t_L g645 ( .A(n_582), .B(n_628), .Y(n_645) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
AND2x2_ASAP7_75t_L g684 ( .A(n_584), .B(n_602), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_585), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_SL g670 ( .A(n_586), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_591), .B1(n_593), .B2(n_600), .C(n_603), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_596), .B1(n_598), .B2(n_599), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OAI22xp33_ASAP7_75t_L g603 ( .A1(n_597), .A2(n_604), .B1(n_606), .B2(n_608), .Y(n_603) );
OR2x2_ASAP7_75t_L g674 ( .A(n_598), .B(n_602), .Y(n_674) );
OR2x2_ASAP7_75t_L g677 ( .A(n_598), .B(n_612), .Y(n_677) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OAI221xp5_ASAP7_75t_L g673 ( .A1(n_619), .A2(n_674), .B1(n_675), .B2(n_677), .C(n_678), .Y(n_673) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVxp67_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND3xp33_ASAP7_75t_SL g629 ( .A(n_630), .B(n_644), .C(n_656), .Y(n_629) );
AOI222xp33_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_635), .B1(n_637), .B2(n_640), .C1(n_642), .C2(n_643), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_634), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_632), .B(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g654 ( .A(n_634), .Y(n_654) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVxp67_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_646), .B1(n_647), .B2(n_649), .C(n_652), .Y(n_644) );
INVx1_ASAP7_75t_L g659 ( .A(n_645), .Y(n_659) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
OAI21xp33_ASAP7_75t_L g678 ( .A1(n_649), .A2(n_679), .B(n_680), .Y(n_678) );
INVx1_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
NOR5xp2_ASAP7_75t_L g656 ( .A(n_657), .B(n_665), .C(n_673), .D(n_682), .E(n_688), .Y(n_656) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OR2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
INVxp67_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
INVx3_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g705 ( .A(n_706), .B(n_708), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_717), .Y(n_716) );
endmodule