module fake_jpeg_2872_n_242 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_242);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_242;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_14),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_58),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_2),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_57),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_48),
.Y(n_73)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_29),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_50),
.Y(n_63)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

AOI21xp33_ASAP7_75t_L g67 ( 
.A1(n_56),
.A2(n_59),
.B(n_60),
.Y(n_67)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx24_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_20),
.B(n_15),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_61),
.B(n_20),
.Y(n_82)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_38),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_27),
.B1(n_25),
.B2(n_30),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_65),
.A2(n_69),
.B1(n_85),
.B2(n_47),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_27),
.B1(n_38),
.B2(n_37),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_66),
.A2(n_86),
.B1(n_93),
.B2(n_43),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_45),
.A2(n_25),
.B1(n_30),
.B2(n_22),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_35),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_87),
.Y(n_95)
);

NOR2x1_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_36),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_81),
.B(n_82),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_41),
.B(n_37),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_89),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_45),
.A2(n_21),
.B1(n_22),
.B2(n_33),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_62),
.A2(n_32),
.B1(n_38),
.B2(n_37),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_36),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_46),
.B(n_35),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_47),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_32),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_32),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_40),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_53),
.A2(n_34),
.B1(n_33),
.B2(n_21),
.Y(n_93)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_78),
.B(n_84),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_100),
.B(n_113),
.Y(n_127)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

AND2x2_ASAP7_75t_SL g104 ( 
.A(n_78),
.B(n_46),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_104),
.B(n_108),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_109),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_34),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_47),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_114),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_111),
.A2(n_115),
.B1(n_121),
.B2(n_124),
.Y(n_135)
);

AOI32xp33_ASAP7_75t_L g112 ( 
.A1(n_89),
.A2(n_60),
.A3(n_39),
.B1(n_28),
.B2(n_31),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_117),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_46),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_83),
.A2(n_51),
.B1(n_48),
.B2(n_58),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_68),
.B1(n_90),
.B2(n_59),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_15),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_125),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_63),
.B(n_13),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_120),
.Y(n_146)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_83),
.A2(n_49),
.B1(n_60),
.B2(n_19),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_63),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_122),
.B(n_123),
.Y(n_139)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_64),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_100),
.A2(n_66),
.B1(n_86),
.B2(n_67),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_130),
.A2(n_140),
.B1(n_145),
.B2(n_149),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_92),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_137),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_72),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_116),
.A2(n_77),
.B1(n_64),
.B2(n_72),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_73),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_133),
.Y(n_166)
);

NOR3xp33_ASAP7_75t_SL g144 ( 
.A(n_110),
.B(n_80),
.C(n_52),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_144),
.B(n_150),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_114),
.A2(n_68),
.B1(n_54),
.B2(n_56),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_148),
.A2(n_150),
.B1(n_123),
.B2(n_120),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_97),
.A2(n_90),
.B1(n_19),
.B2(n_28),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_114),
.A2(n_39),
.B1(n_28),
.B2(n_80),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_96),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_151),
.B(n_160),
.Y(n_179)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_141),
.Y(n_154)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_110),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_155),
.A2(n_156),
.B(n_157),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_128),
.A2(n_97),
.B(n_104),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_128),
.A2(n_96),
.B(n_122),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_95),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_161),
.A2(n_129),
.B1(n_125),
.B2(n_138),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_104),
.Y(n_162)
);

AOI221xp5_ASAP7_75t_L g189 ( 
.A1(n_162),
.A2(n_136),
.B1(n_102),
.B2(n_106),
.C(n_124),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_139),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_167),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_112),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_165),
.B(n_170),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_172),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_99),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_171),
.C(n_129),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_169),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_142),
.B(n_108),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_103),
.C(n_98),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_165),
.A2(n_132),
.B1(n_143),
.B2(n_130),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_176),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_164),
.A2(n_132),
.B1(n_135),
.B2(n_140),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_148),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_188),
.C(n_171),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_169),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_2),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_159),
.A2(n_149),
.B1(n_144),
.B2(n_141),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_182),
.A2(n_186),
.B1(n_155),
.B2(n_159),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_106),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_189),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_174),
.A2(n_156),
.B(n_157),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_191),
.A2(n_187),
.B(n_39),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_195),
.C(n_200),
.Y(n_213)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_180),
.Y(n_194)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_162),
.C(n_166),
.Y(n_195)
);

AOI221xp5_ASAP7_75t_L g196 ( 
.A1(n_184),
.A2(n_170),
.B1(n_163),
.B2(n_155),
.C(n_162),
.Y(n_196)
);

AOI321xp33_ASAP7_75t_L g208 ( 
.A1(n_196),
.A2(n_173),
.A3(n_185),
.B1(n_190),
.B2(n_181),
.C(n_179),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_197),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_183),
.A2(n_168),
.B1(n_172),
.B2(n_158),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_199),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_186),
.A2(n_153),
.B1(n_152),
.B2(n_161),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_136),
.C(n_154),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_180),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_202),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_101),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_205),
.Y(n_211)
);

AOI31xp67_ASAP7_75t_L g222 ( 
.A1(n_208),
.A2(n_209),
.A3(n_210),
.B(n_214),
.Y(n_222)
);

AOI321xp33_ASAP7_75t_L g209 ( 
.A1(n_191),
.A2(n_190),
.A3(n_181),
.B1(n_173),
.B2(n_177),
.C(n_176),
.Y(n_209)
);

AOI321xp33_ASAP7_75t_L g214 ( 
.A1(n_195),
.A2(n_187),
.A3(n_39),
.B1(n_28),
.B2(n_5),
.C(n_6),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_2),
.Y(n_215)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_215),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_212),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_206),
.A2(n_193),
.B(n_203),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_217),
.A2(n_220),
.B1(n_224),
.B2(n_3),
.Y(n_227)
);

AOI21x1_ASAP7_75t_SL g218 ( 
.A1(n_208),
.A2(n_203),
.B(n_193),
.Y(n_218)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_218),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_207),
.A2(n_204),
.B(n_211),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_3),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_202),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_213),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_214),
.A2(n_192),
.B1(n_4),
.B2(n_8),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_213),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_227),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_229),
.Y(n_233)
);

NOR3xp33_ASAP7_75t_SL g230 ( 
.A(n_222),
.B(n_8),
.C(n_10),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_10),
.Y(n_235)
);

OAI21xp33_ASAP7_75t_L g232 ( 
.A1(n_225),
.A2(n_218),
.B(n_223),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_232),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_226),
.A2(n_8),
.B(n_10),
.Y(n_234)
);

OAI221xp5_ASAP7_75t_L g236 ( 
.A1(n_234),
.A2(n_230),
.B1(n_229),
.B2(n_12),
.C(n_11),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_235),
.A2(n_231),
.B1(n_233),
.B2(n_232),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_236),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_237),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_240),
.B(n_238),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_241),
.B(n_239),
.Y(n_242)
);


endmodule