module fake_jpeg_24469_n_221 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_221);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_221;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_43),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_0),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_0),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_1),
.Y(n_51)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_19),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_17),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_31),
.B1(n_27),
.B2(n_30),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_65),
.B1(n_67),
.B2(n_72),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_49),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_64),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_57),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_33),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_59),
.Y(n_74)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_1),
.Y(n_58)
);

OAI21xp33_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_66),
.B(n_2),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_31),
.C(n_17),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_61),
.Y(n_83)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_70),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_26),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_68),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_35),
.A2(n_32),
.B1(n_28),
.B2(n_23),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_35),
.A2(n_26),
.B(n_18),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_34),
.A2(n_30),
.B1(n_27),
.B2(n_20),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_36),
.B(n_26),
.Y(n_68)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_29),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_43),
.A2(n_23),
.B1(n_28),
.B2(n_19),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_22),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_78),
.Y(n_103)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_77),
.B(n_88),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_22),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_51),
.A2(n_22),
.B1(n_21),
.B2(n_18),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_79),
.A2(n_91),
.B1(n_95),
.B2(n_101),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_2),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_82),
.A2(n_85),
.B(n_87),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_21),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_96),
.Y(n_119)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g116 ( 
.A(n_86),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_3),
.Y(n_87)
);

NOR2x1_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_3),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_89),
.Y(n_117)
);

A2O1A1O1Ixp25_ASAP7_75t_L g90 ( 
.A1(n_65),
.A2(n_21),
.B(n_18),
.C(n_16),
.D(n_29),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_97),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_66),
.A2(n_16),
.B1(n_29),
.B2(n_6),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_59),
.B(n_50),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_93),
.B(n_100),
.Y(n_105)
);

AO22x2_ASAP7_75t_L g95 ( 
.A1(n_58),
.A2(n_16),
.B1(n_29),
.B2(n_6),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_4),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_54),
.B(n_4),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_55),
.B(n_4),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_102),
.Y(n_124)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

NAND3xp33_ASAP7_75t_L g100 ( 
.A(n_54),
.B(n_15),
.C(n_12),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_47),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_8),
.Y(n_102)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_110),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_108),
.Y(n_144)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_91),
.A2(n_55),
.B1(n_47),
.B2(n_57),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_111),
.A2(n_115),
.B1(n_120),
.B2(n_122),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_95),
.A2(n_62),
.B1(n_69),
.B2(n_10),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_97),
.B1(n_87),
.B2(n_82),
.Y(n_140)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_121),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_75),
.A2(n_69),
.B1(n_56),
.B2(n_10),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_84),
.A2(n_69),
.B1(n_56),
.B2(n_9),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_78),
.A2(n_8),
.B1(n_73),
.B2(n_90),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_126),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_81),
.A2(n_8),
.B1(n_74),
.B2(n_76),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_125),
.A2(n_74),
.B1(n_82),
.B2(n_87),
.Y(n_141)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_102),
.Y(n_127)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_81),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_130),
.B(n_135),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_109),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_131),
.Y(n_160)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_136),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_88),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_137),
.A2(n_94),
.B(n_121),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_107),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_139),
.A2(n_143),
.B(n_147),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_140),
.A2(n_106),
.B1(n_97),
.B2(n_108),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_125),
.Y(n_155)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_129),
.A2(n_81),
.B(n_74),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

NAND3xp33_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_152),
.C(n_106),
.Y(n_169)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_154),
.B(n_159),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_134),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_119),
.C(n_117),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_158),
.C(n_162),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_122),
.C(n_123),
.Y(n_158)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_164),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_128),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_132),
.A2(n_128),
.B(n_116),
.Y(n_164)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_165),
.Y(n_178)
);

INVxp67_ASAP7_75t_SL g166 ( 
.A(n_133),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_166),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_169),
.B(n_137),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_167),
.A2(n_151),
.B1(n_136),
.B2(n_149),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_170),
.A2(n_180),
.B1(n_183),
.B2(n_168),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_175),
.C(n_165),
.Y(n_185)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_174),
.B(n_177),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_152),
.C(n_150),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_145),
.Y(n_176)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_176),
.Y(n_188)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_168),
.Y(n_180)
);

NAND3xp33_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_135),
.C(n_163),
.Y(n_190)
);

OAI32xp33_ASAP7_75t_L g183 ( 
.A1(n_164),
.A2(n_132),
.A3(n_134),
.B1(n_145),
.B2(n_146),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_142),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_186),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_191),
.C(n_192),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_176),
.Y(n_186)
);

BUFx12_ASAP7_75t_L g187 ( 
.A(n_177),
.Y(n_187)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_187),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_189),
.A2(n_183),
.B1(n_176),
.B2(n_170),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_190),
.A2(n_139),
.B(n_142),
.Y(n_202)
);

MAJx2_ASAP7_75t_L g191 ( 
.A(n_173),
.B(n_162),
.C(n_159),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_158),
.C(n_160),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_178),
.A2(n_145),
.B1(n_154),
.B2(n_143),
.Y(n_194)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_194),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_187),
.Y(n_197)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_197),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_175),
.C(n_172),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_202),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_188),
.A2(n_171),
.B(n_174),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_200),
.B(n_185),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_201),
.A2(n_184),
.B1(n_193),
.B2(n_191),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_205),
.B(n_209),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_203),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_179),
.C(n_187),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_203),
.A2(n_188),
.B(n_194),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_208),
.A2(n_199),
.B(n_197),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_195),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_210),
.B(n_212),
.Y(n_215)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_211),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_208),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_206),
.Y(n_217)
);

AO21x1_ASAP7_75t_L g219 ( 
.A1(n_217),
.A2(n_218),
.B(n_215),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_214),
.A2(n_207),
.B1(n_205),
.B2(n_131),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_219),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_214),
.Y(n_221)
);


endmodule