module real_aes_8265_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g114 ( .A(n_0), .Y(n_114) );
NAND3xp33_ASAP7_75t_SL g745 ( .A(n_0), .B(n_721), .C(n_746), .Y(n_745) );
AOI22xp5_ASAP7_75t_L g724 ( .A1(n_1), .A2(n_725), .B1(n_726), .B2(n_727), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_1), .Y(n_725) );
A2O1A1Ixp33_ASAP7_75t_L g178 ( .A1(n_2), .A2(n_136), .B(n_141), .C(n_179), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_3), .A2(n_131), .B(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_4), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g482 ( .A(n_5), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_6), .B(n_169), .Y(n_235) );
AOI21xp33_ASAP7_75t_L g490 ( .A1(n_7), .A2(n_131), .B(n_491), .Y(n_490) );
AND2x6_ASAP7_75t_L g136 ( .A(n_8), .B(n_137), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_9), .A2(n_266), .B(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g148 ( .A(n_10), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_11), .B(n_43), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_11), .B(n_744), .Y(n_743) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_12), .B(n_146), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_13), .B(n_193), .Y(n_461) );
INVx1_ASAP7_75t_L g495 ( .A(n_14), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_15), .A2(n_33), .B1(n_728), .B2(n_729), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_15), .Y(n_729) );
INVx1_ASAP7_75t_L g129 ( .A(n_16), .Y(n_129) );
INVx1_ASAP7_75t_L g473 ( .A(n_17), .Y(n_473) );
A2O1A1Ixp33_ASAP7_75t_L g162 ( .A1(n_18), .A2(n_149), .B(n_163), .C(n_167), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_19), .B(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_20), .B(n_452), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g447 ( .A(n_21), .B(n_131), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_22), .B(n_275), .Y(n_274) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_23), .A2(n_193), .B(n_194), .C(n_196), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_24), .B(n_169), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_25), .B(n_146), .Y(n_221) );
A2O1A1Ixp33_ASAP7_75t_L g471 ( .A1(n_26), .A2(n_165), .B(n_167), .C(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_27), .B(n_146), .Y(n_207) );
CKINVDCx16_ASAP7_75t_R g217 ( .A(n_28), .Y(n_217) );
INVx1_ASAP7_75t_L g205 ( .A(n_29), .Y(n_205) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_30), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_31), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_32), .B(n_146), .Y(n_483) );
INVx1_ASAP7_75t_L g728 ( .A(n_33), .Y(n_728) );
INVx1_ASAP7_75t_L g271 ( .A(n_34), .Y(n_271) );
INVx1_ASAP7_75t_L g503 ( .A(n_35), .Y(n_503) );
INVx2_ASAP7_75t_L g134 ( .A(n_36), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_37), .Y(n_186) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_38), .A2(n_193), .B(n_231), .C(n_233), .Y(n_230) );
INVxp67_ASAP7_75t_L g272 ( .A(n_39), .Y(n_272) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_40), .A2(n_141), .B(n_204), .C(n_210), .Y(n_203) );
CKINVDCx14_ASAP7_75t_R g229 ( .A(n_41), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g448 ( .A1(n_42), .A2(n_136), .B(n_141), .C(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g744 ( .A(n_43), .Y(n_744) );
INVx1_ASAP7_75t_L g502 ( .A(n_44), .Y(n_502) );
A2O1A1Ixp33_ASAP7_75t_L g144 ( .A1(n_45), .A2(n_145), .B(n_147), .C(n_150), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_46), .B(n_146), .Y(n_537) );
AOI22xp33_ASAP7_75t_SL g103 ( .A1(n_47), .A2(n_104), .B1(n_739), .B2(n_749), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_48), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g268 ( .A(n_49), .Y(n_268) );
INVx1_ASAP7_75t_L g191 ( .A(n_50), .Y(n_191) );
CKINVDCx16_ASAP7_75t_R g504 ( .A(n_51), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_52), .B(n_131), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g500 ( .A1(n_53), .A2(n_141), .B1(n_196), .B2(n_501), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_54), .Y(n_454) );
CKINVDCx16_ASAP7_75t_R g479 ( .A(n_55), .Y(n_479) );
CKINVDCx14_ASAP7_75t_R g139 ( .A(n_56), .Y(n_139) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_57), .A2(n_145), .B(n_233), .C(n_494), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_58), .Y(n_540) );
INVx1_ASAP7_75t_L g492 ( .A(n_59), .Y(n_492) );
INVx1_ASAP7_75t_L g137 ( .A(n_60), .Y(n_137) );
INVx1_ASAP7_75t_L g128 ( .A(n_61), .Y(n_128) );
INVx1_ASAP7_75t_SL g232 ( .A(n_62), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_63), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_64), .B(n_169), .Y(n_198) );
INVx1_ASAP7_75t_L g220 ( .A(n_65), .Y(n_220) );
A2O1A1Ixp33_ASAP7_75t_SL g511 ( .A1(n_66), .A2(n_233), .B(n_452), .C(n_512), .Y(n_511) );
INVxp67_ASAP7_75t_L g513 ( .A(n_67), .Y(n_513) );
AOI222xp33_ASAP7_75t_L g438 ( .A1(n_68), .A2(n_439), .B1(n_724), .B2(n_730), .C1(n_731), .C2(n_735), .Y(n_438) );
INVx1_ASAP7_75t_L g748 ( .A(n_69), .Y(n_748) );
AOI21xp5_ASAP7_75t_L g130 ( .A1(n_70), .A2(n_131), .B(n_138), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_71), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_72), .A2(n_131), .B(n_160), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_73), .Y(n_506) );
INVx1_ASAP7_75t_L g534 ( .A(n_74), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_75), .A2(n_266), .B(n_267), .Y(n_265) );
INVx1_ASAP7_75t_L g161 ( .A(n_76), .Y(n_161) );
CKINVDCx16_ASAP7_75t_R g202 ( .A(n_77), .Y(n_202) );
OAI22xp5_ASAP7_75t_SL g431 ( .A1(n_78), .A2(n_79), .B1(n_432), .B2(n_433), .Y(n_431) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_78), .Y(n_433) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_79), .Y(n_432) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_80), .A2(n_136), .B(n_141), .C(n_536), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_81), .A2(n_131), .B(n_190), .Y(n_189) );
INVx1_ASAP7_75t_L g164 ( .A(n_82), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_83), .B(n_206), .Y(n_450) );
INVx2_ASAP7_75t_L g126 ( .A(n_84), .Y(n_126) );
INVx1_ASAP7_75t_L g180 ( .A(n_85), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_86), .B(n_452), .Y(n_451) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_87), .A2(n_136), .B(n_141), .C(n_481), .Y(n_480) );
OR2x2_ASAP7_75t_L g111 ( .A(n_88), .B(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g721 ( .A(n_88), .Y(n_721) );
OR2x2_ASAP7_75t_L g723 ( .A(n_88), .B(n_113), .Y(n_723) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_89), .A2(n_141), .B(n_219), .C(n_222), .Y(n_218) );
AOI22xp33_ASAP7_75t_L g116 ( .A1(n_90), .A2(n_117), .B1(n_118), .B2(n_434), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_90), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_91), .B(n_125), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_92), .Y(n_486) );
A2O1A1Ixp33_ASAP7_75t_L g458 ( .A1(n_93), .A2(n_136), .B(n_141), .C(n_459), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_94), .Y(n_465) );
INVx1_ASAP7_75t_L g510 ( .A(n_95), .Y(n_510) );
CKINVDCx16_ASAP7_75t_R g470 ( .A(n_96), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_97), .B(n_206), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_98), .B(n_154), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_99), .B(n_154), .Y(n_474) );
INVx2_ASAP7_75t_L g195 ( .A(n_100), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_101), .A2(n_131), .B(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_102), .B(n_748), .Y(n_747) );
OA21x2_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_107), .B(n_437), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g738 ( .A(n_106), .Y(n_738) );
OAI21xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_116), .B(n_435), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_SL g436 ( .A(n_111), .Y(n_436) );
NOR2x2_ASAP7_75t_L g730 ( .A(n_112), .B(n_721), .Y(n_730) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
OR2x2_ASAP7_75t_L g720 ( .A(n_113), .B(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
XOR2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_431), .Y(n_118) );
INVx2_ASAP7_75t_L g722 ( .A(n_119), .Y(n_722) );
OAI22xp5_ASAP7_75t_SL g731 ( .A1(n_119), .A2(n_723), .B1(n_732), .B2(n_733), .Y(n_731) );
OR2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_361), .Y(n_119) );
NAND5xp2_ASAP7_75t_L g120 ( .A(n_121), .B(n_276), .C(n_308), .D(n_325), .E(n_348), .Y(n_120) );
AOI221xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_199), .B1(n_236), .B2(n_240), .C(n_244), .Y(n_121) );
INVx1_ASAP7_75t_L g388 ( .A(n_122), .Y(n_388) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_171), .Y(n_122) );
AND3x2_ASAP7_75t_L g363 ( .A(n_123), .B(n_173), .C(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_156), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_124), .B(n_242), .Y(n_241) );
BUFx3_ASAP7_75t_L g251 ( .A(n_124), .Y(n_251) );
AND2x2_ASAP7_75t_L g255 ( .A(n_124), .B(n_187), .Y(n_255) );
INVx2_ASAP7_75t_L g285 ( .A(n_124), .Y(n_285) );
OR2x2_ASAP7_75t_L g296 ( .A(n_124), .B(n_188), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_124), .B(n_172), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_124), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g375 ( .A(n_124), .B(n_188), .Y(n_375) );
OA21x2_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_130), .B(n_153), .Y(n_124) );
INVx1_ASAP7_75t_L g174 ( .A(n_125), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_L g201 ( .A1(n_125), .A2(n_177), .B(n_202), .C(n_203), .Y(n_201) );
INVx2_ASAP7_75t_L g225 ( .A(n_125), .Y(n_225) );
OA21x2_ASAP7_75t_L g467 ( .A1(n_125), .A2(n_468), .B(n_474), .Y(n_467) );
AND2x2_ASAP7_75t_SL g125 ( .A(n_126), .B(n_127), .Y(n_125) );
AND2x2_ASAP7_75t_L g155 ( .A(n_126), .B(n_127), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
BUFx2_ASAP7_75t_L g266 ( .A(n_131), .Y(n_266) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_136), .Y(n_131) );
NAND2x1p5_ASAP7_75t_L g177 ( .A(n_132), .B(n_136), .Y(n_177) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_135), .Y(n_132) );
INVx1_ASAP7_75t_L g209 ( .A(n_133), .Y(n_209) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g142 ( .A(n_134), .Y(n_142) );
INVx1_ASAP7_75t_L g197 ( .A(n_134), .Y(n_197) );
INVx1_ASAP7_75t_L g143 ( .A(n_135), .Y(n_143) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_135), .Y(n_146) );
INVx3_ASAP7_75t_L g149 ( .A(n_135), .Y(n_149) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_135), .Y(n_166) );
INVx1_ASAP7_75t_L g452 ( .A(n_135), .Y(n_452) );
INVx4_ASAP7_75t_SL g152 ( .A(n_136), .Y(n_152) );
BUFx3_ASAP7_75t_L g210 ( .A(n_136), .Y(n_210) );
O2A1O1Ixp33_ASAP7_75t_SL g138 ( .A1(n_139), .A2(n_140), .B(n_144), .C(n_152), .Y(n_138) );
O2A1O1Ixp33_ASAP7_75t_SL g160 ( .A1(n_140), .A2(n_152), .B(n_161), .C(n_162), .Y(n_160) );
O2A1O1Ixp33_ASAP7_75t_SL g190 ( .A1(n_140), .A2(n_152), .B(n_191), .C(n_192), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_L g228 ( .A1(n_140), .A2(n_152), .B(n_229), .C(n_230), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_SL g267 ( .A1(n_140), .A2(n_152), .B(n_268), .C(n_269), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_140), .A2(n_152), .B(n_470), .C(n_471), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_140), .A2(n_152), .B(n_492), .C(n_493), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_L g509 ( .A1(n_140), .A2(n_152), .B(n_510), .C(n_511), .Y(n_509) );
INVx5_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x6_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
BUFx3_ASAP7_75t_L g151 ( .A(n_142), .Y(n_151) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_142), .Y(n_234) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx4_ASAP7_75t_L g193 ( .A(n_146), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
INVx5_ASAP7_75t_L g206 ( .A(n_149), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_149), .B(n_495), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_149), .B(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g184 ( .A(n_150), .Y(n_184) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g167 ( .A(n_151), .Y(n_167) );
INVx1_ASAP7_75t_L g222 ( .A(n_152), .Y(n_222) );
OAI22xp33_ASAP7_75t_L g499 ( .A1(n_152), .A2(n_177), .B1(n_500), .B2(n_504), .Y(n_499) );
HB1xp67_ASAP7_75t_L g158 ( .A(n_154), .Y(n_158) );
INVx4_ASAP7_75t_L g170 ( .A(n_154), .Y(n_170) );
OA21x2_ASAP7_75t_L g507 ( .A1(n_154), .A2(n_508), .B(n_514), .Y(n_507) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g263 ( .A(n_155), .Y(n_263) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_156), .Y(n_254) );
AND2x2_ASAP7_75t_L g316 ( .A(n_156), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_156), .B(n_172), .Y(n_335) );
INVx1_ASAP7_75t_SL g156 ( .A(n_157), .Y(n_156) );
OR2x2_ASAP7_75t_L g243 ( .A(n_157), .B(n_172), .Y(n_243) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_157), .Y(n_250) );
AND2x2_ASAP7_75t_L g302 ( .A(n_157), .B(n_188), .Y(n_302) );
NAND3xp33_ASAP7_75t_L g327 ( .A(n_157), .B(n_171), .C(n_285), .Y(n_327) );
AND2x2_ASAP7_75t_L g392 ( .A(n_157), .B(n_173), .Y(n_392) );
AND2x2_ASAP7_75t_L g426 ( .A(n_157), .B(n_172), .Y(n_426) );
OA21x2_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_159), .B(n_168), .Y(n_157) );
OA21x2_ASAP7_75t_L g188 ( .A1(n_158), .A2(n_189), .B(n_198), .Y(n_188) );
OA21x2_ASAP7_75t_L g226 ( .A1(n_158), .A2(n_227), .B(n_235), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_165), .B(n_195), .Y(n_194) );
OAI22xp33_ASAP7_75t_L g270 ( .A1(n_165), .A2(n_206), .B1(n_271), .B2(n_272), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_165), .B(n_473), .Y(n_472) );
INVx4_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g182 ( .A(n_166), .Y(n_182) );
OAI22xp5_ASAP7_75t_SL g501 ( .A1(n_166), .A2(n_182), .B1(n_502), .B2(n_503), .Y(n_501) );
OA21x2_ASAP7_75t_L g489 ( .A1(n_169), .A2(n_490), .B(n_496), .Y(n_489) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_170), .B(n_186), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_170), .B(n_212), .Y(n_211) );
AO21x2_ASAP7_75t_L g215 ( .A1(n_170), .A2(n_216), .B(n_223), .Y(n_215) );
NOR2xp33_ASAP7_75t_SL g453 ( .A(n_170), .B(n_454), .Y(n_453) );
INVxp67_ASAP7_75t_L g252 ( .A(n_171), .Y(n_252) );
AND2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_187), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_172), .B(n_285), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_172), .B(n_316), .Y(n_324) );
AND2x2_ASAP7_75t_L g374 ( .A(n_172), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g402 ( .A(n_172), .Y(n_402) );
INVx4_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AND2x2_ASAP7_75t_L g309 ( .A(n_173), .B(n_302), .Y(n_309) );
BUFx3_ASAP7_75t_L g341 ( .A(n_173), .Y(n_341) );
AO21x2_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_185), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_174), .B(n_465), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_174), .B(n_486), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_174), .B(n_540), .Y(n_539) );
OAI21xp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_178), .Y(n_175) );
OAI21xp5_ASAP7_75t_L g216 ( .A1(n_177), .A2(n_217), .B(n_218), .Y(n_216) );
OAI21xp5_ASAP7_75t_L g478 ( .A1(n_177), .A2(n_479), .B(n_480), .Y(n_478) );
OAI21xp5_ASAP7_75t_L g533 ( .A1(n_177), .A2(n_534), .B(n_535), .Y(n_533) );
O2A1O1Ixp5_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B(n_183), .C(n_184), .Y(n_179) );
O2A1O1Ixp33_ASAP7_75t_L g219 ( .A1(n_181), .A2(n_184), .B(n_220), .C(n_221), .Y(n_219) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_184), .A2(n_450), .B(n_451), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_184), .A2(n_537), .B(n_538), .Y(n_536) );
INVx2_ASAP7_75t_L g317 ( .A(n_187), .Y(n_317) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_188), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_193), .B(n_232), .Y(n_231) );
INVx2_ASAP7_75t_L g484 ( .A(n_196), .Y(n_484) );
INVx3_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_199), .A2(n_377), .B1(n_379), .B2(n_380), .Y(n_376) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_213), .Y(n_199) );
AND2x2_ASAP7_75t_L g236 ( .A(n_200), .B(n_237), .Y(n_236) );
INVx3_ASAP7_75t_SL g247 ( .A(n_200), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_200), .B(n_280), .Y(n_312) );
OR2x2_ASAP7_75t_L g331 ( .A(n_200), .B(n_214), .Y(n_331) );
AND2x2_ASAP7_75t_L g336 ( .A(n_200), .B(n_288), .Y(n_336) );
AND2x2_ASAP7_75t_L g339 ( .A(n_200), .B(n_281), .Y(n_339) );
AND2x2_ASAP7_75t_L g351 ( .A(n_200), .B(n_226), .Y(n_351) );
AND2x2_ASAP7_75t_L g367 ( .A(n_200), .B(n_215), .Y(n_367) );
AND2x4_ASAP7_75t_L g370 ( .A(n_200), .B(n_238), .Y(n_370) );
OR2x2_ASAP7_75t_L g387 ( .A(n_200), .B(n_323), .Y(n_387) );
OR2x2_ASAP7_75t_L g418 ( .A(n_200), .B(n_260), .Y(n_418) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_200), .B(n_346), .Y(n_420) );
OR2x6_ASAP7_75t_L g200 ( .A(n_201), .B(n_211), .Y(n_200) );
O2A1O1Ixp33_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_207), .C(n_208), .Y(n_204) );
O2A1O1Ixp33_ASAP7_75t_L g481 ( .A1(n_206), .A2(n_482), .B(n_483), .C(n_484), .Y(n_481) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_209), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g294 ( .A(n_213), .B(n_258), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_213), .B(n_281), .Y(n_413) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_226), .Y(n_213) );
AND2x2_ASAP7_75t_L g246 ( .A(n_214), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g280 ( .A(n_214), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g288 ( .A(n_214), .B(n_260), .Y(n_288) );
AND2x2_ASAP7_75t_L g306 ( .A(n_214), .B(n_238), .Y(n_306) );
OR2x2_ASAP7_75t_L g323 ( .A(n_214), .B(n_281), .Y(n_323) );
INVx2_ASAP7_75t_SL g214 ( .A(n_215), .Y(n_214) );
BUFx2_ASAP7_75t_L g239 ( .A(n_215), .Y(n_239) );
AND2x2_ASAP7_75t_L g346 ( .A(n_215), .B(n_226), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
INVx1_ASAP7_75t_L g275 ( .A(n_225), .Y(n_275) );
AO21x2_ASAP7_75t_L g456 ( .A1(n_225), .A2(n_457), .B(n_464), .Y(n_456) );
INVx2_ASAP7_75t_L g238 ( .A(n_226), .Y(n_238) );
INVx1_ASAP7_75t_L g358 ( .A(n_226), .Y(n_358) );
AND2x2_ASAP7_75t_L g408 ( .A(n_226), .B(n_247), .Y(n_408) );
INVx3_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_234), .Y(n_462) );
AND2x2_ASAP7_75t_L g257 ( .A(n_237), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g292 ( .A(n_237), .B(n_247), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_237), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
AND2x2_ASAP7_75t_L g279 ( .A(n_238), .B(n_247), .Y(n_279) );
OR2x2_ASAP7_75t_L g395 ( .A(n_239), .B(n_369), .Y(n_395) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_242), .B(n_375), .Y(n_381) );
INVx2_ASAP7_75t_SL g242 ( .A(n_243), .Y(n_242) );
OAI32xp33_ASAP7_75t_L g337 ( .A1(n_243), .A2(n_338), .A3(n_340), .B1(n_342), .B2(n_343), .Y(n_337) );
OR2x2_ASAP7_75t_L g354 ( .A(n_243), .B(n_296), .Y(n_354) );
OAI21xp33_ASAP7_75t_SL g379 ( .A1(n_243), .A2(n_253), .B(n_284), .Y(n_379) );
OAI22xp33_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_248), .B1(n_253), .B2(n_256), .Y(n_244) );
INVxp33_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_246), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_247), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g305 ( .A(n_247), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g405 ( .A(n_247), .B(n_346), .Y(n_405) );
OR2x2_ASAP7_75t_L g429 ( .A(n_247), .B(n_323), .Y(n_429) );
AOI21xp33_ASAP7_75t_L g412 ( .A1(n_248), .A2(n_311), .B(n_413), .Y(n_412) );
OR2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_252), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
INVx1_ASAP7_75t_L g289 ( .A(n_250), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_250), .B(n_255), .Y(n_307) );
AND2x2_ASAP7_75t_L g329 ( .A(n_251), .B(n_302), .Y(n_329) );
INVx1_ASAP7_75t_L g342 ( .A(n_251), .Y(n_342) );
OR2x2_ASAP7_75t_L g347 ( .A(n_251), .B(n_281), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_254), .B(n_296), .Y(n_295) );
OAI22xp33_ASAP7_75t_L g277 ( .A1(n_255), .A2(n_278), .B1(n_283), .B2(n_287), .Y(n_277) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
OAI22xp5_ASAP7_75t_L g326 ( .A1(n_258), .A2(n_320), .B1(n_327), .B2(n_328), .Y(n_326) );
AND2x2_ASAP7_75t_L g404 ( .A(n_258), .B(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx1_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_260), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g423 ( .A(n_260), .B(n_306), .Y(n_423) );
AO21x2_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_264), .B(n_273), .Y(n_260) );
INVx1_ASAP7_75t_L g282 ( .A(n_261), .Y(n_282) );
AO21x2_ASAP7_75t_L g532 ( .A1(n_261), .A2(n_533), .B(n_539), .Y(n_532) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AOI21xp5_ASAP7_75t_SL g446 ( .A1(n_262), .A2(n_447), .B(n_448), .Y(n_446) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AO21x2_ASAP7_75t_L g477 ( .A1(n_263), .A2(n_478), .B(n_485), .Y(n_477) );
AO21x2_ASAP7_75t_L g498 ( .A1(n_263), .A2(n_499), .B(n_505), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_263), .B(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
OA21x2_ASAP7_75t_L g281 ( .A1(n_265), .A2(n_274), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AOI221xp5_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_289), .B1(n_290), .B2(n_295), .C(n_297), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_279), .B(n_281), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_279), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g298 ( .A(n_280), .Y(n_298) );
O2A1O1Ixp33_ASAP7_75t_L g385 ( .A1(n_280), .A2(n_386), .B(n_387), .C(n_388), .Y(n_385) );
AND2x2_ASAP7_75t_L g390 ( .A(n_280), .B(n_370), .Y(n_390) );
O2A1O1Ixp33_ASAP7_75t_SL g428 ( .A1(n_280), .A2(n_369), .B(n_429), .C(n_430), .Y(n_428) );
BUFx3_ASAP7_75t_L g320 ( .A(n_281), .Y(n_320) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_284), .B(n_341), .Y(n_384) );
AOI211xp5_ASAP7_75t_L g403 ( .A1(n_284), .A2(n_404), .B(n_406), .C(n_412), .Y(n_403) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVxp67_ASAP7_75t_L g364 ( .A(n_286), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_288), .B(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
AOI211xp5_ASAP7_75t_L g308 ( .A1(n_292), .A2(n_309), .B(n_310), .C(n_318), .Y(n_308) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g393 ( .A(n_296), .Y(n_393) );
OR2x2_ASAP7_75t_L g410 ( .A(n_296), .B(n_340), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_299), .B1(n_304), .B2(n_307), .Y(n_297) );
OAI22xp33_ASAP7_75t_L g310 ( .A1(n_299), .A2(n_311), .B1(n_312), .B2(n_313), .Y(n_310) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
OR2x2_ASAP7_75t_L g397 ( .A(n_301), .B(n_341), .Y(n_397) );
INVx1_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g352 ( .A(n_302), .B(n_342), .Y(n_352) );
INVx1_ASAP7_75t_L g360 ( .A(n_303), .Y(n_360) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_306), .B(n_320), .Y(n_368) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g359 ( .A(n_316), .B(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g425 ( .A(n_317), .Y(n_425) );
AOI21xp33_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_321), .B(n_324), .Y(n_318) );
INVx1_ASAP7_75t_L g355 ( .A(n_319), .Y(n_355) );
NAND2xp5_ASAP7_75t_SL g330 ( .A(n_320), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_320), .B(n_351), .Y(n_350) );
NAND2x1p5_ASAP7_75t_L g371 ( .A(n_320), .B(n_346), .Y(n_371) );
NAND2xp5_ASAP7_75t_SL g378 ( .A(n_320), .B(n_367), .Y(n_378) );
OAI211xp5_ASAP7_75t_L g382 ( .A1(n_320), .A2(n_330), .B(n_370), .C(n_383), .Y(n_382) );
INVx1_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
AOI221xp5_ASAP7_75t_SL g325 ( .A1(n_326), .A2(n_330), .B1(n_332), .B2(n_336), .C(n_337), .Y(n_325) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVxp67_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_334), .B(n_342), .Y(n_416) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
O2A1O1Ixp33_ASAP7_75t_L g427 ( .A1(n_336), .A2(n_351), .B(n_353), .C(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_339), .B(n_346), .Y(n_411) );
NAND2xp5_ASAP7_75t_SL g430 ( .A(n_340), .B(n_393), .Y(n_430) );
CKINVDCx16_ASAP7_75t_R g340 ( .A(n_341), .Y(n_340) );
INVxp33_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_345), .B(n_347), .Y(n_344) );
AOI21xp33_ASAP7_75t_SL g356 ( .A1(n_345), .A2(n_357), .B(n_359), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_345), .B(n_418), .Y(n_417) );
INVx2_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_346), .B(n_400), .Y(n_399) );
AOI221xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_352), .B1(n_353), .B2(n_355), .C(n_356), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_352), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g386 ( .A(n_358), .Y(n_386) );
NAND5xp2_ASAP7_75t_L g361 ( .A(n_362), .B(n_389), .C(n_403), .D(n_414), .E(n_427), .Y(n_361) );
AOI211xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_365), .B(n_372), .C(n_385), .Y(n_362) );
INVx2_ASAP7_75t_SL g409 ( .A(n_363), .Y(n_409) );
NAND4xp25_ASAP7_75t_SL g365 ( .A(n_366), .B(n_368), .C(n_369), .D(n_371), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx3_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OAI211xp5_ASAP7_75t_SL g372 ( .A1(n_371), .A2(n_373), .B(n_376), .C(n_382), .Y(n_372) );
CKINVDCx20_ASAP7_75t_R g373 ( .A(n_374), .Y(n_373) );
AOI221xp5_ASAP7_75t_L g414 ( .A1(n_374), .A2(n_415), .B1(n_417), .B2(n_419), .C(n_421), .Y(n_414) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AOI221xp5_ASAP7_75t_SL g389 ( .A1(n_390), .A2(n_391), .B1(n_394), .B2(n_396), .C(n_398), .Y(n_389) );
AND2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_397), .A2(n_420), .B1(n_422), .B2(n_424), .Y(n_421) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_409), .B1(n_410), .B2(n_411), .Y(n_406) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
NAND3xp33_ASAP7_75t_L g437 ( .A(n_435), .B(n_438), .C(n_736), .Y(n_437) );
OAI22xp5_ASAP7_75t_SL g439 ( .A1(n_440), .A2(n_720), .B1(n_722), .B2(n_723), .Y(n_439) );
INVx2_ASAP7_75t_L g732 ( .A(n_440), .Y(n_732) );
AND2x2_ASAP7_75t_SL g440 ( .A(n_441), .B(n_689), .Y(n_440) );
NOR3xp33_ASAP7_75t_L g441 ( .A(n_442), .B(n_582), .C(n_655), .Y(n_441) );
OAI211xp5_ASAP7_75t_SL g442 ( .A1(n_443), .A2(n_475), .B(n_515), .C(n_566), .Y(n_442) );
INVxp67_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_455), .Y(n_444) );
AND2x2_ASAP7_75t_L g531 ( .A(n_445), .B(n_532), .Y(n_531) );
INVx3_ASAP7_75t_L g549 ( .A(n_445), .Y(n_549) );
INVx2_ASAP7_75t_L g564 ( .A(n_445), .Y(n_564) );
INVx1_ASAP7_75t_L g594 ( .A(n_445), .Y(n_594) );
AND2x2_ASAP7_75t_L g644 ( .A(n_445), .B(n_565), .Y(n_644) );
AOI32xp33_ASAP7_75t_L g671 ( .A1(n_445), .A2(n_599), .A3(n_672), .B1(n_674), .B2(n_675), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_445), .B(n_521), .Y(n_677) );
AND2x2_ASAP7_75t_L g704 ( .A(n_445), .B(n_547), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_445), .B(n_713), .Y(n_712) );
OR2x6_ASAP7_75t_L g445 ( .A(n_446), .B(n_453), .Y(n_445) );
AND2x2_ASAP7_75t_L g593 ( .A(n_455), .B(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g615 ( .A(n_455), .Y(n_615) );
AND2x2_ASAP7_75t_L g700 ( .A(n_455), .B(n_531), .Y(n_700) );
AND2x2_ASAP7_75t_L g703 ( .A(n_455), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_466), .Y(n_455) );
INVx2_ASAP7_75t_L g523 ( .A(n_456), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_456), .B(n_547), .Y(n_553) );
AND2x2_ASAP7_75t_L g563 ( .A(n_456), .B(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g599 ( .A(n_456), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_458), .B(n_463), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_461), .B(n_462), .Y(n_459) );
AND2x2_ASAP7_75t_L g541 ( .A(n_466), .B(n_523), .Y(n_541) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g524 ( .A(n_467), .Y(n_524) );
AND2x2_ASAP7_75t_L g565 ( .A(n_467), .B(n_547), .Y(n_565) );
AND2x2_ASAP7_75t_L g634 ( .A(n_467), .B(n_532), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_487), .Y(n_475) );
OR2x2_ASAP7_75t_L g529 ( .A(n_476), .B(n_498), .Y(n_529) );
INVx1_ASAP7_75t_L g607 ( .A(n_476), .Y(n_607) );
AND2x2_ASAP7_75t_L g621 ( .A(n_476), .B(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_476), .B(n_497), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_476), .B(n_619), .Y(n_673) );
AND2x2_ASAP7_75t_L g681 ( .A(n_476), .B(n_682), .Y(n_681) );
INVx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx3_ASAP7_75t_L g519 ( .A(n_477), .Y(n_519) );
AND2x2_ASAP7_75t_L g588 ( .A(n_477), .B(n_498), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_487), .B(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g715 ( .A(n_487), .Y(n_715) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_497), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_488), .B(n_559), .Y(n_581) );
OR2x2_ASAP7_75t_L g610 ( .A(n_488), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g642 ( .A(n_488), .B(n_622), .Y(n_642) );
INVx1_ASAP7_75t_SL g662 ( .A(n_488), .Y(n_662) );
AND2x2_ASAP7_75t_L g666 ( .A(n_488), .B(n_528), .Y(n_666) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_SL g520 ( .A(n_489), .B(n_497), .Y(n_520) );
AND2x2_ASAP7_75t_L g527 ( .A(n_489), .B(n_507), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_489), .B(n_551), .Y(n_550) );
OR2x2_ASAP7_75t_L g569 ( .A(n_489), .B(n_551), .Y(n_569) );
INVx1_ASAP7_75t_SL g576 ( .A(n_489), .Y(n_576) );
BUFx2_ASAP7_75t_L g587 ( .A(n_489), .Y(n_587) );
AND2x2_ASAP7_75t_L g603 ( .A(n_489), .B(n_519), .Y(n_603) );
AND2x2_ASAP7_75t_L g618 ( .A(n_489), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g682 ( .A(n_489), .B(n_498), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_497), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g606 ( .A(n_497), .B(n_607), .Y(n_606) );
AOI221xp5_ASAP7_75t_L g623 ( .A1(n_497), .A2(n_624), .B1(n_627), .B2(n_630), .C(n_635), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_497), .B(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_507), .Y(n_497) );
INVx3_ASAP7_75t_L g551 ( .A(n_498), .Y(n_551) );
BUFx2_ASAP7_75t_L g561 ( .A(n_507), .Y(n_561) );
AND2x2_ASAP7_75t_L g575 ( .A(n_507), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g592 ( .A(n_507), .Y(n_592) );
OR2x2_ASAP7_75t_L g611 ( .A(n_507), .B(n_551), .Y(n_611) );
INVx3_ASAP7_75t_L g619 ( .A(n_507), .Y(n_619) );
AND2x2_ASAP7_75t_L g622 ( .A(n_507), .B(n_551), .Y(n_622) );
AOI221xp5_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_521), .B1(n_525), .B2(n_530), .C(n_542), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_520), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_518), .B(n_591), .Y(n_716) );
OR2x2_ASAP7_75t_L g719 ( .A(n_518), .B(n_550), .Y(n_719) );
INVx1_ASAP7_75t_SL g518 ( .A(n_519), .Y(n_518) );
OAI221xp5_ASAP7_75t_SL g542 ( .A1(n_519), .A2(n_543), .B1(n_550), .B2(n_552), .C(n_555), .Y(n_542) );
AND2x2_ASAP7_75t_L g559 ( .A(n_519), .B(n_551), .Y(n_559) );
AND2x2_ASAP7_75t_L g567 ( .A(n_519), .B(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_519), .B(n_575), .Y(n_574) );
NAND2x1_ASAP7_75t_L g617 ( .A(n_519), .B(n_618), .Y(n_617) );
OR2x2_ASAP7_75t_L g669 ( .A(n_519), .B(n_611), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_521), .A2(n_629), .B1(n_658), .B2(n_660), .Y(n_657) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AOI322xp5_ASAP7_75t_L g566 ( .A1(n_522), .A2(n_531), .A3(n_567), .B1(n_570), .B2(n_573), .C1(n_577), .C2(n_580), .Y(n_566) );
OR2x2_ASAP7_75t_L g578 ( .A(n_522), .B(n_579), .Y(n_578) );
OR2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_523), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g557 ( .A(n_523), .B(n_532), .Y(n_557) );
INVx1_ASAP7_75t_L g572 ( .A(n_523), .Y(n_572) );
AND2x2_ASAP7_75t_L g638 ( .A(n_523), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g548 ( .A(n_524), .B(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g639 ( .A(n_524), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_524), .B(n_547), .Y(n_713) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_528), .B(n_662), .Y(n_661) );
INVx3_ASAP7_75t_SL g528 ( .A(n_529), .Y(n_528) );
OR2x2_ASAP7_75t_L g613 ( .A(n_529), .B(n_560), .Y(n_613) );
OR2x2_ASAP7_75t_L g710 ( .A(n_529), .B(n_561), .Y(n_710) );
INVx1_ASAP7_75t_L g691 ( .A(n_530), .Y(n_691) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_541), .Y(n_530) );
INVx4_ASAP7_75t_L g579 ( .A(n_531), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_531), .B(n_598), .Y(n_604) );
INVx2_ASAP7_75t_L g547 ( .A(n_532), .Y(n_547) );
INVx1_ASAP7_75t_L g629 ( .A(n_541), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_541), .B(n_601), .Y(n_670) );
AOI21xp33_ASAP7_75t_L g616 ( .A1(n_543), .A2(n_617), .B(n_620), .Y(n_616) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_548), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g601 ( .A(n_547), .Y(n_601) );
INVx1_ASAP7_75t_L g628 ( .A(n_547), .Y(n_628) );
INVx1_ASAP7_75t_L g554 ( .A(n_548), .Y(n_554) );
AND2x2_ASAP7_75t_L g556 ( .A(n_548), .B(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g652 ( .A(n_549), .B(n_638), .Y(n_652) );
AND2x2_ASAP7_75t_L g674 ( .A(n_549), .B(n_634), .Y(n_674) );
BUFx2_ASAP7_75t_L g626 ( .A(n_551), .Y(n_626) );
OR2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
AOI32xp33_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_558), .A3(n_559), .B1(n_560), .B2(n_562), .Y(n_555) );
INVx1_ASAP7_75t_L g636 ( .A(n_556), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_556), .A2(n_684), .B1(n_685), .B2(n_687), .Y(n_683) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_559), .B(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_559), .B(n_618), .Y(n_659) );
AND2x2_ASAP7_75t_L g706 ( .A(n_559), .B(n_591), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_560), .B(n_607), .Y(n_654) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g707 ( .A(n_562), .Y(n_707) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_565), .Y(n_562) );
INVx1_ASAP7_75t_L g632 ( .A(n_563), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_565), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g679 ( .A(n_565), .B(n_599), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_565), .B(n_594), .Y(n_686) );
INVx1_ASAP7_75t_SL g668 ( .A(n_567), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_568), .B(n_619), .Y(n_646) );
NOR4xp25_ASAP7_75t_L g692 ( .A(n_568), .B(n_591), .C(n_693), .D(n_696), .Y(n_692) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_569), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVxp67_ASAP7_75t_L g649 ( .A(n_572), .Y(n_649) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OAI21xp33_ASAP7_75t_L g699 ( .A1(n_575), .A2(n_666), .B(n_700), .Y(n_699) );
AND2x4_ASAP7_75t_L g591 ( .A(n_576), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g640 ( .A(n_579), .Y(n_640) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NAND4xp25_ASAP7_75t_SL g582 ( .A(n_583), .B(n_608), .C(n_623), .D(n_643), .Y(n_582) );
O2A1O1Ixp33_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_589), .B(n_593), .C(n_595), .Y(n_583) );
INVx1_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g675 ( .A(n_588), .B(n_618), .Y(n_675) );
AND2x2_ASAP7_75t_L g684 ( .A(n_588), .B(n_662), .Y(n_684) );
INVx3_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_591), .B(n_626), .Y(n_688) );
AND2x2_ASAP7_75t_L g600 ( .A(n_594), .B(n_601), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_602), .B1(n_604), .B2(n_605), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .Y(n_597) );
AND2x2_ASAP7_75t_L g698 ( .A(n_598), .B(n_644), .Y(n_698) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_600), .B(n_649), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_601), .B(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
O2A1O1Ixp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_612), .B(n_614), .C(n_616), .Y(n_608) );
AOI221xp5_ASAP7_75t_L g643 ( .A1(n_609), .A2(n_644), .B1(n_645), .B2(n_647), .C(n_650), .Y(n_643) );
INVx1_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
OAI221xp5_ASAP7_75t_L g701 ( .A1(n_617), .A2(n_702), .B1(n_705), .B2(n_707), .C(n_708), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_618), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_SL g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_626), .B(n_695), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
INVx1_ASAP7_75t_L g656 ( .A(n_628), .Y(n_656) );
INVx1_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_631), .A2(n_651), .B1(n_653), .B2(n_654), .Y(n_650) );
OR2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AOI21xp33_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_637), .B(n_641), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_640), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
OAI221xp5_ASAP7_75t_L g714 ( .A1(n_651), .A2(n_677), .B1(n_715), .B2(n_716), .C(n_717), .Y(n_714) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g696 ( .A(n_653), .Y(n_696) );
OAI211xp5_ASAP7_75t_SL g655 ( .A1(n_656), .A2(n_657), .B(n_663), .C(n_683), .Y(n_655) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
AOI211xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_666), .B(n_667), .C(n_676), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
A2O1A1Ixp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .B(n_670), .C(n_671), .Y(n_667) );
INVx1_ASAP7_75t_L g695 ( .A(n_673), .Y(n_695) );
OAI21xp5_ASAP7_75t_SL g717 ( .A1(n_674), .A2(n_700), .B(n_718), .Y(n_717) );
AOI21xp33_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_678), .B(n_680), .Y(n_676) );
INVx1_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
INVxp67_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
OAI21xp5_ASAP7_75t_SL g709 ( .A1(n_686), .A2(n_710), .B(n_711), .Y(n_709) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NOR3xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_701), .C(n_714), .Y(n_689) );
OAI211xp5_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_692), .B(n_697), .C(n_699), .Y(n_690) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
CKINVDCx14_ASAP7_75t_R g702 ( .A(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g734 ( .A(n_720), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_724), .Y(n_735) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
CKINVDCx12_ASAP7_75t_R g741 ( .A(n_742), .Y(n_741) );
HB1xp67_ASAP7_75t_L g749 ( .A(n_742), .Y(n_749) );
OR2x2_ASAP7_75t_L g742 ( .A(n_743), .B(n_745), .Y(n_742) );
INVx1_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
endmodule