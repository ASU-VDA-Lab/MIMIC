module real_aes_7842_n_335 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_335);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_335;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_792;
wire n_386;
wire n_503;
wire n_673;
wire n_518;
wire n_635;
wire n_878;
wire n_665;
wire n_991;
wire n_667;
wire n_580;
wire n_577;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_491;
wire n_923;
wire n_894;
wire n_1034;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_353;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_666;
wire n_537;
wire n_551;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_856;
wire n_594;
wire n_983;
wire n_767;
wire n_889;
wire n_696;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1046;
wire n_677;
wire n_958;
wire n_1021;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_815;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_356;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_372;
wire n_528;
wire n_892;
wire n_495;
wire n_994;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_951;
wire n_875;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_1053;
wire n_466;
wire n_559;
wire n_872;
wire n_636;
wire n_976;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_931;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_755;
wire n_656;
wire n_532;
wire n_746;
wire n_1025;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_1049;
wire n_874;
wire n_796;
wire n_801;
wire n_383;
wire n_529;
wire n_725;
wire n_455;
wire n_504;
wire n_960;
wire n_671;
wire n_973;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_345;
wire n_885;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_664;
wire n_367;
wire n_819;
wire n_1017;
wire n_737;
wire n_1013;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_940;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_1006;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_947;
wire n_561;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_769;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_733;
wire n_617;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1037;
wire n_1031;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_488;
wire n_501;
wire n_1041;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1003;
wire n_1000;
wire n_1028;
wire n_366;
wire n_346;
wire n_727;
wire n_1014;
wire n_397;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_354;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_691;
wire n_498;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_1005;
wire n_939;
wire n_831;
wire n_487;
wire n_653;
wire n_365;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_789;
wire n_544;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_741;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_347;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_1045;
wire n_465;
wire n_473;
wire n_566;
wire n_719;
wire n_837;
wire n_967;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_337;
wire n_1024;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_SL g563 ( .A1(n_0), .A2(n_253), .B1(n_564), .B2(n_566), .Y(n_563) );
CKINVDCx20_ASAP7_75t_R g631 ( .A(n_1), .Y(n_631) );
CKINVDCx20_ASAP7_75t_R g819 ( .A(n_2), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_3), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_4), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_5), .A2(n_43), .B1(n_379), .B2(n_729), .Y(n_902) );
CKINVDCx20_ASAP7_75t_R g1027 ( .A(n_6), .Y(n_1027) );
AO22x2_ASAP7_75t_L g368 ( .A1(n_7), .A2(n_194), .B1(n_360), .B2(n_361), .Y(n_368) );
INVx1_ASAP7_75t_L g1018 ( .A(n_7), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_8), .A2(n_133), .B1(n_612), .B2(n_613), .Y(n_611) );
CKINVDCx20_ASAP7_75t_R g914 ( .A(n_9), .Y(n_914) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_10), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g636 ( .A(n_11), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_12), .A2(n_256), .B1(n_478), .B2(n_522), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_13), .A2(n_77), .B1(n_613), .B2(n_984), .Y(n_983) );
CKINVDCx20_ASAP7_75t_R g699 ( .A(n_14), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_15), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_16), .A2(n_130), .B1(n_355), .B2(n_680), .Y(n_810) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_17), .Y(n_557) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_18), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g895 ( .A(n_19), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_20), .A2(n_316), .B1(n_872), .B2(n_929), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_21), .A2(n_319), .B1(n_395), .B2(n_403), .Y(n_394) );
CKINVDCx20_ASAP7_75t_R g665 ( .A(n_22), .Y(n_665) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_23), .Y(n_528) );
AOI222xp33_ASAP7_75t_L g946 ( .A1(n_24), .A2(n_46), .B1(n_302), .B2(n_390), .C1(n_575), .C2(n_947), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_25), .A2(n_105), .B1(n_468), .B2(n_877), .Y(n_1040) );
CKINVDCx20_ASAP7_75t_R g867 ( .A(n_26), .Y(n_867) );
AO22x2_ASAP7_75t_L g364 ( .A1(n_27), .A2(n_90), .B1(n_360), .B2(n_365), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g1043 ( .A1(n_28), .A2(n_330), .B1(n_621), .B2(n_969), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_29), .A2(n_179), .B1(n_420), .B2(n_425), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_30), .A2(n_218), .B1(n_468), .B2(n_533), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_31), .A2(n_44), .B1(n_434), .B2(n_435), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_32), .A2(n_95), .B1(n_412), .B2(n_703), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_33), .A2(n_135), .B1(n_596), .B2(n_889), .Y(n_888) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_34), .A2(n_242), .B1(n_653), .B2(n_654), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_35), .B(n_753), .Y(n_752) );
AOI22xp5_ASAP7_75t_SL g569 ( .A1(n_36), .A2(n_570), .B1(n_571), .B2(n_601), .Y(n_569) );
INVx1_ASAP7_75t_L g601 ( .A(n_36), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_37), .A2(n_260), .B1(n_506), .B2(n_507), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_38), .A2(n_188), .B1(n_506), .B2(n_556), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_39), .A2(n_216), .B1(n_595), .B2(n_596), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_40), .B(n_808), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g629 ( .A(n_41), .Y(n_629) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_42), .Y(n_708) );
CKINVDCx20_ASAP7_75t_R g996 ( .A(n_45), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_47), .A2(n_213), .B1(n_435), .B2(n_619), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g977 ( .A1(n_48), .A2(n_978), .B1(n_1002), .B2(n_1003), .Y(n_977) );
INVx1_ASAP7_75t_L g1002 ( .A(n_48), .Y(n_1002) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_49), .B(n_633), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_50), .A2(n_281), .B1(n_784), .B2(n_891), .Y(n_890) );
AOI22xp33_ASAP7_75t_SL g684 ( .A1(n_51), .A2(n_240), .B1(n_685), .B2(n_686), .Y(n_684) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_52), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_53), .Y(n_727) );
INVx1_ASAP7_75t_L g773 ( .A(n_54), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_55), .A2(n_84), .B1(n_371), .B2(n_468), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_56), .A2(n_301), .B1(n_710), .B2(n_784), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_57), .A2(n_78), .B1(n_872), .B2(n_874), .Y(n_871) );
CKINVDCx20_ASAP7_75t_R g910 ( .A(n_58), .Y(n_910) );
AOI222xp33_ASAP7_75t_L g728 ( .A1(n_59), .A2(n_248), .B1(n_299), .B2(n_575), .C1(n_633), .C2(n_729), .Y(n_728) );
AOI22xp5_ASAP7_75t_L g805 ( .A1(n_60), .A2(n_227), .B1(n_506), .B2(n_507), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_61), .A2(n_259), .B1(n_474), .B2(n_479), .Y(n_945) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_62), .A2(n_183), .B1(n_390), .B2(n_634), .Y(n_748) );
INVx1_ASAP7_75t_L g649 ( .A(n_63), .Y(n_649) );
CKINVDCx20_ASAP7_75t_R g917 ( .A(n_64), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_65), .A2(n_111), .B1(n_586), .B2(n_587), .Y(n_907) );
AO22x2_ASAP7_75t_L g359 ( .A1(n_66), .A2(n_221), .B1(n_360), .B2(n_361), .Y(n_359) );
INVx1_ASAP7_75t_L g1015 ( .A(n_66), .Y(n_1015) );
CKINVDCx20_ASAP7_75t_R g961 ( .A(n_67), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_68), .A2(n_69), .B1(n_478), .B2(n_479), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_70), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_71), .A2(n_88), .B1(n_436), .B2(n_470), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_72), .A2(n_201), .B1(n_381), .B2(n_507), .Y(n_551) );
OA22x2_ASAP7_75t_L g488 ( .A1(n_73), .A2(n_489), .B1(n_490), .B2(n_491), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_73), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g1033 ( .A(n_74), .Y(n_1033) );
CKINVDCx20_ASAP7_75t_R g1001 ( .A(n_75), .Y(n_1001) );
AOI211xp5_ASAP7_75t_L g335 ( .A1(n_76), .A2(n_336), .B(n_345), .C(n_1020), .Y(n_335) );
INVx1_ASAP7_75t_L g638 ( .A(n_79), .Y(n_638) );
AOI221xp5_ASAP7_75t_L g723 ( .A1(n_80), .A2(n_291), .B1(n_395), .B2(n_724), .C(n_725), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_81), .A2(n_120), .B1(n_578), .B2(n_580), .Y(n_577) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_82), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_83), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_85), .A2(n_154), .B1(n_511), .B2(n_680), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g981 ( .A1(n_86), .A2(n_185), .B1(n_619), .B2(n_982), .Y(n_981) );
AOI22xp33_ASAP7_75t_SL g590 ( .A1(n_87), .A2(n_317), .B1(n_591), .B2(n_592), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_89), .A2(n_124), .B1(n_432), .B2(n_686), .Y(n_818) );
INVx1_ASAP7_75t_L g1019 ( .A(n_90), .Y(n_1019) );
AOI22xp33_ASAP7_75t_SL g584 ( .A1(n_91), .A2(n_142), .B1(n_458), .B2(n_511), .Y(n_584) );
CKINVDCx20_ASAP7_75t_R g901 ( .A(n_92), .Y(n_901) );
CKINVDCx20_ASAP7_75t_R g662 ( .A(n_93), .Y(n_662) );
CKINVDCx20_ASAP7_75t_R g1035 ( .A(n_94), .Y(n_1035) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_96), .A2(n_190), .B1(n_621), .B2(n_686), .Y(n_847) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_97), .Y(n_701) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_98), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g672 ( .A(n_99), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_100), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_101), .A2(n_255), .B1(n_474), .B2(n_815), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g986 ( .A1(n_102), .A2(n_239), .B1(n_591), .B2(n_782), .Y(n_986) );
AOI22xp5_ASAP7_75t_L g987 ( .A1(n_103), .A2(n_198), .B1(n_622), .B2(n_784), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_104), .A2(n_112), .B1(n_616), .B2(n_844), .Y(n_843) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_106), .A2(n_273), .B1(n_431), .B2(n_468), .Y(n_560) );
CKINVDCx20_ASAP7_75t_R g1029 ( .A(n_107), .Y(n_1029) );
AOI22xp33_ASAP7_75t_SL g966 ( .A1(n_108), .A2(n_150), .B1(n_355), .B2(n_458), .Y(n_966) );
AOI22xp33_ASAP7_75t_SL g970 ( .A1(n_109), .A2(n_267), .B1(n_478), .B2(n_929), .Y(n_970) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_110), .A2(n_294), .B1(n_381), .B2(n_458), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_113), .A2(n_276), .B1(n_386), .B2(n_556), .Y(n_921) );
AOI22xp33_ASAP7_75t_SL g679 ( .A1(n_114), .A2(n_287), .B1(n_507), .B2(n_680), .Y(n_679) );
AOI22xp33_ASAP7_75t_SL g385 ( .A1(n_115), .A2(n_163), .B1(n_386), .B2(n_390), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_116), .A2(n_292), .B1(n_420), .B2(n_599), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_117), .A2(n_167), .B1(n_689), .B2(n_759), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_118), .A2(n_174), .B1(n_613), .B2(n_656), .Y(n_763) );
CKINVDCx20_ASAP7_75t_R g661 ( .A(n_119), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_121), .B(n_677), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_122), .A2(n_173), .B1(n_530), .B2(n_653), .Y(n_1041) );
AND2x6_ASAP7_75t_L g340 ( .A(n_123), .B(n_341), .Y(n_340) );
HB1xp67_ASAP7_75t_L g1012 ( .A(n_123), .Y(n_1012) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_125), .A2(n_208), .B1(n_782), .B2(n_842), .Y(n_841) );
AOI22xp33_ASAP7_75t_SL g904 ( .A1(n_126), .A2(n_244), .B1(n_580), .B2(n_905), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_127), .A2(n_148), .B1(n_474), .B2(n_476), .Y(n_473) );
INVx1_ASAP7_75t_L g837 ( .A(n_128), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_129), .A2(n_230), .B1(n_470), .B2(n_471), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g856 ( .A(n_131), .Y(n_856) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_132), .A2(n_228), .B1(n_434), .B2(n_519), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_134), .A2(n_155), .B1(n_758), .B2(n_759), .Y(n_757) );
AOI22xp5_ASAP7_75t_SL g765 ( .A1(n_136), .A2(n_766), .B1(n_794), .B2(n_795), .Y(n_765) );
INVx1_ASAP7_75t_L g795 ( .A(n_136), .Y(n_795) );
AOI22xp33_ASAP7_75t_SL g673 ( .A1(n_137), .A2(n_247), .B1(n_506), .B2(n_674), .Y(n_673) );
CKINVDCx20_ASAP7_75t_R g925 ( .A(n_138), .Y(n_925) );
AOI22xp5_ASAP7_75t_L g655 ( .A1(n_139), .A2(n_272), .B1(n_476), .B2(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_SL g965 ( .A(n_140), .B(n_395), .Y(n_965) );
INVx1_ASAP7_75t_L g769 ( .A(n_141), .Y(n_769) );
AO22x2_ASAP7_75t_L g367 ( .A1(n_143), .A2(n_211), .B1(n_360), .B2(n_365), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g1016 ( .A(n_143), .B(n_1017), .Y(n_1016) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_144), .B(n_998), .Y(n_997) );
AOI22xp33_ASAP7_75t_SL g973 ( .A1(n_145), .A2(n_226), .B1(n_527), .B2(n_596), .Y(n_973) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_146), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g930 ( .A1(n_147), .A2(n_315), .B1(n_878), .B2(n_931), .Y(n_930) );
AOI22xp33_ASAP7_75t_SL g962 ( .A1(n_149), .A2(n_236), .B1(n_507), .B2(n_634), .Y(n_962) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_151), .Y(n_804) );
CKINVDCx20_ASAP7_75t_R g858 ( .A(n_152), .Y(n_858) );
CKINVDCx20_ASAP7_75t_R g860 ( .A(n_153), .Y(n_860) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_156), .Y(n_545) );
AOI22xp33_ASAP7_75t_SL g813 ( .A1(n_157), .A2(n_197), .B1(n_429), .B2(n_436), .Y(n_813) );
AOI22xp33_ASAP7_75t_SL g972 ( .A1(n_158), .A2(n_171), .B1(n_436), .B2(n_616), .Y(n_972) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_159), .A2(n_203), .B1(n_415), .B2(n_478), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_160), .A2(n_199), .B1(n_586), .B2(n_587), .Y(n_585) );
AOI22xp33_ASAP7_75t_SL g598 ( .A1(n_161), .A2(n_320), .B1(n_519), .B2(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g576 ( .A(n_162), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_164), .A2(n_279), .B1(n_621), .B2(n_622), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_165), .A2(n_334), .B1(n_429), .B2(n_432), .Y(n_428) );
CKINVDCx20_ASAP7_75t_R g1037 ( .A(n_166), .Y(n_1037) );
CKINVDCx20_ASAP7_75t_R g948 ( .A(n_168), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_169), .A2(n_326), .B1(n_478), .B2(n_522), .Y(n_938) );
CKINVDCx20_ASAP7_75t_R g377 ( .A(n_170), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_172), .A2(n_258), .B1(n_521), .B2(n_522), .Y(n_520) );
AOI22xp33_ASAP7_75t_SL g817 ( .A1(n_175), .A2(n_266), .B1(n_434), .B2(n_685), .Y(n_817) );
AOI22xp33_ASAP7_75t_SL g968 ( .A1(n_176), .A2(n_313), .B1(n_420), .B2(n_969), .Y(n_968) );
CKINVDCx20_ASAP7_75t_R g940 ( .A(n_177), .Y(n_940) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_178), .B(n_633), .Y(n_632) );
AOI22xp33_ASAP7_75t_SL g683 ( .A1(n_180), .A2(n_225), .B1(n_468), .B2(n_474), .Y(n_683) );
CKINVDCx20_ASAP7_75t_R g1032 ( .A(n_181), .Y(n_1032) );
CKINVDCx20_ASAP7_75t_R g627 ( .A(n_182), .Y(n_627) );
CKINVDCx20_ASAP7_75t_R g828 ( .A(n_184), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_186), .A2(n_193), .B1(n_634), .B2(n_863), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_187), .A2(n_293), .B1(n_431), .B2(n_595), .Y(n_932) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_189), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_191), .A2(n_224), .B1(n_479), .B2(n_616), .Y(n_615) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_192), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g924 ( .A(n_195), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_196), .A2(n_305), .B1(n_521), .B2(n_787), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_200), .A2(n_286), .B1(n_478), .B2(n_522), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_202), .A2(n_241), .B1(n_789), .B2(n_792), .Y(n_788) );
OA22x2_ASAP7_75t_L g441 ( .A1(n_204), .A2(n_442), .B1(n_443), .B2(n_480), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_204), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g964 ( .A(n_205), .B(n_724), .Y(n_964) );
XNOR2x2_ASAP7_75t_L g884 ( .A(n_206), .B(n_885), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_207), .A2(n_324), .B1(n_410), .B2(n_415), .Y(n_409) );
INVx2_ASAP7_75t_L g344 ( .A(n_209), .Y(n_344) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_210), .A2(n_608), .B1(n_641), .B2(n_642), .Y(n_607) );
INVx1_ASAP7_75t_L g641 ( .A(n_210), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g876 ( .A1(n_212), .A2(n_223), .B1(n_877), .B2(n_878), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_214), .B(n_587), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g994 ( .A(n_215), .Y(n_994) );
AOI22xp33_ASAP7_75t_SL g690 ( .A1(n_217), .A2(n_332), .B1(n_415), .B2(n_432), .Y(n_690) );
CKINVDCx20_ASAP7_75t_R g893 ( .A(n_219), .Y(n_893) );
AOI22xp33_ASAP7_75t_SL g688 ( .A1(n_220), .A2(n_328), .B1(n_654), .B2(n_689), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_222), .A2(n_307), .B1(n_387), .B2(n_674), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_229), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_231), .A2(n_270), .B1(n_434), .B2(n_435), .Y(n_846) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_232), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_233), .B(n_751), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_234), .A2(n_696), .B1(n_731), .B2(n_732), .Y(n_695) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_234), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_235), .A2(n_329), .B1(n_527), .B2(n_530), .Y(n_870) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_237), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_238), .Y(n_446) );
OA22x2_ASAP7_75t_L g349 ( .A1(n_243), .A2(n_350), .B1(n_351), .B2(n_438), .Y(n_349) );
CKINVDCx20_ASAP7_75t_R g350 ( .A(n_243), .Y(n_350) );
INVx1_ASAP7_75t_L g772 ( .A(n_245), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_246), .A2(n_269), .B1(n_929), .B2(n_1045), .Y(n_1044) );
INVx1_ASAP7_75t_L g776 ( .A(n_249), .Y(n_776) );
INVx1_ASAP7_75t_L g360 ( .A(n_250), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_250), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_251), .A2(n_327), .B1(n_468), .B2(n_470), .Y(n_881) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_252), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g553 ( .A(n_254), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g991 ( .A(n_257), .Y(n_991) );
CKINVDCx20_ASAP7_75t_R g826 ( .A(n_261), .Y(n_826) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_262), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g1054 ( .A(n_263), .Y(n_1054) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_264), .Y(n_369) );
INVx1_ASAP7_75t_L g625 ( .A(n_265), .Y(n_625) );
INVx1_ASAP7_75t_L g990 ( .A(n_268), .Y(n_990) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_271), .B(n_751), .Y(n_941) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_274), .Y(n_496) );
AOI22xp33_ASAP7_75t_SL g762 ( .A1(n_275), .A2(n_323), .B1(n_564), .B2(n_566), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_277), .A2(n_312), .B1(n_415), .B2(n_474), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_278), .A2(n_298), .B1(n_387), .B2(n_582), .Y(n_663) );
INVx1_ASAP7_75t_L g343 ( .A(n_280), .Y(n_343) );
CKINVDCx20_ASAP7_75t_R g830 ( .A(n_282), .Y(n_830) );
CKINVDCx20_ASAP7_75t_R g974 ( .A(n_283), .Y(n_974) );
INVx1_ASAP7_75t_L g341 ( .A(n_284), .Y(n_341) );
CKINVDCx20_ASAP7_75t_R g897 ( .A(n_285), .Y(n_897) );
OA22x2_ASAP7_75t_L g667 ( .A1(n_288), .A2(n_668), .B1(n_669), .B2(n_691), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_288), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_289), .A2(n_318), .B1(n_479), .B2(n_782), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_290), .B(n_396), .Y(n_678) );
CKINVDCx20_ASAP7_75t_R g920 ( .A(n_295), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_296), .B(n_379), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g898 ( .A(n_297), .Y(n_898) );
AOI22xp5_ASAP7_75t_L g1021 ( .A1(n_300), .A2(n_1022), .B1(n_1023), .B2(n_1046), .Y(n_1021) );
CKINVDCx20_ASAP7_75t_R g1046 ( .A(n_300), .Y(n_1046) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_303), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g831 ( .A(n_304), .Y(n_831) );
INVx1_ASAP7_75t_L g882 ( .A(n_306), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g1030 ( .A(n_308), .B(n_580), .Y(n_1030) );
CKINVDCx20_ASAP7_75t_R g1000 ( .A(n_309), .Y(n_1000) );
INVx1_ASAP7_75t_L g770 ( .A(n_310), .Y(n_770) );
CKINVDCx20_ASAP7_75t_R g865 ( .A(n_311), .Y(n_865) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_314), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_321), .Y(n_705) );
INVx1_ASAP7_75t_L g568 ( .A(n_322), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_325), .Y(n_764) );
OA22x2_ASAP7_75t_SL g821 ( .A1(n_331), .A2(n_822), .B1(n_823), .B2(n_848), .Y(n_821) );
INVx1_ASAP7_75t_L g848 ( .A(n_331), .Y(n_848) );
INVx1_ASAP7_75t_L g777 ( .A(n_333), .Y(n_777) );
CKINVDCx20_ASAP7_75t_R g336 ( .A(n_337), .Y(n_336) );
CKINVDCx20_ASAP7_75t_R g337 ( .A(n_338), .Y(n_337) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_340), .B(n_342), .Y(n_339) );
HB1xp67_ASAP7_75t_L g1011 ( .A(n_341), .Y(n_1011) );
OAI21xp5_ASAP7_75t_L g1052 ( .A1(n_342), .A2(n_1010), .B(n_1053), .Y(n_1052) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
AOI221xp5_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_736), .B1(n_1005), .B2(n_1006), .C(n_1007), .Y(n_345) );
INVx1_ASAP7_75t_L g1005 ( .A(n_346), .Y(n_1005) );
AOI22xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_348), .B1(n_483), .B2(n_735), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AOI22xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_439), .B1(n_481), .B2(n_482), .Y(n_348) );
INVx1_ASAP7_75t_L g481 ( .A(n_349), .Y(n_481) );
INVx1_ASAP7_75t_SL g438 ( .A(n_351), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_352), .B(n_407), .Y(n_351) );
NOR2x1_ASAP7_75t_L g352 ( .A(n_353), .B(n_384), .Y(n_352) );
OAI222xp33_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_369), .B1(n_370), .B2(n_377), .C1(n_378), .C2(n_383), .Y(n_353) );
OAI221xp5_ASAP7_75t_L g829 ( .A1(n_354), .A2(n_574), .B1(n_830), .B2(n_831), .C(n_832), .Y(n_829) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx4_ASAP7_75t_L g730 ( .A(n_355), .Y(n_730) );
BUFx2_ASAP7_75t_L g863 ( .A(n_355), .Y(n_863) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx2_ASAP7_75t_L g471 ( .A(n_356), .Y(n_471) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_356), .Y(n_511) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_356), .Y(n_556) );
BUFx4f_ASAP7_75t_SL g674 ( .A(n_356), .Y(n_674) );
AND2x4_ASAP7_75t_L g356 ( .A(n_357), .B(n_366), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_363), .Y(n_357) );
INVx1_ASAP7_75t_L g382 ( .A(n_358), .Y(n_382) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g376 ( .A(n_359), .Y(n_376) );
INVx1_ASAP7_75t_L g393 ( .A(n_359), .Y(n_393) );
AND2x2_ASAP7_75t_L g399 ( .A(n_359), .B(n_375), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_359), .B(n_367), .Y(n_418) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g365 ( .A(n_362), .Y(n_365) );
AND2x2_ASAP7_75t_L g414 ( .A(n_363), .B(n_402), .Y(n_414) );
INVx1_ASAP7_75t_L g515 ( .A(n_363), .Y(n_515) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g373 ( .A(n_364), .B(n_368), .Y(n_373) );
INVx1_ASAP7_75t_L g389 ( .A(n_364), .Y(n_389) );
OR2x2_ASAP7_75t_L g401 ( .A(n_364), .B(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g406 ( .A(n_364), .B(n_402), .Y(n_406) );
AND2x4_ASAP7_75t_L g381 ( .A(n_366), .B(n_382), .Y(n_381) );
AND2x4_ASAP7_75t_L g387 ( .A(n_366), .B(n_388), .Y(n_387) );
NAND2x1p5_ASAP7_75t_L g514 ( .A(n_366), .B(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
INVx2_ASAP7_75t_L g375 ( .A(n_367), .Y(n_375) );
AND2x2_ASAP7_75t_L g424 ( .A(n_367), .B(n_393), .Y(n_424) );
INVx2_ASAP7_75t_L g402 ( .A(n_368), .Y(n_402) );
INVx2_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g747 ( .A(n_371), .Y(n_747) );
BUFx6f_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx3_ASAP7_75t_L g504 ( .A(n_372), .Y(n_504) );
INVx4_ASAP7_75t_L g549 ( .A(n_372), .Y(n_549) );
INVx2_ASAP7_75t_L g803 ( .A(n_372), .Y(n_803) );
INVx2_ASAP7_75t_L g960 ( .A(n_372), .Y(n_960) );
INVx2_ASAP7_75t_SL g993 ( .A(n_372), .Y(n_993) );
AND2x6_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
AND2x4_ASAP7_75t_L g391 ( .A(n_373), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g463 ( .A(n_373), .Y(n_463) );
AND2x2_ASAP7_75t_L g413 ( .A(n_374), .B(n_414), .Y(n_413) );
AND2x6_ASAP7_75t_L g431 ( .A(n_374), .B(n_400), .Y(n_431) );
AND2x4_ASAP7_75t_L g434 ( .A(n_374), .B(n_406), .Y(n_434) );
AND2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
BUFx4f_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g1028 ( .A(n_380), .Y(n_1028) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx12f_ASAP7_75t_L g506 ( .A(n_381), .Y(n_506) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_381), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_394), .Y(n_384) );
BUFx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx2_ASAP7_75t_L g458 ( .A(n_387), .Y(n_458) );
BUFx3_ASAP7_75t_L g680 ( .A(n_387), .Y(n_680) );
INVx1_ASAP7_75t_L g906 ( .A(n_387), .Y(n_906) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OR2x6_ASAP7_75t_L g426 ( .A(n_389), .B(n_418), .Y(n_426) );
BUFx2_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
BUFx2_ASAP7_75t_SL g507 ( .A(n_391), .Y(n_507) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_391), .Y(n_582) );
INVx1_ASAP7_75t_L g464 ( .A(n_392), .Y(n_464) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx5_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g586 ( .A(n_397), .Y(n_586) );
INVx2_ASAP7_75t_L g751 ( .A(n_397), .Y(n_751) );
INVx2_ASAP7_75t_L g808 ( .A(n_397), .Y(n_808) );
INVx4_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AND2x4_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
AND2x6_ASAP7_75t_L g405 ( .A(n_399), .B(n_406), .Y(n_405) );
AND2x4_ASAP7_75t_L g432 ( .A(n_399), .B(n_414), .Y(n_432) );
INVx1_ASAP7_75t_L g449 ( .A(n_399), .Y(n_449) );
NAND2x1p5_ASAP7_75t_L g453 ( .A(n_399), .B(n_406), .Y(n_453) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g448 ( .A(n_401), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_SL g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g677 ( .A(n_404), .Y(n_677) );
INVx1_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
BUFx2_ASAP7_75t_L g587 ( .A(n_405), .Y(n_587) );
BUFx2_ASAP7_75t_L g724 ( .A(n_405), .Y(n_724) );
BUFx4f_ASAP7_75t_L g753 ( .A(n_405), .Y(n_753) );
AND2x2_ASAP7_75t_L g423 ( .A(n_406), .B(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g707 ( .A(n_406), .B(n_424), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_408), .B(n_427), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_419), .Y(n_408) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx3_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx3_ASAP7_75t_L g612 ( .A(n_412), .Y(n_612) );
BUFx3_ASAP7_75t_L g782 ( .A(n_412), .Y(n_782) );
BUFx6f_ASAP7_75t_L g889 ( .A(n_412), .Y(n_889) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g475 ( .A(n_413), .Y(n_475) );
BUFx2_ASAP7_75t_SL g527 ( .A(n_413), .Y(n_527) );
BUFx2_ASAP7_75t_SL g595 ( .A(n_413), .Y(n_595) );
AND2x4_ASAP7_75t_L g416 ( .A(n_414), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g437 ( .A(n_414), .B(n_424), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_414), .B(n_424), .Y(n_538) );
BUFx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx3_ASAP7_75t_L g479 ( .A(n_416), .Y(n_479) );
BUFx2_ASAP7_75t_SL g530 ( .A(n_416), .Y(n_530) );
BUFx2_ASAP7_75t_SL g596 ( .A(n_416), .Y(n_596) );
BUFx3_ASAP7_75t_L g703 ( .A(n_416), .Y(n_703) );
BUFx3_ASAP7_75t_L g815 ( .A(n_416), .Y(n_815) );
BUFx3_ASAP7_75t_L g844 ( .A(n_416), .Y(n_844) );
AND2x2_ASAP7_75t_L g656 ( .A(n_417), .B(n_515), .Y(n_656) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx3_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx3_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx5_ASAP7_75t_L g476 ( .A(n_422), .Y(n_476) );
INVx1_ASAP7_75t_L g519 ( .A(n_422), .Y(n_519) );
INVx3_ASAP7_75t_L g566 ( .A(n_422), .Y(n_566) );
INVx4_ASAP7_75t_L g685 ( .A(n_422), .Y(n_685) );
INVx8_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_426), .A2(n_460), .B1(n_461), .B2(n_462), .Y(n_459) );
INVx6_ASAP7_75t_SL g523 ( .A(n_426), .Y(n_523) );
INVx1_ASAP7_75t_SL g686 ( .A(n_426), .Y(n_686) );
INVx1_ASAP7_75t_L g874 ( .A(n_426), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_433), .Y(n_427) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_429), .Y(n_720) );
INVx1_ASAP7_75t_L g894 ( .A(n_429), .Y(n_894) );
INVx5_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g533 ( .A(n_430), .Y(n_533) );
INVx4_ASAP7_75t_L g758 ( .A(n_430), .Y(n_758) );
INVx2_ASAP7_75t_L g787 ( .A(n_430), .Y(n_787) );
INVx11_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx11_ASAP7_75t_L g455 ( .A(n_431), .Y(n_455) );
BUFx3_ASAP7_75t_L g478 ( .A(n_432), .Y(n_478) );
BUFx3_ASAP7_75t_L g521 ( .A(n_432), .Y(n_521) );
INVx2_ASAP7_75t_L g614 ( .A(n_432), .Y(n_614) );
BUFx6f_ASAP7_75t_L g880 ( .A(n_432), .Y(n_880) );
BUFx3_ASAP7_75t_L g1045 ( .A(n_432), .Y(n_1045) );
BUFx3_ASAP7_75t_L g470 ( .A(n_434), .Y(n_470) );
INVx6_ASAP7_75t_L g565 ( .A(n_434), .Y(n_565) );
BUFx3_ASAP7_75t_L g619 ( .A(n_434), .Y(n_619) );
BUFx3_ASAP7_75t_L g791 ( .A(n_434), .Y(n_791) );
BUFx3_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx3_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx3_ASAP7_75t_L g468 ( .A(n_437), .Y(n_468) );
BUFx3_ASAP7_75t_L g593 ( .A(n_437), .Y(n_593) );
BUFx3_ASAP7_75t_L g759 ( .A(n_437), .Y(n_759) );
INVx1_ASAP7_75t_L g482 ( .A(n_439), .Y(n_482) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g480 ( .A(n_443), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_465), .Y(n_443) );
NOR3xp33_ASAP7_75t_L g444 ( .A(n_445), .B(n_454), .C(n_459), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_447), .B1(n_450), .B2(n_451), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_447), .A2(n_545), .B1(n_546), .B2(n_547), .Y(n_544) );
BUFx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g495 ( .A(n_448), .Y(n_495) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_448), .Y(n_626) );
OAI221xp5_ASAP7_75t_L g660 ( .A1(n_448), .A2(n_499), .B1(n_661), .B2(n_662), .C(n_663), .Y(n_660) );
OA211x2_ASAP7_75t_L g939 ( .A1(n_451), .A2(n_940), .B(n_941), .C(n_942), .Y(n_939) );
OAI22xp5_ASAP7_75t_L g989 ( .A1(n_451), .A2(n_827), .B1(n_990), .B2(n_991), .Y(n_989) );
INVx1_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g547 ( .A(n_452), .Y(n_547) );
INVx2_ASAP7_75t_L g918 ( .A(n_452), .Y(n_918) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx3_ASAP7_75t_L g499 ( .A(n_453), .Y(n_499) );
OAI21xp33_ASAP7_75t_SL g454 ( .A1(n_455), .A2(n_456), .B(n_457), .Y(n_454) );
INVx3_ASAP7_75t_L g591 ( .A(n_455), .Y(n_591) );
INVx4_ASAP7_75t_L g616 ( .A(n_455), .Y(n_616) );
INVx4_ASAP7_75t_L g654 ( .A(n_455), .Y(n_654) );
INVx2_ASAP7_75t_SL g877 ( .A(n_455), .Y(n_877) );
CKINVDCx16_ASAP7_75t_R g640 ( .A(n_462), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_462), .A2(n_514), .B1(n_726), .B2(n_727), .Y(n_725) );
BUFx2_ASAP7_75t_L g838 ( .A(n_462), .Y(n_838) );
OR2x6_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_472), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_469), .Y(n_466) );
BUFx2_ASAP7_75t_L g982 ( .A(n_468), .Y(n_982) );
INVx1_ASAP7_75t_L g630 ( .A(n_471), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_477), .Y(n_472) );
INVx3_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx3_ASAP7_75t_L g653 ( .A(n_475), .Y(n_653) );
BUFx6f_ASAP7_75t_L g621 ( .A(n_476), .Y(n_621) );
INVx1_ASAP7_75t_L g735 ( .A(n_483), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_485), .B1(n_604), .B2(n_734), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_488), .B1(n_539), .B2(n_603), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_516), .Y(n_491) );
NOR3xp33_ASAP7_75t_L g492 ( .A(n_493), .B(n_501), .C(n_508), .Y(n_492) );
OAI22xp5_ASAP7_75t_SL g493 ( .A1(n_494), .A2(n_496), .B1(n_497), .B2(n_500), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_494), .A2(n_547), .B1(n_769), .B2(n_770), .Y(n_768) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g827 ( .A(n_495), .Y(n_827) );
INVx1_ASAP7_75t_SL g857 ( .A(n_495), .Y(n_857) );
OAI22xp5_ASAP7_75t_L g825 ( .A1(n_497), .A2(n_826), .B1(n_827), .B2(n_828), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g855 ( .A1(n_497), .A2(n_856), .B1(n_857), .B2(n_858), .Y(n_855) );
OAI22xp5_ASAP7_75t_L g1031 ( .A1(n_497), .A2(n_915), .B1(n_1032), .B2(n_1033), .Y(n_1031) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_499), .A2(n_625), .B1(n_626), .B2(n_627), .Y(n_624) );
OAI21xp33_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_503), .B(n_505), .Y(n_501) );
OAI21xp5_ASAP7_75t_SL g664 ( .A1(n_503), .A2(n_665), .B(n_666), .Y(n_664) );
OAI21xp5_ASAP7_75t_SL g671 ( .A1(n_503), .A2(n_672), .B(n_673), .Y(n_671) );
INVx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g579 ( .A(n_506), .Y(n_579) );
BUFx4f_ASAP7_75t_SL g947 ( .A(n_506), .Y(n_947) );
OAI22xp33_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_510), .B1(n_512), .B2(n_513), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_511), .Y(n_510) );
OAI22xp5_ASAP7_75t_L g1034 ( .A1(n_513), .A2(n_1035), .B1(n_1036), .B2(n_1037), .Y(n_1034) );
BUFx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_514), .A2(n_553), .B1(n_554), .B2(n_557), .Y(n_552) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_514), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_514), .A2(n_776), .B1(n_777), .B2(n_778), .Y(n_775) );
INVx4_ASAP7_75t_L g836 ( .A(n_514), .Y(n_836) );
NOR3xp33_ASAP7_75t_L g516 ( .A(n_517), .B(n_524), .C(n_531), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_520), .Y(n_517) );
INVx1_ASAP7_75t_L g722 ( .A(n_521), .Y(n_722) );
BUFx2_ASAP7_75t_L g842 ( .A(n_521), .Y(n_842) );
BUFx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
BUFx4f_ASAP7_75t_SL g622 ( .A(n_523), .Y(n_622) );
BUFx2_ASAP7_75t_L g710 ( .A(n_523), .Y(n_710) );
BUFx2_ASAP7_75t_L g891 ( .A(n_523), .Y(n_891) );
BUFx2_ASAP7_75t_L g929 ( .A(n_523), .Y(n_929) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_526), .B1(n_528), .B2(n_529), .Y(n_524) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_534), .B1(n_535), .B2(n_536), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g896 ( .A1(n_536), .A2(n_565), .B1(n_897), .B2(n_898), .Y(n_896) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g716 ( .A(n_537), .Y(n_716) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g603 ( .A(n_539), .Y(n_603) );
OA22x2_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_541), .B1(n_569), .B2(n_602), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_541), .A2(n_606), .B1(n_607), .B2(n_643), .Y(n_605) );
INVx1_ASAP7_75t_L g643 ( .A(n_541), .Y(n_643) );
XOR2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_568), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_558), .Y(n_542) );
NOR3xp33_ASAP7_75t_L g543 ( .A(n_544), .B(n_548), .C(n_552), .Y(n_543) );
OAI21xp5_ASAP7_75t_SL g548 ( .A1(n_549), .A2(n_550), .B(n_551), .Y(n_548) );
INVx4_ASAP7_75t_L g575 ( .A(n_549), .Y(n_575) );
BUFx2_ASAP7_75t_L g861 ( .A(n_549), .Y(n_861) );
INVx2_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_SL g995 ( .A(n_555), .Y(n_995) );
BUFx6f_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g1036 ( .A(n_556), .Y(n_1036) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_559), .B(n_562), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_567), .Y(n_562) );
INVxp67_ASAP7_75t_L g714 ( .A(n_564), .Y(n_714) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g599 ( .A(n_565), .Y(n_599) );
INVx3_ASAP7_75t_L g689 ( .A(n_565), .Y(n_689) );
INVx2_ASAP7_75t_L g969 ( .A(n_565), .Y(n_969) );
INVx1_ASAP7_75t_L g602 ( .A(n_569), .Y(n_602) );
INVx1_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_572), .B(n_588), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_583), .Y(n_572) );
OAI21xp5_ASAP7_75t_SL g573 ( .A1(n_574), .A2(n_576), .B(n_577), .Y(n_573) );
OAI221xp5_ASAP7_75t_SL g628 ( .A1(n_574), .A2(n_629), .B1(n_630), .B2(n_631), .C(n_632), .Y(n_628) );
OAI221xp5_ASAP7_75t_SL g771 ( .A1(n_574), .A2(n_630), .B1(n_772), .B2(n_773), .C(n_774), .Y(n_771) );
OAI21xp33_ASAP7_75t_SL g919 ( .A1(n_574), .A2(n_920), .B(n_921), .Y(n_919) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx3_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_589), .B(n_597), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_594), .Y(n_589) );
BUFx4f_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .Y(n_597) );
INVx1_ASAP7_75t_L g734 ( .A(n_604), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_644), .B1(n_645), .B2(n_733), .Y(n_604) );
INVx1_ASAP7_75t_L g733 ( .A(n_605), .Y(n_733) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g642 ( .A(n_608), .Y(n_642) );
AND2x2_ASAP7_75t_SL g608 ( .A(n_609), .B(n_623), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_610), .B(n_617), .Y(n_609) );
NAND2xp33_ASAP7_75t_SL g610 ( .A(n_611), .B(n_615), .Y(n_610) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
NOR3xp33_ASAP7_75t_L g623 ( .A(n_624), .B(n_628), .C(n_635), .Y(n_623) );
INVx1_ASAP7_75t_L g916 ( .A(n_626), .Y(n_916) );
BUFx3_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g923 ( .A(n_634), .Y(n_923) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_637), .B1(n_638), .B2(n_639), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g999 ( .A1(n_639), .A2(n_835), .B1(n_1000), .B2(n_1001), .Y(n_999) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g778 ( .A(n_640), .Y(n_778) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OAI22xp5_ASAP7_75t_SL g645 ( .A1(n_646), .A2(n_647), .B1(n_694), .B2(n_695), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_667), .B1(n_692), .B2(n_693), .Y(n_647) );
INVx2_ASAP7_75t_SL g692 ( .A(n_648), .Y(n_692) );
XNOR2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
NOR4xp75_ASAP7_75t_L g650 ( .A(n_651), .B(n_657), .C(n_660), .D(n_664), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_652), .B(n_655), .Y(n_651) );
INVxp67_ASAP7_75t_L g700 ( .A(n_653), .Y(n_700) );
NAND2xp5_ASAP7_75t_SL g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx1_ASAP7_75t_L g693 ( .A(n_667), .Y(n_693) );
INVx1_ASAP7_75t_L g691 ( .A(n_669), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_670), .B(n_681), .Y(n_669) );
NOR2xp67_ASAP7_75t_L g670 ( .A(n_671), .B(n_675), .Y(n_670) );
NAND3xp33_ASAP7_75t_L g675 ( .A(n_676), .B(n_678), .C(n_679), .Y(n_675) );
NOR2x1_ASAP7_75t_L g681 ( .A(n_682), .B(n_687), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
BUFx6f_ASAP7_75t_L g784 ( .A(n_685), .Y(n_784) );
INVx2_ASAP7_75t_L g873 ( .A(n_685), .Y(n_873) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_690), .Y(n_687) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g732 ( .A(n_696), .Y(n_732) );
AND4x1_ASAP7_75t_L g696 ( .A(n_697), .B(n_711), .C(n_723), .D(n_728), .Y(n_696) );
NOR2xp33_ASAP7_75t_SL g697 ( .A(n_698), .B(n_704), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_700), .B1(n_701), .B2(n_702), .Y(n_698) );
INVx2_ASAP7_75t_L g931 ( .A(n_702), .Y(n_931) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_706), .B1(n_708), .B2(n_709), .Y(n_704) );
BUFx2_ASAP7_75t_R g706 ( .A(n_707), .Y(n_706) );
INVxp67_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_712), .B(n_717), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_714), .B1(n_715), .B2(n_716), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_719), .B1(n_721), .B2(n_722), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx3_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g1006 ( .A(n_736), .Y(n_1006) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_738), .B1(n_850), .B2(n_1004), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
AOI22xp5_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_796), .B1(n_797), .B2(n_849), .Y(n_738) );
INVx4_ASAP7_75t_L g849 ( .A(n_739), .Y(n_849) );
XOR2x2_ASAP7_75t_L g739 ( .A(n_740), .B(n_765), .Y(n_739) );
INVx2_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
OAI22x1_ASAP7_75t_L g798 ( .A1(n_741), .A2(n_742), .B1(n_799), .B2(n_820), .Y(n_798) );
INVx3_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
XOR2x2_ASAP7_75t_L g742 ( .A(n_743), .B(n_764), .Y(n_742) );
NAND2xp5_ASAP7_75t_SL g743 ( .A(n_744), .B(n_755), .Y(n_743) );
NOR2xp33_ASAP7_75t_L g744 ( .A(n_745), .B(n_749), .Y(n_744) );
OAI21xp5_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_747), .B(n_748), .Y(n_745) );
OAI221xp5_ASAP7_75t_L g1026 ( .A1(n_747), .A2(n_1027), .B1(n_1028), .B2(n_1029), .C(n_1030), .Y(n_1026) );
NAND3xp33_ASAP7_75t_L g749 ( .A(n_750), .B(n_752), .C(n_754), .Y(n_749) );
NOR2x1_ASAP7_75t_L g755 ( .A(n_756), .B(n_761), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_757), .B(n_760), .Y(n_756) );
INVx1_ASAP7_75t_L g793 ( .A(n_759), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_762), .B(n_763), .Y(n_761) );
INVx1_ASAP7_75t_SL g794 ( .A(n_766), .Y(n_794) );
AND2x2_ASAP7_75t_SL g766 ( .A(n_767), .B(n_779), .Y(n_766) );
NOR3xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_771), .C(n_775), .Y(n_767) );
OAI22xp5_ASAP7_75t_L g864 ( .A1(n_778), .A2(n_865), .B1(n_866), .B2(n_867), .Y(n_864) );
NOR2xp33_ASAP7_75t_L g779 ( .A(n_780), .B(n_785), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_781), .B(n_783), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_786), .B(n_788), .Y(n_785) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx3_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx2_ASAP7_75t_SL g796 ( .A(n_797), .Y(n_796) );
XNOR2x2_ASAP7_75t_L g797 ( .A(n_798), .B(n_821), .Y(n_797) );
INVx3_ASAP7_75t_L g820 ( .A(n_799), .Y(n_820) );
XOR2x2_ASAP7_75t_L g799 ( .A(n_800), .B(n_819), .Y(n_799) );
NAND2x1_ASAP7_75t_SL g800 ( .A(n_801), .B(n_811), .Y(n_800) );
NOR2xp33_ASAP7_75t_L g801 ( .A(n_802), .B(n_806), .Y(n_801) );
OAI21xp5_ASAP7_75t_SL g802 ( .A1(n_803), .A2(n_804), .B(n_805), .Y(n_802) );
OAI21xp5_ASAP7_75t_SL g900 ( .A1(n_803), .A2(n_901), .B(n_902), .Y(n_900) );
NAND3xp33_ASAP7_75t_L g806 ( .A(n_807), .B(n_809), .C(n_810), .Y(n_806) );
NOR2x1_ASAP7_75t_L g811 ( .A(n_812), .B(n_816), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .Y(n_812) );
BUFx2_ASAP7_75t_L g984 ( .A(n_815), .Y(n_984) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_817), .B(n_818), .Y(n_816) );
INVx2_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
AND2x2_ASAP7_75t_SL g823 ( .A(n_824), .B(n_839), .Y(n_823) );
NOR3xp33_ASAP7_75t_L g824 ( .A(n_825), .B(n_829), .C(n_833), .Y(n_824) );
OAI22xp5_ASAP7_75t_L g833 ( .A1(n_834), .A2(n_835), .B1(n_837), .B2(n_838), .Y(n_833) );
INVx2_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx3_ASAP7_75t_SL g866 ( .A(n_836), .Y(n_866) );
OAI22xp5_ASAP7_75t_SL g922 ( .A1(n_838), .A2(n_923), .B1(n_924), .B2(n_925), .Y(n_922) );
NOR2xp33_ASAP7_75t_L g839 ( .A(n_840), .B(n_845), .Y(n_839) );
NAND2xp5_ASAP7_75t_SL g840 ( .A(n_841), .B(n_843), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_846), .B(n_847), .Y(n_845) );
INVx1_ASAP7_75t_L g1004 ( .A(n_850), .Y(n_1004) );
XNOR2xp5_ASAP7_75t_SL g850 ( .A(n_851), .B(n_953), .Y(n_850) );
AOI22xp5_ASAP7_75t_L g851 ( .A1(n_852), .A2(n_883), .B1(n_951), .B2(n_952), .Y(n_851) );
INVx1_ASAP7_75t_L g951 ( .A(n_852), .Y(n_951) );
XOR2x2_ASAP7_75t_L g852 ( .A(n_853), .B(n_882), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_854), .B(n_868), .Y(n_853) );
NOR3xp33_ASAP7_75t_L g854 ( .A(n_855), .B(n_859), .C(n_864), .Y(n_854) );
OAI21xp33_ASAP7_75t_L g859 ( .A1(n_860), .A2(n_861), .B(n_862), .Y(n_859) );
NOR2xp33_ASAP7_75t_L g868 ( .A(n_869), .B(n_875), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_870), .B(n_871), .Y(n_869) );
INVx3_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_876), .B(n_881), .Y(n_875) );
INVx4_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
OAI22xp5_ASAP7_75t_L g892 ( .A1(n_879), .A2(n_893), .B1(n_894), .B2(n_895), .Y(n_892) );
INVx4_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g952 ( .A(n_883), .Y(n_952) );
AOI22xp5_ASAP7_75t_L g883 ( .A1(n_884), .A2(n_908), .B1(n_949), .B2(n_950), .Y(n_883) );
INVx2_ASAP7_75t_L g949 ( .A(n_884), .Y(n_949) );
NAND2xp5_ASAP7_75t_SL g885 ( .A(n_886), .B(n_899), .Y(n_885) );
NOR3xp33_ASAP7_75t_L g886 ( .A(n_887), .B(n_892), .C(n_896), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g887 ( .A(n_888), .B(n_890), .Y(n_887) );
NOR2xp33_ASAP7_75t_L g899 ( .A(n_900), .B(n_903), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g903 ( .A(n_904), .B(n_907), .Y(n_903) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx1_ASAP7_75t_L g950 ( .A(n_908), .Y(n_950) );
XNOR2xp5_ASAP7_75t_L g908 ( .A(n_909), .B(n_933), .Y(n_908) );
XNOR2x1_ASAP7_75t_L g909 ( .A(n_910), .B(n_911), .Y(n_909) );
AND2x2_ASAP7_75t_L g911 ( .A(n_912), .B(n_926), .Y(n_911) );
NOR3xp33_ASAP7_75t_L g912 ( .A(n_913), .B(n_919), .C(n_922), .Y(n_912) );
OAI22xp5_ASAP7_75t_L g913 ( .A1(n_914), .A2(n_915), .B1(n_917), .B2(n_918), .Y(n_913) );
INVx2_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
INVx1_ASAP7_75t_L g998 ( .A(n_923), .Y(n_998) );
AND4x1_ASAP7_75t_L g926 ( .A(n_927), .B(n_928), .C(n_930), .D(n_932), .Y(n_926) );
INVx2_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
XOR2x2_ASAP7_75t_L g934 ( .A(n_935), .B(n_948), .Y(n_934) );
NAND4xp75_ASAP7_75t_L g935 ( .A(n_936), .B(n_939), .C(n_943), .D(n_946), .Y(n_935) );
AND2x2_ASAP7_75t_L g936 ( .A(n_937), .B(n_938), .Y(n_936) );
AND2x2_ASAP7_75t_L g943 ( .A(n_944), .B(n_945), .Y(n_943) );
XNOR2xp5_ASAP7_75t_L g953 ( .A(n_954), .B(n_975), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_956), .Y(n_955) );
XOR2x2_ASAP7_75t_L g956 ( .A(n_957), .B(n_974), .Y(n_956) );
NAND3x1_ASAP7_75t_L g957 ( .A(n_958), .B(n_967), .C(n_971), .Y(n_957) );
NOR2xp33_ASAP7_75t_L g958 ( .A(n_959), .B(n_963), .Y(n_958) );
OAI21xp5_ASAP7_75t_SL g959 ( .A1(n_960), .A2(n_961), .B(n_962), .Y(n_959) );
NAND3xp33_ASAP7_75t_L g963 ( .A(n_964), .B(n_965), .C(n_966), .Y(n_963) );
AND2x2_ASAP7_75t_L g967 ( .A(n_968), .B(n_970), .Y(n_967) );
AND2x2_ASAP7_75t_L g971 ( .A(n_972), .B(n_973), .Y(n_971) );
INVx2_ASAP7_75t_L g975 ( .A(n_976), .Y(n_975) );
INVx1_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
INVx1_ASAP7_75t_L g1003 ( .A(n_978), .Y(n_1003) );
AND2x2_ASAP7_75t_SL g978 ( .A(n_979), .B(n_988), .Y(n_978) );
NOR2xp33_ASAP7_75t_SL g979 ( .A(n_980), .B(n_985), .Y(n_979) );
NAND2xp5_ASAP7_75t_L g980 ( .A(n_981), .B(n_983), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g985 ( .A(n_986), .B(n_987), .Y(n_985) );
NOR3xp33_ASAP7_75t_L g988 ( .A(n_989), .B(n_992), .C(n_999), .Y(n_988) );
OAI221xp5_ASAP7_75t_L g992 ( .A1(n_993), .A2(n_994), .B1(n_995), .B2(n_996), .C(n_997), .Y(n_992) );
INVx1_ASAP7_75t_SL g1007 ( .A(n_1008), .Y(n_1007) );
NOR2x1_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1013), .Y(n_1008) );
OR2x2_ASAP7_75t_SL g1058 ( .A(n_1009), .B(n_1014), .Y(n_1058) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1012), .Y(n_1009) );
CKINVDCx20_ASAP7_75t_R g1048 ( .A(n_1010), .Y(n_1048) );
INVx1_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g1053 ( .A(n_1011), .B(n_1050), .Y(n_1053) );
CKINVDCx16_ASAP7_75t_R g1050 ( .A(n_1012), .Y(n_1050) );
CKINVDCx20_ASAP7_75t_R g1013 ( .A(n_1014), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_1015), .B(n_1016), .Y(n_1014) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1019), .Y(n_1017) );
OAI322xp33_ASAP7_75t_L g1020 ( .A1(n_1021), .A2(n_1047), .A3(n_1049), .B1(n_1051), .B2(n_1054), .C1(n_1055), .C2(n_1058), .Y(n_1020) );
CKINVDCx20_ASAP7_75t_R g1022 ( .A(n_1023), .Y(n_1022) );
HB1xp67_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
XOR2x2_ASAP7_75t_L g1057 ( .A(n_1024), .B(n_1054), .Y(n_1057) );
NAND2xp5_ASAP7_75t_L g1024 ( .A(n_1025), .B(n_1038), .Y(n_1024) );
NOR3xp33_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1031), .C(n_1034), .Y(n_1025) );
NOR2xp33_ASAP7_75t_L g1038 ( .A(n_1039), .B(n_1042), .Y(n_1038) );
NAND2xp5_ASAP7_75t_L g1039 ( .A(n_1040), .B(n_1041), .Y(n_1039) );
NAND2xp5_ASAP7_75t_L g1042 ( .A(n_1043), .B(n_1044), .Y(n_1042) );
HB1xp67_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
CKINVDCx20_ASAP7_75t_R g1051 ( .A(n_1052), .Y(n_1051) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
endmodule