module fake_jpeg_25657_n_276 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_276);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_276;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx4f_ASAP7_75t_SL g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_21),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_31),
.B(n_33),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_21),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_40),
.Y(n_43)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_36),
.Y(n_50)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_27),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_36),
.A2(n_15),
.B1(n_25),
.B2(n_19),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_41),
.A2(n_48),
.B1(n_37),
.B2(n_35),
.Y(n_79)
);

NOR2x1_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_29),
.B1(n_23),
.B2(n_25),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_30),
.B1(n_22),
.B2(n_28),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_47),
.A2(n_54),
.B1(n_37),
.B2(n_50),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_36),
.A2(n_15),
.B1(n_19),
.B2(n_27),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_22),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_34),
.Y(n_62)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_30),
.B1(n_22),
.B2(n_28),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

BUFx4f_ASAP7_75t_SL g59 ( 
.A(n_52),
.Y(n_59)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_53),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_60),
.B(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_66),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_64),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_34),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_40),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_40),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_67),
.B(n_71),
.Y(n_90)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

NAND2x1_ASAP7_75t_SL g99 ( 
.A(n_68),
.B(n_70),
.Y(n_99)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_72),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_49),
.A2(n_33),
.B(n_31),
.C(n_24),
.Y(n_73)
);

FAx1_ASAP7_75t_SL g95 ( 
.A(n_73),
.B(n_80),
.CI(n_22),
.CON(n_95),
.SN(n_95)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_46),
.B(n_31),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_78),
.B(n_55),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_79),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_L g80 ( 
.A1(n_48),
.A2(n_33),
.B(n_24),
.Y(n_80)
);

MAJx2_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_41),
.C(n_35),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_71),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_37),
.B1(n_44),
.B2(n_56),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_86),
.A2(n_50),
.B1(n_47),
.B2(n_74),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_59),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_92),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_55),
.B(n_1),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_91),
.A2(n_95),
.B(n_96),
.Y(n_128)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_60),
.A2(n_33),
.B1(n_44),
.B2(n_45),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_94),
.A2(n_50),
.B1(n_72),
.B2(n_77),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_35),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_106),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_65),
.A2(n_51),
.B1(n_56),
.B2(n_44),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_103),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_105),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_54),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_86),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_107),
.B(n_109),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_81),
.A2(n_70),
.B(n_65),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_108),
.A2(n_125),
.B(n_30),
.Y(n_154)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_99),
.Y(n_150)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_114),
.Y(n_133)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_117),
.A2(n_106),
.B1(n_83),
.B2(n_97),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_20),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_118),
.B(n_129),
.Y(n_132)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_120),
.Y(n_146)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_85),
.A2(n_68),
.B1(n_64),
.B2(n_73),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_121),
.A2(n_100),
.B1(n_92),
.B2(n_89),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_93),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_122),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_127),
.B1(n_130),
.B2(n_100),
.Y(n_158)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_85),
.A2(n_0),
.B(n_1),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_30),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_82),
.A2(n_50),
.B1(n_59),
.B2(n_29),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_28),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_85),
.A2(n_32),
.B1(n_39),
.B2(n_38),
.Y(n_130)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_131),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_156),
.Y(n_159)
);

AO22x1_ASAP7_75t_L g135 ( 
.A1(n_126),
.A2(n_121),
.B1(n_112),
.B2(n_99),
.Y(n_135)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_111),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_136),
.B(n_153),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_138),
.A2(n_141),
.B(n_147),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_96),
.C(n_87),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_140),
.C(n_151),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_96),
.C(n_90),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_130),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_116),
.A2(n_119),
.B1(n_108),
.B2(n_128),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_142),
.A2(n_158),
.B1(n_124),
.B2(n_89),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_122),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_144),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_95),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_150),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_112),
.A2(n_95),
.B(n_99),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_83),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_38),
.C(n_32),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_38),
.C(n_32),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_154),
.A2(n_39),
.B(n_38),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_115),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_155),
.B(n_39),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_109),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_58),
.Y(n_185)
);

OA21x2_ASAP7_75t_L g160 ( 
.A1(n_146),
.A2(n_123),
.B(n_114),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_160),
.A2(n_172),
.B(n_58),
.Y(n_204)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_164),
.A2(n_178),
.B1(n_148),
.B2(n_156),
.Y(n_194)
);

A2O1A1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_146),
.A2(n_113),
.B(n_14),
.C(n_9),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_165),
.B(n_183),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_143),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_167),
.A2(n_170),
.B1(n_58),
.B2(n_1),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_158),
.A2(n_20),
.B1(n_16),
.B2(n_26),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

NOR2x1_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_147),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_171),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_149),
.A2(n_57),
.B1(n_32),
.B2(n_39),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

OA21x2_ASAP7_75t_L g172 ( 
.A1(n_135),
.A2(n_39),
.B(n_38),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_133),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_175),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_137),
.B(n_26),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_134),
.A2(n_20),
.B1(n_18),
.B2(n_26),
.Y(n_177)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_177),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_180),
.Y(n_187)
);

XNOR2x1_ASAP7_75t_SL g181 ( 
.A(n_145),
.B(n_18),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_181),
.B(n_153),
.Y(n_192)
);

NOR2x1_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_8),
.Y(n_182)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_182),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_133),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_151),
.Y(n_184)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_184),
.Y(n_196)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_140),
.C(n_139),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_190),
.C(n_193),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_150),
.Y(n_190)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_194),
.A2(n_201),
.B1(n_164),
.B2(n_173),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_141),
.C(n_132),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_198),
.B(n_206),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_163),
.A2(n_141),
.B1(n_58),
.B2(n_18),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_199),
.A2(n_170),
.B1(n_182),
.B2(n_171),
.Y(n_209)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_175),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_205),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_204),
.A2(n_172),
.B(n_178),
.Y(n_214)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_161),
.B(n_7),
.C(n_12),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_195),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_208),
.A2(n_218),
.B(n_185),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_209),
.A2(n_214),
.B1(n_216),
.B2(n_221),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_204),
.A2(n_163),
.B1(n_174),
.B2(n_184),
.Y(n_211)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_211),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_212),
.Y(n_228)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_220),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_199),
.A2(n_169),
.B1(n_181),
.B2(n_160),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_197),
.A2(n_176),
.B(n_160),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_188),
.A2(n_176),
.B1(n_159),
.B2(n_172),
.Y(n_219)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_219),
.Y(n_229)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_201),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_188),
.A2(n_179),
.B1(n_166),
.B2(n_165),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_185),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_200),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_190),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_233),
.C(n_210),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_215),
.B(n_198),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_225),
.Y(n_241)
);

INVx13_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_222),
.B(n_191),
.Y(n_226)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_193),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_216),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_232),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_189),
.C(n_196),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_235),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_226),
.B(n_206),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_236),
.B(n_243),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_242),
.C(n_230),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_221),
.Y(n_238)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_238),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_234),
.B(n_219),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_240),
.B(n_245),
.Y(n_254)
);

AOI21xp33_ASAP7_75t_L g242 ( 
.A1(n_235),
.A2(n_218),
.B(n_207),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_209),
.C(n_207),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_243),
.B(n_223),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_253),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_252),
.C(n_255),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_246),
.B(n_228),
.Y(n_250)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_250),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_241),
.C(n_229),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_244),
.B(n_234),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_229),
.C(n_227),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_251),
.A2(n_244),
.B1(n_227),
.B2(n_225),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_256),
.B(n_257),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_254),
.B(n_186),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_253),
.A2(n_214),
.B1(n_192),
.B2(n_2),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_260),
.A2(n_6),
.B1(n_10),
.B2(n_3),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_247),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_7),
.C(n_11),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_8),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_259),
.A2(n_14),
.B(n_6),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_265),
.B(n_267),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_266),
.A2(n_260),
.B1(n_8),
.B2(n_3),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_7),
.C(n_10),
.Y(n_267)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_268),
.Y(n_272)
);

AOI32xp33_ASAP7_75t_L g271 ( 
.A1(n_269),
.A2(n_263),
.A3(n_261),
.B1(n_4),
.B2(n_5),
.Y(n_271)
);

AOI321xp33_ASAP7_75t_SL g273 ( 
.A1(n_271),
.A2(n_270),
.A3(n_261),
.B1(n_4),
.B2(n_5),
.C(n_9),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_272),
.C(n_4),
.Y(n_274)
);

OAI21xp33_ASAP7_75t_L g275 ( 
.A1(n_274),
.A2(n_14),
.B(n_0),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_1),
.Y(n_276)
);


endmodule