module real_jpeg_27719_n_16 (n_333, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_333;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_0),
.A2(n_31),
.B1(n_33),
.B2(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_0),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_0),
.A2(n_27),
.B1(n_28),
.B2(n_125),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_0),
.A2(n_47),
.B1(n_48),
.B2(n_125),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_0),
.A2(n_63),
.B1(n_65),
.B2(n_125),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_1),
.Y(n_111)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_1),
.Y(n_115)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_1),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_2),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_2),
.B(n_30),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_2),
.B(n_33),
.Y(n_173)
);

AOI21xp33_ASAP7_75t_L g177 ( 
.A1(n_2),
.A2(n_33),
.B(n_173),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_2),
.A2(n_47),
.B1(n_48),
.B2(n_130),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_2),
.A2(n_60),
.B(n_63),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_2),
.B(n_88),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_2),
.A2(n_109),
.B1(n_147),
.B2(n_224),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_3),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_3),
.A2(n_31),
.B1(n_33),
.B2(n_132),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_3),
.A2(n_47),
.B1(n_48),
.B2(n_132),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_3),
.A2(n_63),
.B1(n_65),
.B2(n_132),
.Y(n_224)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_5),
.A2(n_31),
.B1(n_33),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_5),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_53),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_5),
.A2(n_47),
.B1(n_48),
.B2(n_53),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_5),
.A2(n_53),
.B1(n_63),
.B2(n_65),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_8),
.A2(n_35),
.B1(n_47),
.B2(n_48),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_8),
.A2(n_35),
.B1(n_63),
.B2(n_65),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_8),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_280)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_10),
.A2(n_31),
.B1(n_33),
.B2(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_10),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_10),
.A2(n_47),
.B1(n_48),
.B2(n_127),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_10),
.A2(n_63),
.B1(n_65),
.B2(n_127),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_127),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_11),
.A2(n_31),
.B1(n_33),
.B2(n_37),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_11),
.A2(n_37),
.B1(n_63),
.B2(n_65),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_11),
.A2(n_37),
.B1(n_47),
.B2(n_48),
.Y(n_257)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_13),
.A2(n_31),
.B1(n_33),
.B2(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_14),
.A2(n_31),
.B1(n_33),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_14),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_14),
.A2(n_50),
.B1(n_63),
.B2(n_65),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_50),
.Y(n_284)
);

INVx11_ASAP7_75t_SL g64 ( 
.A(n_15),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_95),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_93),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_80),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_19),
.B(n_80),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_70),
.C(n_74),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_20),
.A2(n_21),
.B1(n_70),
.B2(n_319),
.Y(n_323)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_39),
.B1(n_40),
.B2(n_69),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_22),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_23),
.A2(n_38),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_23),
.A2(n_38),
.B1(n_138),
.B2(n_264),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_23),
.A2(n_264),
.B(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_24),
.B(n_72),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_24),
.A2(n_84),
.B(n_85),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_24),
.A2(n_30),
.B1(n_129),
.B2(n_131),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_24),
.A2(n_85),
.B(n_284),
.Y(n_308)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_26),
.B1(n_31),
.B2(n_33),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_25),
.B(n_33),
.Y(n_144)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

HAxp5_ASAP7_75t_SL g129 ( 
.A(n_27),
.B(n_130),
.CON(n_129),
.SN(n_129)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_29),
.A2(n_31),
.B1(n_129),
.B2(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_30),
.B(n_284),
.Y(n_283)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

AOI32xp33_ASAP7_75t_L g171 ( 
.A1(n_31),
.A2(n_47),
.A3(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_171)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_34),
.A2(n_38),
.B(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_36),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_38),
.B(n_73),
.Y(n_85)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_57),
.B2(n_68),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_42),
.B(n_57),
.C(n_69),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_51),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_43),
.A2(n_76),
.B(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_49),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_44),
.B(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_52),
.Y(n_79)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_44),
.A2(n_54),
.B1(n_124),
.B2(n_126),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_44),
.A2(n_54),
.B1(n_124),
.B2(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_44),
.A2(n_54),
.B1(n_156),
.B2(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_44),
.A2(n_54),
.B1(n_78),
.B2(n_302),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_44)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_45),
.Y(n_172)
);

NAND2xp33_ASAP7_75t_SL g174 ( 
.A(n_45),
.B(n_48),
.Y(n_174)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_48),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_48),
.A2(n_61),
.B(n_130),
.C(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_51),
.A2(n_88),
.B(n_280),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_54),
.Y(n_51)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_57),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_57),
.A2(n_68),
.B1(n_75),
.B2(n_317),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_62),
.B(n_66),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_58),
.A2(n_66),
.B(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_58),
.A2(n_62),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_58),
.A2(n_181),
.B(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_58),
.A2(n_62),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_58),
.A2(n_62),
.B1(n_180),
.B2(n_199),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_58),
.A2(n_62),
.B1(n_104),
.B2(n_257),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_58),
.A2(n_120),
.B(n_257),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_62),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_65),
.Y(n_62)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_62),
.A2(n_104),
.B(n_105),
.Y(n_103)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_62),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_62),
.B(n_130),
.Y(n_222)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_65),
.B(n_229),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_67),
.B(n_121),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_70),
.C(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_70),
.A2(n_316),
.B1(n_318),
.B2(n_319),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_70),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_74),
.B(n_323),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_75),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B(n_79),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_76),
.A2(n_88),
.B(n_89),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_76),
.A2(n_79),
.B(n_89),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_81),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_86),
.B2(n_87),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI321xp33_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_312),
.A3(n_324),
.B1(n_330),
.B2(n_331),
.C(n_333),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_294),
.B(n_311),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_270),
.B(n_293),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_162),
.B(n_248),
.C(n_269),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_148),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_100),
.B(n_148),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_133),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_117),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_102),
.B(n_117),
.C(n_133),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_108),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_103),
.B(n_108),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_105),
.B(n_191),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_107),
.B(n_121),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_112),
.B(n_113),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_109),
.A2(n_112),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_109),
.A2(n_209),
.B(n_210),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_109),
.A2(n_216),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_109),
.A2(n_115),
.B(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_110),
.B(n_161),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_110),
.A2(n_114),
.B(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_110),
.A2(n_211),
.B1(n_215),
.B2(n_217),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

INVx11_ASAP7_75t_L g211 ( 
.A(n_115),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_115),
.B(n_130),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_116),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.C(n_128),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_118),
.A2(n_119),
.B1(n_122),
.B2(n_123),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_128),
.B(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_131),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_142),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_139),
.B2(n_140),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_135),
.B(n_140),
.C(n_142),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_145),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_146),
.A2(n_147),
.B(n_160),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.C(n_154),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_149),
.A2(n_150),
.B1(n_243),
.B2(n_245),
.Y(n_242)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_244),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_154),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.C(n_159),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_157),
.A2(n_158),
.B1(n_159),
.B2(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_159),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_160),
.B(n_210),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_247),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_240),
.B(n_246),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_192),
.B(n_239),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_182),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_166),
.B(n_182),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_175),
.C(n_178),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_167),
.A2(n_168),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_171),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_170),
.B(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_170),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_175),
.A2(n_176),
.B1(n_178),
.B2(n_179),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_187),
.B2(n_188),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_183),
.B(n_189),
.C(n_190),
.Y(n_241)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_233),
.B(n_238),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_212),
.B(n_232),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_202),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_195),
.B(n_202),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_200),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_196),
.A2(n_197),
.B1(n_200),
.B2(n_219),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_200),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_208),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_207),
.C(n_208),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_209),
.Y(n_217)
);

INVx11_ASAP7_75t_L g225 ( 
.A(n_211),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_220),
.B(n_231),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_218),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_214),
.B(n_218),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_226),
.B(n_230),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_222),
.B(n_223),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_234),
.B(n_235),
.Y(n_238)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_241),
.B(n_242),
.Y(n_246)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_243),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_249),
.B(n_250),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_267),
.B2(n_268),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_258),
.B2(n_259),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_259),
.C(n_268),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_256),
.Y(n_276)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_262),
.C(n_266),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_265),
.B2(n_266),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_267),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_271),
.B(n_272),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_292),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_285),
.B2(n_286),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_286),
.C(n_292),
.Y(n_295)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_276),
.B(n_279),
.C(n_281),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_281),
.B2(n_282),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_280),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_290),
.B2(n_291),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_287),
.A2(n_288),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_290),
.Y(n_305)
);

AOI21xp33_ASAP7_75t_L g321 ( 
.A1(n_288),
.A2(n_305),
.B(n_308),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_290),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_295),
.B(n_296),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_309),
.B2(n_310),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_304),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_299),
.B(n_304),
.C(n_310),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_301),
.B(n_303),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_301),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_314),
.C(n_320),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_303),
.A2(n_314),
.B1(n_315),
.B2(n_329),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_303),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_308),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_309),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_322),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_313),
.B(n_322),
.Y(n_331)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_316),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_320),
.A2(n_321),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_325),
.B(n_326),
.Y(n_330)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);


endmodule