module real_jpeg_4404_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_1),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_1),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_1),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_1),
.Y(n_143)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_1),
.Y(n_151)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_1),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g202 ( 
.A(n_1),
.Y(n_202)
);

INVx6_ASAP7_75t_L g385 ( 
.A(n_1),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_2),
.A2(n_169),
.B1(n_170),
.B2(n_173),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_2),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_3),
.A2(n_129),
.B1(n_131),
.B2(n_132),
.Y(n_128)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_3),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_3),
.A2(n_131),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_3),
.A2(n_131),
.B1(n_174),
.B2(n_307),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_3),
.A2(n_131),
.B1(n_224),
.B2(n_339),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_4),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_4),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_5),
.A2(n_70),
.B1(n_75),
.B2(n_76),
.Y(n_69)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_5),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_5),
.A2(n_75),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_6),
.A2(n_118),
.B1(n_120),
.B2(n_121),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_6),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_6),
.A2(n_120),
.B1(n_132),
.B2(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_6),
.A2(n_29),
.B1(n_120),
.B2(n_271),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g283 ( 
.A1(n_6),
.A2(n_120),
.B1(n_284),
.B2(n_286),
.Y(n_283)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_7),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_8),
.Y(n_81)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_8),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_8),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_8),
.Y(n_243)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_8),
.Y(n_310)
);

BUFx5_ASAP7_75t_L g345 ( 
.A(n_8),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_9),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_9),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_9),
.A2(n_152),
.B1(n_220),
.B2(n_224),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_9),
.A2(n_87),
.B1(n_152),
.B2(n_280),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_9),
.A2(n_152),
.B1(n_330),
.B2(n_331),
.Y(n_329)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_10),
.Y(n_140)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_10),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_10),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_11),
.A2(n_61),
.B1(n_64),
.B2(n_65),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_11),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_11),
.A2(n_64),
.B1(n_207),
.B2(n_210),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_11),
.A2(n_64),
.B1(n_250),
.B2(n_254),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_12),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_52)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_12),
.A2(n_56),
.B1(n_102),
.B2(n_125),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g343 ( 
.A1(n_12),
.A2(n_56),
.B1(n_77),
.B2(n_344),
.Y(n_343)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_13),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_14),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_14),
.A2(n_53),
.B1(n_199),
.B2(n_239),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_14),
.B(n_42),
.C(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_14),
.B(n_111),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_14),
.B(n_213),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_14),
.B(n_58),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_14),
.B(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_16),
.A2(n_45),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_16),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_16),
.A2(n_86),
.B1(n_236),
.B2(n_238),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_259),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_258),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_230),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_21),
.B(n_230),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_157),
.C(n_177),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_22),
.A2(n_23),
.B1(n_157),
.B2(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_93),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_24),
.B(n_94),
.C(n_156),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_68),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_25),
.B(n_68),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_52),
.B1(n_57),
.B2(n_59),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_26),
.A2(n_268),
.B(n_269),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_26),
.A2(n_57),
.B1(n_290),
.B2(n_329),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_26),
.A2(n_269),
.B(n_329),
.Y(n_360)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_27),
.A2(n_58),
.B1(n_60),
.B2(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_27),
.A2(n_58),
.B1(n_159),
.B2(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_27),
.B(n_270),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_41),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_33),
.B1(n_36),
.B2(n_38),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_30),
.Y(n_160)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_30),
.Y(n_271)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_31),
.Y(n_163)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_32),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g237 ( 
.A(n_32),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_32),
.Y(n_293)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_38),
.Y(n_274)
);

INVx5_ASAP7_75t_SL g332 ( 
.A(n_38),
.Y(n_332)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_41),
.A2(n_290),
.B(n_294),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_41),
.A2(n_52),
.B(n_294),
.Y(n_389)
);

AOI22x1_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_44),
.B1(n_47),
.B2(n_49),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_46),
.Y(n_286)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx11_ASAP7_75t_L g291 ( 
.A(n_55),
.Y(n_291)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_58),
.B(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g347 ( 
.A(n_62),
.Y(n_347)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AO22x2_ASAP7_75t_L g111 ( 
.A1(n_63),
.A2(n_112),
.B1(n_113),
.B2(n_115),
.Y(n_111)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_80),
.B1(n_84),
.B2(n_89),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_69),
.Y(n_216)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_70),
.Y(n_276)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_74),
.Y(n_172)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_78),
.Y(n_308)
);

BUFx8_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g212 ( 
.A(n_79),
.Y(n_212)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_80),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_80),
.B(n_283),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_80),
.A2(n_316),
.B1(n_317),
.B2(n_318),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_80),
.A2(n_206),
.B1(n_242),
.B2(n_343),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_81),
.Y(n_167)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_82),
.Y(n_344)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_85),
.A2(n_165),
.B1(n_166),
.B2(n_168),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_88),
.Y(n_176)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_127),
.B1(n_155),
.B2(n_156),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_94),
.Y(n_155)
);

AOI22x1_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_111),
.B1(n_116),
.B2(n_123),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_95),
.A2(n_218),
.B(n_228),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_95),
.A2(n_228),
.B(n_335),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_95),
.B(n_116),
.Y(n_365)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_96),
.A2(n_124),
.B1(n_229),
.B2(n_249),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_96),
.A2(n_219),
.B1(n_229),
.B2(n_364),
.Y(n_388)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_111),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_102),
.B1(n_107),
.B2(n_109),
.Y(n_97)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_98),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_101),
.Y(n_351)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_103),
.A2(n_146),
.B1(n_147),
.B2(n_149),
.Y(n_145)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_105),
.Y(n_223)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g227 ( 
.A(n_106),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_110),
.Y(n_190)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_110),
.Y(n_197)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_110),
.Y(n_253)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_110),
.Y(n_336)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_111),
.Y(n_229)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_117),
.B(n_229),
.Y(n_228)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx6_ASAP7_75t_SL g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_135),
.B1(n_145),
.B2(n_150),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_128),
.A2(n_180),
.B(n_182),
.Y(n_179)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_133),
.Y(n_192)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_135),
.A2(n_150),
.B(n_257),
.Y(n_256)
);

INVx3_ASAP7_75t_SL g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_136),
.B(n_183),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_136),
.A2(n_383),
.B(n_386),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_145),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_SL g149 ( 
.A(n_140),
.Y(n_149)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_143),
.Y(n_185)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_144),
.Y(n_146)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_145),
.B(n_199),
.Y(n_367)
);

OAI32xp33_ASAP7_75t_L g187 ( 
.A1(n_146),
.A2(n_188),
.A3(n_191),
.B1(n_193),
.B2(n_198),
.Y(n_187)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_157),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_164),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_158),
.B(n_164),
.Y(n_246)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_160),
.Y(n_330)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_165),
.A2(n_205),
.B1(n_213),
.B2(n_216),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_165),
.A2(n_168),
.B(n_241),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_165),
.A2(n_279),
.B(n_282),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_165),
.A2(n_199),
.B(n_282),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_166),
.Y(n_318)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_167),
.B(n_283),
.Y(n_282)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_171),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_172),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_177),
.B(n_404),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_186),
.C(n_217),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_178),
.A2(n_179),
.B1(n_217),
.B2(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_181),
.B(n_183),
.Y(n_257)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_186),
.B(n_398),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_203),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_187),
.A2(n_203),
.B1(n_204),
.B2(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_187),
.Y(n_376)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI21xp33_ASAP7_75t_SL g383 ( 
.A1(n_198),
.A2(n_199),
.B(n_384),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

OAI21xp33_ASAP7_75t_SL g335 ( 
.A1(n_199),
.A2(n_336),
.B(n_337),
.Y(n_335)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_212),
.Y(n_281)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_217),
.Y(n_399)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx4_ASAP7_75t_SL g221 ( 
.A(n_222),
.Y(n_221)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_227),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_229),
.A2(n_364),
.B(n_365),
.Y(n_363)
);

BUFx24_ASAP7_75t_SL g414 ( 
.A(n_230),
.Y(n_414)
);

FAx1_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_232),
.CI(n_245),
.CON(n_230),
.SN(n_230)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_240),
.B2(n_244),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx3_ASAP7_75t_SL g236 ( 
.A(n_237),
.Y(n_236)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_237),
.Y(n_239)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

NAND2xp33_ASAP7_75t_SL g352 ( 
.A(n_239),
.B(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_240),
.Y(n_244)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_256),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_251),
.Y(n_250)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

AOI32xp33_ASAP7_75t_L g346 ( 
.A1(n_254),
.A2(n_338),
.A3(n_347),
.B1(n_348),
.B2(n_352),
.Y(n_346)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_257),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_392),
.B(n_411),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

AOI21x1_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_371),
.B(n_391),
.Y(n_261)
);

AO21x1_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_355),
.B(n_370),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_323),
.B(n_354),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_297),
.B(n_322),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_277),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_266),
.B(n_277),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_272),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_267),
.A2(n_272),
.B1(n_273),
.B2(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_267),
.Y(n_320)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_287),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_278),
.B(n_288),
.C(n_296),
.Y(n_324)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_279),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_284),
.Y(n_301)
);

INVx6_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_295),
.B2(n_296),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx5_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_314),
.B(n_321),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_304),
.B(n_313),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_303),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_312),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_312),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_309),
.B(n_311),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_306),
.Y(n_316)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_311),
.A2(n_342),
.B(n_345),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_319),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_319),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_324),
.B(n_325),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_340),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_328),
.B1(n_333),
.B2(n_334),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_328),
.B(n_333),
.C(n_340),
.Y(n_356)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVxp33_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_346),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_341),
.B(n_346),
.Y(n_361)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx8_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_357),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_356),
.B(n_357),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_358),
.A2(n_359),
.B1(n_362),
.B2(n_369),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_360),
.B(n_361),
.C(n_369),
.Y(n_372)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_362),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g362 ( 
.A(n_363),
.B(n_366),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_363),
.B(n_367),
.C(n_368),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_368),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_372),
.B(n_373),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_380),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_375),
.A2(n_377),
.B1(n_378),
.B2(n_379),
.Y(n_374)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_375),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_377),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_377),
.B(n_378),
.C(n_380),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_381),
.A2(n_382),
.B1(n_387),
.B2(n_390),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_381),
.B(n_388),
.C(n_389),
.Y(n_402)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx8_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_387),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_388),
.B(n_389),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_394),
.B(n_406),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_395),
.A2(n_412),
.B(n_413),
.Y(n_411)
);

NOR2x1_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_403),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_396),
.B(n_403),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_400),
.C(n_402),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_397),
.B(n_409),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_400),
.A2(n_401),
.B1(n_402),
.B2(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_402),
.Y(n_410)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_408),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_407),
.B(n_408),
.Y(n_412)
);


endmodule