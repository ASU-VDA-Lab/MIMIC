module fake_jpeg_29465_n_530 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_530);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_530;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx24_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_SL g37 ( 
.A(n_5),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_45),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_52),
.B(n_64),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_45),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_53),
.B(n_76),
.Y(n_126)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_55),
.Y(n_131)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_26),
.B(n_18),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx11_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_70),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_72),
.Y(n_157)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_73),
.Y(n_150)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_75),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_26),
.B(n_18),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_80),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_85),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_87),
.Y(n_151)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_89),
.Y(n_147)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_91),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_93),
.Y(n_156)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_94),
.Y(n_160)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_99),
.Y(n_108)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_100),
.B(n_101),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_34),
.B(n_48),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_48),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_120),
.B(n_124),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_67),
.A2(n_22),
.B1(n_49),
.B2(n_33),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_121),
.A2(n_127),
.B1(n_129),
.B2(n_146),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_76),
.B(n_34),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_51),
.A2(n_41),
.B1(n_49),
.B2(n_33),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_67),
.A2(n_22),
.B1(n_49),
.B2(n_33),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_63),
.B(n_22),
.C(n_41),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_133),
.B(n_136),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_52),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_82),
.B(n_30),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_137),
.B(n_162),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_55),
.A2(n_49),
.B1(n_36),
.B2(n_47),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_62),
.Y(n_149)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_74),
.A2(n_36),
.B1(n_47),
.B2(n_44),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_158),
.A2(n_159),
.B1(n_161),
.B2(n_83),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_70),
.A2(n_92),
.B1(n_81),
.B2(n_79),
.Y(n_159)
);

OA22x2_ASAP7_75t_L g161 ( 
.A1(n_65),
.A2(n_19),
.B1(n_47),
.B2(n_44),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_82),
.B(n_17),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_100),
.B(n_44),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_163),
.B(n_29),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_36),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_164),
.B(n_169),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_165),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_126),
.A2(n_161),
.B(n_110),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_166),
.A2(n_19),
.B(n_151),
.Y(n_240)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_113),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_167),
.Y(n_252)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_125),
.Y(n_168)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_168),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_126),
.B(n_40),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_145),
.A2(n_84),
.B1(n_68),
.B2(n_23),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_172),
.A2(n_183),
.B1(n_213),
.B2(n_138),
.Y(n_247)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_173),
.Y(n_256)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_128),
.Y(n_174)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_174),
.Y(n_231)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_117),
.Y(n_175)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_175),
.Y(n_225)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_119),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_176),
.Y(n_265)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_177),
.Y(n_263)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_178),
.Y(n_267)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_113),
.Y(n_179)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_179),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_181),
.B(n_191),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_135),
.Y(n_182)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_182),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_145),
.A2(n_42),
.B1(n_28),
.B2(n_23),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_184),
.Y(n_243)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_117),
.Y(n_185)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_185),
.Y(n_245)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

INVx13_ASAP7_75t_L g266 ( 
.A(n_186),
.Y(n_266)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_187),
.Y(n_250)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_122),
.Y(n_188)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_188),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_190),
.A2(n_50),
.B1(n_1),
.B2(n_2),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_42),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_108),
.B(n_42),
.Y(n_192)
);

FAx1_ASAP7_75t_SL g251 ( 
.A(n_192),
.B(n_203),
.CI(n_216),
.CON(n_251),
.SN(n_251)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_132),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_194),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_150),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_115),
.B(n_40),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_196),
.B(n_219),
.Y(n_227)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_123),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_197),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_111),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_198),
.B(n_199),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_109),
.B(n_17),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_150),
.Y(n_200)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_200),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_114),
.B(n_35),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_201),
.B(n_202),
.Y(n_262)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_154),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_107),
.B(n_40),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_111),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_204),
.B(n_205),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_116),
.B(n_24),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_157),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_206),
.Y(n_235)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_149),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_207),
.Y(n_261)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_143),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_218),
.Y(n_242)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_143),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_209),
.Y(n_248)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_130),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_210),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_105),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_211),
.Y(n_232)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_106),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_212),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_152),
.A2(n_23),
.B1(n_28),
.B2(n_29),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_112),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_214),
.A2(n_217),
.B1(n_104),
.B2(n_142),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_118),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_215),
.B(n_222),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_107),
.B(n_29),
.Y(n_216)
);

INVx8_ASAP7_75t_L g217 ( 
.A(n_141),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_121),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_130),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_158),
.B(n_35),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_220),
.B(n_223),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_151),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_221),
.A2(n_152),
.B1(n_104),
.B2(n_19),
.Y(n_226)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_160),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_144),
.B(n_104),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_226),
.B(n_254),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_229),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_191),
.A2(n_129),
.B1(n_71),
.B2(n_102),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_233),
.A2(n_236),
.B1(n_241),
.B2(n_273),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_218),
.A2(n_166),
.B1(n_164),
.B2(n_192),
.Y(n_236)
);

AOI21xp33_ASAP7_75t_L g237 ( 
.A1(n_169),
.A2(n_28),
.B(n_19),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_237),
.B(n_4),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_189),
.A2(n_102),
.B1(n_142),
.B2(n_141),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_238),
.A2(n_260),
.B1(n_264),
.B2(n_270),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_240),
.B(n_35),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_190),
.A2(n_155),
.B1(n_134),
.B2(n_131),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_180),
.B(n_87),
.C(n_86),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_244),
.B(n_249),
.C(n_179),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_247),
.A2(n_175),
.B1(n_212),
.B2(n_217),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_195),
.B(n_155),
.C(n_134),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_215),
.A2(n_32),
.B1(n_103),
.B2(n_131),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_203),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_216),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_171),
.B(n_3),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_272),
.B(n_3),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_222),
.A2(n_32),
.B1(n_35),
.B2(n_24),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_253),
.B(n_188),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_276),
.B(n_270),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_277),
.B(n_282),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_227),
.B(n_197),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_278),
.B(n_281),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_251),
.B(n_177),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_279),
.B(n_286),
.Y(n_330)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_248),
.Y(n_280)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_280),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_259),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_259),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_225),
.Y(n_283)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_283),
.Y(n_324)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_225),
.Y(n_285)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_285),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_251),
.B(n_178),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_287),
.B(n_289),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_227),
.B(n_209),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_288),
.B(n_298),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_251),
.B(n_174),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_250),
.Y(n_290)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_290),
.Y(n_355)
);

INVx8_ASAP7_75t_L g292 ( 
.A(n_239),
.Y(n_292)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_292),
.Y(n_332)
);

OAI32xp33_ASAP7_75t_L g293 ( 
.A1(n_236),
.A2(n_168),
.A3(n_184),
.B1(n_200),
.B2(n_186),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_293),
.B(n_299),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_253),
.B(n_255),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_294),
.B(n_295),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_167),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_248),
.Y(n_296)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_296),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_226),
.Y(n_298)
);

OA21x2_ASAP7_75t_L g300 ( 
.A1(n_240),
.A2(n_210),
.B(n_173),
.Y(n_300)
);

AO21x1_ASAP7_75t_L g353 ( 
.A1(n_300),
.A2(n_305),
.B(n_315),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_241),
.A2(n_214),
.B1(n_165),
.B2(n_170),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_301),
.A2(n_304),
.B1(n_312),
.B2(n_320),
.Y(n_352)
);

INVxp33_ASAP7_75t_SL g302 ( 
.A(n_235),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_302),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_271),
.B(n_32),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_303),
.B(n_307),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_233),
.A2(n_207),
.B1(n_170),
.B2(n_182),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_250),
.Y(n_306)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_306),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_242),
.B(n_32),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_260),
.A2(n_32),
.B1(n_35),
.B2(n_24),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_308),
.A2(n_256),
.B(n_263),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_259),
.Y(n_309)
);

NOR3xp33_ASAP7_75t_L g328 ( 
.A(n_309),
.B(n_232),
.C(n_275),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_242),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_310),
.B(n_318),
.Y(n_354)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_245),
.Y(n_311)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_311),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_269),
.A2(n_258),
.B1(n_262),
.B2(n_249),
.Y(n_312)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_257),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_313),
.Y(n_344)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_230),
.Y(n_316)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_316),
.Y(n_356)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_245),
.Y(n_317)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_317),
.Y(n_360)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_243),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_243),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_319),
.B(n_321),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_244),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_264),
.B(n_32),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_268),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_322),
.A2(n_231),
.B1(n_246),
.B2(n_266),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_284),
.A2(n_265),
.B1(n_232),
.B2(n_275),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_323),
.A2(n_337),
.B1(n_358),
.B2(n_322),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_310),
.A2(n_234),
.B(n_235),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_325),
.B(n_339),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_328),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_336),
.B(n_303),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_314),
.A2(n_235),
.B1(n_254),
.B2(n_268),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_305),
.A2(n_252),
.B(n_272),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_276),
.B(n_274),
.C(n_252),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_341),
.B(n_345),
.C(n_314),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_286),
.B(n_256),
.C(n_224),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_279),
.A2(n_228),
.B(n_224),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_348),
.A2(n_349),
.B(n_362),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_287),
.A2(n_228),
.B(n_257),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_350),
.A2(n_357),
.B1(n_359),
.B2(n_291),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_289),
.B(n_267),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_351),
.B(n_10),
.C(n_11),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_297),
.A2(n_239),
.B1(n_267),
.B2(n_263),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_314),
.A2(n_231),
.B1(n_230),
.B2(n_246),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_297),
.A2(n_298),
.B1(n_277),
.B2(n_304),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_361),
.B(n_282),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_300),
.A2(n_261),
.B(n_266),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_364),
.B(n_388),
.C(n_389),
.Y(n_401)
);

NAND3xp33_ASAP7_75t_L g365 ( 
.A(n_326),
.B(n_295),
.C(n_294),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_365),
.Y(n_410)
);

OAI21xp33_ASAP7_75t_SL g419 ( 
.A1(n_366),
.A2(n_397),
.B(n_342),
.Y(n_419)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_347),
.Y(n_367)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_367),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_368),
.A2(n_373),
.B1(n_374),
.B2(n_375),
.Y(n_424)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_347),
.Y(n_369)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_369),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_370),
.B(n_341),
.Y(n_407)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_360),
.Y(n_371)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_371),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_323),
.A2(n_291),
.B1(n_312),
.B2(n_301),
.Y(n_372)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_372),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_352),
.A2(n_293),
.B1(n_300),
.B2(n_283),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_352),
.A2(n_285),
.B1(n_308),
.B2(n_290),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_359),
.A2(n_311),
.B1(n_317),
.B2(n_307),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_377),
.A2(n_335),
.B1(n_349),
.B2(n_348),
.Y(n_402)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_360),
.Y(n_378)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_378),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_340),
.B(n_320),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_380),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_354),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g409 ( 
.A(n_381),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_333),
.A2(n_346),
.B1(n_357),
.B2(n_350),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_382),
.B(n_383),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_346),
.A2(n_313),
.B1(n_321),
.B2(n_318),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_340),
.B(n_319),
.Y(n_384)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_384),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_346),
.A2(n_292),
.B1(n_296),
.B2(n_280),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_385),
.B(n_386),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_343),
.A2(n_316),
.B1(n_261),
.B2(n_7),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_351),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_387)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_387),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_330),
.B(n_35),
.C(n_24),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_330),
.B(n_24),
.C(n_7),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_335),
.A2(n_24),
.B1(n_8),
.B2(n_9),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_390),
.A2(n_10),
.B(n_11),
.Y(n_428)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_338),
.Y(n_392)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_392),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_336),
.B(n_4),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_393),
.B(n_345),
.C(n_331),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_362),
.A2(n_8),
.B(n_9),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_394),
.A2(n_354),
.B(n_342),
.Y(n_404)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_338),
.Y(n_395)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_395),
.Y(n_416)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_324),
.Y(n_396)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_396),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_331),
.B(n_8),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_398),
.B(n_339),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_402),
.A2(n_411),
.B1(n_421),
.B2(n_422),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_SL g403 ( 
.A1(n_391),
.A2(n_344),
.B1(n_332),
.B2(n_329),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_403),
.A2(n_428),
.B1(n_390),
.B2(n_386),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_404),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_407),
.B(n_375),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_408),
.B(n_427),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_377),
.A2(n_353),
.B1(n_363),
.B2(n_325),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_417),
.B(n_389),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_419),
.A2(n_371),
.B1(n_378),
.B2(n_369),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_379),
.A2(n_353),
.B1(n_363),
.B2(n_337),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_373),
.A2(n_355),
.B1(n_332),
.B2(n_327),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_364),
.B(n_358),
.C(n_356),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_425),
.B(n_388),
.C(n_393),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_370),
.B(n_361),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_415),
.Y(n_429)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_429),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_430),
.B(n_435),
.C(n_443),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_399),
.B(n_397),
.Y(n_432)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_432),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_433),
.B(n_439),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_434),
.A2(n_413),
.B1(n_423),
.B2(n_414),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_407),
.B(n_384),
.C(n_382),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_409),
.B(n_391),
.Y(n_436)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_436),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_427),
.B(n_376),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_415),
.Y(n_440)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_440),
.Y(n_466)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_416),
.Y(n_441)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_441),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_442),
.B(n_445),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_408),
.B(n_376),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_366),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_444),
.B(n_450),
.C(n_400),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_424),
.A2(n_368),
.B1(n_374),
.B2(n_367),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_446),
.A2(n_454),
.B1(n_400),
.B2(n_411),
.Y(n_456)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_416),
.Y(n_447)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_447),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_410),
.B(n_387),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_448),
.B(n_451),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_399),
.B(n_396),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_449),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_421),
.B(n_383),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_426),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_401),
.B(n_398),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_452),
.B(n_453),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_401),
.B(n_385),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_418),
.A2(n_420),
.B1(n_413),
.B2(n_422),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_456),
.A2(n_431),
.B1(n_450),
.B2(n_444),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_459),
.B(n_431),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_453),
.B(n_402),
.C(n_417),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_461),
.B(n_467),
.C(n_472),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_437),
.A2(n_412),
.B(n_428),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_463),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_464),
.A2(n_334),
.B1(n_356),
.B2(n_13),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_438),
.B(n_404),
.C(n_406),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_437),
.B(n_405),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_471),
.B(n_474),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_438),
.B(n_426),
.C(n_412),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_445),
.B(n_394),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_476),
.A2(n_464),
.B1(n_459),
.B2(n_472),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_473),
.B(n_435),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_477),
.B(n_481),
.Y(n_504)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_469),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_478),
.B(n_482),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_473),
.B(n_439),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_457),
.B(n_443),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_483),
.B(n_485),
.Y(n_496)
);

XOR2x1_ASAP7_75t_L g484 ( 
.A(n_460),
.B(n_454),
.Y(n_484)
);

FAx1_ASAP7_75t_SL g500 ( 
.A(n_484),
.B(n_455),
.CI(n_458),
.CON(n_500),
.SN(n_500)
);

AOI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_462),
.A2(n_442),
.B1(n_446),
.B2(n_430),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_457),
.B(n_452),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_486),
.B(n_489),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_461),
.B(n_395),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_488),
.B(n_467),
.C(n_455),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_465),
.A2(n_392),
.B1(n_334),
.B2(n_327),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_490),
.A2(n_475),
.B1(n_468),
.B2(n_466),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_R g491 ( 
.A(n_463),
.B(n_10),
.Y(n_491)
);

NOR2x1_ASAP7_75t_L g501 ( 
.A(n_491),
.B(n_466),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_479),
.A2(n_480),
.B(n_471),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_492),
.A2(n_499),
.B(n_487),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_493),
.B(n_501),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_495),
.B(n_503),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_483),
.A2(n_460),
.B1(n_470),
.B2(n_475),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_497),
.B(n_498),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_491),
.A2(n_474),
.B(n_469),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_500),
.B(n_485),
.Y(n_508)
);

OAI321xp33_ASAP7_75t_L g503 ( 
.A1(n_484),
.A2(n_468),
.A3(n_12),
.B1(n_13),
.B2(n_15),
.C(n_16),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_504),
.B(n_487),
.C(n_488),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_505),
.B(n_511),
.Y(n_517)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_508),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_509),
.B(n_510),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_496),
.B(n_477),
.C(n_481),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_494),
.B(n_500),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_497),
.B(n_502),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_513),
.B(n_496),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_506),
.A2(n_492),
.B(n_501),
.Y(n_514)
);

AOI21x1_ASAP7_75t_L g523 ( 
.A1(n_514),
.A2(n_507),
.B(n_504),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_512),
.A2(n_499),
.B1(n_493),
.B2(n_498),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_518),
.B(n_519),
.Y(n_520)
);

OAI21xp33_ASAP7_75t_L g521 ( 
.A1(n_515),
.A2(n_507),
.B(n_500),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_521),
.B(n_522),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_517),
.B(n_505),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_523),
.B(n_518),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_525),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_526),
.B(n_524),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_527),
.A2(n_520),
.B(n_514),
.Y(n_528)
);

NAND3xp33_ASAP7_75t_L g529 ( 
.A(n_528),
.B(n_516),
.C(n_12),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_529),
.A2(n_10),
.B(n_13),
.Y(n_530)
);


endmodule