module fake_jpeg_21681_n_106 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_106);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_106;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx6_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_7),
.Y(n_11)
);

INVx1_ASAP7_75t_SL g12 ( 
.A(n_9),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_6),
.B(n_5),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx11_ASAP7_75t_SL g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_25),
.Y(n_36)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_12),
.B(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_16),
.C(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_29),
.B(n_24),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_27),
.A2(n_10),
.B1(n_17),
.B2(n_20),
.Y(n_34)
);

OAI32xp33_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_20),
.A3(n_24),
.B1(n_10),
.B2(n_26),
.Y(n_40)
);

O2A1O1Ixp33_ASAP7_75t_L g37 ( 
.A1(n_32),
.A2(n_25),
.B(n_23),
.C(n_15),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_17),
.B1(n_30),
.B2(n_31),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_11),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_11),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_30),
.B1(n_29),
.B2(n_31),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_36),
.B(n_13),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_18),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_26),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_46),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_28),
.B(n_26),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_16),
.C(n_14),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_55),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_30),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_58),
.B(n_59),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_28),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_44),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_67),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_47),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_62),
.C(n_65),
.Y(n_79)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_56),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_70),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_56),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_78),
.Y(n_86)
);

A2O1A1O1Ixp25_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_53),
.B(n_58),
.C(n_51),
.D(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_79),
.Y(n_83)
);

OAI32xp33_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_53),
.A3(n_60),
.B1(n_40),
.B2(n_55),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_46),
.C(n_50),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_63),
.C(n_21),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_75),
.A2(n_71),
.B1(n_68),
.B2(n_43),
.Y(n_81)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_80),
.A2(n_73),
.B1(n_77),
.B2(n_76),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_31),
.B1(n_2),
.B2(n_3),
.Y(n_91)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_85),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_67),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_87),
.B(n_21),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_88),
.B(n_91),
.Y(n_96)
);

MAJx2_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_86),
.C(n_81),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_14),
.Y(n_94)
);

AOI322xp5_ASAP7_75t_L g93 ( 
.A1(n_90),
.A2(n_87),
.A3(n_21),
.B1(n_9),
.B2(n_6),
.C1(n_7),
.C2(n_19),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_93),
.B(n_94),
.Y(n_100)
);

OAI21xp33_ASAP7_75t_L g95 ( 
.A1(n_90),
.A2(n_92),
.B(n_3),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_1),
.B(n_4),
.Y(n_97)
);

NOR3xp33_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_4),
.C(n_98),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_33),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_14),
.C(n_33),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_4),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_99),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_33),
.C(n_101),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_100),
.B(n_33),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_104),
.B(n_105),
.Y(n_106)
);


endmodule