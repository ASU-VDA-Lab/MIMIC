module real_aes_2033_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_250;
wire n_85;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_552;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
AO22x2_ASAP7_75t_L g103 ( .A1(n_0), .A2(n_52), .B1(n_93), .B2(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g192 ( .A(n_1), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_2), .B(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g178 ( .A(n_3), .Y(n_178) );
AO22x2_ASAP7_75t_L g100 ( .A1(n_4), .A2(n_20), .B1(n_93), .B2(n_101), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_5), .Y(n_289) );
AOI22xp33_ASAP7_75t_L g139 ( .A1(n_6), .A2(n_49), .B1(n_140), .B2(n_143), .Y(n_139) );
AOI22xp5_ASAP7_75t_L g118 ( .A1(n_7), .A2(n_14), .B1(n_119), .B2(n_123), .Y(n_118) );
INVx2_ASAP7_75t_L g207 ( .A(n_8), .Y(n_207) );
INVx1_ASAP7_75t_L g253 ( .A(n_9), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g153 ( .A1(n_10), .A2(n_68), .B1(n_154), .B2(n_158), .Y(n_153) );
INVx1_ASAP7_75t_L g172 ( .A(n_11), .Y(n_172) );
AOI22xp5_ASAP7_75t_L g162 ( .A1(n_12), .A2(n_72), .B1(n_163), .B2(n_167), .Y(n_162) );
INVx1_ASAP7_75t_SL g225 ( .A(n_13), .Y(n_225) );
INVx1_ASAP7_75t_L g250 ( .A(n_15), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g333 ( .A(n_16), .B(n_228), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g105 ( .A1(n_17), .A2(n_24), .B1(n_106), .B2(n_113), .Y(n_105) );
AOI33xp33_ASAP7_75t_L g301 ( .A1(n_18), .A2(n_37), .A3(n_213), .B1(n_221), .B2(n_302), .B3(n_303), .Y(n_301) );
INVx1_ASAP7_75t_L g282 ( .A(n_19), .Y(n_282) );
OAI221xp5_ASAP7_75t_L g184 ( .A1(n_20), .A2(n_52), .B1(n_55), .B2(n_185), .C(n_187), .Y(n_184) );
OR2x2_ASAP7_75t_L g208 ( .A(n_21), .B(n_69), .Y(n_208) );
OA21x2_ASAP7_75t_L g238 ( .A1(n_21), .A2(n_69), .B(n_207), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_22), .B(n_211), .Y(n_210) );
INVx3_ASAP7_75t_L g93 ( .A(n_23), .Y(n_93) );
INVx1_ASAP7_75t_SL g94 ( .A(n_25), .Y(n_94) );
INVx1_ASAP7_75t_L g194 ( .A(n_26), .Y(n_194) );
AND2x2_ASAP7_75t_L g216 ( .A(n_26), .B(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g234 ( .A(n_26), .B(n_192), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g284 ( .A(n_27), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_28), .B(n_211), .Y(n_309) );
AOI22xp5_ASAP7_75t_L g326 ( .A1(n_29), .A2(n_237), .B1(n_243), .B2(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_30), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_31), .B(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g85 ( .A(n_32), .B(n_86), .Y(n_85) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_33), .B(n_271), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_34), .B(n_228), .Y(n_274) );
AO22x2_ASAP7_75t_L g96 ( .A1(n_35), .A2(n_55), .B1(n_93), .B2(n_97), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_36), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_38), .B(n_228), .Y(n_313) );
INVx1_ASAP7_75t_L g214 ( .A(n_39), .Y(n_214) );
INVx1_ASAP7_75t_L g230 ( .A(n_39), .Y(n_230) );
AND2x2_ASAP7_75t_L g314 ( .A(n_40), .B(n_205), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g146 ( .A1(n_41), .A2(n_67), .B1(n_147), .B2(n_150), .Y(n_146) );
AOI221xp5_ASAP7_75t_L g272 ( .A1(n_42), .A2(n_57), .B1(n_211), .B2(n_219), .C(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_43), .B(n_211), .Y(n_266) );
INVx1_ASAP7_75t_L g95 ( .A(n_44), .Y(n_95) );
INVx1_ASAP7_75t_L g81 ( .A(n_45), .Y(n_81) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_46), .B(n_237), .Y(n_291) );
AOI21xp5_ASAP7_75t_SL g262 ( .A1(n_47), .A2(n_219), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g246 ( .A(n_48), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_48), .A2(n_82), .B1(n_83), .B2(n_246), .Y(n_559) );
INVx1_ASAP7_75t_L g312 ( .A(n_50), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_51), .A2(n_219), .B(n_311), .Y(n_310) );
INVxp33_ASAP7_75t_L g189 ( .A(n_52), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g129 ( .A1(n_53), .A2(n_66), .B1(n_130), .B2(n_134), .Y(n_129) );
INVx1_ASAP7_75t_L g217 ( .A(n_54), .Y(n_217) );
INVx1_ASAP7_75t_L g232 ( .A(n_54), .Y(n_232) );
INVxp67_ASAP7_75t_L g188 ( .A(n_55), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_56), .B(n_211), .Y(n_304) );
AND2x2_ASAP7_75t_L g235 ( .A(n_58), .B(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g247 ( .A(n_59), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_60), .A2(n_219), .B(n_224), .Y(n_218) );
AOI22xp33_ASAP7_75t_SL g566 ( .A1(n_61), .A2(n_82), .B1(n_83), .B2(n_567), .Y(n_566) );
CKINVDCx20_ASAP7_75t_R g567 ( .A(n_61), .Y(n_567) );
A2O1A1Ixp33_ASAP7_75t_L g331 ( .A1(n_62), .A2(n_219), .B(n_296), .C(n_332), .Y(n_331) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_63), .A2(n_177), .B1(n_178), .B2(n_179), .Y(n_176) );
INVx1_ASAP7_75t_L g179 ( .A(n_63), .Y(n_179) );
AND2x2_ASAP7_75t_SL g260 ( .A(n_64), .B(n_236), .Y(n_260) );
AOI22xp5_ASAP7_75t_L g298 ( .A1(n_65), .A2(n_219), .B1(n_299), .B2(n_300), .Y(n_298) );
INVx1_ASAP7_75t_L g264 ( .A(n_70), .Y(n_264) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_71), .A2(n_172), .B1(n_173), .B2(n_174), .Y(n_171) );
INVx1_ASAP7_75t_L g173 ( .A(n_71), .Y(n_173) );
AND2x2_ASAP7_75t_L g305 ( .A(n_73), .B(n_236), .Y(n_305) );
A2O1A1Ixp33_ASAP7_75t_L g279 ( .A1(n_74), .A2(n_280), .B(n_281), .C(n_283), .Y(n_279) );
BUFx2_ASAP7_75t_SL g186 ( .A(n_75), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_76), .B(n_228), .Y(n_265) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_181), .B1(n_195), .B2(n_555), .C(n_558), .Y(n_77) );
XNOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_170), .Y(n_78) );
AOI22xp33_ASAP7_75t_SL g79 ( .A1(n_80), .A2(n_81), .B1(n_82), .B2(n_83), .Y(n_79) );
CKINVDCx16_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
INVx2_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
OR2x2_ASAP7_75t_L g83 ( .A(n_84), .B(n_138), .Y(n_83) );
NAND4xp25_ASAP7_75t_SL g84 ( .A(n_85), .B(n_105), .C(n_118), .D(n_129), .Y(n_84) );
HB1xp67_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
INVx3_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
INVx6_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
AND2x2_ASAP7_75t_L g89 ( .A(n_90), .B(n_98), .Y(n_89) );
AND2x4_ASAP7_75t_L g115 ( .A(n_90), .B(n_116), .Y(n_115) );
AND2x4_ASAP7_75t_L g136 ( .A(n_90), .B(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g90 ( .A(n_91), .B(n_96), .Y(n_90) );
AND2x2_ASAP7_75t_L g111 ( .A(n_91), .B(n_112), .Y(n_111) );
HB1xp67_ASAP7_75t_L g128 ( .A(n_91), .Y(n_128) );
INVx2_ASAP7_75t_L g133 ( .A(n_91), .Y(n_133) );
OAI22x1_ASAP7_75t_L g91 ( .A1(n_92), .A2(n_93), .B1(n_94), .B2(n_95), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g97 ( .A(n_93), .Y(n_97) );
INVx2_ASAP7_75t_L g101 ( .A(n_93), .Y(n_101) );
INVx1_ASAP7_75t_L g104 ( .A(n_93), .Y(n_104) );
INVx2_ASAP7_75t_L g112 ( .A(n_96), .Y(n_112) );
AND2x2_ASAP7_75t_L g132 ( .A(n_96), .B(n_133), .Y(n_132) );
BUFx2_ASAP7_75t_L g161 ( .A(n_96), .Y(n_161) );
AND2x4_ASAP7_75t_L g142 ( .A(n_98), .B(n_111), .Y(n_142) );
AND2x4_ASAP7_75t_L g149 ( .A(n_98), .B(n_145), .Y(n_149) );
AND2x2_ASAP7_75t_L g166 ( .A(n_98), .B(n_132), .Y(n_166) );
AND2x4_ASAP7_75t_L g98 ( .A(n_99), .B(n_102), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
INVx1_ASAP7_75t_L g110 ( .A(n_100), .Y(n_110) );
AND2x4_ASAP7_75t_L g122 ( .A(n_100), .B(n_102), .Y(n_122) );
AND2x2_ASAP7_75t_L g127 ( .A(n_100), .B(n_103), .Y(n_127) );
INVxp67_ASAP7_75t_L g137 ( .A(n_102), .Y(n_137) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x2_ASAP7_75t_L g109 ( .A(n_103), .B(n_110), .Y(n_109) );
BUFx6f_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
AND2x4_ASAP7_75t_L g152 ( .A(n_109), .B(n_145), .Y(n_152) );
AND2x2_ASAP7_75t_L g157 ( .A(n_109), .B(n_132), .Y(n_157) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_110), .Y(n_117) );
AND2x2_ASAP7_75t_L g121 ( .A(n_111), .B(n_122), .Y(n_121) );
AND2x4_ASAP7_75t_L g145 ( .A(n_112), .B(n_133), .Y(n_145) );
BUFx2_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
BUFx6f_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AND2x4_ASAP7_75t_L g131 ( .A(n_122), .B(n_132), .Y(n_131) );
AND2x4_ASAP7_75t_L g169 ( .A(n_122), .B(n_145), .Y(n_169) );
BUFx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx3_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_128), .Y(n_126) );
AND2x4_ASAP7_75t_L g144 ( .A(n_127), .B(n_145), .Y(n_144) );
AND2x4_ASAP7_75t_L g160 ( .A(n_127), .B(n_161), .Y(n_160) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_SL g134 ( .A(n_135), .Y(n_134) );
INVx6_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
NAND4xp25_ASAP7_75t_L g138 ( .A(n_139), .B(n_146), .C(n_153), .D(n_162), .Y(n_138) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx6_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
BUFx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx4_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx8_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx8_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx5_ASAP7_75t_SL g159 ( .A(n_160), .Y(n_159) );
BUFx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
HB1xp67_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
OAI22xp5_ASAP7_75t_SL g170 ( .A1(n_171), .A2(n_175), .B1(n_176), .B2(n_180), .Y(n_170) );
CKINVDCx16_ASAP7_75t_R g180 ( .A(n_171), .Y(n_180) );
INVx1_ASAP7_75t_L g174 ( .A(n_172), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_SL g273 ( .A1(n_178), .A2(n_226), .B(n_233), .C(n_274), .Y(n_273) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_182), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_183), .Y(n_182) );
AND3x1_ASAP7_75t_SL g183 ( .A(n_184), .B(n_190), .C(n_193), .Y(n_183) );
INVxp67_ASAP7_75t_L g565 ( .A(n_184), .Y(n_565) );
CKINVDCx8_ASAP7_75t_R g185 ( .A(n_186), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_188), .B(n_189), .Y(n_187) );
CKINVDCx16_ASAP7_75t_R g563 ( .A(n_190), .Y(n_563) );
AO21x1_ASAP7_75t_SL g573 ( .A1(n_190), .A2(n_574), .B(n_575), .Y(n_573) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g212 ( .A(n_191), .B(n_213), .Y(n_212) );
OR2x2_ASAP7_75t_SL g570 ( .A(n_191), .B(n_193), .Y(n_570) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_L g223 ( .A(n_192), .B(n_214), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_193), .B(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NOR2x1p5_ASAP7_75t_L g220 ( .A(n_194), .B(n_221), .Y(n_220) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
OR3x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_420), .C(n_491), .Y(n_197) );
NAND3x1_ASAP7_75t_SL g198 ( .A(n_199), .B(n_347), .C(n_369), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_337), .Y(n_199) );
AOI22xp33_ASAP7_75t_SL g200 ( .A1(n_201), .A2(n_267), .B1(n_315), .B2(n_319), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_201), .A2(n_523), .B1(n_524), .B2(n_526), .Y(n_522) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_239), .Y(n_201) );
AND2x2_ASAP7_75t_L g338 ( .A(n_202), .B(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_SL g404 ( .A(n_202), .B(n_385), .Y(n_404) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g322 ( .A(n_203), .Y(n_322) );
AND2x2_ASAP7_75t_L g372 ( .A(n_203), .B(n_241), .Y(n_372) );
INVx1_ASAP7_75t_L g411 ( .A(n_203), .Y(n_411) );
OR2x2_ASAP7_75t_L g448 ( .A(n_203), .B(n_259), .Y(n_448) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_203), .Y(n_460) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_203), .Y(n_484) );
AND2x2_ASAP7_75t_L g541 ( .A(n_203), .B(n_368), .Y(n_541) );
AO21x2_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_209), .B(n_235), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_205), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_SL g206 ( .A(n_207), .B(n_208), .Y(n_206) );
AND2x4_ASAP7_75t_L g243 ( .A(n_207), .B(n_208), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_210), .B(n_218), .Y(n_209) );
INVx1_ASAP7_75t_L g292 ( .A(n_211), .Y(n_292) );
AND2x4_ASAP7_75t_L g211 ( .A(n_212), .B(n_215), .Y(n_211) );
INVx1_ASAP7_75t_L g328 ( .A(n_212), .Y(n_328) );
OR2x6_ASAP7_75t_L g226 ( .A(n_213), .B(n_222), .Y(n_226) );
INVxp33_ASAP7_75t_L g302 ( .A(n_213), .Y(n_302) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_213), .Y(n_575) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AND2x4_ASAP7_75t_L g255 ( .A(n_214), .B(n_231), .Y(n_255) );
INVx1_ASAP7_75t_L g329 ( .A(n_215), .Y(n_329) );
BUFx3_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g222 ( .A(n_217), .Y(n_222) );
AND2x6_ASAP7_75t_L g252 ( .A(n_217), .B(n_229), .Y(n_252) );
INVxp67_ASAP7_75t_L g290 ( .A(n_219), .Y(n_290) );
AND2x4_ASAP7_75t_L g219 ( .A(n_220), .B(n_223), .Y(n_219) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_220), .Y(n_574) );
INVx1_ASAP7_75t_L g303 ( .A(n_221), .Y(n_303) );
INVx3_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_SL g224 ( .A1(n_225), .A2(n_226), .B(n_227), .C(n_233), .Y(n_224) );
OAI22xp5_ASAP7_75t_L g245 ( .A1(n_226), .A2(n_246), .B1(n_247), .B2(n_248), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_L g263 ( .A1(n_226), .A2(n_233), .B(n_264), .C(n_265), .Y(n_263) );
INVxp67_ASAP7_75t_L g280 ( .A(n_226), .Y(n_280) );
O2A1O1Ixp33_ASAP7_75t_L g311 ( .A1(n_226), .A2(n_233), .B(n_312), .C(n_313), .Y(n_311) );
INVx2_ASAP7_75t_L g335 ( .A(n_226), .Y(n_335) );
INVx1_ASAP7_75t_L g248 ( .A(n_228), .Y(n_248) );
AND2x4_ASAP7_75t_L g557 ( .A(n_228), .B(n_234), .Y(n_557) );
AND2x4_ASAP7_75t_L g228 ( .A(n_229), .B(n_231), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_233), .B(n_243), .Y(n_256) );
INVx1_ASAP7_75t_L g299 ( .A(n_233), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g332 ( .A1(n_233), .A2(n_333), .B(n_334), .Y(n_332) );
INVx5_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_234), .Y(n_283) );
OAI22xp5_ASAP7_75t_L g278 ( .A1(n_236), .A2(n_279), .B1(n_284), .B2(n_285), .Y(n_278) );
INVx3_ASAP7_75t_L g285 ( .A(n_236), .Y(n_285) );
INVx4_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_237), .B(n_288), .Y(n_287) );
INVx3_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
BUFx4f_ASAP7_75t_L g271 ( .A(n_238), .Y(n_271) );
NOR2x1_ASAP7_75t_L g239 ( .A(n_240), .B(n_257), .Y(n_239) );
INVx1_ASAP7_75t_L g416 ( .A(n_240), .Y(n_416) );
AND2x2_ASAP7_75t_L g442 ( .A(n_240), .B(n_259), .Y(n_442) );
NAND2x1_ASAP7_75t_L g458 ( .A(n_240), .B(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g339 ( .A(n_241), .B(n_325), .Y(n_339) );
INVx3_ASAP7_75t_L g368 ( .A(n_241), .Y(n_368) );
NOR2x1_ASAP7_75t_SL g487 ( .A(n_241), .B(n_259), .Y(n_487) );
AND2x4_ASAP7_75t_L g241 ( .A(n_242), .B(n_244), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_243), .A2(n_262), .B(n_266), .Y(n_261) );
OAI21xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_249), .B(n_256), .Y(n_244) );
OAI222xp33_ASAP7_75t_L g558 ( .A1(n_247), .A2(n_559), .B1(n_560), .B2(n_566), .C1(n_568), .C2(n_571), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_248), .B(n_282), .Y(n_281) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_251), .B1(n_253), .B2(n_254), .Y(n_249) );
INVxp67_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVxp67_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NOR2x1_ASAP7_75t_L g395 ( .A(n_257), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g366 ( .A(n_258), .B(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx4_ASAP7_75t_L g336 ( .A(n_259), .Y(n_336) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_259), .Y(n_381) );
AND2x2_ASAP7_75t_L g453 ( .A(n_259), .B(n_325), .Y(n_453) );
AND2x4_ASAP7_75t_L g470 ( .A(n_259), .B(n_414), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_259), .B(n_412), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_259), .B(n_321), .Y(n_546) );
OR2x6_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_267), .A2(n_363), .B1(n_434), .B2(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_293), .Y(n_267) );
INVx2_ASAP7_75t_L g436 ( .A(n_268), .Y(n_436) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_276), .Y(n_268) );
BUFx3_ASAP7_75t_L g426 ( .A(n_269), .Y(n_426) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_270), .B(n_295), .Y(n_318) );
INVx2_ASAP7_75t_L g342 ( .A(n_270), .Y(n_342) );
INVx1_ASAP7_75t_L g354 ( .A(n_270), .Y(n_354) );
AND2x4_ASAP7_75t_L g361 ( .A(n_270), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g378 ( .A(n_270), .B(n_277), .Y(n_378) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_270), .Y(n_392) );
INVxp67_ASAP7_75t_L g400 ( .A(n_270), .Y(n_400) );
OA21x2_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_272), .B(n_275), .Y(n_270) );
INVx2_ASAP7_75t_SL g296 ( .A(n_271), .Y(n_296) );
AND2x2_ASAP7_75t_L g429 ( .A(n_276), .B(n_345), .Y(n_429) );
AND2x2_ASAP7_75t_L g445 ( .A(n_276), .B(n_346), .Y(n_445) );
NOR2xp67_ASAP7_75t_L g532 ( .A(n_276), .B(n_345), .Y(n_532) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x4_ASAP7_75t_L g341 ( .A(n_277), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g352 ( .A(n_277), .Y(n_352) );
INVx1_ASAP7_75t_L g365 ( .A(n_277), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_277), .B(n_307), .Y(n_402) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_286), .Y(n_277) );
AO21x2_ASAP7_75t_L g307 ( .A1(n_285), .A2(n_308), .B(n_314), .Y(n_307) );
AO21x2_ASAP7_75t_L g345 ( .A1(n_285), .A2(n_308), .B(n_314), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_290), .B1(n_291), .B2(n_292), .Y(n_286) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g525 ( .A(n_293), .Y(n_525) );
AND2x4_ASAP7_75t_L g293 ( .A(n_294), .B(n_306), .Y(n_293) );
AND2x2_ASAP7_75t_L g399 ( .A(n_294), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g428 ( .A(n_294), .Y(n_428) );
AND2x2_ASAP7_75t_L g530 ( .A(n_294), .B(n_345), .Y(n_530) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_295), .B(n_307), .Y(n_390) );
AO21x2_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_297), .B(n_305), .Y(n_295) );
AO21x2_ASAP7_75t_L g346 ( .A1(n_296), .A2(n_297), .B(n_305), .Y(n_346) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_298), .B(n_304), .Y(n_297) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx3_ASAP7_75t_L g316 ( .A(n_306), .Y(n_316) );
NAND2x1p5_ASAP7_75t_L g505 ( .A(n_306), .B(n_426), .Y(n_505) );
INVx3_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_307), .Y(n_419) );
AND2x2_ASAP7_75t_L g446 ( .A(n_307), .B(n_392), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
AND2x2_ASAP7_75t_L g360 ( .A(n_316), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g376 ( .A(n_316), .Y(n_376) );
AND2x2_ASAP7_75t_L g464 ( .A(n_316), .B(n_341), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_316), .B(n_484), .Y(n_489) );
AND2x2_ASAP7_75t_L g499 ( .A(n_316), .B(n_378), .Y(n_499) );
OR2x2_ASAP7_75t_L g536 ( .A(n_316), .B(n_436), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_317), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g496 ( .A(n_317), .B(n_352), .Y(n_496) );
AND2x2_ASAP7_75t_L g512 ( .A(n_317), .B(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g506 ( .A(n_318), .B(n_402), .Y(n_506) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_323), .Y(n_319) );
INVx1_ASAP7_75t_L g388 ( .A(n_320), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_320), .B(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g486 ( .A(n_320), .B(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_320), .B(n_367), .Y(n_511) );
INVx3_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_321), .Y(n_358) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_322), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_323), .A2(n_356), .B1(n_374), .B2(n_377), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_323), .B(n_458), .Y(n_457) );
INVx2_ASAP7_75t_SL g490 ( .A(n_323), .Y(n_490) );
AND2x4_ASAP7_75t_SL g323 ( .A(n_324), .B(n_336), .Y(n_323) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x4_ASAP7_75t_L g367 ( .A(n_325), .B(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g387 ( .A(n_325), .Y(n_387) );
INVx1_ASAP7_75t_L g414 ( .A(n_325), .Y(n_414) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_331), .Y(n_325) );
NOR3xp33_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .C(n_330), .Y(n_327) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_336), .Y(n_356) );
AND2x4_ASAP7_75t_L g413 ( .A(n_336), .B(n_414), .Y(n_413) );
NOR2x1_ASAP7_75t_L g474 ( .A(n_336), .B(n_443), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_338), .B(n_340), .Y(n_337) );
AND2x2_ASAP7_75t_L g438 ( .A(n_338), .B(n_381), .Y(n_438) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_338), .A2(n_519), .B(n_520), .Y(n_518) );
INVx2_ASAP7_75t_L g396 ( .A(n_339), .Y(n_396) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_340), .A2(n_450), .B1(n_454), .B2(n_457), .Y(n_449) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_343), .Y(n_340) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_341), .Y(n_407) );
AND2x2_ASAP7_75t_L g417 ( .A(n_341), .B(n_418), .Y(n_417) );
INVx3_ASAP7_75t_L g456 ( .A(n_341), .Y(n_456) );
NAND2x1_ASAP7_75t_SL g481 ( .A(n_341), .B(n_350), .Y(n_481) );
AND2x2_ASAP7_75t_L g377 ( .A(n_343), .B(n_378), .Y(n_377) );
AND2x4_ASAP7_75t_L g343 ( .A(n_344), .B(n_346), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NOR2x1_ASAP7_75t_L g353 ( .A(n_345), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g350 ( .A(n_346), .Y(n_350) );
INVx2_ASAP7_75t_L g362 ( .A(n_346), .Y(n_362) );
AOI21xp5_ASAP7_75t_SL g347 ( .A1(n_348), .A2(n_355), .B(n_359), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_350), .B(n_544), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_351), .A2(n_440), .B1(n_444), .B2(n_447), .Y(n_439) );
AND2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
BUFx2_ASAP7_75t_L g544 ( .A(n_352), .Y(n_544) );
INVx1_ASAP7_75t_SL g551 ( .A(n_352), .Y(n_551) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_353), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OA21x2_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_363), .B(n_366), .Y(n_359) );
AND2x2_ASAP7_75t_L g363 ( .A(n_361), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g405 ( .A(n_361), .B(n_401), .Y(n_405) );
AND2x2_ASAP7_75t_L g520 ( .A(n_361), .B(n_418), .Y(n_520) );
AND2x2_ASAP7_75t_L g523 ( .A(n_361), .B(n_429), .Y(n_523) );
AND2x4_ASAP7_75t_L g531 ( .A(n_361), .B(n_532), .Y(n_531) );
OAI21xp33_ASAP7_75t_L g485 ( .A1(n_363), .A2(n_486), .B(n_488), .Y(n_485) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g513 ( .A(n_365), .Y(n_513) );
AND2x2_ASAP7_75t_L g529 ( .A(n_365), .B(n_530), .Y(n_529) );
INVx4_ASAP7_75t_L g443 ( .A(n_367), .Y(n_443) );
INVx1_ASAP7_75t_L g412 ( .A(n_368), .Y(n_412) );
AND2x2_ASAP7_75t_L g434 ( .A(n_368), .B(n_387), .Y(n_434) );
NOR2x1_ASAP7_75t_L g369 ( .A(n_370), .B(n_393), .Y(n_369) );
OAI21xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_373), .B(n_379), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g380 ( .A(n_372), .B(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_SL g533 ( .A(n_372), .B(n_385), .Y(n_533) );
AND2x2_ASAP7_75t_L g554 ( .A(n_372), .B(n_470), .Y(n_554) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g480 ( .A(n_377), .Y(n_480) );
OAI21xp5_ASAP7_75t_SL g379 ( .A1(n_380), .A2(n_382), .B(n_389), .Y(n_379) );
OR2x6_ASAP7_75t_L g432 ( .A(n_381), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_384), .B(n_388), .Y(n_383) );
INVx2_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
OR2x2_ASAP7_75t_L g455 ( .A(n_390), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g552 ( .A(n_390), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_391), .B(n_525), .Y(n_524) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_406), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_397), .B1(n_403), .B2(n_405), .Y(n_394) );
OR2x2_ASAP7_75t_L g466 ( .A(n_396), .B(n_467), .Y(n_466) );
INVx3_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_398), .Y(n_423) );
NAND2x1p5_ASAP7_75t_L g398 ( .A(n_399), .B(n_401), .Y(n_398) );
INVx1_ASAP7_75t_L g472 ( .A(n_401), .Y(n_472) );
INVx2_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
INVxp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_408), .B1(n_415), .B2(n_417), .Y(n_406) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_410), .B(n_413), .Y(n_409) );
AND2x4_ASAP7_75t_SL g410 ( .A(n_411), .B(n_412), .Y(n_410) );
AND2x2_ASAP7_75t_L g415 ( .A(n_413), .B(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g476 ( .A(n_416), .B(n_470), .Y(n_476) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_421), .B(n_461), .Y(n_420) );
NOR2xp67_ASAP7_75t_L g421 ( .A(n_422), .B(n_435), .Y(n_421) );
AOI21xp33_ASAP7_75t_SL g422 ( .A1(n_423), .A2(n_424), .B(n_430), .Y(n_422) );
OR2x2_ASAP7_75t_L g424 ( .A(n_425), .B(n_427), .Y(n_424) );
INVx3_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NAND2x1p5_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OAI22xp33_ASAP7_75t_SL g500 ( .A1(n_432), .A2(n_501), .B1(n_503), .B2(n_506), .Y(n_500) );
NOR2x1_ASAP7_75t_L g447 ( .A(n_433), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g483 ( .A(n_434), .B(n_484), .Y(n_483) );
OAI211xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_437), .B(n_439), .C(n_449), .Y(n_435) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
NAND2xp33_ASAP7_75t_SL g440 ( .A(n_441), .B(n_443), .Y(n_440) );
INVxp33_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g452 ( .A(n_443), .Y(n_452) );
AOI221xp5_ASAP7_75t_L g463 ( .A1(n_444), .A2(n_464), .B1(n_465), .B2(n_468), .C(n_471), .Y(n_463) );
AND2x4_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
INVx1_ASAP7_75t_L g504 ( .A(n_445), .Y(n_504) );
INVx2_ASAP7_75t_SL g502 ( .A(n_448), .Y(n_502) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
NAND2x1_ASAP7_75t_L g501 ( .A(n_452), .B(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g498 ( .A(n_458), .Y(n_498) );
INVx1_ASAP7_75t_L g527 ( .A(n_459), .Y(n_527) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NOR2x1_ASAP7_75t_L g461 ( .A(n_462), .B(n_477), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_463), .B(n_475), .Y(n_462) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g516 ( .A(n_467), .Y(n_516) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g537 ( .A(n_470), .B(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g542 ( .A(n_470), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_472), .B(n_473), .Y(n_471) );
INVxp33_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx2_ASAP7_75t_L g495 ( .A(n_474), .Y(n_495) );
OAI21xp5_ASAP7_75t_SL g477 ( .A1(n_478), .A2(n_482), .B(n_485), .Y(n_477) );
INVxp67_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
BUFx2_ASAP7_75t_L g538 ( .A(n_484), .Y(n_538) );
AND2x2_ASAP7_75t_L g526 ( .A(n_487), .B(n_527), .Y(n_526) );
NOR2xp33_ASAP7_75t_R g488 ( .A(n_489), .B(n_490), .Y(n_488) );
NAND3xp33_ASAP7_75t_L g491 ( .A(n_492), .B(n_507), .C(n_534), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_493), .B(n_500), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_494), .B(n_497), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
OR2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_508), .B(n_521), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_509), .B(n_518), .Y(n_508) );
AOI22xp33_ASAP7_75t_SL g509 ( .A1(n_510), .A2(n_512), .B1(n_514), .B2(n_515), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
NOR2x1_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
INVxp67_ASAP7_75t_SL g519 ( .A(n_517), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_522), .B(n_528), .Y(n_521) );
OAI21xp5_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_531), .B(n_533), .Y(n_528) );
INVx1_ASAP7_75t_L g547 ( .A(n_531), .Y(n_547) );
AOI211xp5_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_537), .B(n_539), .C(n_548), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_543), .B1(n_545), .B2(n_547), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_549), .B(n_553), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
INVxp67_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g560 ( .A(n_561), .Y(n_560) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_562), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
CKINVDCx20_ASAP7_75t_R g568 ( .A(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
CKINVDCx20_ASAP7_75t_R g571 ( .A(n_572), .Y(n_571) );
CKINVDCx20_ASAP7_75t_R g572 ( .A(n_573), .Y(n_572) );
endmodule