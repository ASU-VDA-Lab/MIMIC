module fake_jpeg_10545_n_311 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_311);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_36),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_39),
.Y(n_50)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx5_ASAP7_75t_SL g56 ( 
.A(n_43),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_18),
.B1(n_25),
.B2(n_19),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_49),
.B1(n_59),
.B2(n_26),
.Y(n_65)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_46),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_25),
.B1(n_38),
.B2(n_19),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_41),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_51),
.B(n_32),
.Y(n_83)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_41),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_54),
.Y(n_67)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_58),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_36),
.A2(n_24),
.B1(n_20),
.B2(n_21),
.Y(n_59)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_64),
.Y(n_85)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_65),
.Y(n_105)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_68),
.B(n_69),
.Y(n_104)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_42),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_56),
.Y(n_100)
);

AO22x1_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_52),
.B1(n_60),
.B2(n_56),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_87),
.Y(n_101)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_79),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_35),
.B1(n_40),
.B2(n_53),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_74),
.A2(n_80),
.B1(n_69),
.B2(n_73),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_76),
.A2(n_98),
.B1(n_32),
.B2(n_34),
.Y(n_114)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_77),
.A2(n_93),
.B1(n_94),
.B2(n_32),
.Y(n_115)
);

BUFx8_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_48),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_82),
.Y(n_111)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_84),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_23),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_63),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_46),
.B(n_22),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_89),
.B(n_92),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_36),
.C(n_42),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_43),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_29),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_95),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_51),
.B(n_16),
.Y(n_92)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_56),
.A2(n_22),
.B1(n_16),
.B2(n_33),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_96),
.B(n_97),
.Y(n_99)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_60),
.A2(n_40),
.B1(n_35),
.B2(n_33),
.Y(n_98)
);

NAND2xp33_ASAP7_75t_SL g134 ( 
.A(n_100),
.B(n_43),
.Y(n_134)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_102),
.B(n_107),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_103),
.A2(n_71),
.B(n_27),
.Y(n_155)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_60),
.B1(n_47),
.B2(n_27),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_110),
.A2(n_117),
.B1(n_122),
.B2(n_124),
.Y(n_146)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_112),
.B(n_114),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_87),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_72),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_74),
.A2(n_34),
.B1(n_30),
.B2(n_28),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_120),
.C(n_43),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_37),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_121),
.Y(n_145)
);

AND2x2_ASAP7_75t_SL g120 ( 
.A(n_70),
.B(n_43),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_70),
.B(n_37),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_88),
.A2(n_34),
.B1(n_30),
.B2(n_28),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_90),
.A2(n_43),
.B1(n_30),
.B2(n_28),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_76),
.Y(n_125)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_125),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_88),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_99),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_128),
.B(n_129),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_99),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_113),
.B(n_96),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_131),
.B(n_132),
.Y(n_185)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_135),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_134),
.B(n_153),
.Y(n_176)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_105),
.A2(n_95),
.B1(n_67),
.B2(n_66),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_138),
.A2(n_101),
.B(n_114),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_139),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_111),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_142),
.Y(n_181)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_123),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_121),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_143),
.A2(n_156),
.B1(n_109),
.B2(n_82),
.Y(n_173)
);

AND2x4_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_71),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_144),
.A2(n_154),
.B(n_2),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_105),
.A2(n_97),
.B1(n_66),
.B2(n_77),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_147),
.A2(n_157),
.B1(n_124),
.B2(n_127),
.Y(n_159)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_8),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_119),
.C(n_116),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_68),
.Y(n_151)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_151),
.Y(n_160)
);

A2O1A1O1Ixp25_ASAP7_75t_L g153 ( 
.A1(n_108),
.A2(n_118),
.B(n_120),
.C(n_100),
.D(n_103),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_123),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_155),
.A2(n_122),
.B(n_29),
.Y(n_177)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_110),
.Y(n_156)
);

OAI22x1_ASAP7_75t_SL g157 ( 
.A1(n_120),
.A2(n_37),
.B1(n_29),
.B2(n_75),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_162),
.C(n_164),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_112),
.C(n_102),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_107),
.C(n_101),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_166),
.A2(n_177),
.B(n_189),
.Y(n_208)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_167),
.B(n_170),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_125),
.B1(n_117),
.B2(n_106),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_169),
.A2(n_174),
.B1(n_175),
.B2(n_179),
.Y(n_206)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_146),
.A2(n_106),
.B1(n_115),
.B2(n_113),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_152),
.A2(n_126),
.B1(n_93),
.B2(n_86),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_145),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_178),
.B(n_183),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_152),
.A2(n_86),
.B1(n_37),
.B2(n_78),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_156),
.A2(n_78),
.B1(n_37),
.B2(n_29),
.Y(n_180)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_180),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_0),
.C(n_1),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_182),
.B(n_187),
.C(n_191),
.Y(n_218)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_148),
.Y(n_183)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_130),
.B(n_0),
.Y(n_186)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_0),
.C(n_2),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_138),
.A2(n_144),
.B1(n_130),
.B2(n_157),
.Y(n_188)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_144),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_144),
.A2(n_3),
.B(n_4),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_191),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_181),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_195),
.B(n_198),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_180),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_200),
.A2(n_144),
.B(n_177),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_140),
.Y(n_201)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_201),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_167),
.B(n_149),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_205),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_165),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_203),
.Y(n_239)
);

NOR3xp33_ASAP7_75t_SL g204 ( 
.A(n_185),
.B(n_154),
.C(n_142),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_213),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_129),
.Y(n_205)
);

INVxp33_ASAP7_75t_SL g209 ( 
.A(n_165),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_168),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_214),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_184),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_171),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_179),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_218),
.Y(n_237)
);

INVxp33_ASAP7_75t_L g217 ( 
.A(n_175),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_L g228 ( 
.A1(n_217),
.A2(n_215),
.B1(n_192),
.B2(n_196),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_194),
.A2(n_190),
.B1(n_174),
.B2(n_158),
.Y(n_219)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_176),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_223),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_221),
.A2(n_214),
.B(n_199),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_176),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_161),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_230),
.C(n_210),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_212),
.A2(n_188),
.B1(n_158),
.B2(n_169),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_225),
.A2(n_226),
.B1(n_235),
.B2(n_216),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_212),
.A2(n_135),
.B1(n_159),
.B2(n_163),
.Y(n_226)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_228),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_162),
.C(n_164),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_208),
.A2(n_207),
.B(n_216),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_231),
.A2(n_240),
.B(n_205),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_192),
.A2(n_163),
.B1(n_166),
.B2(n_132),
.Y(n_232)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_206),
.A2(n_187),
.B1(n_133),
.B2(n_160),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_189),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_218),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_201),
.A2(n_172),
.B(n_128),
.Y(n_240)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_242),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_239),
.B(n_202),
.Y(n_244)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_244),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_233),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_245),
.A2(n_246),
.B1(n_234),
.B2(n_226),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_233),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_247),
.A2(n_248),
.B(n_253),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_221),
.A2(n_195),
.B(n_199),
.Y(n_248)
);

AO221x1_ASAP7_75t_L g251 ( 
.A1(n_229),
.A2(n_203),
.B1(n_136),
.B2(n_139),
.C(n_213),
.Y(n_251)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_251),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_227),
.A2(n_203),
.B1(n_197),
.B2(n_210),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_252),
.A2(n_257),
.B1(n_258),
.B2(n_235),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_220),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_237),
.C(n_230),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_197),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_256),
.B(n_222),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_229),
.A2(n_204),
.B1(n_182),
.B2(n_139),
.Y(n_257)
);

NOR3xp33_ASAP7_75t_SL g258 ( 
.A(n_240),
.B(n_10),
.C(n_15),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_260),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_271),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_253),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_250),
.A2(n_225),
.B1(n_236),
.B2(n_237),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_263),
.A2(n_265),
.B1(n_242),
.B2(n_246),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_266),
.C(n_269),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_241),
.A2(n_231),
.B1(n_238),
.B2(n_228),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_223),
.C(n_224),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_136),
.C(n_4),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_9),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_9),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_14),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_275),
.A2(n_276),
.B1(n_282),
.B2(n_283),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_258),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_280),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_267),
.A2(n_243),
.B(n_245),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_278),
.A2(n_3),
.B(n_4),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_256),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_268),
.A2(n_257),
.B1(n_247),
.B2(n_254),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_262),
.A2(n_9),
.B1(n_13),
.B2(n_12),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_285),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_267),
.Y(n_285)
);

MAJx2_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_275),
.C(n_274),
.Y(n_288)
);

AOI21xp33_ASAP7_75t_L g297 ( 
.A1(n_288),
.A2(n_12),
.B(n_10),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_274),
.A2(n_270),
.B1(n_269),
.B2(n_271),
.Y(n_289)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_289),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_264),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_290),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_281),
.A2(n_266),
.B(n_272),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_291),
.A2(n_292),
.B(n_294),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_279),
.C(n_261),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_278),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_295),
.B(n_11),
.Y(n_300)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_297),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_295),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_298),
.Y(n_304)
);

AOI322xp5_ASAP7_75t_L g306 ( 
.A1(n_300),
.A2(n_301),
.A3(n_288),
.B1(n_293),
.B2(n_7),
.C1(n_5),
.C2(n_6),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_11),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_292),
.C(n_287),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_302),
.C(n_7),
.Y(n_308)
);

AOI32xp33_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_298),
.A3(n_7),
.B1(n_5),
.B2(n_296),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_307),
.A2(n_308),
.B(n_303),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_304),
.B(n_305),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_7),
.Y(n_311)
);


endmodule