module fake_jpeg_27413_n_237 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_237);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_237;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_12),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_14),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_12),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_29),
.A2(n_13),
.B1(n_19),
.B2(n_18),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_38),
.A2(n_40),
.B1(n_46),
.B2(n_26),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_29),
.A2(n_13),
.B1(n_19),
.B2(n_24),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_21),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_31),
.Y(n_52)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_24),
.B1(n_25),
.B2(n_22),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_52),
.B(n_56),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_50),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_58),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_39),
.B(n_35),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_47),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_34),
.B1(n_30),
.B2(n_36),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_59),
.A2(n_68),
.B1(n_69),
.B2(n_51),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_65),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_32),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_31),
.Y(n_84)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_48),
.A2(n_20),
.B1(n_33),
.B2(n_26),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_66),
.Y(n_91)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_70),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_28),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_50),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_21),
.Y(n_71)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_21),
.Y(n_72)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_46),
.A2(n_22),
.B1(n_17),
.B2(n_25),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_40),
.B1(n_48),
.B2(n_38),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_79),
.Y(n_119)
);

NAND2x1_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_51),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_81),
.A2(n_37),
.B1(n_23),
.B2(n_3),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_43),
.C(n_45),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_84),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_44),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_88),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_44),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_52),
.A2(n_0),
.B(n_1),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g104 ( 
.A1(n_89),
.A2(n_0),
.B(n_1),
.Y(n_104)
);

AND2x6_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_54),
.Y(n_92)
);

A2O1A1O1Ixp25_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_94),
.B(n_95),
.C(n_97),
.D(n_23),
.Y(n_109)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_67),
.Y(n_99)
);

AND2x6_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_10),
.Y(n_94)
);

A2O1A1O1Ixp25_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_23),
.B(n_26),
.C(n_22),
.D(n_17),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_43),
.C(n_22),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_62),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_56),
.A2(n_23),
.B(n_26),
.C(n_17),
.Y(n_97)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_100),
.B(n_110),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_102),
.B(n_76),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_78),
.A2(n_73),
.B1(n_53),
.B2(n_57),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_103),
.A2(n_111),
.B1(n_95),
.B2(n_86),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_104),
.A2(n_107),
.B(n_109),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_53),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_106),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_55),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_55),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_80),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_108),
.Y(n_123)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_92),
.A2(n_57),
.B1(n_49),
.B2(n_37),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_112),
.B(n_83),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_113),
.A2(n_61),
.B(n_85),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_43),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_116),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_115),
.A2(n_91),
.B1(n_79),
.B2(n_89),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_90),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_62),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_118),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_86),
.B(n_1),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_60),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_93),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_99),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_124),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_125),
.A2(n_129),
.B1(n_131),
.B2(n_138),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_128),
.Y(n_157)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_113),
.A2(n_92),
.B1(n_91),
.B2(n_81),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_82),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_98),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_101),
.A2(n_88),
.B1(n_96),
.B2(n_94),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_134),
.A2(n_109),
.B1(n_117),
.B2(n_118),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_103),
.A2(n_94),
.B1(n_95),
.B2(n_97),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_135),
.A2(n_144),
.B(n_119),
.Y(n_151)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_136),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_139),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_97),
.B1(n_85),
.B2(n_74),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_111),
.A2(n_85),
.B1(n_74),
.B2(n_76),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_140),
.A2(n_110),
.B1(n_100),
.B2(n_108),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_60),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_141),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_107),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_107),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_145),
.B(n_133),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_101),
.C(n_119),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_153),
.C(n_162),
.Y(n_174)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_148),
.B(n_154),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_151),
.A2(n_122),
.B(n_134),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_156),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_119),
.C(n_116),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_112),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_106),
.Y(n_158)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_158),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_159),
.A2(n_125),
.B1(n_135),
.B2(n_121),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_74),
.B1(n_102),
.B2(n_61),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_161),
.A2(n_138),
.B1(n_127),
.B2(n_128),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_61),
.C(n_12),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_144),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_164),
.Y(n_177)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_11),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_166),
.Y(n_181)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_167),
.A2(n_160),
.B1(n_157),
.B2(n_161),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_131),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_171),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_170),
.B(n_178),
.Y(n_188)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_133),
.C(n_122),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_175),
.B(n_176),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_159),
.A2(n_127),
.B1(n_126),
.B2(n_132),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_151),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_142),
.C(n_11),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_179),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_142),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_183),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_163),
.A2(n_150),
.B1(n_166),
.B2(n_148),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_150),
.Y(n_184)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

AOI21x1_ASAP7_75t_L g185 ( 
.A1(n_177),
.A2(n_164),
.B(n_156),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_185),
.A2(n_194),
.B(n_195),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_193),
.Y(n_207)
);

XOR2x1_ASAP7_75t_SL g187 ( 
.A(n_172),
.B(n_178),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_192),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_182),
.B(n_147),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_9),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_147),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_172),
.A2(n_157),
.B(n_149),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_198),
.B(n_203),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_194),
.A2(n_167),
.B1(n_179),
.B2(n_175),
.Y(n_199)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_187),
.A2(n_185),
.B1(n_191),
.B2(n_184),
.Y(n_200)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_200),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_174),
.C(n_169),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_202),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_188),
.A2(n_180),
.B1(n_174),
.B2(n_173),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_162),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_205),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_9),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_206),
.B(n_9),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_196),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_210),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_1),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_216),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_7),
.Y(n_216)
);

OAI21x1_ASAP7_75t_L g217 ( 
.A1(n_208),
.A2(n_204),
.B(n_199),
.Y(n_217)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_217),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_207),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_218),
.B(n_220),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_209),
.B(n_201),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_211),
.B(n_214),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_221),
.B(n_222),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_202),
.C(n_205),
.Y(n_222)
);

NOR2x1_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_215),
.Y(n_226)
);

AOI322xp5_ASAP7_75t_L g230 ( 
.A1(n_226),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_224),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_2),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_2),
.C(n_3),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_2),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_229),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_4),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_3),
.C(n_4),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_233),
.A2(n_226),
.B(n_5),
.Y(n_235)
);

AO21x1_ASAP7_75t_L g236 ( 
.A1(n_235),
.A2(n_234),
.B(n_5),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_236),
.B(n_6),
.Y(n_237)
);


endmodule