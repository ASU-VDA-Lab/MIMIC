module fake_jpeg_3484_n_194 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_194);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_194;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_16),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_14),
.B(n_30),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_6),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_37),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_39),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_9),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_7),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_5),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_69),
.Y(n_80)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

BUFx10_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_76),
.Y(n_87)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_79),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_82),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_79),
.A2(n_58),
.B1(n_68),
.B2(n_64),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_93),
.B1(n_64),
.B2(n_51),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_70),
.Y(n_82)
);

BUFx16f_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_84),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_52),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_89),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_71),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g110 ( 
.A1(n_88),
.A2(n_76),
.B1(n_67),
.B2(n_57),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_52),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_58),
.B1(n_49),
.B2(n_50),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_63),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_96),
.Y(n_119)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

INVxp67_ASAP7_75t_SL g130 ( 
.A(n_98),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_113),
.B1(n_2),
.B2(n_7),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_71),
.Y(n_102)
);

NAND2xp33_ASAP7_75t_SL g129 ( 
.A(n_102),
.B(n_110),
.Y(n_129)
);

AOI32xp33_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_59),
.A3(n_55),
.B1(n_54),
.B2(n_63),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_108),
.Y(n_115)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_93),
.A2(n_66),
.B1(n_65),
.B2(n_60),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_85),
.B1(n_4),
.B2(n_6),
.Y(n_121)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_92),
.B(n_54),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_107),
.B(n_112),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_55),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_91),
.C(n_84),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_111),
.Y(n_120)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_95),
.B(n_1),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_L g114 ( 
.A1(n_84),
.A2(n_23),
.B(n_47),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_114),
.A2(n_26),
.B(n_46),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_94),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_118),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_101),
.A2(n_85),
.B1(n_3),
.B2(n_4),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_117),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_24),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_124),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_122),
.A2(n_22),
.B1(n_27),
.B2(n_36),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_102),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_102),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_127),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_25),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_97),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_17),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_99),
.A2(n_8),
.B(n_10),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_133),
.A2(n_134),
.B(n_114),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_110),
.A2(n_10),
.B(n_11),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_100),
.B(n_11),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_135),
.B(n_32),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_119),
.B(n_113),
.Y(n_136)
);

NAND3xp33_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_141),
.C(n_142),
.Y(n_158)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_120),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_144),
.C(n_148),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_131),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_149),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_33),
.C(n_45),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_38),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_127),
.A2(n_12),
.B1(n_17),
.B2(n_18),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_146),
.A2(n_147),
.B1(n_140),
.B2(n_151),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_34),
.C(n_44),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_18),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_153),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_115),
.B(n_35),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_154),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_132),
.B(n_19),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_20),
.C(n_21),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_123),
.B(n_48),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_157),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_133),
.A2(n_134),
.B1(n_129),
.B2(n_117),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_156),
.A2(n_42),
.B1(n_143),
.B2(n_154),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_167),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_151),
.A2(n_125),
.B(n_123),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_164),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_156),
.A2(n_139),
.B(n_138),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_169),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_137),
.A2(n_131),
.B(n_121),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_170),
.Y(n_176)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_172),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_41),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_166),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_160),
.Y(n_178)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_178),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_169),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_165),
.C(n_168),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_161),
.C(n_164),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_174),
.A2(n_173),
.B1(n_158),
.B2(n_159),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_182),
.A2(n_185),
.B(n_186),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_184),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_163),
.Y(n_186)
);

AOI31xp67_ASAP7_75t_L g188 ( 
.A1(n_184),
.A2(n_176),
.A3(n_167),
.B(n_175),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_188),
.B(n_189),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_190),
.A2(n_191),
.B(n_179),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_187),
.A2(n_179),
.B1(n_183),
.B2(n_177),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_192),
.B(n_191),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_193),
.B(n_165),
.Y(n_194)
);


endmodule