module fake_ariane_204_n_1993 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1993);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1993;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_1083;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_194;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_928;
wire n_253;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_96),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_38),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_85),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_140),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_12),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_9),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_174),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_13),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_12),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_141),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_79),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_173),
.Y(n_205)
);

BUFx5_ASAP7_75t_L g206 ( 
.A(n_14),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_61),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_109),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_39),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_18),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_158),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_51),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_20),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_123),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_154),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_168),
.Y(n_216)
);

BUFx5_ASAP7_75t_L g217 ( 
.A(n_188),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_192),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_64),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_166),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_46),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_24),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_113),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_124),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_164),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_32),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_128),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_60),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_99),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_11),
.Y(n_230)
);

BUFx8_ASAP7_75t_SL g231 ( 
.A(n_161),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_52),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_0),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_121),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_167),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_176),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_61),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_75),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_190),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_31),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_149),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_171),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_146),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_73),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_0),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_179),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_170),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_126),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_93),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_78),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_105),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_32),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_150),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_90),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_77),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_45),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_29),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_106),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_143),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_10),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_104),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_50),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_18),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_191),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_64),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_182),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_95),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_122),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_38),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_91),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_41),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_92),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_186),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_25),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_86),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_84),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_69),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_10),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_181),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_6),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_127),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_131),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_159),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_83),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_17),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_33),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_58),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_89),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_119),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_62),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_71),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_28),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_101),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_162),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_114),
.Y(n_295)
);

BUFx10_ASAP7_75t_L g296 ( 
.A(n_28),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_137),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_31),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_52),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_8),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_9),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_80),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_55),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_142),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_117),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g306 ( 
.A(n_111),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_13),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_139),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_48),
.Y(n_309)
);

BUFx10_ASAP7_75t_L g310 ( 
.A(n_62),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_87),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_48),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_50),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_44),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_151),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_2),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_47),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_40),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_130),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_35),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_58),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_169),
.Y(n_322)
);

BUFx10_ASAP7_75t_L g323 ( 
.A(n_33),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_30),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_76),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_2),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_3),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_16),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_5),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_160),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_152),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_144),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_56),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_36),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_6),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_51),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_53),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_54),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_35),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_156),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_175),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_102),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_49),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_36),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_184),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_37),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_100),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_185),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_74),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_112),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_147),
.Y(n_351)
);

INVx2_ASAP7_75t_SL g352 ( 
.A(n_125),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_136),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_60),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_69),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_59),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_5),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_72),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_108),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_22),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_17),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_178),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_24),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_118),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_132),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_54),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_57),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_110),
.Y(n_368)
);

BUFx2_ASAP7_75t_SL g369 ( 
.A(n_115),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_30),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_53),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_103),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_94),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_15),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_145),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_148),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_172),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_21),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_81),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_47),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_44),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_21),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_41),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_82),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_260),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_231),
.Y(n_386)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_202),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_242),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_194),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_194),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_206),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_206),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_206),
.Y(n_393)
);

INVxp33_ASAP7_75t_SL g394 ( 
.A(n_207),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_206),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_298),
.Y(n_396)
);

INVxp67_ASAP7_75t_SL g397 ( 
.A(n_202),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_328),
.Y(n_398)
);

INVxp67_ASAP7_75t_SL g399 ( 
.A(n_355),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_206),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_203),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_206),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_206),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_234),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_206),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_235),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_355),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_355),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_355),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_355),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_213),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_213),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_242),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_272),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_230),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_230),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_279),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_228),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_302),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_204),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_204),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_296),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_218),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_218),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_304),
.Y(n_425)
);

INVxp67_ASAP7_75t_SL g426 ( 
.A(n_198),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_240),
.Y(n_427)
);

INVxp33_ASAP7_75t_SL g428 ( 
.A(n_207),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_256),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_248),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_201),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_209),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_296),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_219),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_222),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_226),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_248),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_257),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_250),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_250),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_199),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_353),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_353),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_252),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_210),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_262),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_265),
.Y(n_447)
);

CKINVDCx14_ASAP7_75t_R g448 ( 
.A(n_224),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_210),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_277),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g451 ( 
.A(n_296),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_278),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_280),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_263),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_269),
.Y(n_455)
);

INVxp67_ASAP7_75t_SL g456 ( 
.A(n_285),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_212),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_258),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_290),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_237),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_300),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_309),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_313),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_314),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_212),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_318),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_321),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_326),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_327),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_333),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_337),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_338),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_324),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_344),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_354),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_360),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_361),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_271),
.Y(n_478)
);

INVxp33_ASAP7_75t_SL g479 ( 
.A(n_232),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_374),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_445),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_458),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g483 ( 
.A(n_388),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_391),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_388),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_391),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_458),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_393),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_396),
.Y(n_489)
);

NOR2x1_ASAP7_75t_L g490 ( 
.A(n_420),
.B(n_340),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_393),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_395),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_404),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_395),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_399),
.B(n_364),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_400),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_458),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_448),
.B(n_200),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_458),
.Y(n_499)
);

INVx6_ASAP7_75t_L g500 ( 
.A(n_458),
.Y(n_500)
);

OA21x2_ASAP7_75t_L g501 ( 
.A1(n_400),
.A2(n_197),
.B(n_196),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_402),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_413),
.B(n_239),
.Y(n_503)
);

NAND2xp33_ASAP7_75t_SL g504 ( 
.A(n_398),
.B(n_228),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_392),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_402),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_387),
.B(n_288),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_403),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_403),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_392),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_413),
.B(n_340),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_405),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_405),
.Y(n_513)
);

OR2x2_ASAP7_75t_L g514 ( 
.A(n_385),
.B(n_221),
.Y(n_514)
);

BUFx8_ASAP7_75t_L g515 ( 
.A(n_386),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_407),
.Y(n_516)
);

OA21x2_ASAP7_75t_L g517 ( 
.A1(n_420),
.A2(n_215),
.B(n_211),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_421),
.B(n_229),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_421),
.B(n_238),
.Y(n_519)
);

AND2x6_ASAP7_75t_L g520 ( 
.A(n_423),
.B(n_258),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_407),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_417),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_449),
.Y(n_523)
);

NOR2x1_ASAP7_75t_L g524 ( 
.A(n_423),
.B(n_369),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_408),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_424),
.B(n_241),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_408),
.Y(n_527)
);

NOR2x1_ASAP7_75t_L g528 ( 
.A(n_424),
.B(n_214),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_397),
.B(n_310),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_419),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_409),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_409),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_394),
.B(n_291),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_410),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_R g535 ( 
.A(n_427),
.B(n_236),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_410),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_430),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_430),
.B(n_437),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_437),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_439),
.Y(n_540)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_429),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_428),
.A2(n_383),
.B1(n_382),
.B2(n_381),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_439),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_440),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_440),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_438),
.B(n_306),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_442),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_401),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_442),
.B(n_283),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_443),
.B(n_243),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_443),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_426),
.B(n_283),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_454),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_441),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_456),
.B(n_310),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_411),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_389),
.B(n_390),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_457),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_411),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_418),
.B(n_444),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_510),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_513),
.Y(n_562)
);

NOR3xp33_ASAP7_75t_L g563 ( 
.A(n_542),
.B(n_478),
.C(n_455),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_513),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_493),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_513),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_505),
.Y(n_567)
);

OR2x6_ASAP7_75t_L g568 ( 
.A(n_541),
.B(n_538),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_535),
.B(n_479),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_514),
.B(n_422),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_507),
.B(n_552),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_505),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_505),
.Y(n_573)
);

INVxp33_ASAP7_75t_L g574 ( 
.A(n_514),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_533),
.B(n_433),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_507),
.B(n_451),
.Y(n_576)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_557),
.B(n_465),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_505),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_512),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_512),
.Y(n_580)
);

INVxp67_ASAP7_75t_SL g581 ( 
.A(n_485),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_522),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_512),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_530),
.Y(n_584)
);

AND2x6_ASAP7_75t_L g585 ( 
.A(n_528),
.B(n_258),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_552),
.B(n_444),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_483),
.B(n_431),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_512),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_527),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_542),
.A2(n_245),
.B1(n_233),
.B2(n_232),
.Y(n_590)
);

INVxp67_ASAP7_75t_SL g591 ( 
.A(n_485),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_541),
.B(n_193),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_527),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_483),
.B(n_432),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_485),
.Y(n_595)
);

INVx1_ASAP7_75t_SL g596 ( 
.A(n_554),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_484),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_510),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_484),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_527),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_531),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_531),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_531),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_486),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_510),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_521),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_552),
.B(n_538),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_510),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_555),
.B(n_193),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_521),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_525),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_552),
.B(n_446),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_498),
.B(n_434),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_525),
.Y(n_614)
);

OR2x6_ASAP7_75t_L g615 ( 
.A(n_538),
.B(n_446),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_528),
.B(n_447),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_555),
.B(n_195),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_532),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_510),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_486),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_549),
.A2(n_378),
.B1(n_435),
.B2(n_436),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_538),
.B(n_447),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_532),
.Y(n_623)
);

INVx5_ASAP7_75t_L g624 ( 
.A(n_520),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_536),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_536),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_488),
.Y(n_627)
);

INVx1_ASAP7_75t_SL g628 ( 
.A(n_548),
.Y(n_628)
);

AND3x2_ASAP7_75t_L g629 ( 
.A(n_489),
.B(n_452),
.C(n_450),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_488),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_557),
.Y(n_631)
);

AO21x2_ASAP7_75t_L g632 ( 
.A1(n_491),
.A2(n_494),
.B(n_492),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_510),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_491),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_492),
.Y(n_635)
);

NAND2xp33_ASAP7_75t_SL g636 ( 
.A(n_553),
.B(n_233),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_494),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_496),
.Y(n_638)
);

INVxp67_ASAP7_75t_SL g639 ( 
.A(n_524),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_496),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_502),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_529),
.B(n_450),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_502),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_506),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_506),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_508),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_529),
.B(n_452),
.Y(n_647)
);

INVx2_ASAP7_75t_SL g648 ( 
.A(n_560),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_495),
.B(n_453),
.Y(n_649)
);

INVxp67_ASAP7_75t_SL g650 ( 
.A(n_524),
.Y(n_650)
);

NAND3xp33_ASAP7_75t_L g651 ( 
.A(n_508),
.B(n_254),
.C(n_251),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_495),
.B(n_453),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_509),
.B(n_459),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_516),
.Y(n_654)
);

AO21x2_ASAP7_75t_L g655 ( 
.A1(n_509),
.A2(n_268),
.B(n_255),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_516),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_501),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_539),
.Y(n_658)
);

OAI22xp33_ASAP7_75t_L g659 ( 
.A1(n_481),
.A2(n_558),
.B1(n_523),
.B2(n_336),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_560),
.B(n_195),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_516),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_546),
.A2(n_335),
.B1(n_370),
.B2(n_371),
.Y(n_662)
);

BUFx2_ASAP7_75t_L g663 ( 
.A(n_515),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_516),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_516),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_516),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_504),
.B(n_205),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_534),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_511),
.B(n_459),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_534),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_534),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_549),
.B(n_205),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_539),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_534),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_503),
.B(n_461),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_534),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_539),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_549),
.B(n_208),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_544),
.Y(n_679)
);

INVx2_ASAP7_75t_SL g680 ( 
.A(n_511),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_544),
.Y(n_681)
);

INVx5_ASAP7_75t_L g682 ( 
.A(n_520),
.Y(n_682)
);

NAND2xp33_ASAP7_75t_L g683 ( 
.A(n_537),
.B(n_208),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_534),
.Y(n_684)
);

INVx1_ASAP7_75t_SL g685 ( 
.A(n_503),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_544),
.Y(n_686)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_511),
.B(n_480),
.Y(n_687)
);

NAND2xp33_ASAP7_75t_SL g688 ( 
.A(n_549),
.B(n_335),
.Y(n_688)
);

AND2x4_ASAP7_75t_L g689 ( 
.A(n_511),
.B(n_461),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_518),
.B(n_216),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_490),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_518),
.Y(n_692)
);

CKINVDCx20_ASAP7_75t_R g693 ( 
.A(n_515),
.Y(n_693)
);

NAND2xp33_ASAP7_75t_SL g694 ( 
.A(n_519),
.B(n_336),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_559),
.Y(n_695)
);

NAND3xp33_ASAP7_75t_L g696 ( 
.A(n_501),
.B(n_276),
.C(n_270),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_559),
.Y(n_697)
);

OAI21xp33_ASAP7_75t_SL g698 ( 
.A1(n_537),
.A2(n_463),
.B(n_462),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_519),
.B(n_216),
.Y(n_699)
);

NAND3xp33_ASAP7_75t_L g700 ( 
.A(n_501),
.B(n_308),
.C(n_297),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_500),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_526),
.B(n_220),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_540),
.B(n_462),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_540),
.B(n_543),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_543),
.B(n_463),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_545),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_559),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_490),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_545),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_517),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_487),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_487),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_501),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_692),
.B(n_547),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_685),
.B(n_547),
.Y(n_715)
);

NOR2xp67_ASAP7_75t_L g716 ( 
.A(n_565),
.B(n_551),
.Y(n_716)
);

INVxp67_ASAP7_75t_L g717 ( 
.A(n_570),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_692),
.B(n_551),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_685),
.B(n_526),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_606),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_649),
.B(n_556),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_SL g722 ( 
.A(n_565),
.B(n_582),
.Y(n_722)
);

AO221x1_ASAP7_75t_L g723 ( 
.A1(n_659),
.A2(n_663),
.B1(n_590),
.B2(n_563),
.C(n_605),
.Y(n_723)
);

NAND3xp33_ASAP7_75t_L g724 ( 
.A(n_613),
.B(n_515),
.C(n_343),
.Y(n_724)
);

O2A1O1Ixp33_ASAP7_75t_L g725 ( 
.A1(n_698),
.A2(n_556),
.B(n_550),
.C(n_469),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_652),
.B(n_550),
.Y(n_726)
);

NAND2xp33_ASAP7_75t_L g727 ( 
.A(n_630),
.B(n_220),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_571),
.B(n_225),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_597),
.B(n_225),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_675),
.B(n_517),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_607),
.B(n_517),
.Y(n_731)
);

OAI22xp33_ASAP7_75t_SL g732 ( 
.A1(n_590),
.A2(n_357),
.B1(n_339),
.B2(n_363),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_570),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_576),
.B(n_274),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_597),
.B(n_227),
.Y(n_735)
);

INVxp67_ASAP7_75t_L g736 ( 
.A(n_596),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_609),
.B(n_286),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_574),
.B(n_406),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_617),
.B(n_287),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_607),
.B(n_586),
.Y(n_740)
);

NOR2xp67_ASAP7_75t_SL g741 ( 
.A(n_569),
.B(n_339),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_562),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_562),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_564),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_597),
.B(n_227),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_586),
.B(n_517),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_610),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_612),
.B(n_587),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_612),
.B(n_594),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_642),
.B(n_223),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_631),
.B(n_414),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_647),
.B(n_315),
.Y(n_752)
);

OR2x2_ASAP7_75t_L g753 ( 
.A(n_596),
.B(n_425),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_564),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_655),
.A2(n_306),
.B1(n_310),
.B2(n_323),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_611),
.Y(n_756)
);

O2A1O1Ixp5_ASAP7_75t_L g757 ( 
.A1(n_690),
.A2(n_362),
.B(n_311),
.C(n_372),
.Y(n_757)
);

BUFx3_ASAP7_75t_L g758 ( 
.A(n_663),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_691),
.B(n_292),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_611),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_631),
.B(n_515),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_604),
.Y(n_762)
);

INVxp67_ASAP7_75t_SL g763 ( 
.A(n_599),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_577),
.B(n_460),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_639),
.B(n_650),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_622),
.B(n_376),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_604),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_620),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_622),
.B(n_342),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_616),
.B(n_342),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_691),
.B(n_348),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_614),
.Y(n_772)
);

NAND2xp33_ASAP7_75t_L g773 ( 
.A(n_630),
.B(n_348),
.Y(n_773)
);

O2A1O1Ixp33_ASAP7_75t_L g774 ( 
.A1(n_698),
.A2(n_469),
.B(n_464),
.C(n_480),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_708),
.B(n_648),
.Y(n_775)
);

OAI22xp33_ASAP7_75t_L g776 ( 
.A1(n_568),
.A2(n_343),
.B1(n_346),
.B2(n_356),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_599),
.B(n_349),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_620),
.Y(n_778)
);

INVx2_ASAP7_75t_SL g779 ( 
.A(n_577),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_708),
.B(n_299),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_634),
.A2(n_640),
.B(n_638),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_614),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_648),
.B(n_301),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_618),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_615),
.B(n_349),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_618),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_623),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_599),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_615),
.B(n_351),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_634),
.B(n_351),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_615),
.B(n_358),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_615),
.B(n_358),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_623),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_615),
.B(n_359),
.Y(n_794)
);

O2A1O1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_638),
.A2(n_472),
.B(n_477),
.C(n_464),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_655),
.A2(n_306),
.B1(n_323),
.B2(n_352),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_568),
.B(n_466),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_628),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_689),
.B(n_359),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_625),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_627),
.Y(n_801)
);

O2A1O1Ixp5_ASAP7_75t_L g802 ( 
.A1(n_699),
.A2(n_350),
.B(n_325),
.C(n_345),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_625),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_689),
.B(n_680),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_689),
.B(n_365),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_640),
.B(n_365),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_627),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_689),
.B(n_368),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_680),
.B(n_706),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_641),
.B(n_368),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_706),
.B(n_373),
.Y(n_811)
);

AND2x4_ASAP7_75t_L g812 ( 
.A(n_568),
.B(n_687),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_635),
.Y(n_813)
);

NAND2xp33_ASAP7_75t_L g814 ( 
.A(n_641),
.B(n_373),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_709),
.B(n_375),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_626),
.Y(n_816)
);

BUFx12f_ASAP7_75t_SL g817 ( 
.A(n_568),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_643),
.B(n_375),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_568),
.A2(n_356),
.B1(n_357),
.B2(n_363),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_635),
.Y(n_820)
);

OR2x6_ASAP7_75t_L g821 ( 
.A(n_687),
.B(n_466),
.Y(n_821)
);

NOR2xp67_ASAP7_75t_L g822 ( 
.A(n_582),
.B(n_467),
.Y(n_822)
);

NAND2xp33_ASAP7_75t_L g823 ( 
.A(n_643),
.B(n_377),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_660),
.B(n_592),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_709),
.B(n_377),
.Y(n_825)
);

INVx2_ASAP7_75t_SL g826 ( 
.A(n_629),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_595),
.B(n_379),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_595),
.B(n_653),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_626),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_702),
.B(n_303),
.Y(n_830)
);

INVxp67_ASAP7_75t_L g831 ( 
.A(n_628),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_644),
.B(n_379),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_644),
.B(n_467),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_584),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_575),
.B(n_307),
.Y(n_835)
);

AOI22xp5_ASAP7_75t_L g836 ( 
.A1(n_688),
.A2(n_352),
.B1(n_341),
.B2(n_322),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_672),
.B(n_312),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_646),
.B(n_217),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_646),
.B(n_217),
.Y(n_839)
);

OR2x2_ASAP7_75t_L g840 ( 
.A(n_584),
.B(n_473),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_581),
.B(n_468),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_567),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_662),
.B(n_474),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_637),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_591),
.B(n_468),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_669),
.B(n_470),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_637),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_704),
.B(n_470),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_567),
.Y(n_849)
);

OR2x2_ASAP7_75t_L g850 ( 
.A(n_636),
.B(n_471),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_572),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_572),
.Y(n_852)
);

INVx2_ASAP7_75t_SL g853 ( 
.A(n_703),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_678),
.B(n_316),
.Y(n_854)
);

AND2x4_ASAP7_75t_L g855 ( 
.A(n_667),
.B(n_471),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_693),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_573),
.B(n_472),
.Y(n_857)
);

OAI22xp5_ASAP7_75t_L g858 ( 
.A1(n_662),
.A2(n_380),
.B1(n_383),
.B2(n_382),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_683),
.B(n_573),
.Y(n_859)
);

NOR2x1p5_ASAP7_75t_L g860 ( 
.A(n_705),
.B(n_346),
.Y(n_860)
);

INVx5_ASAP7_75t_L g861 ( 
.A(n_598),
.Y(n_861)
);

OR2x2_ASAP7_75t_L g862 ( 
.A(n_621),
.B(n_475),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_598),
.B(n_217),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_645),
.Y(n_864)
);

NAND2xp33_ASAP7_75t_L g865 ( 
.A(n_645),
.B(n_317),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_SL g866 ( 
.A(n_651),
.B(n_323),
.Y(n_866)
);

BUFx3_ASAP7_75t_L g867 ( 
.A(n_605),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_579),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_566),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_579),
.B(n_475),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_694),
.A2(n_319),
.B1(n_244),
.B2(n_246),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_658),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_585),
.B(n_476),
.Y(n_873)
);

INVxp33_ASAP7_75t_L g874 ( 
.A(n_651),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_598),
.B(n_217),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_658),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_585),
.B(n_476),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_561),
.B(n_320),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_686),
.Y(n_879)
);

OR2x2_ASAP7_75t_L g880 ( 
.A(n_578),
.B(n_477),
.Y(n_880)
);

AND2x2_ASAP7_75t_SL g881 ( 
.A(n_561),
.B(n_673),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_561),
.B(n_329),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_673),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_723),
.A2(n_655),
.B1(n_585),
.B2(n_713),
.Y(n_884)
);

INVxp67_ASAP7_75t_L g885 ( 
.A(n_798),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_719),
.B(n_726),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_742),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_720),
.Y(n_888)
);

NAND2x1p5_ASAP7_75t_L g889 ( 
.A(n_881),
.B(n_657),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_719),
.B(n_715),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_881),
.B(n_812),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_742),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_861),
.Y(n_893)
);

AOI22xp5_ASAP7_75t_L g894 ( 
.A1(n_812),
.A2(n_585),
.B1(n_632),
.B2(n_681),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_874),
.B(n_561),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_743),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_715),
.B(n_585),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_748),
.A2(n_657),
.B1(n_713),
.B2(n_583),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_779),
.B(n_412),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_812),
.B(n_598),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_749),
.B(n_585),
.Y(n_901)
);

INVx4_ASAP7_75t_L g902 ( 
.A(n_834),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_747),
.Y(n_903)
);

NAND2xp33_ASAP7_75t_L g904 ( 
.A(n_788),
.B(n_598),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_781),
.A2(n_632),
.B(n_605),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_740),
.B(n_578),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_743),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_744),
.Y(n_908)
);

OR2x6_ASAP7_75t_L g909 ( 
.A(n_831),
.B(n_657),
.Y(n_909)
);

INVx2_ASAP7_75t_SL g910 ( 
.A(n_840),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_817),
.B(n_580),
.Y(n_911)
);

INVx2_ASAP7_75t_SL g912 ( 
.A(n_753),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_758),
.Y(n_913)
);

OR2x6_ASAP7_75t_L g914 ( 
.A(n_736),
.B(n_713),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_821),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_756),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_760),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_772),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_782),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_751),
.Y(n_920)
);

INVxp67_ASAP7_75t_L g921 ( 
.A(n_738),
.Y(n_921)
);

INVx4_ASAP7_75t_L g922 ( 
.A(n_861),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_717),
.B(n_412),
.Y(n_923)
);

AND2x6_ASAP7_75t_SL g924 ( 
.A(n_843),
.B(n_415),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_867),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_714),
.B(n_585),
.Y(n_926)
);

AOI22xp33_ASAP7_75t_SL g927 ( 
.A1(n_866),
.A2(n_367),
.B1(n_370),
.B2(n_371),
.Y(n_927)
);

BUFx12f_ASAP7_75t_L g928 ( 
.A(n_856),
.Y(n_928)
);

AND2x6_ASAP7_75t_L g929 ( 
.A(n_797),
.B(n_677),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_718),
.B(n_677),
.Y(n_930)
);

AO22x1_ASAP7_75t_L g931 ( 
.A1(n_733),
.A2(n_366),
.B1(n_381),
.B2(n_367),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_853),
.B(n_679),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_784),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_721),
.B(n_679),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_797),
.B(n_681),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_788),
.B(n_608),
.Y(n_936)
);

INVx2_ASAP7_75t_SL g937 ( 
.A(n_758),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_786),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_787),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_821),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_867),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_828),
.A2(n_632),
.B(n_583),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_793),
.Y(n_943)
);

NOR3xp33_ASAP7_75t_SL g944 ( 
.A(n_858),
.B(n_380),
.C(n_366),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_734),
.B(n_580),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_744),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_861),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_754),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_754),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_879),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_797),
.B(n_588),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_763),
.A2(n_588),
.B1(n_710),
.B2(n_654),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_800),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_879),
.Y(n_954)
);

OR2x6_ASAP7_75t_L g955 ( 
.A(n_821),
.B(n_710),
.Y(n_955)
);

INVx4_ASAP7_75t_L g956 ( 
.A(n_861),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_SL g957 ( 
.A1(n_859),
.A2(n_676),
.B(n_674),
.C(n_654),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_803),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_750),
.B(n_686),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_716),
.B(n_695),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_816),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_829),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_880),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_752),
.B(n_695),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_764),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_850),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_847),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_826),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_869),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_761),
.B(n_697),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_809),
.A2(n_654),
.B(n_674),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_847),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_766),
.B(n_697),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_734),
.B(n_707),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_859),
.B(n_608),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_869),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_848),
.B(n_707),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_762),
.Y(n_978)
);

OR2x6_ASAP7_75t_L g979 ( 
.A(n_822),
.B(n_804),
.Y(n_979)
);

AOI22xp33_ASAP7_75t_L g980 ( 
.A1(n_746),
.A2(n_696),
.B1(n_700),
.B2(n_603),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_855),
.Y(n_981)
);

BUFx2_ASAP7_75t_L g982 ( 
.A(n_785),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_762),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_759),
.B(n_589),
.Y(n_984)
);

NOR3xp33_ASAP7_75t_SL g985 ( 
.A(n_776),
.B(n_334),
.C(n_284),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_855),
.B(n_674),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_775),
.B(n_676),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_842),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_759),
.B(n_589),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_849),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_767),
.B(n_608),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_767),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_780),
.B(n_593),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_780),
.B(n_593),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_860),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_768),
.Y(n_996)
);

AND2x6_ASAP7_75t_L g997 ( 
.A(n_731),
.B(n_608),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_768),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_778),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_722),
.B(n_415),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_851),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_783),
.B(n_416),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_852),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_778),
.B(n_608),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_841),
.B(n_600),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_868),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_845),
.B(n_600),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_855),
.B(n_601),
.Y(n_1008)
);

AOI22xp33_ASAP7_75t_L g1009 ( 
.A1(n_862),
.A2(n_700),
.B1(n_696),
.B2(n_601),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_801),
.B(n_619),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_801),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_835),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_783),
.B(n_416),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_872),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_769),
.B(n_602),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_807),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_876),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_883),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_807),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_765),
.B(n_602),
.Y(n_1020)
);

NOR3xp33_ASAP7_75t_SL g1021 ( 
.A(n_819),
.B(n_724),
.C(n_790),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_846),
.B(n_603),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_SL g1023 ( 
.A(n_741),
.Y(n_1023)
);

NAND2x1p5_ASAP7_75t_L g1024 ( 
.A(n_813),
.B(n_820),
.Y(n_1024)
);

BUFx8_ASAP7_75t_L g1025 ( 
.A(n_813),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_824),
.B(n_676),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_820),
.Y(n_1027)
);

AND2x4_ASAP7_75t_L g1028 ( 
.A(n_824),
.B(n_701),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_833),
.B(n_619),
.Y(n_1029)
);

INVx2_ASAP7_75t_SL g1030 ( 
.A(n_799),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_770),
.B(n_619),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_844),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_844),
.B(n_864),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_864),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_857),
.Y(n_1035)
);

OR2x2_ASAP7_75t_L g1036 ( 
.A(n_835),
.B(n_701),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_873),
.Y(n_1037)
);

NAND2x2_ASAP7_75t_L g1038 ( 
.A(n_732),
.B(n_1),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_730),
.B(n_619),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_870),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_878),
.B(n_619),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_729),
.B(n_701),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_877),
.Y(n_1043)
);

BUFx8_ASAP7_75t_L g1044 ( 
.A(n_774),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_838),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_811),
.B(n_633),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_725),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_795),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_815),
.Y(n_1049)
);

AOI22xp33_ASAP7_75t_L g1050 ( 
.A1(n_796),
.A2(n_712),
.B1(n_711),
.B2(n_664),
.Y(n_1050)
);

NOR2x1_ASAP7_75t_L g1051 ( 
.A(n_789),
.B(n_656),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_838),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_878),
.B(n_633),
.Y(n_1053)
);

BUFx12f_ASAP7_75t_L g1054 ( 
.A(n_755),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_728),
.B(n_790),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_825),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_737),
.B(n_656),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_882),
.B(n_633),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_839),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_882),
.B(n_633),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_832),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_839),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_805),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_808),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_827),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_728),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_791),
.B(n_633),
.Y(n_1067)
);

AOI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_727),
.A2(n_661),
.B1(n_664),
.B2(n_666),
.Y(n_1068)
);

HB1xp67_ASAP7_75t_L g1069 ( 
.A(n_792),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_794),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_771),
.B(n_661),
.Y(n_1071)
);

BUFx2_ASAP7_75t_L g1072 ( 
.A(n_836),
.Y(n_1072)
);

NAND2xp33_ASAP7_75t_R g1073 ( 
.A(n_1012),
.B(n_968),
.Y(n_1073)
);

INVx3_ASAP7_75t_L g1074 ( 
.A(n_955),
.Y(n_1074)
);

NOR2x1_ASAP7_75t_L g1075 ( 
.A(n_902),
.B(n_729),
.Y(n_1075)
);

BUFx4f_ASAP7_75t_L g1076 ( 
.A(n_928),
.Y(n_1076)
);

BUFx8_ASAP7_75t_L g1077 ( 
.A(n_928),
.Y(n_1077)
);

O2A1O1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_890),
.A2(n_830),
.B(n_806),
.C(n_810),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_886),
.A2(n_830),
.B(n_818),
.C(n_810),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_886),
.A2(n_818),
.B1(n_854),
.B2(n_837),
.Y(n_1080)
);

AOI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_965),
.A2(n_739),
.B1(n_737),
.B2(n_837),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_888),
.Y(n_1082)
);

BUFx4f_ASAP7_75t_L g1083 ( 
.A(n_909),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_1055),
.A2(n_739),
.B(n_854),
.C(n_823),
.Y(n_1084)
);

INVx4_ASAP7_75t_L g1085 ( 
.A(n_955),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_905),
.A2(n_875),
.B(n_863),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_1049),
.A2(n_814),
.B(n_773),
.C(n_745),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1002),
.B(n_735),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_934),
.A2(n_865),
.B(n_745),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_904),
.A2(n_735),
.B(n_777),
.Y(n_1090)
);

OAI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_942),
.A2(n_875),
.B(n_863),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_893),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_1055),
.A2(n_777),
.B1(n_871),
.B2(n_668),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_1041),
.A2(n_666),
.B(n_668),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_1054),
.A2(n_670),
.B1(n_671),
.B2(n_712),
.Y(n_1095)
);

O2A1O1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_1056),
.A2(n_802),
.B(n_757),
.C(n_670),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_893),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_920),
.B(n_671),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1013),
.B(n_665),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_1072),
.B(n_665),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_893),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1041),
.A2(n_684),
.B(n_665),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_945),
.A2(n_711),
.B(n_684),
.C(n_665),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_966),
.B(n_665),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_885),
.B(n_684),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_963),
.B(n_684),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_903),
.Y(n_1107)
);

NOR2xp67_ASAP7_75t_L g1108 ( 
.A(n_902),
.B(n_684),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_915),
.B(n_247),
.Y(n_1109)
);

AND2x2_ASAP7_75t_SL g1110 ( 
.A(n_915),
.B(n_258),
.Y(n_1110)
);

NOR3xp33_ASAP7_75t_SL g1111 ( 
.A(n_995),
.B(n_253),
.C(n_249),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1035),
.B(n_520),
.Y(n_1112)
);

CKINVDCx11_ASAP7_75t_R g1113 ( 
.A(n_1038),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1053),
.A2(n_294),
.B(n_259),
.Y(n_1114)
);

AND2x4_ASAP7_75t_SL g1115 ( 
.A(n_940),
.B(n_258),
.Y(n_1115)
);

INVxp67_ASAP7_75t_L g1116 ( 
.A(n_1000),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_945),
.A2(n_487),
.B(n_497),
.C(n_499),
.Y(n_1117)
);

O2A1O1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_1061),
.A2(n_497),
.B(n_499),
.C(n_4),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_940),
.B(n_1),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_913),
.Y(n_1120)
);

AOI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_891),
.A2(n_332),
.B1(n_282),
.B2(n_289),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1053),
.A2(n_261),
.B(n_264),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_916),
.Y(n_1123)
);

NAND2xp33_ASAP7_75t_SL g1124 ( 
.A(n_1021),
.B(n_266),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_895),
.A2(n_497),
.B(n_499),
.C(n_273),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1058),
.A2(n_330),
.B(n_275),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1058),
.A2(n_331),
.B(n_281),
.Y(n_1127)
);

O2A1O1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_1065),
.A2(n_3),
.B(n_4),
.C(n_7),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_937),
.B(n_267),
.Y(n_1129)
);

O2A1O1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_1064),
.A2(n_7),
.B(n_8),
.C(n_11),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1060),
.A2(n_293),
.B(n_295),
.Y(n_1131)
);

O2A1O1Ixp5_ASAP7_75t_SL g1132 ( 
.A1(n_1067),
.A2(n_520),
.B(n_500),
.C(n_217),
.Y(n_1132)
);

NOR3xp33_ASAP7_75t_SL g1133 ( 
.A(n_1066),
.B(n_384),
.C(n_15),
.Y(n_1133)
);

INVx6_ASAP7_75t_L g1134 ( 
.A(n_1025),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_910),
.B(n_14),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1040),
.B(n_520),
.Y(n_1136)
);

NOR2xp67_ASAP7_75t_L g1137 ( 
.A(n_912),
.B(n_682),
.Y(n_1137)
);

O2A1O1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_1063),
.A2(n_16),
.B(n_19),
.C(n_20),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_921),
.B(n_982),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_981),
.B(n_1063),
.Y(n_1140)
);

BUFx4f_ASAP7_75t_L g1141 ( 
.A(n_909),
.Y(n_1141)
);

O2A1O1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_1030),
.A2(n_19),
.B(n_22),
.C(n_23),
.Y(n_1142)
);

OAI22x1_ASAP7_75t_L g1143 ( 
.A1(n_1070),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_1143)
);

AND2x4_ASAP7_75t_L g1144 ( 
.A(n_913),
.B(n_981),
.Y(n_1144)
);

AOI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1060),
.A2(n_500),
.B(n_482),
.Y(n_1145)
);

OR2x6_ASAP7_75t_L g1146 ( 
.A(n_955),
.B(n_347),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_895),
.A2(n_347),
.B(n_305),
.C(n_682),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1039),
.A2(n_1029),
.B(n_974),
.Y(n_1148)
);

CKINVDCx16_ASAP7_75t_R g1149 ( 
.A(n_1023),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_906),
.A2(n_347),
.B(n_305),
.C(n_682),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1039),
.A2(n_682),
.B(n_624),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1069),
.B(n_923),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1046),
.A2(n_682),
.B(n_624),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_906),
.B(n_520),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_R g1155 ( 
.A(n_924),
.B(n_893),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_1069),
.B(n_26),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_897),
.A2(n_347),
.B(n_305),
.C(n_624),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_969),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_891),
.B(n_624),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_917),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1031),
.A2(n_624),
.B(n_347),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_918),
.Y(n_1162)
);

HB1xp67_ASAP7_75t_L g1163 ( 
.A(n_909),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_957),
.A2(n_624),
.B(n_305),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_1023),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_944),
.Y(n_1166)
);

A2O1A1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_1047),
.A2(n_901),
.B(n_984),
.C(n_989),
.Y(n_1167)
);

AOI21x1_ASAP7_75t_L g1168 ( 
.A1(n_975),
.A2(n_1067),
.B(n_1004),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1054),
.B(n_27),
.Y(n_1169)
);

OAI21xp33_ASAP7_75t_L g1170 ( 
.A1(n_927),
.A2(n_985),
.B(n_1048),
.Y(n_1170)
);

O2A1O1Ixp5_ASAP7_75t_L g1171 ( 
.A1(n_957),
.A2(n_27),
.B(n_29),
.C(n_34),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_977),
.A2(n_305),
.B(n_482),
.Y(n_1172)
);

O2A1O1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_1026),
.A2(n_34),
.B(n_37),
.C(n_39),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_919),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1028),
.B(n_40),
.Y(n_1175)
);

BUFx2_ASAP7_75t_L g1176 ( 
.A(n_914),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1028),
.B(n_42),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_993),
.A2(n_482),
.B(n_153),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_914),
.Y(n_1179)
);

INVx3_ASAP7_75t_L g1180 ( 
.A(n_922),
.Y(n_1180)
);

BUFx3_ASAP7_75t_L g1181 ( 
.A(n_899),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_930),
.B(n_520),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_933),
.Y(n_1183)
);

OAI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_898),
.A2(n_520),
.B(n_217),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_938),
.B(n_42),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_986),
.B(n_43),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_939),
.B(n_43),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_914),
.Y(n_1188)
);

BUFx2_ASAP7_75t_L g1189 ( 
.A(n_1044),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_994),
.A2(n_482),
.B(n_217),
.C(n_49),
.Y(n_1190)
);

INVx8_ASAP7_75t_L g1191 ( 
.A(n_929),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_960),
.B(n_482),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_943),
.B(n_45),
.Y(n_1193)
);

AND2x6_ASAP7_75t_L g1194 ( 
.A(n_947),
.B(n_482),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_931),
.Y(n_1195)
);

A2O1A1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_987),
.A2(n_217),
.B(n_55),
.C(n_56),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_969),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_953),
.B(n_46),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_975),
.A2(n_129),
.B(n_189),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1015),
.A2(n_120),
.B(n_187),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_958),
.Y(n_1201)
);

CKINVDCx10_ASAP7_75t_R g1202 ( 
.A(n_979),
.Y(n_1202)
);

O2A1O1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_1014),
.A2(n_57),
.B(n_59),
.C(n_63),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_1044),
.Y(n_1204)
);

BUFx2_ASAP7_75t_L g1205 ( 
.A(n_929),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_986),
.B(n_63),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_976),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_936),
.A2(n_1022),
.B(n_971),
.Y(n_1208)
);

AND3x1_ASAP7_75t_SL g1209 ( 
.A(n_961),
.B(n_65),
.C(n_66),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_962),
.B(n_65),
.Y(n_1210)
);

OR2x2_ASAP7_75t_L g1211 ( 
.A(n_986),
.B(n_66),
.Y(n_1211)
);

O2A1O1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1017),
.A2(n_67),
.B(n_68),
.C(n_500),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_988),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_900),
.B(n_67),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_960),
.B(n_68),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_936),
.A2(n_1005),
.B(n_1007),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_929),
.B(n_500),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1018),
.A2(n_70),
.B1(n_88),
.B2(n_97),
.Y(n_1218)
);

BUFx2_ASAP7_75t_L g1219 ( 
.A(n_929),
.Y(n_1219)
);

AOI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_929),
.A2(n_98),
.B1(n_107),
.B2(n_116),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_979),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_952),
.A2(n_133),
.B(n_134),
.Y(n_1222)
);

NAND2x1p5_ASAP7_75t_L g1223 ( 
.A(n_922),
.B(n_135),
.Y(n_1223)
);

O2A1O1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_990),
.A2(n_138),
.B(n_155),
.C(n_157),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_900),
.B(n_163),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_911),
.B(n_165),
.Y(n_1226)
);

AOI21xp33_ASAP7_75t_L g1227 ( 
.A1(n_884),
.A2(n_177),
.B(n_180),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_987),
.A2(n_1057),
.B(n_960),
.C(n_1062),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1080),
.A2(n_889),
.B(n_991),
.Y(n_1229)
);

NOR2xp67_ASAP7_75t_SL g1230 ( 
.A(n_1134),
.B(n_947),
.Y(n_1230)
);

NAND2x1p5_ASAP7_75t_L g1231 ( 
.A(n_1083),
.B(n_956),
.Y(n_1231)
);

BUFx4f_ASAP7_75t_SL g1232 ( 
.A(n_1077),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1080),
.A2(n_889),
.B(n_991),
.Y(n_1233)
);

A2O1A1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_1079),
.A2(n_1036),
.B(n_970),
.C(n_932),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1084),
.B(n_1006),
.Y(n_1235)
);

OR2x2_ASAP7_75t_L g1236 ( 
.A(n_1152),
.B(n_935),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1167),
.A2(n_1010),
.B(n_1004),
.Y(n_1237)
);

AO31x2_ASAP7_75t_L g1238 ( 
.A1(n_1148),
.A2(n_1045),
.A3(n_1052),
.B(n_1059),
.Y(n_1238)
);

BUFx2_ASAP7_75t_SL g1239 ( 
.A(n_1181),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1086),
.A2(n_1010),
.B(n_1024),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1208),
.A2(n_1145),
.B(n_1091),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_1092),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_1092),
.Y(n_1243)
);

CKINVDCx20_ASAP7_75t_R g1244 ( 
.A(n_1077),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1081),
.A2(n_1001),
.B1(n_1003),
.B2(n_1038),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1091),
.A2(n_1024),
.B(n_1033),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1216),
.A2(n_1020),
.B(n_926),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1168),
.A2(n_1033),
.B(n_1051),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1172),
.A2(n_1045),
.B(n_1052),
.Y(n_1249)
);

HB1xp67_ASAP7_75t_L g1250 ( 
.A(n_1144),
.Y(n_1250)
);

OA22x2_ASAP7_75t_L g1251 ( 
.A1(n_1195),
.A2(n_894),
.B1(n_970),
.B2(n_1042),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1094),
.A2(n_1059),
.B(n_983),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1088),
.B(n_973),
.Y(n_1253)
);

INVxp67_ASAP7_75t_SL g1254 ( 
.A(n_1140),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1170),
.B(n_911),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1099),
.A2(n_1071),
.B(n_964),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_1144),
.B(n_972),
.Y(n_1257)
);

OAI21xp33_ASAP7_75t_L g1258 ( 
.A1(n_1196),
.A2(n_1042),
.B(n_959),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1116),
.B(n_1008),
.Y(n_1259)
);

INVx3_ASAP7_75t_L g1260 ( 
.A(n_1191),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1102),
.A2(n_1011),
.B(n_1016),
.Y(n_1261)
);

BUFx2_ASAP7_75t_L g1262 ( 
.A(n_1120),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_1092),
.Y(n_1263)
);

OAI22x1_ASAP7_75t_L g1264 ( 
.A1(n_1169),
.A2(n_1042),
.B1(n_1019),
.B2(n_1032),
.Y(n_1264)
);

AO22x2_ASAP7_75t_L g1265 ( 
.A1(n_1093),
.A2(n_1027),
.B1(n_1034),
.B2(n_978),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_L g1266 ( 
.A(n_1097),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1089),
.A2(n_941),
.B(n_925),
.Y(n_1267)
);

OAI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1078),
.A2(n_884),
.B(n_1068),
.Y(n_1268)
);

OAI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1093),
.A2(n_951),
.B(n_980),
.Y(n_1269)
);

AND2x4_ASAP7_75t_L g1270 ( 
.A(n_1085),
.B(n_941),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1161),
.A2(n_992),
.B(n_983),
.Y(n_1271)
);

INVx5_ASAP7_75t_L g1272 ( 
.A(n_1194),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1175),
.B(n_972),
.Y(n_1273)
);

AOI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1073),
.A2(n_997),
.B1(n_967),
.B2(n_925),
.Y(n_1274)
);

BUFx5_ASAP7_75t_L g1275 ( 
.A(n_1194),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1090),
.A2(n_980),
.B(n_997),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1164),
.A2(n_998),
.B(n_992),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1139),
.B(n_998),
.Y(n_1278)
);

OAI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1154),
.A2(n_997),
.B(n_1009),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1178),
.A2(n_978),
.B(n_999),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1103),
.A2(n_947),
.B(n_956),
.Y(n_1281)
);

A2O1A1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_1087),
.A2(n_1043),
.B(n_996),
.C(n_1037),
.Y(n_1282)
);

NOR4xp25_ASAP7_75t_L g1283 ( 
.A(n_1138),
.B(n_996),
.C(n_1016),
.D(n_1011),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1222),
.A2(n_947),
.B(n_967),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1100),
.B(n_999),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1228),
.A2(n_967),
.B(n_1009),
.Y(n_1286)
);

AOI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1186),
.A2(n_1177),
.B1(n_1156),
.B2(n_1124),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1107),
.Y(n_1288)
);

BUFx8_ASAP7_75t_SL g1289 ( 
.A(n_1076),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1132),
.A2(n_887),
.B(n_892),
.Y(n_1290)
);

A2O1A1Ixp33_ASAP7_75t_L g1291 ( 
.A1(n_1214),
.A2(n_1037),
.B(n_967),
.C(n_1050),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1123),
.B(n_887),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1184),
.A2(n_892),
.B(n_896),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1160),
.Y(n_1294)
);

INVxp67_ASAP7_75t_SL g1295 ( 
.A(n_1105),
.Y(n_1295)
);

AO31x2_ASAP7_75t_L g1296 ( 
.A1(n_1157),
.A2(n_896),
.A3(n_907),
.B(n_908),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1162),
.B(n_907),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1154),
.A2(n_908),
.B(n_946),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1200),
.A2(n_946),
.B(n_948),
.Y(n_1299)
);

OR2x6_ASAP7_75t_L g1300 ( 
.A(n_1191),
.B(n_948),
.Y(n_1300)
);

BUFx3_ASAP7_75t_L g1301 ( 
.A(n_1076),
.Y(n_1301)
);

OAI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1171),
.A2(n_997),
.B(n_1050),
.Y(n_1302)
);

AOI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1184),
.A2(n_949),
.B(n_950),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1098),
.B(n_949),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1206),
.A2(n_950),
.B1(n_954),
.B2(n_997),
.Y(n_1305)
);

AOI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1109),
.A2(n_954),
.B1(n_1206),
.B2(n_1135),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1174),
.B(n_1183),
.Y(n_1307)
);

AO21x2_ASAP7_75t_L g1308 ( 
.A1(n_1227),
.A2(n_1125),
.B(n_1150),
.Y(n_1308)
);

OR2x6_ASAP7_75t_L g1309 ( 
.A(n_1191),
.B(n_1205),
.Y(n_1309)
);

AOI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1192),
.A2(n_1163),
.B(n_1179),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1119),
.B(n_1211),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1201),
.B(n_1213),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1199),
.A2(n_1151),
.B(n_1153),
.Y(n_1313)
);

NAND3xp33_ASAP7_75t_L g1314 ( 
.A(n_1173),
.B(n_1130),
.C(n_1128),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_1165),
.Y(n_1315)
);

INVx3_ASAP7_75t_L g1316 ( 
.A(n_1085),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1110),
.B(n_1155),
.Y(n_1317)
);

OR2x2_ASAP7_75t_L g1318 ( 
.A(n_1185),
.B(n_1187),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1189),
.B(n_1204),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1182),
.A2(n_1136),
.B(n_1112),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1223),
.A2(n_1074),
.B(n_1112),
.Y(n_1321)
);

INVx3_ASAP7_75t_L g1322 ( 
.A(n_1097),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_SL g1323 ( 
.A(n_1083),
.B(n_1141),
.Y(n_1323)
);

AOI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1176),
.A2(n_1188),
.B(n_1122),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1223),
.A2(n_1074),
.B(n_1136),
.Y(n_1325)
);

NAND2xp33_ASAP7_75t_L g1326 ( 
.A(n_1194),
.B(n_1075),
.Y(n_1326)
);

AOI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1114),
.A2(n_1131),
.B(n_1127),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1221),
.B(n_1115),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1166),
.B(n_1143),
.Y(n_1329)
);

AO31x2_ASAP7_75t_L g1330 ( 
.A1(n_1147),
.A2(n_1190),
.A3(n_1197),
.B(n_1158),
.Y(n_1330)
);

BUFx3_ASAP7_75t_L g1331 ( 
.A(n_1134),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1182),
.A2(n_1218),
.B(n_1146),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1193),
.A2(n_1198),
.B1(n_1210),
.B2(n_1141),
.Y(n_1333)
);

OA21x2_ASAP7_75t_L g1334 ( 
.A1(n_1227),
.A2(n_1117),
.B(n_1207),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1106),
.B(n_1226),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1217),
.A2(n_1096),
.B(n_1224),
.Y(n_1336)
);

NAND2x1p5_ASAP7_75t_L g1337 ( 
.A(n_1219),
.B(n_1101),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1202),
.B(n_1149),
.Y(n_1338)
);

AO21x2_ASAP7_75t_L g1339 ( 
.A1(n_1126),
.A2(n_1118),
.B(n_1217),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1104),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1180),
.B(n_1159),
.Y(n_1341)
);

AO31x2_ASAP7_75t_L g1342 ( 
.A1(n_1218),
.A2(n_1225),
.A3(n_1209),
.B(n_1095),
.Y(n_1342)
);

BUFx10_ASAP7_75t_L g1343 ( 
.A(n_1101),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_SL g1344 ( 
.A(n_1101),
.B(n_1180),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1159),
.B(n_1194),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1220),
.A2(n_1212),
.B(n_1215),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1133),
.B(n_1111),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1146),
.Y(n_1348)
);

AO21x1_ASAP7_75t_L g1349 ( 
.A1(n_1203),
.A2(n_1142),
.B(n_1129),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1146),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1108),
.A2(n_1137),
.B(n_1121),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1113),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1152),
.B(n_886),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1086),
.A2(n_1208),
.B(n_1145),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1080),
.A2(n_843),
.B1(n_1054),
.B2(n_401),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1152),
.B(n_886),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1152),
.B(n_886),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1152),
.B(n_886),
.Y(n_1358)
);

O2A1O1Ixp33_ASAP7_75t_SL g1359 ( 
.A1(n_1084),
.A2(n_890),
.B(n_1080),
.C(n_886),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1152),
.B(n_886),
.Y(n_1360)
);

INVx1_ASAP7_75t_SL g1361 ( 
.A(n_1144),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1082),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1080),
.A2(n_890),
.B(n_904),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1152),
.B(n_886),
.Y(n_1364)
);

NAND2x1p5_ASAP7_75t_L g1365 ( 
.A(n_1083),
.B(n_1141),
.Y(n_1365)
);

NAND3xp33_ASAP7_75t_L g1366 ( 
.A(n_1080),
.B(n_890),
.C(n_886),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1081),
.B(n_1012),
.Y(n_1367)
);

NAND3x1_ASAP7_75t_L g1368 ( 
.A(n_1081),
.B(n_1169),
.C(n_1075),
.Y(n_1368)
);

OAI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1081),
.A2(n_1012),
.B1(n_890),
.B2(n_1080),
.Y(n_1369)
);

A2O1A1Ixp33_ASAP7_75t_L g1370 ( 
.A1(n_1079),
.A2(n_886),
.B(n_1080),
.C(n_1078),
.Y(n_1370)
);

AOI211x1_ASAP7_75t_L g1371 ( 
.A1(n_1080),
.A2(n_1170),
.B(n_776),
.C(n_1185),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1080),
.A2(n_890),
.B(n_904),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1082),
.Y(n_1373)
);

OAI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1080),
.A2(n_886),
.B(n_890),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1080),
.B(n_886),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1181),
.Y(n_1376)
);

INVxp67_ASAP7_75t_SL g1377 ( 
.A(n_1140),
.Y(n_1377)
);

AND2x4_ASAP7_75t_L g1378 ( 
.A(n_1085),
.B(n_1144),
.Y(n_1378)
);

BUFx2_ASAP7_75t_L g1379 ( 
.A(n_1120),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1080),
.A2(n_890),
.B(n_904),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1080),
.A2(n_890),
.B1(n_886),
.B2(n_1081),
.Y(n_1381)
);

INVx4_ASAP7_75t_L g1382 ( 
.A(n_1191),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1086),
.A2(n_1208),
.B(n_1145),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1080),
.A2(n_890),
.B1(n_886),
.B2(n_1081),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1080),
.A2(n_890),
.B(n_904),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1080),
.A2(n_890),
.B(n_904),
.Y(n_1386)
);

AO21x1_ASAP7_75t_L g1387 ( 
.A1(n_1080),
.A2(n_890),
.B(n_1079),
.Y(n_1387)
);

AO31x2_ASAP7_75t_L g1388 ( 
.A1(n_1167),
.A2(n_1148),
.A3(n_1228),
.B(n_1103),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1080),
.A2(n_890),
.B(n_904),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1238),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1238),
.Y(n_1391)
);

OR2x2_ASAP7_75t_L g1392 ( 
.A(n_1254),
.B(n_1377),
.Y(n_1392)
);

OR2x2_ASAP7_75t_L g1393 ( 
.A(n_1307),
.B(n_1361),
.Y(n_1393)
);

INVx6_ASAP7_75t_L g1394 ( 
.A(n_1343),
.Y(n_1394)
);

AOI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1333),
.A2(n_1332),
.B(n_1324),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1354),
.A2(n_1383),
.B(n_1313),
.Y(n_1396)
);

AOI222xp33_ASAP7_75t_L g1397 ( 
.A1(n_1355),
.A2(n_1381),
.B1(n_1384),
.B2(n_1374),
.C1(n_1375),
.C2(n_1369),
.Y(n_1397)
);

OAI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1366),
.A2(n_1384),
.B(n_1381),
.Y(n_1398)
);

INVx8_ASAP7_75t_L g1399 ( 
.A(n_1289),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1375),
.A2(n_1366),
.B1(n_1374),
.B2(n_1367),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1238),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1265),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1241),
.A2(n_1247),
.B(n_1277),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1307),
.Y(n_1404)
);

AND2x4_ASAP7_75t_L g1405 ( 
.A(n_1378),
.B(n_1309),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1336),
.A2(n_1303),
.B(n_1321),
.Y(n_1406)
);

AND2x2_ASAP7_75t_SL g1407 ( 
.A(n_1323),
.B(n_1283),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1287),
.A2(n_1370),
.B1(n_1357),
.B2(n_1353),
.Y(n_1408)
);

BUFx2_ASAP7_75t_L g1409 ( 
.A(n_1262),
.Y(n_1409)
);

BUFx8_ASAP7_75t_L g1410 ( 
.A(n_1301),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1325),
.A2(n_1237),
.B(n_1261),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1311),
.B(n_1250),
.Y(n_1412)
);

BUFx3_ASAP7_75t_L g1413 ( 
.A(n_1331),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1255),
.A2(n_1251),
.B1(n_1387),
.B2(n_1314),
.Y(n_1414)
);

BUFx2_ASAP7_75t_L g1415 ( 
.A(n_1379),
.Y(n_1415)
);

OA21x2_ASAP7_75t_L g1416 ( 
.A1(n_1276),
.A2(n_1268),
.B(n_1302),
.Y(n_1416)
);

AOI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1333),
.A2(n_1372),
.B(n_1363),
.Y(n_1417)
);

AND2x4_ASAP7_75t_L g1418 ( 
.A(n_1378),
.B(n_1309),
.Y(n_1418)
);

INVxp67_ASAP7_75t_L g1419 ( 
.A(n_1376),
.Y(n_1419)
);

AOI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1380),
.A2(n_1389),
.B(n_1386),
.Y(n_1420)
);

A2O1A1Ixp33_ASAP7_75t_L g1421 ( 
.A1(n_1385),
.A2(n_1268),
.B(n_1258),
.C(n_1314),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1240),
.A2(n_1249),
.B(n_1280),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1293),
.A2(n_1246),
.B(n_1252),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1356),
.B(n_1358),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1320),
.A2(n_1271),
.B(n_1248),
.Y(n_1425)
);

A2O1A1Ixp33_ASAP7_75t_L g1426 ( 
.A1(n_1302),
.A2(n_1276),
.B(n_1269),
.C(n_1229),
.Y(n_1426)
);

AOI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1267),
.A2(n_1235),
.B(n_1233),
.Y(n_1427)
);

OAI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1290),
.A2(n_1299),
.B(n_1298),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1286),
.A2(n_1284),
.B(n_1279),
.Y(n_1429)
);

AO21x1_ASAP7_75t_L g1430 ( 
.A1(n_1245),
.A2(n_1235),
.B(n_1295),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1360),
.B(n_1364),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1312),
.Y(n_1432)
);

OAI221xp5_ASAP7_75t_L g1433 ( 
.A1(n_1245),
.A2(n_1306),
.B1(n_1318),
.B2(n_1359),
.C(n_1283),
.Y(n_1433)
);

AO21x2_ASAP7_75t_L g1434 ( 
.A1(n_1279),
.A2(n_1269),
.B(n_1308),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1281),
.A2(n_1327),
.B(n_1256),
.Y(n_1435)
);

NAND3xp33_ASAP7_75t_SL g1436 ( 
.A(n_1347),
.B(n_1349),
.C(n_1329),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1265),
.Y(n_1437)
);

CKINVDCx20_ASAP7_75t_R g1438 ( 
.A(n_1244),
.Y(n_1438)
);

AO21x1_ASAP7_75t_L g1439 ( 
.A1(n_1305),
.A2(n_1335),
.B(n_1346),
.Y(n_1439)
);

AOI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1368),
.A2(n_1273),
.B1(n_1317),
.B2(n_1239),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1305),
.A2(n_1334),
.B(n_1351),
.Y(n_1441)
);

AOI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1285),
.A2(n_1310),
.B(n_1264),
.Y(n_1442)
);

AOI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1323),
.A2(n_1361),
.B1(n_1257),
.B2(n_1230),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1371),
.A2(n_1272),
.B1(n_1274),
.B2(n_1236),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1341),
.B(n_1253),
.Y(n_1445)
);

INVx3_ASAP7_75t_L g1446 ( 
.A(n_1242),
.Y(n_1446)
);

NOR2x1_ASAP7_75t_SL g1447 ( 
.A(n_1300),
.B(n_1345),
.Y(n_1447)
);

NAND3xp33_ASAP7_75t_L g1448 ( 
.A(n_1234),
.B(n_1253),
.C(n_1291),
.Y(n_1448)
);

AO32x2_ASAP7_75t_L g1449 ( 
.A1(n_1251),
.A2(n_1388),
.A3(n_1382),
.B1(n_1296),
.B2(n_1334),
.Y(n_1449)
);

AOI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1285),
.A2(n_1345),
.B(n_1344),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1341),
.B(n_1278),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1292),
.A2(n_1297),
.B(n_1337),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1292),
.A2(n_1297),
.B(n_1337),
.Y(n_1453)
);

AOI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1319),
.A2(n_1270),
.B1(n_1326),
.B2(n_1348),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1340),
.A2(n_1316),
.B(n_1260),
.Y(n_1455)
);

BUFx2_ASAP7_75t_L g1456 ( 
.A(n_1242),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1316),
.A2(n_1260),
.B(n_1373),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1288),
.A2(n_1362),
.B(n_1294),
.Y(n_1458)
);

AOI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1304),
.A2(n_1300),
.B(n_1350),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1365),
.B(n_1231),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1296),
.Y(n_1461)
);

O2A1O1Ixp33_ASAP7_75t_L g1462 ( 
.A1(n_1282),
.A2(n_1352),
.B(n_1259),
.C(n_1308),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1242),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_SL g1464 ( 
.A1(n_1382),
.A2(n_1328),
.B(n_1342),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1296),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_SL g1466 ( 
.A1(n_1342),
.A2(n_1275),
.B(n_1339),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1300),
.A2(n_1365),
.B1(n_1339),
.B2(n_1270),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1330),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1330),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_SL g1470 ( 
.A1(n_1342),
.A2(n_1275),
.B(n_1343),
.Y(n_1470)
);

OAI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1322),
.A2(n_1231),
.B(n_1388),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_SL g1472 ( 
.A(n_1275),
.B(n_1243),
.Y(n_1472)
);

OAI21x1_ASAP7_75t_L g1473 ( 
.A1(n_1322),
.A2(n_1388),
.B(n_1275),
.Y(n_1473)
);

AO31x2_ASAP7_75t_L g1474 ( 
.A1(n_1330),
.A2(n_1275),
.A3(n_1243),
.B(n_1263),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1263),
.Y(n_1475)
);

AO31x2_ASAP7_75t_L g1476 ( 
.A1(n_1266),
.A2(n_1387),
.A3(n_1247),
.B(n_1167),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1232),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1354),
.A2(n_1383),
.B(n_1313),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1353),
.B(n_1356),
.Y(n_1479)
);

NAND3xp33_ASAP7_75t_L g1480 ( 
.A(n_1381),
.B(n_1384),
.C(n_1081),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1375),
.A2(n_890),
.B1(n_1366),
.B2(n_1381),
.Y(n_1481)
);

INVx1_ASAP7_75t_SL g1482 ( 
.A(n_1239),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1238),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1378),
.B(n_1309),
.Y(n_1484)
);

AOI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1333),
.A2(n_1145),
.B(n_1332),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1262),
.Y(n_1486)
);

INVx3_ASAP7_75t_L g1487 ( 
.A(n_1272),
.Y(n_1487)
);

NAND2xp33_ASAP7_75t_R g1488 ( 
.A(n_1375),
.B(n_1374),
.Y(n_1488)
);

NAND3xp33_ASAP7_75t_SL g1489 ( 
.A(n_1287),
.B(n_1081),
.C(n_1012),
.Y(n_1489)
);

NAND2x1p5_ASAP7_75t_L g1490 ( 
.A(n_1272),
.B(n_1083),
.Y(n_1490)
);

A2O1A1Ixp33_ASAP7_75t_L g1491 ( 
.A1(n_1374),
.A2(n_886),
.B(n_1375),
.C(n_1366),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1311),
.B(n_1181),
.Y(n_1492)
);

INVx3_ASAP7_75t_L g1493 ( 
.A(n_1272),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1354),
.A2(n_1383),
.B(n_1313),
.Y(n_1494)
);

OA21x2_ASAP7_75t_L g1495 ( 
.A1(n_1241),
.A2(n_1354),
.B(n_1383),
.Y(n_1495)
);

AOI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1375),
.A2(n_1374),
.B(n_1359),
.Y(n_1496)
);

CKINVDCx20_ASAP7_75t_R g1497 ( 
.A(n_1244),
.Y(n_1497)
);

NOR2x1_ASAP7_75t_R g1498 ( 
.A(n_1315),
.B(n_834),
.Y(n_1498)
);

OAI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1366),
.A2(n_1384),
.B(n_1381),
.Y(n_1499)
);

OAI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1366),
.A2(n_1384),
.B(n_1381),
.Y(n_1500)
);

INVx8_ASAP7_75t_L g1501 ( 
.A(n_1289),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1375),
.A2(n_890),
.B1(n_1366),
.B2(n_1381),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1311),
.B(n_1181),
.Y(n_1503)
);

BUFx3_ASAP7_75t_L g1504 ( 
.A(n_1331),
.Y(n_1504)
);

OA21x2_ASAP7_75t_L g1505 ( 
.A1(n_1241),
.A2(n_1354),
.B(n_1383),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1238),
.Y(n_1506)
);

INVx3_ASAP7_75t_L g1507 ( 
.A(n_1272),
.Y(n_1507)
);

BUFx3_ASAP7_75t_L g1508 ( 
.A(n_1331),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1238),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1311),
.B(n_1181),
.Y(n_1510)
);

INVx8_ASAP7_75t_L g1511 ( 
.A(n_1289),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1307),
.Y(n_1512)
);

OAI21x1_ASAP7_75t_SL g1513 ( 
.A1(n_1374),
.A2(n_1375),
.B(n_1387),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1307),
.Y(n_1514)
);

AND2x4_ASAP7_75t_L g1515 ( 
.A(n_1378),
.B(n_1309),
.Y(n_1515)
);

OAI21x1_ASAP7_75t_L g1516 ( 
.A1(n_1354),
.A2(n_1383),
.B(n_1313),
.Y(n_1516)
);

AO21x2_ASAP7_75t_L g1517 ( 
.A1(n_1268),
.A2(n_1302),
.B(n_1276),
.Y(n_1517)
);

BUFx10_ASAP7_75t_L g1518 ( 
.A(n_1338),
.Y(n_1518)
);

NAND2x1p5_ASAP7_75t_L g1519 ( 
.A(n_1272),
.B(n_1083),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1381),
.B(n_1384),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1311),
.B(n_1181),
.Y(n_1521)
);

NAND2x1p5_ASAP7_75t_L g1522 ( 
.A(n_1272),
.B(n_1083),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1355),
.A2(n_1384),
.B1(n_1381),
.B2(n_1080),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1238),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1254),
.B(n_1377),
.Y(n_1525)
);

OAI21x1_ASAP7_75t_L g1526 ( 
.A1(n_1354),
.A2(n_1383),
.B(n_1313),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1307),
.Y(n_1527)
);

AOI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1375),
.A2(n_1374),
.B(n_1359),
.Y(n_1528)
);

AOI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1375),
.A2(n_1374),
.B(n_1359),
.Y(n_1529)
);

AO21x2_ASAP7_75t_L g1530 ( 
.A1(n_1268),
.A2(n_1302),
.B(n_1276),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1355),
.A2(n_1384),
.B1(n_1381),
.B2(n_1080),
.Y(n_1531)
);

AO31x2_ASAP7_75t_L g1532 ( 
.A1(n_1387),
.A2(n_1247),
.A3(n_1167),
.B(n_1228),
.Y(n_1532)
);

AOI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1375),
.A2(n_1374),
.B(n_1359),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1412),
.B(n_1492),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1393),
.B(n_1392),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1503),
.B(n_1510),
.Y(n_1536)
);

O2A1O1Ixp5_ASAP7_75t_L g1537 ( 
.A1(n_1520),
.A2(n_1499),
.B(n_1500),
.C(n_1398),
.Y(n_1537)
);

A2O1A1Ixp33_ASAP7_75t_L g1538 ( 
.A1(n_1523),
.A2(n_1531),
.B(n_1520),
.C(n_1480),
.Y(n_1538)
);

OA21x2_ASAP7_75t_L g1539 ( 
.A1(n_1435),
.A2(n_1441),
.B(n_1406),
.Y(n_1539)
);

BUFx3_ASAP7_75t_L g1540 ( 
.A(n_1413),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1521),
.B(n_1409),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1523),
.A2(n_1531),
.B1(n_1400),
.B2(n_1491),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1525),
.Y(n_1543)
);

AOI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1481),
.A2(n_1502),
.B(n_1421),
.Y(n_1544)
);

AOI21xp5_ASAP7_75t_SL g1545 ( 
.A1(n_1462),
.A2(n_1491),
.B(n_1421),
.Y(n_1545)
);

BUFx6f_ASAP7_75t_L g1546 ( 
.A(n_1413),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1415),
.B(n_1486),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1445),
.B(n_1400),
.Y(n_1548)
);

NOR2xp67_ASAP7_75t_L g1549 ( 
.A(n_1436),
.B(n_1489),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1408),
.A2(n_1414),
.B1(n_1433),
.B2(n_1426),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1445),
.B(n_1451),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1451),
.B(n_1404),
.Y(n_1552)
);

NOR2xp67_ASAP7_75t_L g1553 ( 
.A(n_1440),
.B(n_1448),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1414),
.A2(n_1528),
.B1(n_1533),
.B2(n_1496),
.Y(n_1554)
);

AOI21xp5_ASAP7_75t_L g1555 ( 
.A1(n_1529),
.A2(n_1397),
.B(n_1430),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1431),
.B(n_1419),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1424),
.B(n_1479),
.Y(n_1557)
);

AND2x4_ASAP7_75t_L g1558 ( 
.A(n_1405),
.B(n_1418),
.Y(n_1558)
);

O2A1O1Ixp5_ASAP7_75t_L g1559 ( 
.A1(n_1439),
.A2(n_1417),
.B(n_1471),
.C(n_1395),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1512),
.B(n_1514),
.Y(n_1560)
);

O2A1O1Ixp33_ASAP7_75t_L g1561 ( 
.A1(n_1513),
.A2(n_1482),
.B(n_1464),
.C(n_1466),
.Y(n_1561)
);

BUFx12f_ASAP7_75t_L g1562 ( 
.A(n_1518),
.Y(n_1562)
);

AOI21xp5_ASAP7_75t_L g1563 ( 
.A1(n_1517),
.A2(n_1530),
.B(n_1416),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1416),
.A2(n_1407),
.B1(n_1488),
.B2(n_1527),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1432),
.B(n_1517),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1407),
.B(n_1530),
.Y(n_1566)
);

OA21x2_ASAP7_75t_L g1567 ( 
.A1(n_1428),
.A2(n_1494),
.B(n_1478),
.Y(n_1567)
);

AOI21x1_ASAP7_75t_SL g1568 ( 
.A1(n_1399),
.A2(n_1511),
.B(n_1501),
.Y(n_1568)
);

AOI221xp5_ASAP7_75t_L g1569 ( 
.A1(n_1402),
.A2(n_1437),
.B1(n_1444),
.B2(n_1434),
.C(n_1467),
.Y(n_1569)
);

O2A1O1Ixp33_ASAP7_75t_L g1570 ( 
.A1(n_1477),
.A2(n_1463),
.B(n_1475),
.C(n_1470),
.Y(n_1570)
);

AOI21xp5_ASAP7_75t_SL g1571 ( 
.A1(n_1490),
.A2(n_1519),
.B(n_1522),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1456),
.B(n_1405),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1452),
.B(n_1453),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1402),
.B(n_1437),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1488),
.A2(n_1454),
.B1(n_1443),
.B2(n_1484),
.Y(n_1575)
);

OA21x2_ASAP7_75t_L g1576 ( 
.A1(n_1428),
.A2(n_1478),
.B(n_1526),
.Y(n_1576)
);

AOI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1472),
.A2(n_1429),
.B(n_1411),
.Y(n_1577)
);

OA21x2_ASAP7_75t_L g1578 ( 
.A1(n_1396),
.A2(n_1526),
.B(n_1516),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1532),
.B(n_1476),
.Y(n_1579)
);

BUFx2_ASAP7_75t_L g1580 ( 
.A(n_1410),
.Y(n_1580)
);

A2O1A1Ixp33_ASAP7_75t_L g1581 ( 
.A1(n_1429),
.A2(n_1460),
.B(n_1473),
.C(n_1455),
.Y(n_1581)
);

AOI221xp5_ASAP7_75t_L g1582 ( 
.A1(n_1483),
.A2(n_1468),
.B1(n_1469),
.B2(n_1504),
.C(n_1508),
.Y(n_1582)
);

INVx3_ASAP7_75t_SL g1583 ( 
.A(n_1399),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1532),
.B(n_1476),
.Y(n_1584)
);

A2O1A1Ixp33_ASAP7_75t_L g1585 ( 
.A1(n_1473),
.A2(n_1455),
.B(n_1484),
.C(n_1515),
.Y(n_1585)
);

OAI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1484),
.A2(n_1420),
.B1(n_1522),
.B2(n_1519),
.Y(n_1586)
);

AOI21x1_ASAP7_75t_SL g1587 ( 
.A1(n_1399),
.A2(n_1511),
.B(n_1501),
.Y(n_1587)
);

AOI21x1_ASAP7_75t_SL g1588 ( 
.A1(n_1501),
.A2(n_1511),
.B(n_1498),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1446),
.B(n_1450),
.Y(n_1589)
);

O2A1O1Ixp5_ASAP7_75t_L g1590 ( 
.A1(n_1485),
.A2(n_1427),
.B(n_1442),
.C(n_1493),
.Y(n_1590)
);

O2A1O1Ixp33_ASAP7_75t_L g1591 ( 
.A1(n_1487),
.A2(n_1507),
.B(n_1483),
.C(n_1468),
.Y(n_1591)
);

AND2x4_ASAP7_75t_L g1592 ( 
.A(n_1447),
.B(n_1474),
.Y(n_1592)
);

OAI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1394),
.A2(n_1497),
.B1(n_1438),
.B2(n_1507),
.Y(n_1593)
);

AOI21xp5_ASAP7_75t_SL g1594 ( 
.A1(n_1469),
.A2(n_1495),
.B(n_1505),
.Y(n_1594)
);

O2A1O1Ixp5_ASAP7_75t_L g1595 ( 
.A1(n_1459),
.A2(n_1461),
.B(n_1465),
.C(n_1390),
.Y(n_1595)
);

OA21x2_ASAP7_75t_L g1596 ( 
.A1(n_1396),
.A2(n_1516),
.B(n_1494),
.Y(n_1596)
);

INVx4_ASAP7_75t_L g1597 ( 
.A(n_1518),
.Y(n_1597)
);

OA21x2_ASAP7_75t_L g1598 ( 
.A1(n_1411),
.A2(n_1403),
.B(n_1422),
.Y(n_1598)
);

O2A1O1Ixp33_ASAP7_75t_L g1599 ( 
.A1(n_1438),
.A2(n_1497),
.B(n_1465),
.C(n_1461),
.Y(n_1599)
);

OAI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1532),
.A2(n_1390),
.B1(n_1391),
.B2(n_1401),
.Y(n_1600)
);

OAI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1391),
.A2(n_1401),
.B1(n_1509),
.B2(n_1506),
.Y(n_1601)
);

INVx3_ASAP7_75t_SL g1602 ( 
.A(n_1518),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1476),
.B(n_1474),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1474),
.B(n_1457),
.Y(n_1604)
);

OAI22xp5_ASAP7_75t_SL g1605 ( 
.A1(n_1410),
.A2(n_1449),
.B1(n_1505),
.B2(n_1495),
.Y(n_1605)
);

CKINVDCx20_ASAP7_75t_R g1606 ( 
.A(n_1410),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1457),
.B(n_1524),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1506),
.A2(n_1509),
.B1(n_1505),
.B2(n_1495),
.Y(n_1608)
);

OAI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1449),
.A2(n_1403),
.B1(n_1425),
.B2(n_1423),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1425),
.B(n_1423),
.Y(n_1610)
);

HB1xp67_ASAP7_75t_L g1611 ( 
.A(n_1422),
.Y(n_1611)
);

INVx5_ASAP7_75t_L g1612 ( 
.A(n_1449),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1449),
.Y(n_1613)
);

OA21x2_ASAP7_75t_L g1614 ( 
.A1(n_1435),
.A2(n_1441),
.B(n_1406),
.Y(n_1614)
);

AOI21x1_ASAP7_75t_SL g1615 ( 
.A1(n_1424),
.A2(n_1347),
.B(n_1375),
.Y(n_1615)
);

CKINVDCx16_ASAP7_75t_R g1616 ( 
.A(n_1438),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1393),
.B(n_1392),
.Y(n_1617)
);

A2O1A1Ixp33_ASAP7_75t_L g1618 ( 
.A1(n_1523),
.A2(n_1081),
.B(n_1367),
.C(n_1080),
.Y(n_1618)
);

NOR2xp67_ASAP7_75t_L g1619 ( 
.A(n_1436),
.B(n_1489),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1393),
.B(n_1392),
.Y(n_1620)
);

AOI21xp5_ASAP7_75t_SL g1621 ( 
.A1(n_1462),
.A2(n_1375),
.B(n_1381),
.Y(n_1621)
);

AOI21xp5_ASAP7_75t_SL g1622 ( 
.A1(n_1462),
.A2(n_1375),
.B(n_1381),
.Y(n_1622)
);

AOI21x1_ASAP7_75t_SL g1623 ( 
.A1(n_1424),
.A2(n_1347),
.B(n_1375),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1458),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1458),
.Y(n_1625)
);

AOI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1481),
.A2(n_1375),
.B(n_1374),
.Y(n_1626)
);

AOI21xp5_ASAP7_75t_SL g1627 ( 
.A1(n_1462),
.A2(n_1375),
.B(n_1381),
.Y(n_1627)
);

O2A1O1Ixp33_ASAP7_75t_L g1628 ( 
.A1(n_1489),
.A2(n_1369),
.B(n_1384),
.C(n_1381),
.Y(n_1628)
);

O2A1O1Ixp33_ASAP7_75t_L g1629 ( 
.A1(n_1489),
.A2(n_1369),
.B(n_1384),
.C(n_1381),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1520),
.B(n_1445),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1393),
.B(n_1392),
.Y(n_1631)
);

AOI21xp5_ASAP7_75t_L g1632 ( 
.A1(n_1481),
.A2(n_1375),
.B(n_1374),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1393),
.B(n_1392),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_SL g1634 ( 
.A1(n_1523),
.A2(n_1367),
.B1(n_1531),
.B2(n_1497),
.Y(n_1634)
);

OA21x2_ASAP7_75t_L g1635 ( 
.A1(n_1435),
.A2(n_1441),
.B(n_1406),
.Y(n_1635)
);

AOI21xp5_ASAP7_75t_SL g1636 ( 
.A1(n_1462),
.A2(n_1375),
.B(n_1381),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1626),
.B(n_1632),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1565),
.Y(n_1638)
);

AND2x4_ASAP7_75t_L g1639 ( 
.A(n_1592),
.B(n_1585),
.Y(n_1639)
);

XNOR2xp5_ASAP7_75t_L g1640 ( 
.A(n_1634),
.B(n_1550),
.Y(n_1640)
);

AO21x2_ASAP7_75t_L g1641 ( 
.A1(n_1563),
.A2(n_1608),
.B(n_1594),
.Y(n_1641)
);

BUFx6f_ASAP7_75t_L g1642 ( 
.A(n_1610),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1566),
.B(n_1612),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1566),
.B(n_1543),
.Y(n_1644)
);

INVx2_ASAP7_75t_SL g1645 ( 
.A(n_1589),
.Y(n_1645)
);

INVxp67_ASAP7_75t_L g1646 ( 
.A(n_1604),
.Y(n_1646)
);

NOR2x1_ASAP7_75t_L g1647 ( 
.A(n_1621),
.B(n_1622),
.Y(n_1647)
);

AO21x2_ASAP7_75t_L g1648 ( 
.A1(n_1579),
.A2(n_1584),
.B(n_1609),
.Y(n_1648)
);

NAND3xp33_ASAP7_75t_L g1649 ( 
.A(n_1618),
.B(n_1544),
.C(n_1550),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1613),
.B(n_1535),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1581),
.B(n_1624),
.Y(n_1651)
);

OAI21x1_ASAP7_75t_L g1652 ( 
.A1(n_1559),
.A2(n_1590),
.B(n_1577),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1560),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1625),
.Y(n_1654)
);

INVxp67_ASAP7_75t_L g1655 ( 
.A(n_1604),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1560),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1612),
.B(n_1610),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_1616),
.Y(n_1658)
);

HB1xp67_ASAP7_75t_L g1659 ( 
.A(n_1573),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1573),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1630),
.B(n_1548),
.Y(n_1661)
);

INVxp67_ASAP7_75t_L g1662 ( 
.A(n_1607),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1612),
.B(n_1564),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1564),
.B(n_1611),
.Y(n_1664)
);

AOI221xp5_ASAP7_75t_L g1665 ( 
.A1(n_1542),
.A2(n_1555),
.B1(n_1545),
.B2(n_1636),
.C(n_1627),
.Y(n_1665)
);

BUFx3_ASAP7_75t_L g1666 ( 
.A(n_1558),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1539),
.Y(n_1667)
);

OA21x2_ASAP7_75t_L g1668 ( 
.A1(n_1603),
.A2(n_1537),
.B(n_1609),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_L g1669 ( 
.A(n_1548),
.B(n_1630),
.Y(n_1669)
);

AO21x2_ASAP7_75t_L g1670 ( 
.A1(n_1600),
.A2(n_1554),
.B(n_1601),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1617),
.B(n_1620),
.Y(n_1671)
);

AO21x2_ASAP7_75t_L g1672 ( 
.A1(n_1600),
.A2(n_1554),
.B(n_1601),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1614),
.B(n_1635),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1614),
.B(n_1635),
.Y(n_1674)
);

INVx3_ASAP7_75t_L g1675 ( 
.A(n_1578),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1556),
.B(n_1567),
.Y(n_1676)
);

OA21x2_ASAP7_75t_L g1677 ( 
.A1(n_1595),
.A2(n_1569),
.B(n_1582),
.Y(n_1677)
);

OR2x6_ASAP7_75t_L g1678 ( 
.A(n_1571),
.B(n_1591),
.Y(n_1678)
);

BUFx2_ASAP7_75t_L g1679 ( 
.A(n_1605),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1574),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1552),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1567),
.B(n_1576),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1598),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1552),
.Y(n_1684)
);

OA21x2_ASAP7_75t_L g1685 ( 
.A1(n_1538),
.A2(n_1542),
.B(n_1586),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1598),
.Y(n_1686)
);

BUFx2_ASAP7_75t_L g1687 ( 
.A(n_1576),
.Y(n_1687)
);

OR2x2_ASAP7_75t_SL g1688 ( 
.A(n_1649),
.B(n_1551),
.Y(n_1688)
);

INVx3_ASAP7_75t_L g1689 ( 
.A(n_1642),
.Y(n_1689)
);

AO31x2_ASAP7_75t_L g1690 ( 
.A1(n_1637),
.A2(n_1679),
.A3(n_1638),
.B(n_1687),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1683),
.Y(n_1691)
);

INVxp67_ASAP7_75t_SL g1692 ( 
.A(n_1667),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1640),
.A2(n_1649),
.B1(n_1685),
.B2(n_1665),
.Y(n_1693)
);

BUFx2_ASAP7_75t_SL g1694 ( 
.A(n_1657),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1676),
.B(n_1596),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1644),
.B(n_1633),
.Y(n_1696)
);

OAI21xp5_ASAP7_75t_L g1697 ( 
.A1(n_1640),
.A2(n_1628),
.B(n_1629),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1669),
.B(n_1551),
.Y(n_1698)
);

NOR2xp33_ASAP7_75t_L g1699 ( 
.A(n_1669),
.B(n_1549),
.Y(n_1699)
);

AO21x2_ASAP7_75t_L g1700 ( 
.A1(n_1641),
.A2(n_1686),
.B(n_1670),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1644),
.B(n_1631),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1659),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_L g1703 ( 
.A(n_1661),
.B(n_1619),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1676),
.B(n_1547),
.Y(n_1704)
);

BUFx12f_ASAP7_75t_L g1705 ( 
.A(n_1658),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1644),
.B(n_1557),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1675),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1650),
.B(n_1534),
.Y(n_1708)
);

CKINVDCx20_ASAP7_75t_R g1709 ( 
.A(n_1666),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1661),
.B(n_1561),
.Y(n_1710)
);

HB1xp67_ASAP7_75t_L g1711 ( 
.A(n_1659),
.Y(n_1711)
);

NOR4xp25_ASAP7_75t_SL g1712 ( 
.A(n_1679),
.B(n_1580),
.C(n_1615),
.D(n_1623),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1676),
.B(n_1541),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1657),
.B(n_1663),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1654),
.Y(n_1715)
);

INVxp67_ASAP7_75t_SL g1716 ( 
.A(n_1667),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1660),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1682),
.B(n_1536),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1663),
.B(n_1572),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1654),
.Y(n_1720)
);

OAI21x1_ASAP7_75t_L g1721 ( 
.A1(n_1652),
.A2(n_1575),
.B(n_1599),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_SL g1722 ( 
.A(n_1647),
.B(n_1553),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1675),
.Y(n_1723)
);

AOI22xp33_ASAP7_75t_SL g1724 ( 
.A1(n_1721),
.A2(n_1679),
.B1(n_1685),
.B2(n_1670),
.Y(n_1724)
);

OAI22xp33_ASAP7_75t_L g1725 ( 
.A1(n_1697),
.A2(n_1685),
.B1(n_1665),
.B2(n_1647),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_R g1726 ( 
.A(n_1705),
.B(n_1606),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1696),
.Y(n_1727)
);

NAND3xp33_ASAP7_75t_L g1728 ( 
.A(n_1693),
.B(n_1640),
.C(n_1646),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1714),
.B(n_1639),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1713),
.B(n_1718),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1696),
.Y(n_1731)
);

HB1xp67_ASAP7_75t_L g1732 ( 
.A(n_1702),
.Y(n_1732)
);

AOI211xp5_ASAP7_75t_L g1733 ( 
.A1(n_1697),
.A2(n_1664),
.B(n_1593),
.C(n_1639),
.Y(n_1733)
);

NAND3xp33_ASAP7_75t_L g1734 ( 
.A(n_1693),
.B(n_1646),
.C(n_1655),
.Y(n_1734)
);

INVxp67_ASAP7_75t_SL g1735 ( 
.A(n_1702),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1696),
.Y(n_1736)
);

INVx3_ASAP7_75t_L g1737 ( 
.A(n_1689),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1710),
.B(n_1698),
.Y(n_1738)
);

NAND4xp75_ASAP7_75t_L g1739 ( 
.A(n_1722),
.B(n_1685),
.C(n_1703),
.D(n_1677),
.Y(n_1739)
);

INVx3_ASAP7_75t_L g1740 ( 
.A(n_1689),
.Y(n_1740)
);

A2O1A1Ixp33_ASAP7_75t_L g1741 ( 
.A1(n_1722),
.A2(n_1639),
.B(n_1664),
.C(n_1643),
.Y(n_1741)
);

AND4x1_ASAP7_75t_L g1742 ( 
.A(n_1699),
.B(n_1703),
.C(n_1688),
.D(n_1710),
.Y(n_1742)
);

NOR2x1_ASAP7_75t_L g1743 ( 
.A(n_1699),
.B(n_1681),
.Y(n_1743)
);

BUFx2_ASAP7_75t_L g1744 ( 
.A(n_1709),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1698),
.B(n_1681),
.Y(n_1745)
);

AOI22xp33_ASAP7_75t_SL g1746 ( 
.A1(n_1721),
.A2(n_1685),
.B1(n_1672),
.B2(n_1670),
.Y(n_1746)
);

AOI22xp33_ASAP7_75t_L g1747 ( 
.A1(n_1700),
.A2(n_1685),
.B1(n_1672),
.B2(n_1670),
.Y(n_1747)
);

OAI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1688),
.A2(n_1678),
.B1(n_1677),
.B2(n_1671),
.Y(n_1748)
);

INVx2_ASAP7_75t_SL g1749 ( 
.A(n_1705),
.Y(n_1749)
);

OR2x2_ASAP7_75t_L g1750 ( 
.A(n_1701),
.B(n_1650),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1713),
.B(n_1645),
.Y(n_1751)
);

AOI22xp33_ASAP7_75t_L g1752 ( 
.A1(n_1700),
.A2(n_1672),
.B1(n_1670),
.B2(n_1677),
.Y(n_1752)
);

OAI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1688),
.A2(n_1593),
.B1(n_1684),
.B2(n_1597),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1691),
.Y(n_1754)
);

OAI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1712),
.A2(n_1684),
.B1(n_1597),
.B2(n_1664),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1701),
.Y(n_1756)
);

INVxp67_ASAP7_75t_L g1757 ( 
.A(n_1706),
.Y(n_1757)
);

OAI221xp5_ASAP7_75t_L g1758 ( 
.A1(n_1706),
.A2(n_1677),
.B1(n_1655),
.B2(n_1662),
.C(n_1668),
.Y(n_1758)
);

INVx2_ASAP7_75t_SL g1759 ( 
.A(n_1705),
.Y(n_1759)
);

AOI221xp5_ASAP7_75t_L g1760 ( 
.A1(n_1695),
.A2(n_1672),
.B1(n_1653),
.B2(n_1656),
.C(n_1648),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1711),
.Y(n_1761)
);

NAND4xp25_ASAP7_75t_SL g1762 ( 
.A(n_1714),
.B(n_1588),
.C(n_1568),
.D(n_1587),
.Y(n_1762)
);

BUFx3_ASAP7_75t_L g1763 ( 
.A(n_1705),
.Y(n_1763)
);

AOI222xp33_ASAP7_75t_L g1764 ( 
.A1(n_1721),
.A2(n_1643),
.B1(n_1639),
.B2(n_1638),
.C1(n_1680),
.C2(n_1651),
.Y(n_1764)
);

OA21x2_ASAP7_75t_L g1765 ( 
.A1(n_1707),
.A2(n_1687),
.B(n_1682),
.Y(n_1765)
);

OAI211xp5_ASAP7_75t_SL g1766 ( 
.A1(n_1715),
.A2(n_1720),
.B(n_1716),
.C(n_1692),
.Y(n_1766)
);

OR2x2_ASAP7_75t_L g1767 ( 
.A(n_1701),
.B(n_1650),
.Y(n_1767)
);

NAND3xp33_ASAP7_75t_L g1768 ( 
.A(n_1711),
.B(n_1660),
.C(n_1668),
.Y(n_1768)
);

OAI31xp33_ASAP7_75t_L g1769 ( 
.A1(n_1695),
.A2(n_1639),
.A3(n_1643),
.B(n_1651),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1691),
.Y(n_1770)
);

NAND4xp25_ASAP7_75t_L g1771 ( 
.A(n_1715),
.B(n_1687),
.C(n_1673),
.D(n_1674),
.Y(n_1771)
);

OAI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1708),
.A2(n_1678),
.B1(n_1677),
.B2(n_1671),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1715),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1763),
.B(n_1583),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1727),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1731),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1738),
.B(n_1690),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1765),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1773),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1765),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1765),
.Y(n_1781)
);

OAI21x1_ASAP7_75t_L g1782 ( 
.A1(n_1752),
.A2(n_1707),
.B(n_1723),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1736),
.Y(n_1783)
);

INVx4_ASAP7_75t_SL g1784 ( 
.A(n_1763),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1756),
.B(n_1690),
.Y(n_1785)
);

AO21x1_ASAP7_75t_L g1786 ( 
.A1(n_1725),
.A2(n_1716),
.B(n_1692),
.Y(n_1786)
);

INVx4_ASAP7_75t_SL g1787 ( 
.A(n_1749),
.Y(n_1787)
);

INVx4_ASAP7_75t_SL g1788 ( 
.A(n_1759),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1750),
.Y(n_1789)
);

HB1xp67_ASAP7_75t_L g1790 ( 
.A(n_1732),
.Y(n_1790)
);

NOR2x1_ASAP7_75t_L g1791 ( 
.A(n_1762),
.B(n_1743),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1729),
.B(n_1714),
.Y(n_1792)
);

OR2x2_ASAP7_75t_L g1793 ( 
.A(n_1757),
.B(n_1690),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1745),
.B(n_1690),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1767),
.Y(n_1795)
);

INVxp67_ASAP7_75t_L g1796 ( 
.A(n_1744),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1742),
.B(n_1690),
.Y(n_1797)
);

INVx1_ASAP7_75t_SL g1798 ( 
.A(n_1726),
.Y(n_1798)
);

NAND3xp33_ASAP7_75t_L g1799 ( 
.A(n_1746),
.B(n_1668),
.C(n_1717),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1732),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1761),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1761),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1735),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1754),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1733),
.B(n_1690),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1734),
.Y(n_1806)
);

OAI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1725),
.A2(n_1739),
.B(n_1724),
.Y(n_1807)
);

INVx3_ASAP7_75t_L g1808 ( 
.A(n_1729),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1770),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1741),
.B(n_1690),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_R g1811 ( 
.A(n_1726),
.B(n_1562),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1770),
.Y(n_1812)
);

OAI21xp5_ASAP7_75t_SL g1813 ( 
.A1(n_1771),
.A2(n_1695),
.B(n_1718),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1779),
.Y(n_1814)
);

BUFx3_ASAP7_75t_L g1815 ( 
.A(n_1798),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_SL g1816 ( 
.A(n_1786),
.B(n_1741),
.Y(n_1816)
);

INVxp67_ASAP7_75t_L g1817 ( 
.A(n_1806),
.Y(n_1817)
);

BUFx2_ASAP7_75t_L g1818 ( 
.A(n_1786),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1792),
.B(n_1791),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1808),
.B(n_1730),
.Y(n_1820)
);

OAI211xp5_ASAP7_75t_SL g1821 ( 
.A1(n_1807),
.A2(n_1797),
.B(n_1813),
.C(n_1805),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1779),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1775),
.Y(n_1823)
);

INVx1_ASAP7_75t_SL g1824 ( 
.A(n_1811),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1806),
.B(n_1690),
.Y(n_1825)
);

NAND4xp25_ASAP7_75t_L g1826 ( 
.A(n_1799),
.B(n_1768),
.C(n_1747),
.D(n_1760),
.Y(n_1826)
);

NAND3xp33_ASAP7_75t_L g1827 ( 
.A(n_1810),
.B(n_1758),
.C(n_1747),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1787),
.B(n_1718),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1787),
.B(n_1751),
.Y(n_1829)
);

INVx1_ASAP7_75t_SL g1830 ( 
.A(n_1784),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1778),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1776),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_1790),
.Y(n_1833)
);

HB1xp67_ASAP7_75t_L g1834 ( 
.A(n_1800),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1783),
.Y(n_1835)
);

OAI33xp33_ASAP7_75t_L g1836 ( 
.A1(n_1810),
.A2(n_1748),
.A3(n_1772),
.B1(n_1728),
.B2(n_1766),
.B3(n_1753),
.Y(n_1836)
);

AOI21xp5_ASAP7_75t_SL g1837 ( 
.A1(n_1774),
.A2(n_1748),
.B(n_1772),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1787),
.B(n_1713),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_SL g1839 ( 
.A(n_1787),
.B(n_1769),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1794),
.B(n_1789),
.Y(n_1840)
);

INVx2_ASAP7_75t_SL g1841 ( 
.A(n_1778),
.Y(n_1841)
);

AND2x4_ASAP7_75t_L g1842 ( 
.A(n_1788),
.B(n_1700),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_SL g1843 ( 
.A(n_1788),
.B(n_1764),
.Y(n_1843)
);

INVx2_ASAP7_75t_SL g1844 ( 
.A(n_1780),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1784),
.B(n_1704),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1795),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1784),
.B(n_1694),
.Y(n_1847)
);

INVxp67_ASAP7_75t_SL g1848 ( 
.A(n_1780),
.Y(n_1848)
);

AOI211x1_ASAP7_75t_L g1849 ( 
.A1(n_1777),
.A2(n_1755),
.B(n_1719),
.C(n_1720),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1781),
.Y(n_1850)
);

INVx1_ASAP7_75t_SL g1851 ( 
.A(n_1784),
.Y(n_1851)
);

NOR3xp33_ASAP7_75t_L g1852 ( 
.A(n_1793),
.B(n_1570),
.C(n_1652),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1818),
.B(n_1801),
.Y(n_1853)
);

AOI21xp33_ASAP7_75t_L g1854 ( 
.A1(n_1818),
.A2(n_1700),
.B(n_1793),
.Y(n_1854)
);

OR2x2_ASAP7_75t_L g1855 ( 
.A(n_1817),
.B(n_1802),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1834),
.Y(n_1856)
);

OR2x6_ASAP7_75t_L g1857 ( 
.A(n_1837),
.B(n_1678),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1817),
.B(n_1816),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1815),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1819),
.B(n_1803),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1815),
.B(n_1796),
.Y(n_1861)
);

NOR2x1_ASAP7_75t_L g1862 ( 
.A(n_1815),
.B(n_1540),
.Y(n_1862)
);

O2A1O1Ixp33_ASAP7_75t_L g1863 ( 
.A1(n_1836),
.A2(n_1781),
.B(n_1785),
.C(n_1700),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1841),
.Y(n_1864)
);

OAI21xp33_ASAP7_75t_L g1865 ( 
.A1(n_1821),
.A2(n_1785),
.B(n_1782),
.Y(n_1865)
);

AOI22xp5_ASAP7_75t_L g1866 ( 
.A1(n_1836),
.A2(n_1672),
.B1(n_1677),
.B2(n_1641),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1834),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1819),
.B(n_1737),
.Y(n_1868)
);

NAND2x1p5_ASAP7_75t_L g1869 ( 
.A(n_1830),
.B(n_1851),
.Y(n_1869)
);

NOR4xp25_ASAP7_75t_L g1870 ( 
.A(n_1821),
.B(n_1812),
.C(n_1809),
.D(n_1804),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1846),
.B(n_1717),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1833),
.B(n_1720),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1845),
.B(n_1740),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1814),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1845),
.B(n_1694),
.Y(n_1875)
);

NAND2x1p5_ASAP7_75t_L g1876 ( 
.A(n_1830),
.B(n_1546),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1841),
.Y(n_1877)
);

OR2x2_ASAP7_75t_L g1878 ( 
.A(n_1846),
.B(n_1708),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1814),
.Y(n_1879)
);

OAI22xp5_ASAP7_75t_L g1880 ( 
.A1(n_1837),
.A2(n_1709),
.B1(n_1694),
.B2(n_1712),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1822),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1829),
.B(n_1847),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1833),
.B(n_1656),
.Y(n_1883)
);

HB1xp67_ASAP7_75t_L g1884 ( 
.A(n_1823),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1822),
.Y(n_1885)
);

O2A1O1Ixp33_ASAP7_75t_L g1886 ( 
.A1(n_1826),
.A2(n_1843),
.B(n_1825),
.C(n_1827),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1823),
.Y(n_1887)
);

OR2x2_ASAP7_75t_L g1888 ( 
.A(n_1858),
.B(n_1825),
.Y(n_1888)
);

AO21x2_ASAP7_75t_L g1889 ( 
.A1(n_1870),
.A2(n_1827),
.B(n_1848),
.Y(n_1889)
);

AND2x4_ASAP7_75t_L g1890 ( 
.A(n_1859),
.B(n_1851),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1858),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1878),
.B(n_1826),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1859),
.B(n_1847),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1860),
.B(n_1832),
.Y(n_1894)
);

OR2x2_ASAP7_75t_L g1895 ( 
.A(n_1878),
.B(n_1832),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1884),
.Y(n_1896)
);

NAND2x1_ASAP7_75t_SL g1897 ( 
.A(n_1862),
.B(n_1828),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1874),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1879),
.Y(n_1899)
);

AND2x4_ASAP7_75t_L g1900 ( 
.A(n_1882),
.B(n_1841),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1860),
.B(n_1835),
.Y(n_1901)
);

INVx2_ASAP7_75t_SL g1902 ( 
.A(n_1869),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1882),
.B(n_1829),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1886),
.B(n_1835),
.Y(n_1904)
);

HB1xp67_ASAP7_75t_L g1905 ( 
.A(n_1861),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1869),
.B(n_1828),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1881),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1885),
.Y(n_1908)
);

INVxp67_ASAP7_75t_L g1909 ( 
.A(n_1855),
.Y(n_1909)
);

INVx3_ASAP7_75t_L g1910 ( 
.A(n_1857),
.Y(n_1910)
);

BUFx3_ASAP7_75t_L g1911 ( 
.A(n_1856),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1857),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1853),
.Y(n_1913)
);

INVx1_ASAP7_75t_SL g1914 ( 
.A(n_1853),
.Y(n_1914)
);

NAND3xp33_ASAP7_75t_L g1915 ( 
.A(n_1904),
.B(n_1866),
.C(n_1867),
.Y(n_1915)
);

NAND3xp33_ASAP7_75t_L g1916 ( 
.A(n_1891),
.B(n_1865),
.C(n_1855),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1898),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1898),
.Y(n_1918)
);

INVxp67_ASAP7_75t_L g1919 ( 
.A(n_1902),
.Y(n_1919)
);

OAI211xp5_ASAP7_75t_SL g1920 ( 
.A1(n_1914),
.A2(n_1877),
.B(n_1864),
.C(n_1839),
.Y(n_1920)
);

AOI21xp5_ASAP7_75t_L g1921 ( 
.A1(n_1889),
.A2(n_1857),
.B(n_1880),
.Y(n_1921)
);

INVx2_ASAP7_75t_SL g1922 ( 
.A(n_1903),
.Y(n_1922)
);

AOI22xp33_ASAP7_75t_SL g1923 ( 
.A1(n_1889),
.A2(n_1857),
.B1(n_1848),
.B2(n_1844),
.Y(n_1923)
);

OR2x2_ASAP7_75t_L g1924 ( 
.A(n_1892),
.B(n_1883),
.Y(n_1924)
);

XNOR2xp5_ASAP7_75t_L g1925 ( 
.A(n_1903),
.B(n_1824),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1889),
.B(n_1864),
.Y(n_1926)
);

OAI21xp5_ASAP7_75t_SL g1927 ( 
.A1(n_1892),
.A2(n_1824),
.B(n_1868),
.Y(n_1927)
);

OAI22xp5_ASAP7_75t_L g1928 ( 
.A1(n_1914),
.A2(n_1849),
.B1(n_1838),
.B2(n_1876),
.Y(n_1928)
);

AOI21xp33_ASAP7_75t_L g1929 ( 
.A1(n_1889),
.A2(n_1877),
.B(n_1863),
.Y(n_1929)
);

AND2x4_ASAP7_75t_L g1930 ( 
.A(n_1890),
.B(n_1868),
.Y(n_1930)
);

AOI22xp5_ASAP7_75t_L g1931 ( 
.A1(n_1891),
.A2(n_1852),
.B1(n_1844),
.B2(n_1831),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1899),
.Y(n_1932)
);

AOI322xp5_ASAP7_75t_L g1933 ( 
.A1(n_1891),
.A2(n_1854),
.A3(n_1844),
.B1(n_1852),
.B2(n_1887),
.C1(n_1831),
.C2(n_1850),
.Y(n_1933)
);

INVx1_ASAP7_75t_SL g1934 ( 
.A(n_1893),
.Y(n_1934)
);

NOR2xp33_ASAP7_75t_L g1935 ( 
.A(n_1905),
.B(n_1876),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1906),
.B(n_1820),
.Y(n_1936)
);

NOR2xp33_ASAP7_75t_L g1937 ( 
.A(n_1934),
.B(n_1925),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1922),
.B(n_1890),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1930),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1936),
.B(n_1906),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1930),
.B(n_1893),
.Y(n_1941)
);

OR2x2_ASAP7_75t_L g1942 ( 
.A(n_1924),
.B(n_1894),
.Y(n_1942)
);

INVxp67_ASAP7_75t_L g1943 ( 
.A(n_1926),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1919),
.B(n_1890),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1927),
.B(n_1890),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1935),
.B(n_1900),
.Y(n_1946)
);

INVxp67_ASAP7_75t_L g1947 ( 
.A(n_1917),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1918),
.Y(n_1948)
);

NAND4xp25_ASAP7_75t_L g1949 ( 
.A(n_1937),
.B(n_1923),
.C(n_1916),
.D(n_1915),
.Y(n_1949)
);

CKINVDCx5p33_ASAP7_75t_R g1950 ( 
.A(n_1937),
.Y(n_1950)
);

NAND3xp33_ASAP7_75t_L g1951 ( 
.A(n_1945),
.B(n_1921),
.C(n_1929),
.Y(n_1951)
);

AO21x1_ASAP7_75t_L g1952 ( 
.A1(n_1944),
.A2(n_1913),
.B(n_1932),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1942),
.Y(n_1953)
);

O2A1O1Ixp33_ASAP7_75t_L g1954 ( 
.A1(n_1943),
.A2(n_1920),
.B(n_1909),
.C(n_1913),
.Y(n_1954)
);

NAND4xp25_ASAP7_75t_SL g1955 ( 
.A(n_1940),
.B(n_1931),
.C(n_1933),
.D(n_1896),
.Y(n_1955)
);

NAND3xp33_ASAP7_75t_L g1956 ( 
.A(n_1939),
.B(n_1933),
.C(n_1902),
.Y(n_1956)
);

AOI221x1_ASAP7_75t_SL g1957 ( 
.A1(n_1938),
.A2(n_1896),
.B1(n_1928),
.B2(n_1900),
.C(n_1899),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1941),
.B(n_1911),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1947),
.B(n_1911),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1959),
.Y(n_1960)
);

AOI221xp5_ASAP7_75t_L g1961 ( 
.A1(n_1955),
.A2(n_1943),
.B1(n_1947),
.B2(n_1888),
.C(n_1948),
.Y(n_1961)
);

OAI31xp33_ASAP7_75t_L g1962 ( 
.A1(n_1951),
.A2(n_1910),
.A3(n_1888),
.B(n_1912),
.Y(n_1962)
);

AOI211xp5_ASAP7_75t_L g1963 ( 
.A1(n_1949),
.A2(n_1946),
.B(n_1911),
.C(n_1900),
.Y(n_1963)
);

OAI21xp33_ASAP7_75t_L g1964 ( 
.A1(n_1950),
.A2(n_1897),
.B(n_1900),
.Y(n_1964)
);

NOR2xp33_ASAP7_75t_L g1965 ( 
.A(n_1958),
.B(n_1901),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1963),
.B(n_1953),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1965),
.B(n_1952),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1960),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1961),
.B(n_1954),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1962),
.B(n_1957),
.Y(n_1970)
);

NOR2x1p5_ASAP7_75t_L g1971 ( 
.A(n_1964),
.B(n_1956),
.Y(n_1971)
);

AOI22xp5_ASAP7_75t_SL g1972 ( 
.A1(n_1967),
.A2(n_1908),
.B1(n_1907),
.B2(n_1910),
.Y(n_1972)
);

OAI221xp5_ASAP7_75t_L g1973 ( 
.A1(n_1969),
.A2(n_1897),
.B1(n_1910),
.B2(n_1912),
.C(n_1907),
.Y(n_1973)
);

INVxp33_ASAP7_75t_L g1974 ( 
.A(n_1966),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1968),
.Y(n_1975)
);

OR2x2_ASAP7_75t_L g1976 ( 
.A(n_1969),
.B(n_1895),
.Y(n_1976)
);

OR2x6_ASAP7_75t_L g1977 ( 
.A(n_1975),
.B(n_1971),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1976),
.Y(n_1978)
);

INVxp67_ASAP7_75t_L g1979 ( 
.A(n_1972),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1978),
.Y(n_1980)
);

OAI322xp33_ASAP7_75t_L g1981 ( 
.A1(n_1980),
.A2(n_1970),
.A3(n_1979),
.B1(n_1973),
.B2(n_1974),
.C1(n_1977),
.C2(n_1908),
.Y(n_1981)
);

A2O1A1Ixp33_ASAP7_75t_L g1982 ( 
.A1(n_1981),
.A2(n_1910),
.B(n_1912),
.C(n_1895),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1981),
.Y(n_1983)
);

INVxp67_ASAP7_75t_L g1984 ( 
.A(n_1983),
.Y(n_1984)
);

AOI22xp5_ASAP7_75t_L g1985 ( 
.A1(n_1982),
.A2(n_1831),
.B1(n_1850),
.B2(n_1842),
.Y(n_1985)
);

HB1xp67_ASAP7_75t_L g1986 ( 
.A(n_1984),
.Y(n_1986)
);

OAI22xp33_ASAP7_75t_SL g1987 ( 
.A1(n_1985),
.A2(n_1850),
.B1(n_1871),
.B2(n_1872),
.Y(n_1987)
);

AOI221xp5_ASAP7_75t_L g1988 ( 
.A1(n_1986),
.A2(n_1849),
.B1(n_1842),
.B2(n_1871),
.C(n_1840),
.Y(n_1988)
);

AOI21x1_ASAP7_75t_L g1989 ( 
.A1(n_1988),
.A2(n_1987),
.B(n_1873),
.Y(n_1989)
);

NAND2x1p5_ASAP7_75t_L g1990 ( 
.A(n_1989),
.B(n_1546),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1990),
.B(n_1842),
.Y(n_1991)
);

OA22x2_ASAP7_75t_L g1992 ( 
.A1(n_1991),
.A2(n_1842),
.B1(n_1602),
.B2(n_1873),
.Y(n_1992)
);

AOI211xp5_ASAP7_75t_L g1993 ( 
.A1(n_1992),
.A2(n_1546),
.B(n_1840),
.C(n_1875),
.Y(n_1993)
);


endmodule