module real_aes_6441_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_527;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g111 ( .A(n_0), .Y(n_111) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_1), .A2(n_162), .B(n_165), .C(n_245), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_2), .A2(n_191), .B(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g492 ( .A(n_3), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_4), .B(n_221), .Y(n_220) );
AOI21xp33_ASAP7_75t_L g475 ( .A1(n_5), .A2(n_191), .B(n_476), .Y(n_475) );
AND2x6_ASAP7_75t_L g162 ( .A(n_6), .B(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g258 ( .A(n_7), .Y(n_258) );
INVx1_ASAP7_75t_L g109 ( .A(n_8), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_8), .B(n_41), .Y(n_127) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_9), .A2(n_190), .B(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_10), .B(n_174), .Y(n_247) );
INVx1_ASAP7_75t_L g480 ( .A(n_11), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_12), .B(n_215), .Y(n_515) );
INVx1_ASAP7_75t_L g154 ( .A(n_13), .Y(n_154) );
INVx1_ASAP7_75t_L g527 ( .A(n_14), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g134 ( .A1(n_15), .A2(n_78), .B1(n_135), .B2(n_136), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_15), .Y(n_135) );
A2O1A1Ixp33_ASAP7_75t_L g279 ( .A1(n_16), .A2(n_199), .B(n_280), .C(n_282), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_17), .B(n_221), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_18), .B(n_458), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_19), .B(n_191), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_20), .B(n_205), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g265 ( .A1(n_21), .A2(n_215), .B(n_266), .C(n_268), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_22), .B(n_221), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_23), .B(n_174), .Y(n_173) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_24), .A2(n_201), .B(n_282), .C(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_25), .B(n_174), .Y(n_229) );
CKINVDCx16_ASAP7_75t_R g156 ( .A(n_26), .Y(n_156) );
INVx1_ASAP7_75t_L g228 ( .A(n_27), .Y(n_228) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_28), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g243 ( .A(n_29), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_30), .B(n_174), .Y(n_493) );
INVx1_ASAP7_75t_L g197 ( .A(n_31), .Y(n_197) );
INVx1_ASAP7_75t_L g470 ( .A(n_32), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g131 ( .A1(n_33), .A2(n_132), .B1(n_133), .B2(n_134), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_33), .Y(n_132) );
INVx2_ASAP7_75t_L g160 ( .A(n_34), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_35), .Y(n_249) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_36), .A2(n_215), .B(n_216), .C(n_218), .Y(n_214) );
INVxp67_ASAP7_75t_L g200 ( .A(n_37), .Y(n_200) );
CKINVDCx14_ASAP7_75t_R g213 ( .A(n_38), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g226 ( .A1(n_39), .A2(n_165), .B(n_227), .C(n_231), .Y(n_226) );
A2O1A1Ixp33_ASAP7_75t_L g502 ( .A1(n_40), .A2(n_162), .B(n_165), .C(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_41), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g469 ( .A(n_42), .Y(n_469) );
A2O1A1Ixp33_ASAP7_75t_L g255 ( .A1(n_43), .A2(n_176), .B(n_256), .C(n_257), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_44), .B(n_174), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_45), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g193 ( .A(n_46), .Y(n_193) );
INVx1_ASAP7_75t_L g264 ( .A(n_47), .Y(n_264) );
CKINVDCx16_ASAP7_75t_R g471 ( .A(n_48), .Y(n_471) );
OAI22xp5_ASAP7_75t_SL g740 ( .A1(n_49), .A2(n_58), .B1(n_741), .B2(n_742), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_49), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_50), .B(n_191), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_51), .A2(n_165), .B1(n_268), .B2(n_468), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_52), .Y(n_507) );
CKINVDCx16_ASAP7_75t_R g489 ( .A(n_53), .Y(n_489) );
CKINVDCx14_ASAP7_75t_R g254 ( .A(n_54), .Y(n_254) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_55), .A2(n_218), .B(n_256), .C(n_479), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_56), .Y(n_539) );
INVx1_ASAP7_75t_L g477 ( .A(n_57), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_58), .Y(n_742) );
INVx1_ASAP7_75t_L g163 ( .A(n_59), .Y(n_163) );
INVx1_ASAP7_75t_L g153 ( .A(n_60), .Y(n_153) );
INVx1_ASAP7_75t_SL g217 ( .A(n_61), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_62), .Y(n_121) );
OAI22xp5_ASAP7_75t_SL g739 ( .A1(n_63), .A2(n_740), .B1(n_743), .B2(n_744), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_63), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_64), .B(n_221), .Y(n_270) );
INVx1_ASAP7_75t_L g169 ( .A(n_65), .Y(n_169) );
AOI222xp33_ASAP7_75t_SL g129 ( .A1(n_66), .A2(n_130), .B1(n_131), .B2(n_137), .C1(n_731), .C2(n_733), .Y(n_129) );
A2O1A1Ixp33_ASAP7_75t_SL g457 ( .A1(n_67), .A2(n_218), .B(n_458), .C(n_459), .Y(n_457) );
INVxp67_ASAP7_75t_L g460 ( .A(n_68), .Y(n_460) );
INVx1_ASAP7_75t_L g114 ( .A(n_69), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_70), .A2(n_191), .B(n_253), .Y(n_252) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_71), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_72), .A2(n_191), .B(n_277), .Y(n_276) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_73), .Y(n_473) );
INVx1_ASAP7_75t_L g533 ( .A(n_74), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_75), .A2(n_190), .B(n_192), .Y(n_189) );
CKINVDCx16_ASAP7_75t_R g225 ( .A(n_76), .Y(n_225) );
INVx1_ASAP7_75t_L g278 ( .A(n_77), .Y(n_278) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_78), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_79), .A2(n_162), .B(n_165), .C(n_535), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_80), .A2(n_191), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g281 ( .A(n_81), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_82), .B(n_198), .Y(n_504) );
INVx2_ASAP7_75t_L g151 ( .A(n_83), .Y(n_151) );
INVx1_ASAP7_75t_L g246 ( .A(n_84), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_85), .B(n_458), .Y(n_505) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_86), .A2(n_162), .B(n_165), .C(n_491), .Y(n_490) );
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_87), .B(n_111), .C(n_112), .Y(n_110) );
OR2x2_ASAP7_75t_L g124 ( .A(n_87), .B(n_125), .Y(n_124) );
OR2x2_ASAP7_75t_L g444 ( .A(n_87), .B(n_126), .Y(n_444) );
INVx2_ASAP7_75t_L g730 ( .A(n_87), .Y(n_730) );
A2O1A1Ixp33_ASAP7_75t_L g164 ( .A1(n_88), .A2(n_165), .B(n_168), .C(n_178), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_89), .B(n_183), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_90), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_91), .A2(n_104), .B1(n_115), .B2(n_746), .Y(n_103) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_92), .A2(n_162), .B(n_165), .C(n_513), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_93), .Y(n_519) );
INVx1_ASAP7_75t_L g456 ( .A(n_94), .Y(n_456) );
CKINVDCx16_ASAP7_75t_R g524 ( .A(n_95), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_96), .B(n_198), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_97), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_98), .B(n_149), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_99), .B(n_149), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_100), .B(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g267 ( .A(n_101), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_102), .A2(n_191), .B(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx5_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
CKINVDCx9p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
BUFx2_ASAP7_75t_L g746 ( .A(n_107), .Y(n_746) );
OR2x4_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
AND2x2_ASAP7_75t_L g126 ( .A(n_111), .B(n_127), .Y(n_126) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AOI22xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_129), .B1(n_736), .B2(n_737), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_118), .B(n_122), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_SL g736 ( .A(n_120), .Y(n_736) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AOI21xp5_ASAP7_75t_L g737 ( .A1(n_122), .A2(n_738), .B(n_745), .Y(n_737) );
NOR2xp33_ASAP7_75t_SL g122 ( .A(n_123), .B(n_128), .Y(n_122) );
HB1xp67_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_124), .Y(n_745) );
NOR2x2_ASAP7_75t_L g735 ( .A(n_125), .B(n_730), .Y(n_735) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OR2x2_ASAP7_75t_L g729 ( .A(n_126), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OAI22xp5_ASAP7_75t_SL g137 ( .A1(n_138), .A2(n_444), .B1(n_445), .B2(n_727), .Y(n_137) );
INVx2_ASAP7_75t_L g732 ( .A(n_138), .Y(n_732) );
XOR2xp5_ASAP7_75t_L g738 ( .A(n_138), .B(n_739), .Y(n_738) );
OR2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_378), .Y(n_138) );
NAND5xp2_ASAP7_75t_L g139 ( .A(n_140), .B(n_307), .C(n_337), .D(n_358), .E(n_364), .Y(n_139) );
AOI221xp5_ASAP7_75t_SL g140 ( .A1(n_141), .A2(n_237), .B1(n_271), .B2(n_273), .C(n_284), .Y(n_140) );
INVxp67_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g142 ( .A(n_143), .B(n_234), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_144), .B(n_206), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
A2O1A1Ixp33_ASAP7_75t_SL g358 ( .A1(n_145), .A2(n_222), .B(n_359), .C(n_362), .Y(n_358) );
AND2x2_ASAP7_75t_L g428 ( .A(n_145), .B(n_223), .Y(n_428) );
AND2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_184), .Y(n_145) );
AND2x2_ASAP7_75t_L g286 ( .A(n_146), .B(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g290 ( .A(n_146), .B(n_287), .Y(n_290) );
OR2x2_ASAP7_75t_L g316 ( .A(n_146), .B(n_223), .Y(n_316) );
AND2x2_ASAP7_75t_L g318 ( .A(n_146), .B(n_209), .Y(n_318) );
AND2x2_ASAP7_75t_L g336 ( .A(n_146), .B(n_208), .Y(n_336) );
INVx1_ASAP7_75t_L g369 ( .A(n_146), .Y(n_369) );
INVx2_ASAP7_75t_SL g146 ( .A(n_147), .Y(n_146) );
BUFx2_ASAP7_75t_L g236 ( .A(n_147), .Y(n_236) );
AND2x2_ASAP7_75t_L g272 ( .A(n_147), .B(n_209), .Y(n_272) );
AND2x2_ASAP7_75t_L g425 ( .A(n_147), .B(n_223), .Y(n_425) );
AO21x2_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_155), .B(n_180), .Y(n_147) );
INVx3_ASAP7_75t_L g221 ( .A(n_148), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_148), .B(n_233), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_148), .B(n_249), .Y(n_248) );
NOR2xp33_ASAP7_75t_SL g506 ( .A(n_148), .B(n_507), .Y(n_506) );
INVx4_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
HB1xp67_ASAP7_75t_L g210 ( .A(n_149), .Y(n_210) );
OA21x2_ASAP7_75t_L g453 ( .A1(n_149), .A2(n_454), .B(n_461), .Y(n_453) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g187 ( .A(n_150), .Y(n_187) );
AND2x2_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
AND2x2_ASAP7_75t_SL g183 ( .A(n_151), .B(n_152), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
OAI21xp5_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_157), .B(n_164), .Y(n_155) );
O2A1O1Ixp33_ASAP7_75t_L g224 ( .A1(n_157), .A2(n_183), .B(n_225), .C(n_226), .Y(n_224) );
OAI21xp5_ASAP7_75t_L g242 ( .A1(n_157), .A2(n_243), .B(n_244), .Y(n_242) );
OAI22xp33_ASAP7_75t_L g466 ( .A1(n_157), .A2(n_179), .B1(n_467), .B2(n_471), .Y(n_466) );
OAI21xp5_ASAP7_75t_L g488 ( .A1(n_157), .A2(n_489), .B(n_490), .Y(n_488) );
OAI21xp5_ASAP7_75t_L g532 ( .A1(n_157), .A2(n_533), .B(n_534), .Y(n_532) );
NAND2x1p5_ASAP7_75t_L g157 ( .A(n_158), .B(n_162), .Y(n_157) );
AND2x4_ASAP7_75t_L g191 ( .A(n_158), .B(n_162), .Y(n_191) );
AND2x2_ASAP7_75t_L g158 ( .A(n_159), .B(n_161), .Y(n_158) );
INVx1_ASAP7_75t_L g202 ( .A(n_159), .Y(n_202) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g166 ( .A(n_160), .Y(n_166) );
INVx1_ASAP7_75t_L g269 ( .A(n_160), .Y(n_269) );
INVx1_ASAP7_75t_L g167 ( .A(n_161), .Y(n_167) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_161), .Y(n_172) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_161), .Y(n_174) );
INVx3_ASAP7_75t_L g199 ( .A(n_161), .Y(n_199) );
INVx1_ASAP7_75t_L g458 ( .A(n_161), .Y(n_458) );
INVx4_ASAP7_75t_SL g179 ( .A(n_162), .Y(n_179) );
BUFx3_ASAP7_75t_L g231 ( .A(n_162), .Y(n_231) );
INVx5_ASAP7_75t_L g194 ( .A(n_165), .Y(n_194) );
AND2x6_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
BUFx3_ASAP7_75t_L g177 ( .A(n_166), .Y(n_177) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_166), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B(n_173), .C(n_175), .Y(n_168) );
O2A1O1Ixp5_ASAP7_75t_L g245 ( .A1(n_170), .A2(n_175), .B(n_246), .C(n_247), .Y(n_245) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
OAI22xp5_ASAP7_75t_SL g468 ( .A1(n_171), .A2(n_172), .B1(n_469), .B2(n_470), .Y(n_468) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx4_ASAP7_75t_L g201 ( .A(n_172), .Y(n_201) );
INVx4_ASAP7_75t_L g215 ( .A(n_174), .Y(n_215) );
INVx2_ASAP7_75t_L g256 ( .A(n_174), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_175), .A2(n_504), .B(n_505), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_175), .A2(n_536), .B(n_537), .Y(n_535) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g282 ( .A(n_177), .Y(n_282) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
O2A1O1Ixp33_ASAP7_75t_SL g192 ( .A1(n_179), .A2(n_193), .B(n_194), .C(n_195), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g212 ( .A1(n_179), .A2(n_194), .B(n_213), .C(n_214), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_SL g253 ( .A1(n_179), .A2(n_194), .B(n_254), .C(n_255), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_SL g263 ( .A1(n_179), .A2(n_194), .B(n_264), .C(n_265), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_SL g277 ( .A1(n_179), .A2(n_194), .B(n_278), .C(n_279), .Y(n_277) );
O2A1O1Ixp33_ASAP7_75t_L g455 ( .A1(n_179), .A2(n_194), .B(n_456), .C(n_457), .Y(n_455) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_179), .A2(n_194), .B(n_477), .C(n_478), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g523 ( .A1(n_179), .A2(n_194), .B(n_524), .C(n_525), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
INVx1_ASAP7_75t_L g205 ( .A(n_182), .Y(n_205) );
AO21x2_ASAP7_75t_L g510 ( .A1(n_182), .A2(n_511), .B(n_518), .Y(n_510) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g241 ( .A(n_183), .Y(n_241) );
OA21x2_ASAP7_75t_L g251 ( .A1(n_183), .A2(n_252), .B(n_259), .Y(n_251) );
OA21x2_ASAP7_75t_L g521 ( .A1(n_183), .A2(n_522), .B(n_528), .Y(n_521) );
AND2x2_ASAP7_75t_L g306 ( .A(n_184), .B(n_207), .Y(n_306) );
OR2x2_ASAP7_75t_L g310 ( .A(n_184), .B(n_223), .Y(n_310) );
AND2x2_ASAP7_75t_L g335 ( .A(n_184), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_SL g382 ( .A(n_184), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_184), .B(n_344), .Y(n_430) );
AO21x2_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_188), .B(n_203), .Y(n_184) );
INVx1_ASAP7_75t_L g288 ( .A(n_185), .Y(n_288) );
AO21x2_ASAP7_75t_L g531 ( .A1(n_185), .A2(n_532), .B(n_538), .Y(n_531) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AOI21xp5_ASAP7_75t_SL g500 ( .A1(n_186), .A2(n_501), .B(n_502), .Y(n_500) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AO21x2_ASAP7_75t_L g465 ( .A1(n_187), .A2(n_466), .B(n_472), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_187), .B(n_473), .Y(n_472) );
AO21x2_ASAP7_75t_L g487 ( .A1(n_187), .A2(n_488), .B(n_495), .Y(n_487) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
OA21x2_ASAP7_75t_L g287 ( .A1(n_189), .A2(n_204), .B(n_288), .Y(n_287) );
BUFx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_196), .B(n_202), .Y(n_195) );
OAI22xp33_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B1(n_200), .B2(n_201), .Y(n_196) );
O2A1O1Ixp33_ASAP7_75t_L g227 ( .A1(n_198), .A2(n_228), .B(n_229), .C(n_230), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_198), .A2(n_492), .B(n_493), .C(n_494), .Y(n_491) );
INVx5_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_199), .B(n_258), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_199), .B(n_460), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_199), .B(n_480), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_201), .B(n_267), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_201), .B(n_281), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_201), .B(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g230 ( .A(n_202), .Y(n_230) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
OAI322xp33_ASAP7_75t_L g431 ( .A1(n_206), .A2(n_367), .A3(n_390), .B1(n_411), .B2(n_432), .C1(n_434), .C2(n_435), .Y(n_431) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_207), .B(n_287), .Y(n_434) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_222), .Y(n_207) );
AND2x2_ASAP7_75t_L g235 ( .A(n_208), .B(n_236), .Y(n_235) );
AND2x4_ASAP7_75t_L g303 ( .A(n_208), .B(n_223), .Y(n_303) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g344 ( .A(n_209), .B(n_223), .Y(n_344) );
AND2x2_ASAP7_75t_L g388 ( .A(n_209), .B(n_222), .Y(n_388) );
OA21x2_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_220), .Y(n_209) );
OA21x2_ASAP7_75t_L g261 ( .A1(n_210), .A2(n_262), .B(n_270), .Y(n_261) );
OA21x2_ASAP7_75t_L g275 ( .A1(n_210), .A2(n_276), .B(n_283), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_215), .B(n_217), .Y(n_216) );
INVx3_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_219), .Y(n_516) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_221), .A2(n_475), .B(n_481), .Y(n_474) );
AND2x2_ASAP7_75t_L g271 ( .A(n_222), .B(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g289 ( .A(n_222), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_222), .B(n_318), .Y(n_442) );
INVx3_ASAP7_75t_SL g222 ( .A(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g234 ( .A(n_223), .B(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_223), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g356 ( .A(n_223), .B(n_287), .Y(n_356) );
AND2x2_ASAP7_75t_L g383 ( .A(n_223), .B(n_318), .Y(n_383) );
OR2x2_ASAP7_75t_L g439 ( .A(n_223), .B(n_290), .Y(n_439) );
OR2x6_ASAP7_75t_L g223 ( .A(n_224), .B(n_232), .Y(n_223) );
INVx1_ASAP7_75t_SL g325 ( .A(n_234), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_235), .B(n_356), .Y(n_357) );
AND2x2_ASAP7_75t_L g391 ( .A(n_235), .B(n_381), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_235), .B(n_314), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_235), .B(n_436), .Y(n_435) );
OAI31xp33_ASAP7_75t_L g409 ( .A1(n_237), .A2(n_271), .A3(n_410), .B(n_412), .Y(n_409) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_250), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g376 ( .A(n_238), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g392 ( .A(n_238), .B(n_327), .Y(n_392) );
OR2x2_ASAP7_75t_L g399 ( .A(n_238), .B(n_400), .Y(n_399) );
OR2x2_ASAP7_75t_L g411 ( .A(n_238), .B(n_300), .Y(n_411) );
CKINVDCx16_ASAP7_75t_R g238 ( .A(n_239), .Y(n_238) );
OR2x2_ASAP7_75t_L g345 ( .A(n_239), .B(n_346), .Y(n_345) );
BUFx3_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g273 ( .A(n_240), .B(n_274), .Y(n_273) );
INVx4_ASAP7_75t_L g294 ( .A(n_240), .Y(n_294) );
AND2x2_ASAP7_75t_L g331 ( .A(n_240), .B(n_275), .Y(n_331) );
AO21x2_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_242), .B(n_248), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_241), .B(n_496), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_241), .B(n_519), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_241), .B(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g330 ( .A(n_250), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_SL g400 ( .A(n_250), .Y(n_400) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_260), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_251), .B(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g300 ( .A(n_251), .B(n_261), .Y(n_300) );
INVx2_ASAP7_75t_L g320 ( .A(n_251), .Y(n_320) );
AND2x2_ASAP7_75t_L g334 ( .A(n_251), .B(n_261), .Y(n_334) );
AND2x2_ASAP7_75t_L g341 ( .A(n_251), .B(n_297), .Y(n_341) );
BUFx3_ASAP7_75t_L g351 ( .A(n_251), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_251), .B(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g296 ( .A(n_260), .Y(n_296) );
AND2x2_ASAP7_75t_L g304 ( .A(n_260), .B(n_294), .Y(n_304) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g274 ( .A(n_261), .B(n_275), .Y(n_274) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_261), .Y(n_328) );
INVx2_ASAP7_75t_L g494 ( .A(n_268), .Y(n_494) );
INVx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx2_ASAP7_75t_SL g311 ( .A(n_272), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_272), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_272), .B(n_381), .Y(n_402) );
NAND2xp5_ASAP7_75t_SL g404 ( .A(n_273), .B(n_351), .Y(n_404) );
INVx1_ASAP7_75t_SL g438 ( .A(n_273), .Y(n_438) );
INVx1_ASAP7_75t_SL g346 ( .A(n_274), .Y(n_346) );
INVx1_ASAP7_75t_SL g297 ( .A(n_275), .Y(n_297) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_275), .Y(n_308) );
OR2x2_ASAP7_75t_L g319 ( .A(n_275), .B(n_294), .Y(n_319) );
AND2x2_ASAP7_75t_L g333 ( .A(n_275), .B(n_294), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_275), .B(n_323), .Y(n_385) );
A2O1A1Ixp33_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_289), .B(n_291), .C(n_302), .Y(n_284) );
AOI31xp33_ASAP7_75t_L g401 ( .A1(n_285), .A2(n_402), .A3(n_403), .B(n_404), .Y(n_401) );
AND2x2_ASAP7_75t_L g374 ( .A(n_286), .B(n_303), .Y(n_374) );
BUFx3_ASAP7_75t_L g314 ( .A(n_287), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_287), .B(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g350 ( .A(n_287), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_287), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_SL g305 ( .A(n_290), .Y(n_305) );
OAI222xp33_ASAP7_75t_L g414 ( .A1(n_290), .A2(n_415), .B1(n_418), .B2(n_419), .C1(n_420), .C2(n_421), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_292), .B(n_298), .Y(n_291) );
INVx1_ASAP7_75t_L g420 ( .A(n_292), .Y(n_420) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_294), .B(n_297), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_294), .B(n_320), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_294), .B(n_295), .Y(n_390) );
INVx1_ASAP7_75t_L g441 ( .A(n_294), .Y(n_441) );
NAND2xp5_ASAP7_75t_SL g371 ( .A(n_295), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g443 ( .A(n_295), .Y(n_443) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
INVx2_ASAP7_75t_L g323 ( .A(n_296), .Y(n_323) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_297), .Y(n_366) );
AOI32xp33_ASAP7_75t_L g302 ( .A1(n_298), .A2(n_303), .A3(n_304), .B1(n_305), .B2(n_306), .Y(n_302) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_300), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g377 ( .A(n_300), .Y(n_377) );
OR2x2_ASAP7_75t_L g418 ( .A(n_300), .B(n_319), .Y(n_418) );
INVx1_ASAP7_75t_L g354 ( .A(n_301), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_303), .B(n_314), .Y(n_339) );
INVx3_ASAP7_75t_L g348 ( .A(n_303), .Y(n_348) );
AOI322xp5_ASAP7_75t_L g364 ( .A1(n_303), .A2(n_348), .A3(n_365), .B1(n_367), .B2(n_370), .C1(n_374), .C2(n_375), .Y(n_364) );
AND2x2_ASAP7_75t_L g340 ( .A(n_304), .B(n_341), .Y(n_340) );
INVxp67_ASAP7_75t_L g417 ( .A(n_304), .Y(n_417) );
A2O1A1O1Ixp25_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_309), .B(n_312), .C(n_320), .D(n_321), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_308), .B(n_351), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
OAI221xp5_ASAP7_75t_L g321 ( .A1(n_310), .A2(n_322), .B1(n_325), .B2(n_326), .C(n_329), .Y(n_321) );
INVx1_ASAP7_75t_SL g436 ( .A(n_310), .Y(n_436) );
AOI21xp33_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_317), .B(n_319), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
NAND2xp5_ASAP7_75t_SL g424 ( .A(n_314), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OAI221xp5_ASAP7_75t_SL g406 ( .A1(n_316), .A2(n_400), .B1(n_407), .B2(n_408), .C(n_409), .Y(n_406) );
OAI222xp33_ASAP7_75t_L g437 ( .A1(n_317), .A2(n_438), .B1(n_439), .B2(n_440), .C1(n_442), .C2(n_443), .Y(n_437) );
AND2x2_ASAP7_75t_L g395 ( .A(n_318), .B(n_381), .Y(n_395) );
AOI21xp5_ASAP7_75t_L g407 ( .A1(n_318), .A2(n_333), .B(n_380), .Y(n_407) );
INVx1_ASAP7_75t_L g421 ( .A(n_318), .Y(n_421) );
INVx2_ASAP7_75t_SL g324 ( .A(n_319), .Y(n_324) );
AND2x2_ASAP7_75t_L g327 ( .A(n_320), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx1_ASAP7_75t_SL g361 ( .A(n_323), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_323), .B(n_333), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_324), .B(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_324), .B(n_334), .Y(n_363) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OAI21xp5_ASAP7_75t_SL g329 ( .A1(n_330), .A2(n_332), .B(n_335), .Y(n_329) );
INVx1_ASAP7_75t_SL g347 ( .A(n_331), .Y(n_347) );
AND2x2_ASAP7_75t_L g394 ( .A(n_331), .B(n_377), .Y(n_394) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
AND2x2_ASAP7_75t_L g433 ( .A(n_333), .B(n_351), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_334), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_SL g419 ( .A(n_335), .Y(n_419) );
AOI221xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_340), .B1(n_342), .B2(n_349), .C(n_352), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OAI22xp5_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_345), .B1(n_347), .B2(n_348), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
OAI22xp33_ASAP7_75t_L g352 ( .A1(n_346), .A2(n_353), .B1(n_355), .B2(n_357), .Y(n_352) );
OR2x2_ASAP7_75t_L g423 ( .A(n_347), .B(n_351), .Y(n_423) );
OR2x2_ASAP7_75t_L g426 ( .A(n_347), .B(n_361), .Y(n_426) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OAI221xp5_ASAP7_75t_L g422 ( .A1(n_368), .A2(n_423), .B1(n_424), .B2(n_426), .C(n_427), .Y(n_422) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVxp67_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND3xp33_ASAP7_75t_SL g378 ( .A(n_379), .B(n_393), .C(n_405), .Y(n_378) );
AOI222xp33_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_384), .B1(n_386), .B2(n_389), .C1(n_391), .C2(n_392), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_381), .B(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g403 ( .A(n_383), .Y(n_403) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVxp67_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AOI221xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_395), .B1(n_396), .B2(n_398), .C(n_401), .Y(n_393) );
INVx1_ASAP7_75t_L g408 ( .A(n_394), .Y(n_408) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OAI21xp33_ASAP7_75t_L g427 ( .A1(n_398), .A2(n_428), .B(n_429), .Y(n_427) );
INVx1_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
NOR5xp2_ASAP7_75t_L g405 ( .A(n_406), .B(n_414), .C(n_422), .D(n_431), .E(n_437), .Y(n_405) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
OR2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
INVxp67_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OAI22xp5_ASAP7_75t_SL g731 ( .A1(n_444), .A2(n_446), .B1(n_727), .B2(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_SL g446 ( .A(n_447), .B(n_664), .Y(n_446) );
NOR4xp25_ASAP7_75t_L g447 ( .A(n_448), .B(n_594), .C(n_625), .D(n_644), .Y(n_447) );
NAND4xp25_ASAP7_75t_L g448 ( .A(n_449), .B(n_552), .C(n_567), .D(n_585), .Y(n_448) );
AOI222xp33_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_497), .B1(n_529), .B2(n_540), .C1(n_545), .C2(n_547), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_482), .Y(n_450) );
INVx1_ASAP7_75t_L g608 ( .A(n_451), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_462), .Y(n_451) );
AND2x2_ASAP7_75t_L g483 ( .A(n_452), .B(n_474), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_452), .B(n_486), .Y(n_637) );
INVx3_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
OR2x2_ASAP7_75t_L g544 ( .A(n_453), .B(n_464), .Y(n_544) );
AND2x2_ASAP7_75t_L g553 ( .A(n_453), .B(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g579 ( .A(n_453), .Y(n_579) );
AND2x2_ASAP7_75t_L g600 ( .A(n_453), .B(n_464), .Y(n_600) );
BUFx2_ASAP7_75t_L g623 ( .A(n_453), .Y(n_623) );
AND2x2_ASAP7_75t_L g647 ( .A(n_453), .B(n_465), .Y(n_647) );
AND2x2_ASAP7_75t_L g711 ( .A(n_453), .B(n_474), .Y(n_711) );
AND2x2_ASAP7_75t_L g612 ( .A(n_462), .B(n_543), .Y(n_612) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_463), .B(n_637), .Y(n_636) );
OR2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_474), .Y(n_463) );
OR2x2_ASAP7_75t_L g572 ( .A(n_464), .B(n_487), .Y(n_572) );
AND2x2_ASAP7_75t_L g584 ( .A(n_464), .B(n_543), .Y(n_584) );
BUFx2_ASAP7_75t_L g716 ( .A(n_464), .Y(n_716) );
INVx3_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
OR2x2_ASAP7_75t_L g485 ( .A(n_465), .B(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g566 ( .A(n_465), .B(n_487), .Y(n_566) );
AND2x2_ASAP7_75t_L g619 ( .A(n_465), .B(n_474), .Y(n_619) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_465), .Y(n_655) );
AND2x2_ASAP7_75t_L g542 ( .A(n_474), .B(n_543), .Y(n_542) );
INVx1_ASAP7_75t_SL g554 ( .A(n_474), .Y(n_554) );
INVx2_ASAP7_75t_L g565 ( .A(n_474), .Y(n_565) );
BUFx2_ASAP7_75t_L g589 ( .A(n_474), .Y(n_589) );
AND2x2_ASAP7_75t_SL g646 ( .A(n_474), .B(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_484), .Y(n_482) );
AOI332xp33_ASAP7_75t_L g567 ( .A1(n_483), .A2(n_568), .A3(n_572), .B1(n_573), .B2(n_577), .B3(n_580), .C1(n_581), .C2(n_583), .Y(n_567) );
NAND2x1_ASAP7_75t_L g652 ( .A(n_483), .B(n_543), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_483), .B(n_557), .Y(n_703) );
A2O1A1Ixp33_ASAP7_75t_SL g585 ( .A1(n_484), .A2(n_586), .B(n_589), .C(n_590), .Y(n_585) );
AND2x2_ASAP7_75t_L g724 ( .A(n_484), .B(n_565), .Y(n_724) );
INVx3_ASAP7_75t_SL g484 ( .A(n_485), .Y(n_484) );
OR2x2_ASAP7_75t_L g621 ( .A(n_485), .B(n_622), .Y(n_621) );
OR2x2_ASAP7_75t_L g626 ( .A(n_485), .B(n_623), .Y(n_626) );
INVx1_ASAP7_75t_L g557 ( .A(n_486), .Y(n_557) );
AND2x2_ASAP7_75t_L g660 ( .A(n_486), .B(n_619), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_486), .B(n_600), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_486), .B(n_671), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_486), .B(n_578), .Y(n_686) );
INVx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx3_ASAP7_75t_L g543 ( .A(n_487), .Y(n_543) );
OAI31xp33_ASAP7_75t_L g725 ( .A1(n_497), .A2(n_646), .A3(n_653), .B(n_726), .Y(n_725) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_508), .Y(n_497) );
AND2x2_ASAP7_75t_L g529 ( .A(n_498), .B(n_530), .Y(n_529) );
NAND2x1_ASAP7_75t_SL g548 ( .A(n_498), .B(n_549), .Y(n_548) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_498), .Y(n_635) );
AND2x2_ASAP7_75t_L g640 ( .A(n_498), .B(n_551), .Y(n_640) );
INVx3_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g552 ( .A1(n_499), .A2(n_553), .B(n_555), .C(n_558), .Y(n_552) );
OR2x2_ASAP7_75t_L g569 ( .A(n_499), .B(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g582 ( .A(n_499), .Y(n_582) );
AND2x2_ASAP7_75t_L g588 ( .A(n_499), .B(n_531), .Y(n_588) );
INVx2_ASAP7_75t_L g606 ( .A(n_499), .Y(n_606) );
AND2x2_ASAP7_75t_L g617 ( .A(n_499), .B(n_571), .Y(n_617) );
AND2x2_ASAP7_75t_L g649 ( .A(n_499), .B(n_607), .Y(n_649) );
AND2x2_ASAP7_75t_L g653 ( .A(n_499), .B(n_576), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_499), .B(n_508), .Y(n_658) );
AND2x2_ASAP7_75t_L g692 ( .A(n_499), .B(n_693), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_499), .B(n_595), .Y(n_726) );
OR2x6_ASAP7_75t_L g499 ( .A(n_500), .B(n_506), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_508), .B(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g634 ( .A(n_508), .Y(n_634) );
AND2x2_ASAP7_75t_L g696 ( .A(n_508), .B(n_617), .Y(n_696) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_520), .Y(n_508) );
OR2x2_ASAP7_75t_L g550 ( .A(n_509), .B(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g560 ( .A(n_509), .B(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_509), .B(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g668 ( .A(n_509), .Y(n_668) );
AND2x2_ASAP7_75t_L g685 ( .A(n_509), .B(n_531), .Y(n_685) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g576 ( .A(n_510), .B(n_520), .Y(n_576) );
AND2x2_ASAP7_75t_L g605 ( .A(n_510), .B(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g616 ( .A(n_510), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_510), .B(n_571), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_512), .B(n_517), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B(n_516), .Y(n_513) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g530 ( .A(n_521), .B(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g551 ( .A(n_521), .Y(n_551) );
AND2x2_ASAP7_75t_L g607 ( .A(n_521), .B(n_571), .Y(n_607) );
INVx1_ASAP7_75t_L g709 ( .A(n_529), .Y(n_709) );
INVx1_ASAP7_75t_L g713 ( .A(n_530), .Y(n_713) );
INVx2_ASAP7_75t_L g571 ( .A(n_531), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_541), .B(n_544), .Y(n_540) );
INVx1_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_542), .B(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_542), .B(n_647), .Y(n_705) );
OR2x2_ASAP7_75t_L g546 ( .A(n_543), .B(n_544), .Y(n_546) );
INVx1_ASAP7_75t_SL g598 ( .A(n_543), .Y(n_598) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AOI221xp5_ASAP7_75t_L g601 ( .A1(n_549), .A2(n_602), .B1(n_604), .B2(n_608), .C(n_609), .Y(n_601) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
OR2x2_ASAP7_75t_L g629 ( .A(n_550), .B(n_593), .Y(n_629) );
INVx2_ASAP7_75t_L g561 ( .A(n_551), .Y(n_561) );
INVx1_ASAP7_75t_L g587 ( .A(n_551), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_551), .B(n_571), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_551), .B(n_574), .Y(n_681) );
INVx1_ASAP7_75t_L g689 ( .A(n_551), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_553), .B(n_557), .Y(n_603) );
AND2x4_ASAP7_75t_L g578 ( .A(n_554), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g691 ( .A(n_557), .B(n_647), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_559), .B(n_562), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_560), .B(n_592), .Y(n_591) );
INVxp67_ASAP7_75t_L g699 ( .A(n_561), .Y(n_699) );
INVxp67_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_566), .Y(n_563) );
INVx1_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g599 ( .A(n_565), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g671 ( .A(n_565), .B(n_647), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_565), .B(n_584), .Y(n_677) );
AOI322xp5_ASAP7_75t_L g631 ( .A1(n_566), .A2(n_600), .A3(n_607), .B1(n_632), .B2(n_635), .C1(n_636), .C2(n_638), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_566), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
OR2x2_ASAP7_75t_L g697 ( .A(n_569), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g643 ( .A(n_570), .Y(n_643) );
INVx2_ASAP7_75t_L g574 ( .A(n_571), .Y(n_574) );
INVx1_ASAP7_75t_L g633 ( .A(n_571), .Y(n_633) );
CKINVDCx16_ASAP7_75t_R g580 ( .A(n_572), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
AND2x2_ASAP7_75t_L g669 ( .A(n_574), .B(n_582), .Y(n_669) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g581 ( .A(n_576), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g624 ( .A(n_576), .B(n_617), .Y(n_624) );
AND2x2_ASAP7_75t_L g628 ( .A(n_576), .B(n_588), .Y(n_628) );
OAI21xp33_ASAP7_75t_SL g638 ( .A1(n_577), .A2(n_639), .B(n_641), .Y(n_638) );
OAI22xp33_ASAP7_75t_L g708 ( .A1(n_577), .A2(n_709), .B1(n_710), .B2(n_712), .Y(n_708) );
INVx3_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g583 ( .A(n_578), .B(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_578), .B(n_598), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_580), .B(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx1_ASAP7_75t_L g720 ( .A(n_587), .Y(n_720) );
INVx4_ASAP7_75t_L g593 ( .A(n_588), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_588), .B(n_615), .Y(n_663) );
INVx1_ASAP7_75t_SL g675 ( .A(n_589), .Y(n_675) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NOR2xp67_ASAP7_75t_L g688 ( .A(n_593), .B(n_689), .Y(n_688) );
OAI211xp5_ASAP7_75t_SL g594 ( .A1(n_595), .A2(n_596), .B(n_601), .C(n_618), .Y(n_594) );
OAI221xp5_ASAP7_75t_SL g714 ( .A1(n_596), .A2(n_634), .B1(n_713), .B2(n_715), .C(n_717), .Y(n_714) );
INVx1_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_598), .B(n_711), .Y(n_710) );
OAI31xp33_ASAP7_75t_L g690 ( .A1(n_599), .A2(n_676), .A3(n_691), .B(n_692), .Y(n_690) );
INVx1_ASAP7_75t_L g630 ( .A(n_600), .Y(n_630) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_607), .Y(n_604) );
INVx1_ASAP7_75t_L g680 ( .A(n_605), .Y(n_680) );
AND2x2_ASAP7_75t_L g693 ( .A(n_607), .B(n_616), .Y(n_693) );
AOI21xp33_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_611), .B(n_613), .Y(n_609) );
INVx1_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
INVxp67_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_617), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_617), .B(n_720), .Y(n_719) );
OAI21xp33_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_620), .B(n_624), .Y(n_618) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OAI221xp5_ASAP7_75t_SL g625 ( .A1(n_626), .A2(n_627), .B1(n_629), .B2(n_630), .C(n_631), .Y(n_625) );
A2O1A1Ixp33_ASAP7_75t_L g694 ( .A1(n_626), .A2(n_695), .B(n_697), .C(n_700), .Y(n_694) );
CKINVDCx16_ASAP7_75t_R g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_629), .B(n_679), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
INVx1_ASAP7_75t_L g656 ( .A(n_637), .Y(n_656) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g642 ( .A(n_640), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g684 ( .A(n_640), .B(n_685), .Y(n_684) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OAI211xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_648), .B(n_650), .C(n_659), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
OAI221xp5_ASAP7_75t_L g721 ( .A1(n_648), .A2(n_658), .B1(n_722), .B2(n_723), .C(n_725), .Y(n_721) );
INVx1_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_653), .B1(n_654), .B2(n_657), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
OAI21xp5_ASAP7_75t_SL g659 ( .A1(n_660), .A2(n_661), .B(n_662), .Y(n_659) );
INVx1_ASAP7_75t_SL g722 ( .A(n_661), .Y(n_722) );
INVxp67_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NOR4xp25_ASAP7_75t_L g664 ( .A(n_665), .B(n_694), .C(n_714), .D(n_721), .Y(n_664) );
OAI211xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_670), .B(n_672), .C(n_690), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_667), .B(n_669), .Y(n_666) );
INVxp67_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
O2A1O1Ixp33_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_676), .B(n_678), .C(n_682), .Y(n_672) );
INVx1_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_SL g701 ( .A(n_679), .Y(n_701) );
OR2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
OR2x2_ASAP7_75t_L g712 ( .A(n_680), .B(n_713), .Y(n_712) );
OAI21xp33_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_686), .B(n_687), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AOI221xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_702), .B1(n_704), .B2(n_706), .C(n_708), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVxp67_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_711), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_740), .Y(n_744) );
endmodule