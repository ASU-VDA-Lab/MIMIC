module real_jpeg_25098_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_9;
wire n_72;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

OAI22xp33_ASAP7_75t_SL g14 ( 
.A1(n_2),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_14)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_2),
.A2(n_17),
.B1(n_24),
.B2(n_25),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_2),
.A2(n_17),
.B1(n_46),
.B2(n_48),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_5),
.A2(n_15),
.B1(n_18),
.B2(n_28),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_5),
.B(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_5),
.A2(n_28),
.B1(n_46),
.B2(n_48),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_5),
.B(n_15),
.C(n_40),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_5),
.B(n_21),
.C(n_24),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_5),
.B(n_61),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_5),
.B(n_26),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_7),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_29)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_68),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_67),
.Y(n_9)
);

INVxp67_ASAP7_75t_L g10 ( 
.A(n_11),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_41),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_12),
.B(n_41),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_29),
.C(n_36),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_13),
.A2(n_36),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_13),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_19),
.B1(n_26),
.B2(n_27),
.Y(n_13)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

INVx5_ASAP7_75t_SL g18 ( 
.A(n_15),
.Y(n_18)
);

OAI22xp33_ASAP7_75t_L g20 ( 
.A1(n_15),
.A2(n_18),
.B1(n_21),
.B2(n_22),
.Y(n_20)
);

OA22x2_ASAP7_75t_SL g38 ( 
.A1(n_15),
.A2(n_18),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_15),
.B(n_77),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_19),
.B(n_27),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_23),
.Y(n_19)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_21),
.Y(n_22)
);

OA22x2_ASAP7_75t_L g23 ( 
.A1(n_21),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_23)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_23),
.A2(n_54),
.B(n_55),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_24),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_24),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_29),
.B(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_29),
.B(n_84),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_29),
.A2(n_90),
.B1(n_91),
.B2(n_94),
.Y(n_89)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_31),
.B(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_31),
.B(n_35),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_33),
.A2(n_73),
.B(n_74),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_36),
.Y(n_93)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_45),
.B(n_49),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_40),
.B1(n_46),
.B2(n_48),
.Y(n_51)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_57),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_53),
.B2(n_56),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g48 ( 
.A(n_46),
.Y(n_48)
);

CKINVDCx6p67_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_52),
.Y(n_49)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_53),
.A2(n_56),
.B1(n_76),
.B2(n_78),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_78),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_58),
.Y(n_66)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_87),
.B(n_95),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_79),
.B(n_86),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_75),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_71),
.B(n_75),
.Y(n_86)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_72),
.B(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_76),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_83),
.B(n_85),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_88),
.B(n_89),
.Y(n_95)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);


endmodule