module fake_jpeg_16495_n_119 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_119);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_119;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_27),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_54),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_43),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_0),
.B(n_1),
.Y(n_66)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_48),
.Y(n_54)
);

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_45),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_55),
.Y(n_63)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_53),
.A2(n_40),
.B1(n_42),
.B2(n_46),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_64),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_37),
.Y(n_61)
);

OR2x2_ASAP7_75t_SL g75 ( 
.A(n_61),
.B(n_65),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_56),
.A2(n_49),
.B1(n_47),
.B2(n_50),
.Y(n_64)
);

CKINVDCx12_ASAP7_75t_R g65 ( 
.A(n_55),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_66),
.A2(n_4),
.B1(n_5),
.B2(n_49),
.Y(n_73)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_3),
.Y(n_69)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_74),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_73),
.A2(n_76),
.B1(n_71),
.B2(n_5),
.Y(n_85)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_81),
.B(n_82),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_58),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_63),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_83),
.A2(n_84),
.B1(n_85),
.B2(n_87),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_63),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_77),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_47),
.Y(n_88)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_76),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_90)
);

AOI22x1_ASAP7_75t_L g95 ( 
.A1(n_90),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_91),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_93),
.B(n_97),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_44),
.C(n_39),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_89),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_95),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_98),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_101),
.C(n_94),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g101 ( 
.A(n_96),
.B(n_86),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_102),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_103),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_19),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_100),
.A2(n_86),
.B1(n_39),
.B2(n_21),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_106),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_99),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_109),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_110),
.A2(n_107),
.B(n_22),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_108),
.B1(n_24),
.B2(n_25),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_113),
.A2(n_111),
.B1(n_26),
.B2(n_28),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_114),
.A2(n_20),
.B(n_30),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_116),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_34),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_35),
.Y(n_119)
);


endmodule