module fake_netlist_5_965_n_1854 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1854);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1854;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_798;
wire n_196;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_1809;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_677;
wire n_293;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_334;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_102),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_109),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_155),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_100),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_110),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_74),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_127),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_83),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_6),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_98),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g191 ( 
.A(n_117),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_16),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_150),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_58),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_75),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_21),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_76),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_6),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_119),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_138),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_90),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_156),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_121),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_96),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_49),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_58),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_140),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_54),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_173),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_125),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_62),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_47),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_64),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_47),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_114),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_123),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_162),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_131),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_0),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_63),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_7),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_10),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_59),
.Y(n_223)
);

BUFx8_ASAP7_75t_SL g224 ( 
.A(n_169),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_3),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_69),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_52),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_161),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_139),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_77),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_11),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_14),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_60),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_142),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_60),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_115),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_108),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_2),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_37),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_134),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_45),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_73),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_89),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_167),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_136),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_38),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_36),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_157),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_12),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_105),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_29),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_22),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_153),
.Y(n_253)
);

BUFx10_ASAP7_75t_L g254 ( 
.A(n_84),
.Y(n_254)
);

BUFx10_ASAP7_75t_L g255 ( 
.A(n_148),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_20),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_92),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_72),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_179),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_177),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_67),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_118),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_18),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_1),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_39),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_130),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_50),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_37),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_86),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_8),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_53),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_116),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_52),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_81),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_3),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_34),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_93),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_120),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_56),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_16),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_28),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_94),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_78),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_163),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_106),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_9),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_112),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_45),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_132),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_68),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_19),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_101),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_26),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_61),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_57),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_8),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_53),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_166),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_46),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_154),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_85),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_70),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_164),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_50),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_87),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_0),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_48),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_20),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_82),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_137),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_172),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_40),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_56),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_180),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_13),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_15),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_129),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_44),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_22),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_59),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_122),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g322 ( 
.A(n_158),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_128),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_104),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_44),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_88),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_33),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_91),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_38),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_17),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_66),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_46),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_143),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_48),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_171),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_55),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_1),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_165),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_170),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_151),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_36),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_51),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_35),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_152),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_43),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_39),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_21),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_124),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_51),
.Y(n_349)
);

BUFx10_ASAP7_75t_L g350 ( 
.A(n_17),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_99),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_135),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_57),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_65),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_5),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_7),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_49),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_41),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_11),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_159),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_224),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_186),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_317),
.B(n_2),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_214),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_182),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_221),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_222),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_222),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_183),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_184),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_187),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_221),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_185),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_188),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_313),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_190),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_313),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_234),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_336),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_193),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_336),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_195),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_201),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_294),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_197),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_317),
.B(n_4),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_263),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g388 ( 
.A(n_211),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_199),
.Y(n_389)
);

INVxp33_ASAP7_75t_SL g390 ( 
.A(n_312),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_202),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_341),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_341),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_352),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_189),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_263),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_200),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_209),
.Y(n_398)
);

INVxp33_ASAP7_75t_SL g399 ( 
.A(n_327),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_327),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_213),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_189),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_192),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_215),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_216),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_217),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_192),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_228),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_194),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_194),
.Y(n_410)
);

NOR2xp67_ASAP7_75t_L g411 ( 
.A(n_232),
.B(n_4),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_232),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_191),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_218),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_311),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_238),
.Y(n_416)
);

NOR2xp67_ASAP7_75t_L g417 ( 
.A(n_233),
.B(n_5),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_233),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_320),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_229),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_235),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_235),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_246),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_236),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_322),
.B(n_9),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_246),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_247),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_242),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_355),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_244),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_322),
.B(n_10),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_247),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_245),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_191),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_248),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_251),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_196),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_257),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_326),
.B(n_12),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_251),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g441 ( 
.A(n_254),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_264),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_260),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_264),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_266),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_274),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_277),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_234),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_326),
.B(n_13),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_431),
.B(n_278),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_395),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_395),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_402),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_439),
.B(n_282),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_429),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_437),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_378),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_413),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_367),
.Y(n_459)
);

AND2x6_ASAP7_75t_L g460 ( 
.A(n_413),
.B(n_181),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_402),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_403),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_378),
.B(n_284),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_413),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_403),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_425),
.B(n_261),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_378),
.B(n_243),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_407),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_434),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_448),
.B(n_366),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_434),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_434),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_366),
.Y(n_473)
);

AND2x6_ASAP7_75t_L g474 ( 
.A(n_449),
.B(n_181),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_448),
.B(n_285),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_448),
.B(n_243),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_372),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_407),
.B(n_289),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_409),
.B(n_292),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_409),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_372),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_375),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_375),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_377),
.B(n_379),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_410),
.B(n_301),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_377),
.B(n_262),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_379),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_381),
.Y(n_488)
);

OA21x2_ASAP7_75t_L g489 ( 
.A1(n_381),
.A2(n_204),
.B(n_203),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_367),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_410),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_412),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_412),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_418),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_418),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_392),
.Y(n_496)
);

CKINVDCx6p67_ASAP7_75t_R g497 ( 
.A(n_364),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_421),
.B(n_303),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_399),
.A2(n_223),
.B1(n_357),
.B2(n_353),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_421),
.B(n_422),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_422),
.Y(n_501)
);

NAND2xp33_ASAP7_75t_SL g502 ( 
.A(n_416),
.B(n_419),
.Y(n_502)
);

NAND2xp33_ASAP7_75t_L g503 ( 
.A(n_423),
.B(n_181),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_423),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_426),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_368),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_411),
.B(n_262),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_426),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_392),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_393),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_393),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_427),
.B(n_310),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_427),
.Y(n_513)
);

NAND2xp33_ASAP7_75t_L g514 ( 
.A(n_432),
.B(n_181),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_432),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_387),
.Y(n_516)
);

NAND2xp33_ASAP7_75t_L g517 ( 
.A(n_436),
.B(n_181),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_436),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_440),
.Y(n_519)
);

NAND2xp33_ASAP7_75t_L g520 ( 
.A(n_440),
.B(n_240),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_442),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_442),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_444),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_444),
.Y(n_524)
);

INVx4_ASAP7_75t_L g525 ( 
.A(n_365),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_411),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_369),
.Y(n_527)
);

INVx4_ASAP7_75t_L g528 ( 
.A(n_464),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_466),
.A2(n_435),
.B1(n_424),
.B2(n_430),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_464),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_469),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_470),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_466),
.B(n_370),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_457),
.B(n_373),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_464),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_470),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_457),
.B(n_374),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_469),
.Y(n_538)
);

OR2x2_ASAP7_75t_L g539 ( 
.A(n_459),
.B(n_364),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_457),
.B(n_376),
.Y(n_540)
);

INVx4_ASAP7_75t_L g541 ( 
.A(n_464),
.Y(n_541)
);

NAND3xp33_ASAP7_75t_L g542 ( 
.A(n_456),
.B(n_386),
.C(n_363),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_450),
.B(n_380),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_450),
.B(n_382),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_470),
.Y(n_545)
);

OAI22xp33_ASAP7_75t_L g546 ( 
.A1(n_459),
.A2(n_441),
.B1(n_388),
.B2(n_279),
.Y(n_546)
);

AND3x4_ASAP7_75t_L g547 ( 
.A(n_499),
.B(n_417),
.C(n_307),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_457),
.B(n_417),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_464),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_454),
.B(n_385),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g551 ( 
.A1(n_454),
.A2(n_438),
.B1(n_433),
.B2(n_390),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_SL g552 ( 
.A(n_497),
.B(n_361),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_451),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_469),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_471),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_490),
.B(n_362),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_451),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_452),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_527),
.B(n_250),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_463),
.B(n_389),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_452),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_464),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_464),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_527),
.B(n_250),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_458),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_453),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_497),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_471),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_453),
.Y(n_569)
);

BUFx10_ASAP7_75t_L g570 ( 
.A(n_507),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_463),
.B(n_391),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_458),
.Y(n_572)
);

INVx1_ASAP7_75t_SL g573 ( 
.A(n_490),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_461),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_471),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_461),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_526),
.B(n_396),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_458),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_462),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_474),
.A2(n_400),
.B1(n_212),
.B2(n_307),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_526),
.B(n_441),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_462),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_472),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_465),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_458),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_472),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_467),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_458),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_497),
.Y(n_589)
);

OR2x6_ASAP7_75t_L g590 ( 
.A(n_527),
.B(n_212),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_458),
.Y(n_591)
);

OAI22xp33_ASAP7_75t_L g592 ( 
.A1(n_456),
.A2(n_208),
.B1(n_359),
.B2(n_288),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_458),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_465),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_458),
.Y(n_595)
);

INVx8_ASAP7_75t_L g596 ( 
.A(n_474),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_472),
.Y(n_597)
);

INVx4_ASAP7_75t_L g598 ( 
.A(n_460),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_477),
.Y(n_599)
);

INVx4_ASAP7_75t_L g600 ( 
.A(n_460),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_475),
.B(n_398),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_474),
.A2(n_315),
.B1(n_267),
.B2(n_286),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_467),
.B(n_401),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_SL g604 ( 
.A(n_467),
.B(n_337),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_477),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_R g606 ( 
.A(n_527),
.B(n_404),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_476),
.Y(n_607)
);

INVx1_ASAP7_75t_SL g608 ( 
.A(n_476),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_468),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_475),
.B(n_405),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_525),
.B(n_406),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_507),
.B(n_408),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_502),
.Y(n_613)
);

OR2x6_ASAP7_75t_L g614 ( 
.A(n_527),
.B(n_315),
.Y(n_614)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_460),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_476),
.B(n_420),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_477),
.Y(n_617)
);

INVx1_ASAP7_75t_SL g618 ( 
.A(n_502),
.Y(n_618)
);

INVx1_ASAP7_75t_SL g619 ( 
.A(n_506),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_468),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_507),
.B(n_428),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_474),
.A2(n_349),
.B1(n_267),
.B2(n_286),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_477),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_474),
.A2(n_347),
.B1(n_295),
.B2(n_356),
.Y(n_624)
);

INVx4_ASAP7_75t_L g625 ( 
.A(n_460),
.Y(n_625)
);

OR2x6_ASAP7_75t_L g626 ( 
.A(n_525),
.B(n_295),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_486),
.B(n_443),
.Y(n_627)
);

OAI22xp33_ASAP7_75t_L g628 ( 
.A1(n_516),
.A2(n_455),
.B1(n_205),
.B2(n_206),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_480),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_477),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_507),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_474),
.A2(n_318),
.B1(n_297),
.B2(n_356),
.Y(n_632)
);

INVxp67_ASAP7_75t_L g633 ( 
.A(n_506),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_480),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_491),
.Y(n_635)
);

BUFx2_ASAP7_75t_L g636 ( 
.A(n_455),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_491),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_492),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_477),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_516),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_525),
.B(n_445),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_525),
.B(n_446),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_507),
.B(n_447),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_478),
.B(n_272),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_477),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_486),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_525),
.B(n_478),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_496),
.Y(n_648)
);

CKINVDCx16_ASAP7_75t_R g649 ( 
.A(n_499),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_492),
.Y(n_650)
);

OR2x6_ASAP7_75t_L g651 ( 
.A(n_479),
.B(n_297),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_496),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_486),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_489),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_479),
.Y(n_655)
);

AO22x2_ASAP7_75t_L g656 ( 
.A1(n_485),
.A2(n_347),
.B1(n_304),
.B2(n_308),
.Y(n_656)
);

AND2x6_ASAP7_75t_L g657 ( 
.A(n_485),
.B(n_259),
.Y(n_657)
);

AO21x2_ASAP7_75t_L g658 ( 
.A1(n_498),
.A2(n_204),
.B(n_203),
.Y(n_658)
);

INVx4_ASAP7_75t_L g659 ( 
.A(n_460),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_498),
.B(n_259),
.Y(n_660)
);

AND2x6_ASAP7_75t_L g661 ( 
.A(n_512),
.B(n_333),
.Y(n_661)
);

CKINVDCx6p67_ASAP7_75t_R g662 ( 
.A(n_512),
.Y(n_662)
);

AND2x6_ASAP7_75t_L g663 ( 
.A(n_493),
.B(n_333),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_493),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_494),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_494),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_474),
.A2(n_304),
.B1(n_308),
.B2(n_316),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_513),
.B(n_348),
.Y(n_668)
);

BUFx2_ASAP7_75t_L g669 ( 
.A(n_474),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_496),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_474),
.A2(n_330),
.B1(n_316),
.B2(n_318),
.Y(n_671)
);

BUFx2_ASAP7_75t_L g672 ( 
.A(n_474),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_495),
.B(n_314),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_484),
.B(n_207),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_496),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_495),
.B(n_397),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_501),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_489),
.A2(n_330),
.B1(n_342),
.B2(n_349),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_513),
.B(n_348),
.Y(n_679)
);

NAND3xp33_ASAP7_75t_L g680 ( 
.A(n_533),
.B(n_219),
.C(n_198),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_531),
.Y(n_681)
);

BUFx6f_ASAP7_75t_SL g682 ( 
.A(n_626),
.Y(n_682)
);

OAI221xp5_ASAP7_75t_L g683 ( 
.A1(n_580),
.A2(n_646),
.B1(n_542),
.B2(n_532),
.C(n_545),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_573),
.B(n_371),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_539),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_587),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_SL g687 ( 
.A(n_567),
.B(n_589),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_587),
.Y(n_688)
);

NOR2xp67_ASAP7_75t_L g689 ( 
.A(n_529),
.B(n_501),
.Y(n_689)
);

NAND3xp33_ASAP7_75t_L g690 ( 
.A(n_655),
.B(n_227),
.C(n_225),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_607),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_538),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_607),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_655),
.B(n_608),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_647),
.B(n_240),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_536),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_653),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_SL g698 ( 
.A(n_567),
.B(n_383),
.Y(n_698)
);

NOR2xp67_ASAP7_75t_L g699 ( 
.A(n_611),
.B(n_504),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_653),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_543),
.B(n_544),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_631),
.B(n_240),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_610),
.B(n_487),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_550),
.B(n_487),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_631),
.B(n_240),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_646),
.A2(n_414),
.B1(n_415),
.B2(n_384),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_538),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_644),
.B(n_487),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_581),
.B(n_231),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_554),
.Y(n_710)
);

INVxp67_ASAP7_75t_L g711 ( 
.A(n_640),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_539),
.Y(n_712)
);

A2O1A1Ixp33_ASAP7_75t_L g713 ( 
.A1(n_654),
.A2(n_351),
.B(n_258),
.C(n_269),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_560),
.B(n_487),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_581),
.B(n_239),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_627),
.B(n_394),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_554),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_553),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_557),
.Y(n_719)
);

BUFx5_ASAP7_75t_L g720 ( 
.A(n_654),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_558),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_612),
.A2(n_500),
.B(n_503),
.Y(n_722)
);

NOR2x1p5_ASAP7_75t_L g723 ( 
.A(n_589),
.B(n_241),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_571),
.B(n_487),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_627),
.B(n_603),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_603),
.Y(n_726)
);

NOR3xp33_ASAP7_75t_L g727 ( 
.A(n_604),
.B(n_210),
.C(n_207),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_561),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_570),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_566),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_555),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_555),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_568),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_601),
.B(n_548),
.Y(n_734)
);

AND2x6_ASAP7_75t_L g735 ( 
.A(n_674),
.B(n_210),
.Y(n_735)
);

NAND2xp33_ASAP7_75t_L g736 ( 
.A(n_657),
.B(n_191),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_569),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_574),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_576),
.Y(n_739)
);

OR2x2_ASAP7_75t_L g740 ( 
.A(n_619),
.B(n_500),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_579),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_548),
.B(n_511),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_621),
.A2(n_514),
.B(n_503),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_548),
.B(n_511),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_570),
.B(n_240),
.Y(n_745)
);

O2A1O1Ixp33_ASAP7_75t_L g746 ( 
.A1(n_660),
.A2(n_524),
.B(n_508),
.C(n_522),
.Y(n_746)
);

INVx8_ASAP7_75t_L g747 ( 
.A(n_590),
.Y(n_747)
);

NOR3xp33_ASAP7_75t_SL g748 ( 
.A(n_649),
.B(n_252),
.C(n_249),
.Y(n_748)
);

O2A1O1Ixp33_ASAP7_75t_L g749 ( 
.A1(n_660),
.A2(n_524),
.B(n_508),
.C(n_522),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_616),
.B(n_321),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_582),
.B(n_511),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_584),
.B(n_511),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_594),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_662),
.B(n_256),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_609),
.B(n_511),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_620),
.B(n_489),
.Y(n_756)
);

INVxp33_ASAP7_75t_L g757 ( 
.A(n_556),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_640),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_629),
.B(n_634),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_635),
.B(n_489),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_636),
.B(n_484),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_637),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_638),
.B(n_489),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_650),
.B(n_513),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_568),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_570),
.B(n_283),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_598),
.B(n_283),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_636),
.B(n_484),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_575),
.Y(n_769)
);

AOI22xp5_ASAP7_75t_L g770 ( 
.A1(n_662),
.A2(n_323),
.B1(n_328),
.B2(n_331),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_664),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_643),
.A2(n_514),
.B(n_520),
.Y(n_772)
);

INVxp67_ASAP7_75t_SL g773 ( 
.A(n_665),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_616),
.B(n_265),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_577),
.B(n_268),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_666),
.B(n_515),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_565),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_677),
.B(n_674),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_598),
.B(n_283),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_606),
.A2(n_340),
.B1(n_335),
.B2(n_338),
.Y(n_780)
);

INVx2_ASAP7_75t_SL g781 ( 
.A(n_577),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_641),
.B(n_515),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_676),
.B(n_270),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_626),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_575),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_583),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_642),
.B(n_515),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_559),
.B(n_518),
.Y(n_788)
);

BUFx10_ASAP7_75t_L g789 ( 
.A(n_613),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_633),
.B(n_651),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_600),
.B(n_283),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_600),
.B(n_191),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_586),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_559),
.B(n_518),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_564),
.B(n_518),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_564),
.B(n_523),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_534),
.B(n_523),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_537),
.B(n_540),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_586),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_669),
.Y(n_800)
);

BUFx5_ASAP7_75t_L g801 ( 
.A(n_663),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_597),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_600),
.B(n_191),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_615),
.B(n_191),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_673),
.B(n_658),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_658),
.B(n_523),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_658),
.B(n_496),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_669),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_546),
.B(n_344),
.Y(n_809)
);

OR2x6_ASAP7_75t_L g810 ( 
.A(n_590),
.B(n_342),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_551),
.B(n_628),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_651),
.B(n_496),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_597),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_668),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_668),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_604),
.B(n_354),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_679),
.Y(n_817)
);

INVxp67_ASAP7_75t_L g818 ( 
.A(n_651),
.Y(n_818)
);

O2A1O1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_651),
.A2(n_521),
.B(n_519),
.C(n_505),
.Y(n_819)
);

AOI22xp5_ASAP7_75t_L g820 ( 
.A1(n_590),
.A2(n_253),
.B1(n_360),
.B2(n_351),
.Y(n_820)
);

INVx2_ASAP7_75t_SL g821 ( 
.A(n_626),
.Y(n_821)
);

BUFx6f_ASAP7_75t_SL g822 ( 
.A(n_626),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_613),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_679),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_590),
.B(n_271),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_678),
.B(n_496),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_591),
.B(n_496),
.Y(n_827)
);

AOI22xp5_ASAP7_75t_L g828 ( 
.A1(n_614),
.A2(n_237),
.B1(n_360),
.B2(n_339),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_623),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_591),
.B(n_220),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_672),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_591),
.B(n_220),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_623),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_595),
.B(n_226),
.Y(n_834)
);

NOR3xp33_ASAP7_75t_L g835 ( 
.A(n_592),
.B(n_237),
.C(n_339),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_615),
.B(n_191),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_R g837 ( 
.A(n_552),
.B(n_273),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_595),
.B(n_226),
.Y(n_838)
);

OAI22xp33_ASAP7_75t_L g839 ( 
.A1(n_614),
.A2(n_230),
.B1(n_324),
.B2(n_309),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_639),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_639),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_648),
.Y(n_842)
);

NAND2xp33_ASAP7_75t_L g843 ( 
.A(n_657),
.B(n_191),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_596),
.A2(n_517),
.B(n_520),
.Y(n_844)
);

INVxp67_ASAP7_75t_L g845 ( 
.A(n_656),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_615),
.B(n_230),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_L g847 ( 
.A1(n_701),
.A2(n_614),
.B1(n_672),
.B2(n_547),
.Y(n_847)
);

NOR3xp33_ASAP7_75t_L g848 ( 
.A(n_811),
.B(n_618),
.C(n_258),
.Y(n_848)
);

NOR2x1_ASAP7_75t_L g849 ( 
.A(n_740),
.B(n_547),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_734),
.A2(n_797),
.B(n_744),
.Y(n_850)
);

NAND2xp33_ASAP7_75t_L g851 ( 
.A(n_800),
.B(n_808),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_773),
.B(n_657),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_798),
.B(n_657),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_720),
.B(n_625),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_800),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_800),
.Y(n_856)
);

INVx5_ASAP7_75t_L g857 ( 
.A(n_800),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_742),
.A2(n_596),
.B(n_528),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_703),
.A2(n_596),
.B(n_528),
.Y(n_859)
);

BUFx2_ASAP7_75t_L g860 ( 
.A(n_684),
.Y(n_860)
);

OAI21xp5_ASAP7_75t_L g861 ( 
.A1(n_805),
.A2(n_595),
.B(n_549),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_699),
.B(n_657),
.Y(n_862)
);

INVx4_ASAP7_75t_L g863 ( 
.A(n_808),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_714),
.A2(n_596),
.B(n_528),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_720),
.B(n_625),
.Y(n_865)
);

INVx11_ASAP7_75t_L g866 ( 
.A(n_735),
.Y(n_866)
);

BUFx2_ASAP7_75t_L g867 ( 
.A(n_711),
.Y(n_867)
);

NOR2x1_ASAP7_75t_L g868 ( 
.A(n_694),
.B(n_625),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_778),
.B(n_657),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_720),
.B(n_659),
.Y(n_870)
);

INVx3_ASAP7_75t_L g871 ( 
.A(n_808),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_720),
.B(n_808),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_831),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_691),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_782),
.B(n_787),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_711),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_761),
.B(n_656),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_720),
.B(n_831),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_691),
.B(n_661),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_831),
.B(n_661),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_831),
.B(n_661),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_783),
.B(n_661),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_724),
.A2(n_541),
.B(n_593),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_783),
.B(n_661),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_694),
.B(n_530),
.Y(n_885)
);

OAI21x1_ASAP7_75t_L g886 ( 
.A1(n_827),
.A2(n_530),
.B(n_535),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_696),
.B(n_661),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_704),
.B(n_656),
.Y(n_888)
);

OAI21xp5_ASAP7_75t_L g889 ( 
.A1(n_807),
.A2(n_563),
.B(n_549),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_697),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_708),
.A2(n_541),
.B(n_593),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_758),
.B(n_530),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_700),
.Y(n_893)
);

INVx2_ASAP7_75t_SL g894 ( 
.A(n_781),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_686),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_718),
.B(n_656),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_826),
.A2(n_541),
.B(n_593),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_688),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_693),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_722),
.A2(n_659),
.B(n_562),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_768),
.B(n_350),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_719),
.B(n_535),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_844),
.A2(n_659),
.B(n_562),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_721),
.B(n_535),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_728),
.B(n_730),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_720),
.B(n_565),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_745),
.A2(n_562),
.B(n_572),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_801),
.B(n_565),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_738),
.B(n_549),
.Y(n_909)
);

INVxp67_ASAP7_75t_L g910 ( 
.A(n_790),
.Y(n_910)
);

INVx4_ASAP7_75t_L g911 ( 
.A(n_747),
.Y(n_911)
);

AOI22xp5_ASAP7_75t_L g912 ( 
.A1(n_725),
.A2(n_663),
.B1(n_563),
.B2(n_602),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_739),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_741),
.B(n_563),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_758),
.B(n_562),
.Y(n_915)
);

NOR2x1_ASAP7_75t_L g916 ( 
.A(n_690),
.B(n_823),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_753),
.B(n_565),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_762),
.B(n_565),
.Y(n_918)
);

INVx3_ASAP7_75t_L g919 ( 
.A(n_777),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_745),
.A2(n_562),
.B(n_572),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_L g921 ( 
.A1(n_756),
.A2(n_652),
.B(n_671),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_683),
.A2(n_622),
.B1(n_624),
.B2(n_667),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_685),
.B(n_712),
.Y(n_923)
);

O2A1O1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_845),
.A2(n_713),
.B(n_818),
.C(n_835),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_771),
.B(n_572),
.Y(n_925)
);

INVxp67_ASAP7_75t_L g926 ( 
.A(n_775),
.Y(n_926)
);

AOI33xp33_ASAP7_75t_L g927 ( 
.A1(n_726),
.A2(n_504),
.A3(n_521),
.B1(n_519),
.B2(n_505),
.B3(n_632),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_759),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_775),
.B(n_572),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_818),
.B(n_572),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_764),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_766),
.A2(n_578),
.B(n_585),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_737),
.B(n_253),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_776),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_774),
.B(n_350),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_774),
.B(n_350),
.Y(n_936)
);

AOI21xp33_ASAP7_75t_L g937 ( 
.A1(n_709),
.A2(n_324),
.B(n_309),
.Y(n_937)
);

BUFx6f_ASAP7_75t_SL g938 ( 
.A(n_789),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_709),
.B(n_578),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_715),
.B(n_578),
.Y(n_940)
);

A2O1A1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_819),
.A2(n_269),
.B(n_305),
.C(n_287),
.Y(n_941)
);

BUFx8_ASAP7_75t_SL g942 ( 
.A(n_682),
.Y(n_942)
);

O2A1O1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_845),
.A2(n_287),
.B(n_302),
.C(n_300),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_715),
.B(n_578),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_760),
.A2(n_670),
.B(n_645),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_785),
.Y(n_946)
);

INVxp67_ASAP7_75t_L g947 ( 
.A(n_689),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_766),
.A2(n_578),
.B(n_585),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_735),
.B(n_729),
.Y(n_949)
);

BUFx12f_ASAP7_75t_L g950 ( 
.A(n_789),
.Y(n_950)
);

INVx5_ASAP7_75t_L g951 ( 
.A(n_735),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_763),
.A2(n_585),
.B(n_588),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_729),
.A2(n_585),
.B(n_588),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_735),
.B(n_814),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_846),
.A2(n_585),
.B(n_588),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_793),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_801),
.B(n_588),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_806),
.A2(n_670),
.B(n_645),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_716),
.B(n_588),
.Y(n_959)
);

NOR2xp67_ASAP7_75t_L g960 ( 
.A(n_680),
.B(n_599),
.Y(n_960)
);

AOI21x1_ASAP7_75t_L g961 ( 
.A1(n_792),
.A2(n_483),
.B(n_473),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_846),
.A2(n_675),
.B(n_617),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_735),
.B(n_663),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_799),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_777),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_815),
.B(n_663),
.Y(n_966)
);

AOI22xp33_ASAP7_75t_L g967 ( 
.A1(n_835),
.A2(n_663),
.B1(n_305),
.B2(n_298),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_747),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_801),
.B(n_599),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_817),
.B(n_663),
.Y(n_970)
);

NAND2x1p5_ASAP7_75t_L g971 ( 
.A(n_784),
.B(n_599),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_839),
.A2(n_302),
.B(n_300),
.C(n_298),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_813),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_751),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_824),
.B(n_695),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_767),
.A2(n_675),
.B(n_617),
.Y(n_976)
);

OAI21xp5_ASAP7_75t_L g977 ( 
.A1(n_695),
.A2(n_670),
.B(n_645),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_723),
.Y(n_978)
);

BUFx4f_ASAP7_75t_L g979 ( 
.A(n_747),
.Y(n_979)
);

AOI21x1_ASAP7_75t_L g980 ( 
.A1(n_792),
.A2(n_483),
.B(n_482),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_746),
.B(n_605),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_752),
.Y(n_982)
);

AND2x2_ASAP7_75t_SL g983 ( 
.A(n_727),
.B(n_290),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_810),
.Y(n_984)
);

AOI21x1_ASAP7_75t_L g985 ( 
.A1(n_803),
.A2(n_483),
.B(n_482),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_821),
.B(n_290),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_779),
.A2(n_675),
.B(n_617),
.Y(n_987)
);

AOI21x1_ASAP7_75t_L g988 ( 
.A1(n_803),
.A2(n_488),
.B(n_482),
.Y(n_988)
);

NOR2xp67_ASAP7_75t_L g989 ( 
.A(n_780),
.B(n_605),
.Y(n_989)
);

NAND2x1p5_ASAP7_75t_L g990 ( 
.A(n_829),
.B(n_605),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_754),
.B(n_275),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_812),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_779),
.A2(n_791),
.B(n_804),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_791),
.A2(n_675),
.B(n_617),
.Y(n_994)
);

AOI22x1_ASAP7_75t_L g995 ( 
.A1(n_743),
.A2(n_630),
.B1(n_332),
.B2(n_329),
.Y(n_995)
);

AOI21x1_ASAP7_75t_L g996 ( 
.A1(n_804),
.A2(n_481),
.B(n_473),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_749),
.B(n_630),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_755),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_836),
.A2(n_630),
.B(n_517),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_772),
.A2(n_510),
.B(n_509),
.Y(n_1000)
);

NAND2xp33_ASAP7_75t_L g1001 ( 
.A(n_801),
.B(n_460),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_754),
.Y(n_1002)
);

INVx2_ASAP7_75t_SL g1003 ( 
.A(n_750),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_R g1004 ( 
.A(n_698),
.B(n_687),
.Y(n_1004)
);

O2A1O1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_839),
.A2(n_510),
.B(n_509),
.C(n_488),
.Y(n_1005)
);

NOR2xp67_ASAP7_75t_L g1006 ( 
.A(n_770),
.B(n_71),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_842),
.B(n_510),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_681),
.B(n_473),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_810),
.B(n_481),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_788),
.A2(n_460),
.B(n_481),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_702),
.A2(n_488),
.B(n_460),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_702),
.A2(n_705),
.B(n_796),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_705),
.A2(n_460),
.B(n_358),
.Y(n_1013)
);

AND2x4_ASAP7_75t_L g1014 ( 
.A(n_810),
.B(n_113),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_794),
.A2(n_346),
.B(n_345),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_795),
.A2(n_343),
.B(n_334),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_801),
.B(n_254),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_825),
.B(n_325),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_833),
.A2(n_319),
.B(n_306),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_840),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_841),
.A2(n_299),
.B(n_296),
.Y(n_1021)
);

AOI22xp33_ASAP7_75t_L g1022 ( 
.A1(n_727),
.A2(n_255),
.B1(n_254),
.B2(n_281),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_830),
.A2(n_293),
.B(n_291),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_692),
.B(n_280),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_832),
.A2(n_276),
.B(n_79),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_707),
.Y(n_1026)
);

AOI22xp33_ASAP7_75t_L g1027 ( 
.A1(n_736),
.A2(n_843),
.B1(n_786),
.B2(n_769),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_710),
.B(n_255),
.Y(n_1028)
);

AOI21x1_ASAP7_75t_L g1029 ( 
.A1(n_834),
.A2(n_255),
.B(n_178),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_825),
.B(n_14),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_717),
.B(n_15),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_731),
.B(n_18),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_857),
.Y(n_1033)
);

O2A1O1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_937),
.A2(n_809),
.B(n_816),
.C(n_748),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_928),
.B(n_828),
.Y(n_1035)
);

NOR3xp33_ASAP7_75t_L g1036 ( 
.A(n_991),
.B(n_706),
.C(n_820),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_855),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_913),
.Y(n_1038)
);

A2O1A1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_991),
.A2(n_748),
.B(n_838),
.C(n_765),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_926),
.A2(n_732),
.B(n_802),
.C(n_733),
.Y(n_1040)
);

NOR3xp33_ASAP7_75t_L g1041 ( 
.A(n_926),
.B(n_947),
.C(n_849),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_857),
.B(n_837),
.Y(n_1042)
);

O2A1O1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_947),
.A2(n_757),
.B(n_837),
.C(n_822),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_875),
.B(n_801),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_946),
.Y(n_1045)
);

OAI22x1_ASAP7_75t_L g1046 ( 
.A1(n_910),
.A2(n_822),
.B1(n_682),
.B2(n_24),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_851),
.A2(n_176),
.B(n_175),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_922),
.A2(n_19),
.B1(n_23),
.B2(n_24),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_931),
.B(n_174),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_857),
.B(n_168),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_1002),
.B(n_23),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_855),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_847),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_857),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_850),
.A2(n_160),
.B(n_149),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_1004),
.B(n_147),
.Y(n_1056)
);

OA21x2_ASAP7_75t_L g1057 ( 
.A1(n_861),
.A2(n_146),
.B(n_145),
.Y(n_1057)
);

AO21x1_ASAP7_75t_L g1058 ( 
.A1(n_944),
.A2(n_25),
.B(n_27),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_867),
.B(n_28),
.Y(n_1059)
);

INVx3_ASAP7_75t_L g1060 ( 
.A(n_855),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_876),
.B(n_29),
.Y(n_1061)
);

AOI221xp5_ASAP7_75t_L g1062 ( 
.A1(n_1022),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.C(n_33),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_901),
.B(n_30),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_924),
.A2(n_959),
.B(n_935),
.C(n_936),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_934),
.B(n_31),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_959),
.A2(n_32),
.B(n_34),
.C(n_35),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_855),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_876),
.B(n_860),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_910),
.B(n_40),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_885),
.B(n_848),
.Y(n_1070)
);

O2A1O1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_848),
.A2(n_41),
.B(n_42),
.C(n_43),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_886),
.A2(n_103),
.B(n_141),
.Y(n_1072)
);

CKINVDCx8_ASAP7_75t_R g1073 ( 
.A(n_968),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_854),
.A2(n_97),
.B(n_133),
.Y(n_1074)
);

INVx3_ASAP7_75t_L g1075 ( 
.A(n_863),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_1018),
.B(n_42),
.Y(n_1076)
);

AOI22xp33_ASAP7_75t_L g1077 ( 
.A1(n_983),
.A2(n_54),
.B1(n_55),
.B2(n_80),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_854),
.A2(n_95),
.B(n_107),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_865),
.A2(n_111),
.B(n_126),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_950),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_865),
.A2(n_144),
.B(n_870),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_870),
.A2(n_903),
.B(n_859),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_864),
.A2(n_878),
.B(n_872),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_896),
.A2(n_888),
.B1(n_967),
.B2(n_877),
.Y(n_1084)
);

CKINVDCx20_ASAP7_75t_R g1085 ( 
.A(n_1004),
.Y(n_1085)
);

NOR3xp33_ASAP7_75t_SL g1086 ( 
.A(n_923),
.B(n_899),
.C(n_890),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_863),
.Y(n_1087)
);

INVx8_ASAP7_75t_L g1088 ( 
.A(n_968),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_1003),
.B(n_1030),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_942),
.Y(n_1090)
);

O2A1O1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_972),
.A2(n_943),
.B(n_941),
.C(n_905),
.Y(n_1091)
);

A2O1A1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_944),
.A2(n_853),
.B(n_954),
.C(n_993),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_933),
.B(n_923),
.Y(n_1093)
);

INVx2_ASAP7_75t_SL g1094 ( 
.A(n_894),
.Y(n_1094)
);

OR2x6_ASAP7_75t_L g1095 ( 
.A(n_968),
.B(n_911),
.Y(n_1095)
);

OA22x2_ASAP7_75t_L g1096 ( 
.A1(n_984),
.A2(n_978),
.B1(n_1014),
.B2(n_933),
.Y(n_1096)
);

BUFx4f_ASAP7_75t_L g1097 ( 
.A(n_968),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_986),
.B(n_893),
.Y(n_1098)
);

NAND2x1p5_ASAP7_75t_L g1099 ( 
.A(n_856),
.B(n_871),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_885),
.B(n_974),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_952),
.A2(n_961),
.B(n_996),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_982),
.B(n_998),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_979),
.Y(n_1103)
);

OR2x2_ASAP7_75t_L g1104 ( 
.A(n_895),
.B(n_898),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_992),
.B(n_929),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_992),
.B(n_939),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_992),
.B(n_856),
.Y(n_1107)
);

OAI21xp33_ASAP7_75t_L g1108 ( 
.A1(n_1022),
.A2(n_983),
.B(n_986),
.Y(n_1108)
);

O2A1O1Ixp5_ASAP7_75t_SL g1109 ( 
.A1(n_1017),
.A2(n_884),
.B(n_882),
.C(n_964),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_940),
.A2(n_906),
.B(n_881),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_906),
.A2(n_880),
.B(n_883),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_979),
.Y(n_1112)
);

OAI21xp33_ASAP7_75t_L g1113 ( 
.A1(n_916),
.A2(n_1024),
.B(n_967),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_1028),
.A2(n_1032),
.B(n_1031),
.C(n_869),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_911),
.Y(n_1115)
);

OR2x6_ASAP7_75t_SL g1116 ( 
.A(n_874),
.B(n_956),
.Y(n_1116)
);

OAI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_945),
.A2(n_958),
.B(n_889),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_858),
.A2(n_908),
.B(n_957),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_992),
.B(n_975),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_915),
.B(n_892),
.Y(n_1120)
);

INVx3_ASAP7_75t_L g1121 ( 
.A(n_871),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_1012),
.A2(n_887),
.B(n_852),
.C(n_927),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_908),
.A2(n_957),
.B(n_900),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_892),
.B(n_915),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_891),
.A2(n_897),
.B(n_949),
.Y(n_1125)
);

NOR2xp67_ASAP7_75t_L g1126 ( 
.A(n_1015),
.B(n_1016),
.Y(n_1126)
);

INVx2_ASAP7_75t_SL g1127 ( 
.A(n_1009),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_951),
.A2(n_912),
.B1(n_873),
.B2(n_1027),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_953),
.A2(n_862),
.B(n_969),
.Y(n_1129)
);

INVxp67_ASAP7_75t_SL g1130 ( 
.A(n_873),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_930),
.B(n_1009),
.Y(n_1131)
);

INVx5_ASAP7_75t_L g1132 ( 
.A(n_951),
.Y(n_1132)
);

BUFx10_ASAP7_75t_L g1133 ( 
.A(n_938),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_930),
.B(n_973),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_969),
.A2(n_921),
.B(n_879),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_868),
.B(n_1026),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_919),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_951),
.A2(n_966),
.B(n_970),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_951),
.B(n_1014),
.Y(n_1139)
);

AOI22x1_ASAP7_75t_L g1140 ( 
.A1(n_999),
.A2(n_1000),
.B1(n_948),
.B2(n_932),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_971),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_1006),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_938),
.B(n_925),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_902),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_971),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_919),
.Y(n_1146)
);

AOI22xp33_ASAP7_75t_L g1147 ( 
.A1(n_995),
.A2(n_1017),
.B1(n_989),
.B2(n_904),
.Y(n_1147)
);

O2A1O1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_1023),
.A2(n_1019),
.B(n_1021),
.C(n_909),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_914),
.Y(n_1149)
);

INVx3_ASAP7_75t_L g1150 ( 
.A(n_965),
.Y(n_1150)
);

BUFx2_ASAP7_75t_L g1151 ( 
.A(n_965),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1007),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_917),
.Y(n_1153)
);

NOR3xp33_ASAP7_75t_SL g1154 ( 
.A(n_1025),
.B(n_1013),
.C(n_918),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_963),
.A2(n_1001),
.B(n_955),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_990),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_990),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_960),
.B(n_1027),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1010),
.B(n_1029),
.Y(n_1159)
);

NAND2x1p5_ASAP7_75t_L g1160 ( 
.A(n_980),
.B(n_985),
.Y(n_1160)
);

INVx1_ASAP7_75t_SL g1161 ( 
.A(n_1008),
.Y(n_1161)
);

CKINVDCx14_ASAP7_75t_R g1162 ( 
.A(n_981),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_866),
.A2(n_997),
.B1(n_977),
.B2(n_962),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1005),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_988),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1011),
.Y(n_1166)
);

BUFx2_ASAP7_75t_L g1167 ( 
.A(n_907),
.Y(n_1167)
);

BUFx3_ASAP7_75t_L g1168 ( 
.A(n_920),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_976),
.B(n_987),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_994),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_851),
.A2(n_631),
.B(n_850),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_851),
.A2(n_631),
.B(n_850),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_875),
.B(n_701),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1020),
.Y(n_1174)
);

AOI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_926),
.A2(n_701),
.B1(n_991),
.B2(n_849),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_937),
.A2(n_701),
.B(n_811),
.C(n_926),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_901),
.B(n_459),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_851),
.A2(n_631),
.B(n_850),
.Y(n_1178)
);

NAND3xp33_ASAP7_75t_L g1179 ( 
.A(n_991),
.B(n_701),
.C(n_926),
.Y(n_1179)
);

INVxp67_ASAP7_75t_L g1180 ( 
.A(n_867),
.Y(n_1180)
);

INVxp33_ASAP7_75t_L g1181 ( 
.A(n_860),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_875),
.A2(n_701),
.B1(n_928),
.B2(n_926),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_875),
.B(n_701),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_937),
.A2(n_701),
.B(n_811),
.C(n_926),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_928),
.B(n_701),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_901),
.B(n_459),
.Y(n_1186)
);

INVx3_ASAP7_75t_L g1187 ( 
.A(n_1146),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1176),
.A2(n_1184),
.B(n_1179),
.C(n_1183),
.Y(n_1188)
);

OAI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1064),
.A2(n_1179),
.B(n_1173),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1102),
.Y(n_1190)
);

OAI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1173),
.A2(n_1183),
.B(n_1185),
.Y(n_1191)
);

AO31x2_ASAP7_75t_L g1192 ( 
.A1(n_1092),
.A2(n_1163),
.A3(n_1128),
.B(n_1122),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_1180),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1171),
.A2(n_1178),
.B(n_1172),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1102),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_SL g1196 ( 
.A(n_1090),
.B(n_1085),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1101),
.A2(n_1082),
.B(n_1125),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1111),
.A2(n_1123),
.B(n_1129),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1083),
.A2(n_1140),
.B(n_1160),
.Y(n_1199)
);

O2A1O1Ixp33_ASAP7_75t_SL g1200 ( 
.A1(n_1049),
.A2(n_1039),
.B(n_1070),
.C(n_1158),
.Y(n_1200)
);

AO31x2_ASAP7_75t_L g1201 ( 
.A1(n_1163),
.A2(n_1128),
.A3(n_1058),
.B(n_1110),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1044),
.A2(n_1117),
.B(n_1132),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1175),
.A2(n_1182),
.B1(n_1131),
.B2(n_1035),
.Y(n_1203)
);

INVxp67_ASAP7_75t_SL g1204 ( 
.A(n_1119),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1038),
.Y(n_1205)
);

A2O1A1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1036),
.A2(n_1034),
.B(n_1108),
.C(n_1113),
.Y(n_1206)
);

AOI221x1_ASAP7_75t_L g1207 ( 
.A1(n_1053),
.A2(n_1048),
.B1(n_1066),
.B2(n_1124),
.C(n_1041),
.Y(n_1207)
);

INVxp67_ASAP7_75t_L g1208 ( 
.A(n_1068),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1045),
.Y(n_1209)
);

O2A1O1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_1182),
.A2(n_1053),
.B(n_1089),
.C(n_1048),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_L g1211 ( 
.A(n_1103),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_1181),
.B(n_1177),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1186),
.B(n_1093),
.Y(n_1213)
);

INVx2_ASAP7_75t_SL g1214 ( 
.A(n_1094),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_1103),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1160),
.A2(n_1118),
.B(n_1155),
.Y(n_1216)
);

AO21x2_ASAP7_75t_L g1217 ( 
.A1(n_1117),
.A2(n_1169),
.B(n_1135),
.Y(n_1217)
);

AO21x1_ASAP7_75t_L g1218 ( 
.A1(n_1120),
.A2(n_1114),
.B(n_1100),
.Y(n_1218)
);

CKINVDCx20_ASAP7_75t_R g1219 ( 
.A(n_1162),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1119),
.Y(n_1220)
);

NOR2x1_ASAP7_75t_L g1221 ( 
.A(n_1095),
.B(n_1033),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1138),
.A2(n_1072),
.B(n_1081),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1104),
.Y(n_1223)
);

AOI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1159),
.A2(n_1167),
.B(n_1105),
.Y(n_1224)
);

AO22x2_ASAP7_75t_L g1225 ( 
.A1(n_1084),
.A2(n_1076),
.B1(n_1065),
.B2(n_1164),
.Y(n_1225)
);

AO31x2_ASAP7_75t_L g1226 ( 
.A1(n_1084),
.A2(n_1165),
.A3(n_1170),
.B(n_1040),
.Y(n_1226)
);

BUFx2_ASAP7_75t_L g1227 ( 
.A(n_1116),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1161),
.B(n_1134),
.Y(n_1228)
);

AOI21xp33_ASAP7_75t_L g1229 ( 
.A1(n_1091),
.A2(n_1142),
.B(n_1098),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1063),
.B(n_1061),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1127),
.B(n_1069),
.Y(n_1231)
);

AO32x2_ASAP7_75t_L g1232 ( 
.A1(n_1109),
.A2(n_1086),
.A3(n_1071),
.B1(n_1062),
.B2(n_1057),
.Y(n_1232)
);

NOR2x1_ASAP7_75t_L g1233 ( 
.A(n_1095),
.B(n_1033),
.Y(n_1233)
);

BUFx3_ASAP7_75t_L g1234 ( 
.A(n_1103),
.Y(n_1234)
);

AOI221xp5_ASAP7_75t_SL g1235 ( 
.A1(n_1077),
.A2(n_1051),
.B1(n_1043),
.B2(n_1046),
.C(n_1059),
.Y(n_1235)
);

NAND3xp33_ASAP7_75t_L g1236 ( 
.A(n_1143),
.B(n_1056),
.C(n_1049),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_1112),
.Y(n_1237)
);

BUFx2_ASAP7_75t_L g1238 ( 
.A(n_1096),
.Y(n_1238)
);

BUFx6f_ASAP7_75t_L g1239 ( 
.A(n_1112),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1132),
.A2(n_1106),
.B(n_1147),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1139),
.A2(n_1132),
.B1(n_1096),
.B2(n_1144),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1166),
.A2(n_1055),
.B(n_1148),
.Y(n_1242)
);

OA21x2_ASAP7_75t_L g1243 ( 
.A1(n_1154),
.A2(n_1136),
.B(n_1149),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1126),
.A2(n_1152),
.B(n_1107),
.Y(n_1244)
);

AOI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1042),
.A2(n_1112),
.B1(n_1050),
.B2(n_1153),
.Y(n_1245)
);

HB1xp67_ASAP7_75t_L g1246 ( 
.A(n_1151),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1074),
.A2(n_1079),
.B(n_1078),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1132),
.A2(n_1168),
.B(n_1057),
.Y(n_1248)
);

AO21x2_ASAP7_75t_L g1249 ( 
.A1(n_1047),
.A2(n_1156),
.B(n_1130),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1054),
.A2(n_1087),
.B(n_1075),
.Y(n_1250)
);

AO31x2_ASAP7_75t_L g1251 ( 
.A1(n_1174),
.A2(n_1153),
.A3(n_1099),
.B(n_1150),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1054),
.A2(n_1087),
.B(n_1075),
.Y(n_1252)
);

INVx5_ASAP7_75t_L g1253 ( 
.A(n_1037),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1153),
.A2(n_1095),
.B1(n_1097),
.B2(n_1073),
.Y(n_1254)
);

BUFx2_ASAP7_75t_SL g1255 ( 
.A(n_1115),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1137),
.B(n_1121),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1157),
.A2(n_1137),
.B(n_1099),
.Y(n_1257)
);

INVx5_ASAP7_75t_L g1258 ( 
.A(n_1037),
.Y(n_1258)
);

OAI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1060),
.A2(n_1067),
.B(n_1145),
.Y(n_1259)
);

AO31x2_ASAP7_75t_L g1260 ( 
.A1(n_1141),
.A2(n_1145),
.A3(n_1060),
.B(n_1067),
.Y(n_1260)
);

AOI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1080),
.A2(n_1115),
.B1(n_1088),
.B2(n_1141),
.Y(n_1261)
);

AND2x2_ASAP7_75t_SL g1262 ( 
.A(n_1052),
.B(n_1141),
.Y(n_1262)
);

AO21x2_ASAP7_75t_L g1263 ( 
.A1(n_1133),
.A2(n_1117),
.B(n_1125),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1171),
.A2(n_701),
.B(n_851),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1171),
.A2(n_701),
.B(n_851),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1171),
.A2(n_701),
.B(n_851),
.Y(n_1266)
);

NOR2xp67_ASAP7_75t_SL g1267 ( 
.A(n_1132),
.B(n_857),
.Y(n_1267)
);

OAI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1064),
.A2(n_701),
.B(n_1176),
.Y(n_1268)
);

INVx3_ASAP7_75t_L g1269 ( 
.A(n_1146),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1101),
.A2(n_886),
.B(n_1082),
.Y(n_1270)
);

AOI221xp5_ASAP7_75t_L g1271 ( 
.A1(n_1036),
.A2(n_811),
.B1(n_459),
.B2(n_937),
.C(n_592),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1171),
.A2(n_701),
.B(n_851),
.Y(n_1272)
);

A2O1A1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1176),
.A2(n_701),
.B(n_1184),
.C(n_1179),
.Y(n_1273)
);

AO32x2_ASAP7_75t_L g1274 ( 
.A1(n_1053),
.A2(n_1084),
.A3(n_1048),
.B1(n_1182),
.B2(n_1163),
.Y(n_1274)
);

OR2x2_ASAP7_75t_L g1275 ( 
.A(n_1177),
.B(n_573),
.Y(n_1275)
);

A2O1A1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_1176),
.A2(n_701),
.B(n_1184),
.C(n_1179),
.Y(n_1276)
);

OR2x2_ASAP7_75t_L g1277 ( 
.A(n_1177),
.B(n_573),
.Y(n_1277)
);

A2O1A1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1176),
.A2(n_701),
.B(n_1184),
.C(n_1179),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1101),
.A2(n_886),
.B(n_1082),
.Y(n_1279)
);

INVxp67_ASAP7_75t_SL g1280 ( 
.A(n_1119),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1102),
.Y(n_1281)
);

A2O1A1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_1176),
.A2(n_701),
.B(n_1184),
.C(n_1179),
.Y(n_1282)
);

AO31x2_ASAP7_75t_L g1283 ( 
.A1(n_1092),
.A2(n_1064),
.A3(n_1163),
.B(n_1128),
.Y(n_1283)
);

AND2x6_ASAP7_75t_L g1284 ( 
.A(n_1157),
.B(n_855),
.Y(n_1284)
);

AOI221xp5_ASAP7_75t_L g1285 ( 
.A1(n_1036),
.A2(n_811),
.B1(n_459),
.B2(n_937),
.C(n_592),
.Y(n_1285)
);

O2A1O1Ixp33_ASAP7_75t_L g1286 ( 
.A1(n_1036),
.A2(n_701),
.B(n_811),
.C(n_783),
.Y(n_1286)
);

O2A1O1Ixp33_ASAP7_75t_L g1287 ( 
.A1(n_1036),
.A2(n_701),
.B(n_811),
.C(n_783),
.Y(n_1287)
);

INVx2_ASAP7_75t_SL g1288 ( 
.A(n_1094),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1102),
.Y(n_1289)
);

A2O1A1Ixp33_ASAP7_75t_L g1290 ( 
.A1(n_1176),
.A2(n_701),
.B(n_1184),
.C(n_1179),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1102),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1171),
.A2(n_701),
.B(n_851),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1171),
.A2(n_701),
.B(n_851),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1175),
.B(n_701),
.Y(n_1294)
);

INVx2_ASAP7_75t_SL g1295 ( 
.A(n_1094),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1171),
.A2(n_701),
.B(n_851),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1171),
.A2(n_701),
.B(n_851),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1064),
.A2(n_701),
.B(n_1176),
.Y(n_1298)
);

AO31x2_ASAP7_75t_L g1299 ( 
.A1(n_1092),
.A2(n_1064),
.A3(n_1163),
.B(n_1128),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1101),
.A2(n_886),
.B(n_1082),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_SL g1301 ( 
.A(n_1175),
.B(n_701),
.Y(n_1301)
);

AOI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1036),
.A2(n_701),
.B1(n_991),
.B2(n_783),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1102),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1102),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1173),
.A2(n_701),
.B1(n_1183),
.B2(n_1185),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1171),
.A2(n_701),
.B(n_851),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1038),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1173),
.B(n_1183),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1038),
.Y(n_1309)
);

O2A1O1Ixp33_ASAP7_75t_L g1310 ( 
.A1(n_1036),
.A2(n_701),
.B(n_811),
.C(n_783),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_1179),
.B(n_701),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1171),
.A2(n_701),
.B(n_851),
.Y(n_1312)
);

AO21x2_ASAP7_75t_L g1313 ( 
.A1(n_1117),
.A2(n_1125),
.B(n_1082),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1173),
.B(n_1183),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1171),
.A2(n_701),
.B(n_851),
.Y(n_1315)
);

A2O1A1Ixp33_ASAP7_75t_L g1316 ( 
.A1(n_1176),
.A2(n_701),
.B(n_1184),
.C(n_1179),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_SL g1317 ( 
.A(n_1175),
.B(n_701),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1173),
.A2(n_701),
.B1(n_1183),
.B2(n_1185),
.Y(n_1318)
);

BUFx8_ASAP7_75t_L g1319 ( 
.A(n_1103),
.Y(n_1319)
);

BUFx2_ASAP7_75t_L g1320 ( 
.A(n_1180),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1101),
.A2(n_886),
.B(n_1082),
.Y(n_1321)
);

NOR2xp67_ASAP7_75t_L g1322 ( 
.A(n_1142),
.B(n_947),
.Y(n_1322)
);

OA21x2_ASAP7_75t_L g1323 ( 
.A1(n_1117),
.A2(n_861),
.B(n_1092),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1173),
.B(n_1183),
.Y(n_1324)
);

NAND3xp33_ASAP7_75t_SL g1325 ( 
.A(n_1036),
.B(n_701),
.C(n_459),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1102),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1177),
.B(n_1186),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1171),
.A2(n_701),
.B(n_851),
.Y(n_1328)
);

OR2x6_ASAP7_75t_L g1329 ( 
.A(n_1088),
.B(n_1103),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_1090),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_SL g1331 ( 
.A1(n_1064),
.A2(n_701),
.B(n_1128),
.Y(n_1331)
);

OR2x2_ASAP7_75t_L g1332 ( 
.A(n_1177),
.B(n_573),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1101),
.A2(n_886),
.B(n_1082),
.Y(n_1333)
);

OAI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1064),
.A2(n_701),
.B(n_1176),
.Y(n_1334)
);

AO31x2_ASAP7_75t_L g1335 ( 
.A1(n_1092),
.A2(n_1064),
.A3(n_1163),
.B(n_1128),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_L g1336 ( 
.A(n_1262),
.Y(n_1336)
);

INVx3_ASAP7_75t_SL g1337 ( 
.A(n_1330),
.Y(n_1337)
);

INVx4_ASAP7_75t_L g1338 ( 
.A(n_1329),
.Y(n_1338)
);

INVx2_ASAP7_75t_R g1339 ( 
.A(n_1190),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1308),
.A2(n_1324),
.B1(n_1314),
.B2(n_1302),
.Y(n_1340)
);

INVx1_ASAP7_75t_SL g1341 ( 
.A(n_1193),
.Y(n_1341)
);

INVx6_ASAP7_75t_L g1342 ( 
.A(n_1319),
.Y(n_1342)
);

BUFx2_ASAP7_75t_L g1343 ( 
.A(n_1227),
.Y(n_1343)
);

BUFx3_ASAP7_75t_L g1344 ( 
.A(n_1319),
.Y(n_1344)
);

BUFx2_ASAP7_75t_L g1345 ( 
.A(n_1320),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_SL g1346 ( 
.A1(n_1311),
.A2(n_1230),
.B1(n_1203),
.B2(n_1268),
.Y(n_1346)
);

OAI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1207),
.A2(n_1285),
.B1(n_1271),
.B2(n_1228),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1305),
.B(n_1318),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1234),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1205),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1307),
.Y(n_1351)
);

INVx1_ASAP7_75t_SL g1352 ( 
.A(n_1213),
.Y(n_1352)
);

OAI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1325),
.A2(n_1191),
.B1(n_1304),
.B2(n_1195),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1190),
.B(n_1195),
.Y(n_1354)
);

AOI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1235),
.A2(n_1219),
.B1(n_1327),
.B2(n_1212),
.Y(n_1355)
);

AOI21xp33_ASAP7_75t_L g1356 ( 
.A1(n_1286),
.A2(n_1310),
.B(n_1287),
.Y(n_1356)
);

BUFx8_ASAP7_75t_L g1357 ( 
.A(n_1211),
.Y(n_1357)
);

BUFx8_ASAP7_75t_SL g1358 ( 
.A(n_1211),
.Y(n_1358)
);

BUFx2_ASAP7_75t_L g1359 ( 
.A(n_1246),
.Y(n_1359)
);

OAI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1281),
.A2(n_1303),
.B1(n_1304),
.B2(n_1289),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1309),
.Y(n_1361)
);

INVx4_ASAP7_75t_L g1362 ( 
.A(n_1329),
.Y(n_1362)
);

NAND2x1p5_ASAP7_75t_L g1363 ( 
.A(n_1267),
.B(n_1221),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_SL g1364 ( 
.A1(n_1298),
.A2(n_1334),
.B1(n_1189),
.B2(n_1225),
.Y(n_1364)
);

AOI22x1_ASAP7_75t_SL g1365 ( 
.A1(n_1281),
.A2(n_1289),
.B1(n_1326),
.B2(n_1303),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_SL g1366 ( 
.A1(n_1225),
.A2(n_1238),
.B1(n_1326),
.B2(n_1291),
.Y(n_1366)
);

BUFx3_ASAP7_75t_L g1367 ( 
.A(n_1215),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1294),
.A2(n_1301),
.B1(n_1317),
.B2(n_1229),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1291),
.A2(n_1208),
.B1(n_1236),
.B2(n_1332),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1218),
.A2(n_1204),
.B1(n_1280),
.B2(n_1220),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1275),
.A2(n_1277),
.B1(n_1322),
.B2(n_1206),
.Y(n_1371)
);

INVx6_ASAP7_75t_L g1372 ( 
.A(n_1253),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1231),
.B(n_1223),
.Y(n_1373)
);

CKINVDCx20_ASAP7_75t_R g1374 ( 
.A(n_1261),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1331),
.A2(n_1245),
.B1(n_1188),
.B2(n_1273),
.Y(n_1375)
);

CKINVDCx16_ASAP7_75t_R g1376 ( 
.A(n_1196),
.Y(n_1376)
);

BUFx10_ASAP7_75t_L g1377 ( 
.A(n_1215),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1323),
.A2(n_1217),
.B1(n_1243),
.B2(n_1241),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1276),
.B(n_1278),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1251),
.Y(n_1380)
);

BUFx6f_ASAP7_75t_L g1381 ( 
.A(n_1253),
.Y(n_1381)
);

INVx1_ASAP7_75t_SL g1382 ( 
.A(n_1214),
.Y(n_1382)
);

OAI22xp33_ASAP7_75t_SL g1383 ( 
.A1(n_1240),
.A2(n_1254),
.B1(n_1224),
.B2(n_1244),
.Y(n_1383)
);

BUFx8_ASAP7_75t_L g1384 ( 
.A(n_1237),
.Y(n_1384)
);

NAND2x1p5_ASAP7_75t_L g1385 ( 
.A(n_1233),
.B(n_1258),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1226),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_1288),
.Y(n_1387)
);

INVx6_ASAP7_75t_L g1388 ( 
.A(n_1258),
.Y(n_1388)
);

BUFx4f_ASAP7_75t_SL g1389 ( 
.A(n_1237),
.Y(n_1389)
);

AOI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1295),
.A2(n_1200),
.B1(n_1316),
.B2(n_1290),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1260),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1260),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1260),
.Y(n_1393)
);

OAI22xp33_ASAP7_75t_SL g1394 ( 
.A1(n_1210),
.A2(n_1274),
.B1(n_1328),
.B2(n_1315),
.Y(n_1394)
);

AOI22x1_ASAP7_75t_SL g1395 ( 
.A1(n_1187),
.A2(n_1269),
.B1(n_1255),
.B2(n_1274),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_SL g1396 ( 
.A1(n_1274),
.A2(n_1293),
.B1(n_1264),
.B2(n_1265),
.Y(n_1396)
);

INVx3_ASAP7_75t_SL g1397 ( 
.A(n_1237),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1239),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_SL g1399 ( 
.A1(n_1266),
.A2(n_1292),
.B1(n_1296),
.B2(n_1272),
.Y(n_1399)
);

BUFx10_ASAP7_75t_L g1400 ( 
.A(n_1239),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_SL g1401 ( 
.A1(n_1297),
.A2(n_1312),
.B1(n_1306),
.B2(n_1263),
.Y(n_1401)
);

CKINVDCx8_ASAP7_75t_R g1402 ( 
.A(n_1239),
.Y(n_1402)
);

BUFx12f_ASAP7_75t_L g1403 ( 
.A(n_1284),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1263),
.A2(n_1313),
.B1(n_1202),
.B2(n_1249),
.Y(n_1404)
);

OAI21xp33_ASAP7_75t_L g1405 ( 
.A1(n_1282),
.A2(n_1256),
.B(n_1259),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1313),
.A2(n_1249),
.B1(n_1247),
.B2(n_1248),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1226),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1284),
.A2(n_1194),
.B1(n_1257),
.B2(n_1242),
.Y(n_1408)
);

CKINVDCx11_ASAP7_75t_R g1409 ( 
.A(n_1232),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1198),
.A2(n_1216),
.B1(n_1192),
.B2(n_1199),
.Y(n_1410)
);

CKINVDCx11_ASAP7_75t_R g1411 ( 
.A(n_1232),
.Y(n_1411)
);

CKINVDCx11_ASAP7_75t_R g1412 ( 
.A(n_1232),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1250),
.A2(n_1252),
.B1(n_1335),
.B2(n_1299),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1283),
.A2(n_1299),
.B1(n_1335),
.B2(n_1201),
.Y(n_1414)
);

CKINVDCx20_ASAP7_75t_R g1415 ( 
.A(n_1283),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1201),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1283),
.Y(n_1417)
);

BUFx3_ASAP7_75t_L g1418 ( 
.A(n_1222),
.Y(n_1418)
);

BUFx8_ASAP7_75t_L g1419 ( 
.A(n_1299),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1335),
.A2(n_1197),
.B1(n_1270),
.B2(n_1279),
.Y(n_1420)
);

NAND2x1p5_ASAP7_75t_L g1421 ( 
.A(n_1300),
.B(n_1321),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1333),
.A2(n_1271),
.B1(n_1285),
.B2(n_701),
.Y(n_1422)
);

INVx1_ASAP7_75t_SL g1423 ( 
.A(n_1193),
.Y(n_1423)
);

INVxp33_ASAP7_75t_L g1424 ( 
.A(n_1212),
.Y(n_1424)
);

CKINVDCx20_ASAP7_75t_R g1425 ( 
.A(n_1330),
.Y(n_1425)
);

INVx5_ASAP7_75t_L g1426 ( 
.A(n_1284),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1209),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1271),
.A2(n_1285),
.B1(n_701),
.B2(n_1036),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1209),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1220),
.Y(n_1430)
);

BUFx3_ASAP7_75t_L g1431 ( 
.A(n_1319),
.Y(n_1431)
);

BUFx4f_ASAP7_75t_SL g1432 ( 
.A(n_1319),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1209),
.Y(n_1433)
);

BUFx12f_ASAP7_75t_L g1434 ( 
.A(n_1319),
.Y(n_1434)
);

BUFx3_ASAP7_75t_L g1435 ( 
.A(n_1319),
.Y(n_1435)
);

INVx6_ASAP7_75t_L g1436 ( 
.A(n_1319),
.Y(n_1436)
);

CKINVDCx20_ASAP7_75t_R g1437 ( 
.A(n_1330),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1271),
.A2(n_1285),
.B1(n_701),
.B2(n_1036),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1308),
.A2(n_701),
.B1(n_1324),
.B2(n_1314),
.Y(n_1439)
);

INVx2_ASAP7_75t_SL g1440 ( 
.A(n_1319),
.Y(n_1440)
);

BUFx12f_ASAP7_75t_L g1441 ( 
.A(n_1319),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1271),
.A2(n_1285),
.B1(n_701),
.B2(n_1036),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1271),
.A2(n_1285),
.B1(n_701),
.B2(n_1036),
.Y(n_1443)
);

CKINVDCx11_ASAP7_75t_R g1444 ( 
.A(n_1219),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1209),
.Y(n_1445)
);

AOI21xp33_ASAP7_75t_L g1446 ( 
.A1(n_1302),
.A2(n_701),
.B(n_1286),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1271),
.A2(n_1285),
.B1(n_701),
.B2(n_1036),
.Y(n_1447)
);

BUFx12f_ASAP7_75t_L g1448 ( 
.A(n_1319),
.Y(n_1448)
);

INVx2_ASAP7_75t_SL g1449 ( 
.A(n_1319),
.Y(n_1449)
);

INVx3_ASAP7_75t_SL g1450 ( 
.A(n_1330),
.Y(n_1450)
);

CKINVDCx11_ASAP7_75t_R g1451 ( 
.A(n_1219),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1308),
.A2(n_701),
.B1(n_1324),
.B2(n_1314),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1308),
.A2(n_701),
.B1(n_1324),
.B2(n_1314),
.Y(n_1453)
);

OAI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1302),
.A2(n_701),
.B1(n_649),
.B2(n_1308),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_1444),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1415),
.B(n_1417),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1421),
.A2(n_1406),
.B(n_1410),
.Y(n_1457)
);

INVx2_ASAP7_75t_SL g1458 ( 
.A(n_1372),
.Y(n_1458)
);

INVx3_ASAP7_75t_L g1459 ( 
.A(n_1380),
.Y(n_1459)
);

BUFx2_ASAP7_75t_L g1460 ( 
.A(n_1419),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1364),
.B(n_1366),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1407),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1359),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1430),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1424),
.B(n_1352),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1386),
.Y(n_1466)
);

OAI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1421),
.A2(n_1406),
.B(n_1410),
.Y(n_1467)
);

AND2x4_ASAP7_75t_L g1468 ( 
.A(n_1350),
.B(n_1351),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1430),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1420),
.A2(n_1408),
.B(n_1404),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1386),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1391),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1361),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1392),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1393),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1414),
.B(n_1416),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1339),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1339),
.Y(n_1478)
);

BUFx3_ASAP7_75t_L g1479 ( 
.A(n_1357),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1428),
.A2(n_1438),
.B1(n_1447),
.B2(n_1442),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1428),
.A2(n_1438),
.B1(n_1447),
.B2(n_1442),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1360),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1360),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1354),
.Y(n_1484)
);

BUFx2_ASAP7_75t_L g1485 ( 
.A(n_1419),
.Y(n_1485)
);

NAND2x1_ASAP7_75t_L g1486 ( 
.A(n_1390),
.B(n_1408),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1379),
.Y(n_1487)
);

NAND2x1_ASAP7_75t_L g1488 ( 
.A(n_1375),
.B(n_1413),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1348),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1420),
.A2(n_1404),
.B(n_1413),
.Y(n_1490)
);

INVxp67_ASAP7_75t_L g1491 ( 
.A(n_1345),
.Y(n_1491)
);

AO21x2_ASAP7_75t_L g1492 ( 
.A1(n_1353),
.A2(n_1356),
.B(n_1446),
.Y(n_1492)
);

OR2x6_ASAP7_75t_L g1493 ( 
.A(n_1418),
.B(n_1363),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1394),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1427),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1429),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1433),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1378),
.A2(n_1368),
.B(n_1422),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1445),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1370),
.B(n_1353),
.Y(n_1500)
);

OAI22x1_ASAP7_75t_L g1501 ( 
.A1(n_1355),
.A2(n_1412),
.B1(n_1411),
.B2(n_1409),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1366),
.Y(n_1502)
);

AOI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1340),
.A2(n_1369),
.B(n_1453),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1365),
.Y(n_1504)
);

BUFx6f_ASAP7_75t_L g1505 ( 
.A(n_1426),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1370),
.B(n_1378),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1346),
.B(n_1422),
.Y(n_1507)
);

BUFx2_ASAP7_75t_L g1508 ( 
.A(n_1343),
.Y(n_1508)
);

CKINVDCx6p67_ASAP7_75t_R g1509 ( 
.A(n_1337),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1443),
.A2(n_1454),
.B1(n_1347),
.B2(n_1346),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1395),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1439),
.B(n_1452),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1383),
.Y(n_1513)
);

OR2x6_ASAP7_75t_L g1514 ( 
.A(n_1363),
.B(n_1342),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1396),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1373),
.Y(n_1516)
);

OR2x6_ASAP7_75t_SL g1517 ( 
.A(n_1371),
.B(n_1387),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1454),
.B(n_1347),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1405),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1401),
.Y(n_1520)
);

AOI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1399),
.A2(n_1443),
.B(n_1426),
.Y(n_1521)
);

BUFx3_ASAP7_75t_L g1522 ( 
.A(n_1357),
.Y(n_1522)
);

INVx2_ASAP7_75t_SL g1523 ( 
.A(n_1372),
.Y(n_1523)
);

INVxp33_ASAP7_75t_L g1524 ( 
.A(n_1451),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1341),
.B(n_1423),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1336),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1385),
.Y(n_1527)
);

BUFx2_ASAP7_75t_SL g1528 ( 
.A(n_1381),
.Y(n_1528)
);

BUFx3_ASAP7_75t_L g1529 ( 
.A(n_1384),
.Y(n_1529)
);

INVxp67_ASAP7_75t_L g1530 ( 
.A(n_1382),
.Y(n_1530)
);

INVx3_ASAP7_75t_L g1531 ( 
.A(n_1403),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1376),
.B(n_1374),
.Y(n_1532)
);

INVx1_ASAP7_75t_SL g1533 ( 
.A(n_1349),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1338),
.B(n_1362),
.Y(n_1534)
);

BUFx3_ASAP7_75t_L g1535 ( 
.A(n_1384),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1397),
.B(n_1338),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1362),
.B(n_1398),
.Y(n_1537)
);

BUFx2_ASAP7_75t_L g1538 ( 
.A(n_1508),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1466),
.Y(n_1539)
);

OAI21xp5_ASAP7_75t_L g1540 ( 
.A1(n_1510),
.A2(n_1440),
.B(n_1449),
.Y(n_1540)
);

OR2x6_ASAP7_75t_L g1541 ( 
.A(n_1488),
.B(n_1342),
.Y(n_1541)
);

NAND3xp33_ASAP7_75t_L g1542 ( 
.A(n_1480),
.B(n_1402),
.C(n_1367),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1456),
.B(n_1337),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1489),
.B(n_1450),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1493),
.B(n_1468),
.Y(n_1545)
);

OAI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1481),
.A2(n_1437),
.B(n_1425),
.Y(n_1546)
);

AOI21xp5_ASAP7_75t_L g1547 ( 
.A1(n_1521),
.A2(n_1388),
.B(n_1344),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1473),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1519),
.B(n_1342),
.Y(n_1549)
);

A2O1A1Ixp33_ASAP7_75t_SL g1550 ( 
.A1(n_1513),
.A2(n_1389),
.B(n_1388),
.C(n_1432),
.Y(n_1550)
);

AND2x4_ASAP7_75t_L g1551 ( 
.A(n_1493),
.B(n_1431),
.Y(n_1551)
);

A2O1A1Ixp33_ASAP7_75t_L g1552 ( 
.A1(n_1486),
.A2(n_1435),
.B(n_1389),
.C(n_1436),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1507),
.A2(n_1436),
.B1(n_1448),
.B2(n_1434),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_L g1554 ( 
.A(n_1519),
.B(n_1432),
.Y(n_1554)
);

A2O1A1Ixp33_ASAP7_75t_L g1555 ( 
.A1(n_1486),
.A2(n_1358),
.B(n_1441),
.C(n_1400),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1512),
.B(n_1377),
.Y(n_1556)
);

OA21x2_ASAP7_75t_L g1557 ( 
.A1(n_1490),
.A2(n_1470),
.B(n_1498),
.Y(n_1557)
);

AND2x4_ASAP7_75t_L g1558 ( 
.A(n_1493),
.B(n_1468),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1526),
.B(n_1516),
.Y(n_1559)
);

NOR2x1_ASAP7_75t_SL g1560 ( 
.A(n_1514),
.B(n_1503),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1464),
.B(n_1494),
.Y(n_1561)
);

BUFx2_ASAP7_75t_L g1562 ( 
.A(n_1508),
.Y(n_1562)
);

AND2x4_ASAP7_75t_L g1563 ( 
.A(n_1477),
.B(n_1478),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1464),
.B(n_1494),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1517),
.B(n_1518),
.Y(n_1565)
);

O2A1O1Ixp33_ASAP7_75t_SL g1566 ( 
.A1(n_1518),
.A2(n_1504),
.B(n_1511),
.C(n_1500),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1469),
.B(n_1513),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1517),
.B(n_1504),
.Y(n_1568)
);

OAI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1503),
.A2(n_1507),
.B(n_1500),
.Y(n_1569)
);

A2O1A1Ixp33_ASAP7_75t_L g1570 ( 
.A1(n_1461),
.A2(n_1498),
.B(n_1506),
.C(n_1515),
.Y(n_1570)
);

OAI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1461),
.A2(n_1485),
.B1(n_1460),
.B2(n_1530),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_L g1572 ( 
.A(n_1487),
.B(n_1502),
.Y(n_1572)
);

OA21x2_ASAP7_75t_L g1573 ( 
.A1(n_1490),
.A2(n_1470),
.B(n_1457),
.Y(n_1573)
);

AOI221xp5_ASAP7_75t_L g1574 ( 
.A1(n_1501),
.A2(n_1492),
.B1(n_1520),
.B2(n_1502),
.C(n_1515),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1477),
.B(n_1478),
.Y(n_1575)
);

NOR2xp67_ASAP7_75t_L g1576 ( 
.A(n_1531),
.B(n_1534),
.Y(n_1576)
);

OA21x2_ASAP7_75t_L g1577 ( 
.A1(n_1457),
.A2(n_1467),
.B(n_1520),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_1487),
.B(n_1492),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1463),
.B(n_1460),
.Y(n_1579)
);

A2O1A1Ixp33_ASAP7_75t_L g1580 ( 
.A1(n_1506),
.A2(n_1483),
.B(n_1482),
.C(n_1484),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1501),
.A2(n_1465),
.B1(n_1525),
.B2(n_1483),
.Y(n_1581)
);

OAI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1532),
.A2(n_1491),
.B(n_1527),
.Y(n_1582)
);

A2O1A1Ixp33_ASAP7_75t_L g1583 ( 
.A1(n_1482),
.A2(n_1484),
.B(n_1505),
.C(n_1476),
.Y(n_1583)
);

INVx2_ASAP7_75t_SL g1584 ( 
.A(n_1525),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1496),
.B(n_1497),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1557),
.B(n_1462),
.Y(n_1586)
);

BUFx2_ASAP7_75t_L g1587 ( 
.A(n_1563),
.Y(n_1587)
);

NOR2xp67_ASAP7_75t_L g1588 ( 
.A(n_1578),
.B(n_1495),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1539),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1561),
.B(n_1564),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1567),
.B(n_1476),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1548),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1557),
.B(n_1472),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1573),
.B(n_1474),
.Y(n_1594)
);

INVx3_ASAP7_75t_L g1595 ( 
.A(n_1573),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1577),
.B(n_1471),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1578),
.B(n_1471),
.Y(n_1597)
);

BUFx3_ASAP7_75t_L g1598 ( 
.A(n_1541),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1577),
.B(n_1475),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1575),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_1538),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1585),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1575),
.Y(n_1603)
);

INVx3_ASAP7_75t_L g1604 ( 
.A(n_1545),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1565),
.B(n_1534),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1570),
.B(n_1562),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1570),
.B(n_1459),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1569),
.B(n_1499),
.Y(n_1608)
);

NAND4xp25_ASAP7_75t_SL g1609 ( 
.A(n_1606),
.B(n_1581),
.C(n_1574),
.D(n_1546),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1597),
.B(n_1584),
.Y(n_1610)
);

BUFx2_ASAP7_75t_L g1611 ( 
.A(n_1586),
.Y(n_1611)
);

BUFx3_ASAP7_75t_L g1612 ( 
.A(n_1598),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1600),
.B(n_1545),
.Y(n_1613)
);

BUFx3_ASAP7_75t_L g1614 ( 
.A(n_1598),
.Y(n_1614)
);

AOI31xp33_ASAP7_75t_L g1615 ( 
.A1(n_1606),
.A2(n_1581),
.A3(n_1565),
.B(n_1553),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1594),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1592),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1592),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1597),
.B(n_1580),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1602),
.B(n_1580),
.Y(n_1620)
);

HB1xp67_ASAP7_75t_L g1621 ( 
.A(n_1589),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1594),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1606),
.A2(n_1542),
.B1(n_1583),
.B2(n_1553),
.Y(n_1623)
);

AND2x2_ASAP7_75t_SL g1624 ( 
.A(n_1607),
.B(n_1558),
.Y(n_1624)
);

BUFx2_ASAP7_75t_L g1625 ( 
.A(n_1586),
.Y(n_1625)
);

BUFx2_ASAP7_75t_L g1626 ( 
.A(n_1586),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1602),
.B(n_1572),
.Y(n_1627)
);

INVxp67_ASAP7_75t_L g1628 ( 
.A(n_1589),
.Y(n_1628)
);

AND2x4_ASAP7_75t_L g1629 ( 
.A(n_1604),
.B(n_1558),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1596),
.B(n_1559),
.Y(n_1630)
);

OAI221xp5_ASAP7_75t_L g1631 ( 
.A1(n_1608),
.A2(n_1540),
.B1(n_1555),
.B2(n_1544),
.C(n_1568),
.Y(n_1631)
);

INVx3_ASAP7_75t_L g1632 ( 
.A(n_1595),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1600),
.B(n_1558),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1603),
.B(n_1560),
.Y(n_1634)
);

AOI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1605),
.A2(n_1568),
.B1(n_1571),
.B2(n_1566),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1586),
.B(n_1593),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1596),
.B(n_1591),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1587),
.B(n_1583),
.Y(n_1638)
);

BUFx2_ASAP7_75t_L g1639 ( 
.A(n_1593),
.Y(n_1639)
);

BUFx2_ASAP7_75t_L g1640 ( 
.A(n_1624),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1621),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1616),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1619),
.B(n_1590),
.Y(n_1643)
);

INVx1_ASAP7_75t_SL g1644 ( 
.A(n_1620),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1619),
.B(n_1590),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1636),
.B(n_1611),
.Y(n_1646)
);

INVx2_ASAP7_75t_SL g1647 ( 
.A(n_1624),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1619),
.B(n_1590),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1621),
.Y(n_1649)
);

NAND2x1p5_ASAP7_75t_L g1650 ( 
.A(n_1624),
.B(n_1598),
.Y(n_1650)
);

INVx3_ASAP7_75t_L g1651 ( 
.A(n_1632),
.Y(n_1651)
);

HB1xp67_ASAP7_75t_L g1652 ( 
.A(n_1628),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1628),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1636),
.B(n_1607),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1629),
.B(n_1599),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1637),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1636),
.B(n_1607),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1616),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1611),
.B(n_1607),
.Y(n_1659)
);

AND2x4_ASAP7_75t_L g1660 ( 
.A(n_1629),
.B(n_1599),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1620),
.B(n_1602),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1637),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1627),
.B(n_1608),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1637),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1627),
.B(n_1588),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1610),
.B(n_1588),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1617),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1617),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1611),
.B(n_1599),
.Y(n_1669)
);

AND2x4_ASAP7_75t_SL g1670 ( 
.A(n_1638),
.B(n_1551),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1617),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1610),
.B(n_1588),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1616),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1616),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1618),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1652),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1644),
.B(n_1605),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1640),
.B(n_1624),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1652),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1644),
.B(n_1630),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1653),
.Y(n_1681)
);

AOI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1640),
.A2(n_1609),
.B1(n_1623),
.B2(n_1635),
.Y(n_1682)
);

INVx2_ASAP7_75t_SL g1683 ( 
.A(n_1650),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1653),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1647),
.B(n_1638),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1641),
.Y(n_1686)
);

NAND2x1p5_ASAP7_75t_L g1687 ( 
.A(n_1647),
.B(n_1612),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1641),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1663),
.B(n_1610),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1663),
.B(n_1635),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1643),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1649),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1643),
.B(n_1630),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1661),
.B(n_1635),
.Y(n_1694)
);

INVx2_ASAP7_75t_SL g1695 ( 
.A(n_1650),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1647),
.B(n_1638),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1650),
.B(n_1613),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1650),
.B(n_1613),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1670),
.B(n_1613),
.Y(n_1699)
);

INVxp67_ASAP7_75t_SL g1700 ( 
.A(n_1661),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1670),
.B(n_1633),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1670),
.B(n_1633),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1645),
.B(n_1630),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1649),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1645),
.B(n_1622),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1667),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1648),
.Y(n_1707)
);

BUFx2_ASAP7_75t_L g1708 ( 
.A(n_1646),
.Y(n_1708)
);

OAI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1648),
.A2(n_1631),
.B1(n_1615),
.B2(n_1623),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1667),
.Y(n_1710)
);

HB1xp67_ASAP7_75t_L g1711 ( 
.A(n_1659),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1646),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1668),
.Y(n_1713)
);

INVxp67_ASAP7_75t_L g1714 ( 
.A(n_1666),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1668),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1654),
.B(n_1633),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1665),
.B(n_1615),
.Y(n_1717)
);

AOI32xp33_ASAP7_75t_L g1718 ( 
.A1(n_1659),
.A2(n_1631),
.A3(n_1634),
.B1(n_1609),
.B2(n_1614),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1676),
.Y(n_1719)
);

HB1xp67_ASAP7_75t_L g1720 ( 
.A(n_1708),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1678),
.B(n_1654),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1690),
.B(n_1665),
.Y(n_1722)
);

NOR2xp67_ASAP7_75t_L g1723 ( 
.A(n_1678),
.B(n_1659),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1706),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1708),
.B(n_1699),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1694),
.B(n_1666),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1716),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1676),
.Y(n_1728)
);

OAI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1682),
.A2(n_1552),
.B1(n_1555),
.B2(n_1612),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1706),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1716),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1680),
.B(n_1656),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1710),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1692),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1709),
.B(n_1524),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1677),
.B(n_1672),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1699),
.B(n_1701),
.Y(n_1737)
);

INVxp67_ASAP7_75t_L g1738 ( 
.A(n_1679),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1701),
.B(n_1702),
.Y(n_1739)
);

NAND3xp33_ASAP7_75t_L g1740 ( 
.A(n_1718),
.B(n_1556),
.C(n_1547),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1680),
.B(n_1656),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1702),
.B(n_1654),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1689),
.B(n_1662),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1681),
.B(n_1662),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1685),
.B(n_1657),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1717),
.B(n_1672),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1710),
.Y(n_1747)
);

INVx1_ASAP7_75t_SL g1748 ( 
.A(n_1691),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1684),
.B(n_1657),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1700),
.B(n_1657),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1711),
.B(n_1664),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1707),
.B(n_1664),
.Y(n_1752)
);

INVx1_ASAP7_75t_SL g1753 ( 
.A(n_1685),
.Y(n_1753)
);

OAI322xp33_ASAP7_75t_L g1754 ( 
.A1(n_1714),
.A2(n_1712),
.A3(n_1693),
.B1(n_1703),
.B2(n_1688),
.C1(n_1704),
.C2(n_1686),
.Y(n_1754)
);

OAI21xp33_ASAP7_75t_L g1755 ( 
.A1(n_1726),
.A2(n_1696),
.B(n_1695),
.Y(n_1755)
);

AOI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1740),
.A2(n_1683),
.B1(n_1695),
.B2(n_1696),
.Y(n_1756)
);

AOI211x1_ASAP7_75t_L g1757 ( 
.A1(n_1729),
.A2(n_1698),
.B(n_1697),
.C(n_1646),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1720),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1724),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1748),
.B(n_1692),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1738),
.B(n_1722),
.Y(n_1761)
);

INVx1_ASAP7_75t_SL g1762 ( 
.A(n_1725),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1724),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1735),
.B(n_1712),
.Y(n_1764)
);

NOR2xp33_ASAP7_75t_L g1765 ( 
.A(n_1754),
.B(n_1455),
.Y(n_1765)
);

AOI21xp33_ASAP7_75t_L g1766 ( 
.A1(n_1746),
.A2(n_1753),
.B(n_1736),
.Y(n_1766)
);

OAI21xp5_ASAP7_75t_L g1767 ( 
.A1(n_1723),
.A2(n_1687),
.B(n_1683),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1725),
.B(n_1693),
.Y(n_1768)
);

AOI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1737),
.A2(n_1697),
.B1(n_1698),
.B2(n_1687),
.Y(n_1769)
);

INVxp33_ASAP7_75t_L g1770 ( 
.A(n_1737),
.Y(n_1770)
);

NOR2xp33_ASAP7_75t_R g1771 ( 
.A(n_1719),
.B(n_1455),
.Y(n_1771)
);

INVxp67_ASAP7_75t_SL g1772 ( 
.A(n_1730),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1721),
.B(n_1703),
.Y(n_1773)
);

AOI32xp33_ASAP7_75t_L g1774 ( 
.A1(n_1739),
.A2(n_1669),
.A3(n_1614),
.B1(n_1612),
.B2(n_1634),
.Y(n_1774)
);

OAI32xp33_ASAP7_75t_SL g1775 ( 
.A1(n_1749),
.A2(n_1687),
.A3(n_1705),
.B1(n_1625),
.B2(n_1639),
.Y(n_1775)
);

INVx1_ASAP7_75t_SL g1776 ( 
.A(n_1739),
.Y(n_1776)
);

AOI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1721),
.A2(n_1612),
.B1(n_1614),
.B2(n_1556),
.Y(n_1777)
);

OAI322xp33_ASAP7_75t_L g1778 ( 
.A1(n_1728),
.A2(n_1705),
.A3(n_1715),
.B1(n_1713),
.B2(n_1642),
.C1(n_1674),
.C2(n_1673),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1730),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_SL g1780 ( 
.A(n_1750),
.B(n_1614),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1772),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1768),
.B(n_1743),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1772),
.Y(n_1783)
);

NOR2xp33_ASAP7_75t_L g1784 ( 
.A(n_1765),
.B(n_1509),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1762),
.B(n_1745),
.Y(n_1785)
);

O2A1O1Ixp33_ASAP7_75t_L g1786 ( 
.A1(n_1765),
.A2(n_1734),
.B(n_1752),
.C(n_1744),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1759),
.Y(n_1787)
);

OAI22xp33_ASAP7_75t_L g1788 ( 
.A1(n_1756),
.A2(n_1727),
.B1(n_1731),
.B2(n_1601),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1763),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1776),
.B(n_1745),
.Y(n_1790)
);

INVxp67_ASAP7_75t_L g1791 ( 
.A(n_1758),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1779),
.Y(n_1792)
);

NOR2xp33_ASAP7_75t_SL g1793 ( 
.A(n_1766),
.B(n_1509),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1760),
.Y(n_1794)
);

OAI21xp33_ASAP7_75t_L g1795 ( 
.A1(n_1770),
.A2(n_1731),
.B(n_1727),
.Y(n_1795)
);

OAI32xp33_ASAP7_75t_L g1796 ( 
.A1(n_1775),
.A2(n_1751),
.A3(n_1732),
.B1(n_1741),
.B2(n_1744),
.Y(n_1796)
);

AOI21xp33_ASAP7_75t_L g1797 ( 
.A1(n_1761),
.A2(n_1741),
.B(n_1732),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1771),
.B(n_1742),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1757),
.B(n_1742),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1769),
.B(n_1743),
.Y(n_1800)
);

OAI21xp33_ASAP7_75t_L g1801 ( 
.A1(n_1793),
.A2(n_1755),
.B(n_1764),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1791),
.B(n_1773),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1781),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1783),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1798),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1785),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1791),
.B(n_1780),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1790),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1800),
.B(n_1767),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1786),
.B(n_1794),
.Y(n_1810)
);

INVxp67_ASAP7_75t_L g1811 ( 
.A(n_1784),
.Y(n_1811)
);

NAND3xp33_ASAP7_75t_SL g1812 ( 
.A(n_1784),
.B(n_1774),
.C(n_1777),
.Y(n_1812)
);

AOI21xp5_ASAP7_75t_L g1813 ( 
.A1(n_1810),
.A2(n_1788),
.B(n_1797),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1805),
.B(n_1808),
.Y(n_1814)
);

NOR2xp67_ASAP7_75t_L g1815 ( 
.A(n_1805),
.B(n_1782),
.Y(n_1815)
);

OAI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1811),
.A2(n_1788),
.B(n_1795),
.Y(n_1816)
);

NOR3x1_ASAP7_75t_L g1817 ( 
.A(n_1807),
.B(n_1799),
.C(n_1789),
.Y(n_1817)
);

OR2x2_ASAP7_75t_L g1818 ( 
.A(n_1808),
.B(n_1787),
.Y(n_1818)
);

INVxp67_ASAP7_75t_L g1819 ( 
.A(n_1809),
.Y(n_1819)
);

NAND2xp33_ASAP7_75t_SL g1820 ( 
.A(n_1802),
.B(n_1792),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1811),
.B(n_1796),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1803),
.Y(n_1822)
);

AOI221xp5_ASAP7_75t_L g1823 ( 
.A1(n_1813),
.A2(n_1801),
.B1(n_1812),
.B2(n_1804),
.C(n_1806),
.Y(n_1823)
);

OAI211xp5_ASAP7_75t_SL g1824 ( 
.A1(n_1816),
.A2(n_1747),
.B(n_1733),
.C(n_1533),
.Y(n_1824)
);

O2A1O1Ixp33_ASAP7_75t_SL g1825 ( 
.A1(n_1822),
.A2(n_1733),
.B(n_1747),
.C(n_1751),
.Y(n_1825)
);

OAI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1815),
.A2(n_1554),
.B(n_1552),
.Y(n_1826)
);

AOI221xp5_ASAP7_75t_L g1827 ( 
.A1(n_1821),
.A2(n_1778),
.B1(n_1715),
.B2(n_1713),
.C(n_1554),
.Y(n_1827)
);

OAI211xp5_ASAP7_75t_SL g1828 ( 
.A1(n_1819),
.A2(n_1543),
.B(n_1531),
.C(n_1582),
.Y(n_1828)
);

AOI221xp5_ASAP7_75t_L g1829 ( 
.A1(n_1823),
.A2(n_1820),
.B1(n_1814),
.B2(n_1818),
.C(n_1817),
.Y(n_1829)
);

AOI222xp33_ASAP7_75t_L g1830 ( 
.A1(n_1827),
.A2(n_1669),
.B1(n_1625),
.B2(n_1626),
.C1(n_1639),
.C2(n_1579),
.Y(n_1830)
);

OAI221xp5_ASAP7_75t_L g1831 ( 
.A1(n_1826),
.A2(n_1550),
.B1(n_1531),
.B2(n_1529),
.C(n_1535),
.Y(n_1831)
);

AOI21xp5_ASAP7_75t_SL g1832 ( 
.A1(n_1825),
.A2(n_1522),
.B(n_1479),
.Y(n_1832)
);

A2O1A1Ixp33_ASAP7_75t_L g1833 ( 
.A1(n_1824),
.A2(n_1479),
.B(n_1529),
.C(n_1522),
.Y(n_1833)
);

OAI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1828),
.A2(n_1601),
.B1(n_1669),
.B2(n_1625),
.Y(n_1834)
);

HB1xp67_ASAP7_75t_L g1835 ( 
.A(n_1829),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1834),
.B(n_1833),
.Y(n_1836)
);

NAND4xp75_ASAP7_75t_L g1837 ( 
.A(n_1832),
.B(n_1549),
.C(n_1536),
.D(n_1576),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1830),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1831),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1835),
.Y(n_1840)
);

XNOR2xp5_ASAP7_75t_L g1841 ( 
.A(n_1835),
.B(n_1838),
.Y(n_1841)
);

AOI221x1_ASAP7_75t_L g1842 ( 
.A1(n_1839),
.A2(n_1651),
.B1(n_1549),
.B2(n_1675),
.C(n_1671),
.Y(n_1842)
);

XNOR2xp5_ASAP7_75t_L g1843 ( 
.A(n_1841),
.B(n_1836),
.Y(n_1843)
);

INVxp67_ASAP7_75t_L g1844 ( 
.A(n_1843),
.Y(n_1844)
);

OAI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1844),
.A2(n_1840),
.B1(n_1837),
.B2(n_1842),
.Y(n_1845)
);

OAI22xp5_ASAP7_75t_SL g1846 ( 
.A1(n_1844),
.A2(n_1535),
.B1(n_1528),
.B2(n_1523),
.Y(n_1846)
);

AOI22xp5_ASAP7_75t_L g1847 ( 
.A1(n_1845),
.A2(n_1651),
.B1(n_1660),
.B2(n_1655),
.Y(n_1847)
);

INVxp67_ASAP7_75t_SL g1848 ( 
.A(n_1846),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1848),
.Y(n_1849)
);

AOI31xp33_ASAP7_75t_L g1850 ( 
.A1(n_1849),
.A2(n_1847),
.A3(n_1458),
.B(n_1523),
.Y(n_1850)
);

OA21x2_ASAP7_75t_L g1851 ( 
.A1(n_1850),
.A2(n_1658),
.B(n_1642),
.Y(n_1851)
);

INVxp67_ASAP7_75t_L g1852 ( 
.A(n_1851),
.Y(n_1852)
);

AOI221xp5_ASAP7_75t_L g1853 ( 
.A1(n_1852),
.A2(n_1651),
.B1(n_1675),
.B2(n_1671),
.C(n_1673),
.Y(n_1853)
);

AOI211xp5_ASAP7_75t_L g1854 ( 
.A1(n_1853),
.A2(n_1550),
.B(n_1551),
.C(n_1537),
.Y(n_1854)
);


endmodule