module fake_jpeg_16909_n_364 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_364);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_364;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_18),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_54),
.Y(n_70)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_22),
.B(n_19),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_22),
.B(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_63),
.Y(n_86)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_56),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_84),
.Y(n_111)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_59),
.A2(n_33),
.B1(n_20),
.B2(n_22),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_76),
.A2(n_58),
.B1(n_51),
.B2(n_42),
.Y(n_116)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_57),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_36),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_0),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_59),
.A2(n_33),
.B1(n_20),
.B2(n_23),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_87),
.A2(n_50),
.B1(n_62),
.B2(n_61),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_50),
.Y(n_88)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_36),
.Y(n_89)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_30),
.Y(n_90)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

BUFx12_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_91),
.B(n_102),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_72),
.A2(n_33),
.B1(n_49),
.B2(n_52),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_93),
.A2(n_100),
.B1(n_122),
.B2(n_82),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_70),
.B(n_30),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_94),
.B(n_97),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_84),
.A2(n_23),
.B1(n_27),
.B2(n_55),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_96),
.A2(n_120),
.B1(n_75),
.B2(n_81),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_25),
.B(n_40),
.C(n_42),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_51),
.B1(n_52),
.B2(n_55),
.Y(n_100)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_105),
.Y(n_137)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_106),
.A2(n_116),
.B1(n_66),
.B2(n_74),
.Y(n_147)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_107),
.B(n_88),
.Y(n_153)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_109),
.Y(n_152)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_114),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_77),
.Y(n_114)
);

BUFx4f_ASAP7_75t_SL g115 ( 
.A(n_73),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_115),
.Y(n_127)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_119),
.Y(n_146)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_118),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_25),
.Y(n_119)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_31),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_L g122 ( 
.A1(n_66),
.A2(n_63),
.B1(n_60),
.B2(n_46),
.Y(n_122)
);

AOI21xp33_ASAP7_75t_L g123 ( 
.A1(n_111),
.A2(n_83),
.B(n_86),
.Y(n_123)
);

BUFx24_ASAP7_75t_SL g174 ( 
.A(n_123),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_125),
.A2(n_142),
.B1(n_150),
.B2(n_120),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_126),
.B(n_108),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_121),
.A2(n_81),
.B1(n_75),
.B2(n_71),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_128),
.A2(n_130),
.B1(n_64),
.B2(n_62),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_98),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_129),
.A2(n_147),
.B1(n_149),
.B2(n_95),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_121),
.A2(n_100),
.B1(n_82),
.B2(n_74),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_78),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_139),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_109),
.A2(n_40),
.B1(n_79),
.B2(n_78),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_135),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_97),
.B(n_79),
.Y(n_139)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_122),
.Y(n_144)
);

INVxp33_ASAP7_75t_L g171 ( 
.A(n_144),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_64),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_80),
.Y(n_173)
);

OR2x4_ASAP7_75t_L g148 ( 
.A(n_103),
.B(n_26),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_148),
.A2(n_61),
.B(n_53),
.Y(n_170)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_92),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

INVx5_ASAP7_75t_SL g163 ( 
.A(n_151),
.Y(n_163)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_153),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_132),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_157),
.B(n_160),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_145),
.Y(n_161)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_88),
.C(n_101),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_164),
.C(n_167),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_77),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_148),
.A2(n_112),
.B1(n_95),
.B2(n_107),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_165),
.A2(n_152),
.B1(n_150),
.B2(n_142),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_139),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_166),
.A2(n_170),
.B(n_173),
.Y(n_184)
);

MAJx2_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_91),
.C(n_104),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_149),
.A2(n_102),
.B1(n_118),
.B2(n_80),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_73),
.C(n_44),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_172),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_44),
.C(n_47),
.Y(n_172)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_173),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_146),
.Y(n_175)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_133),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_31),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_R g198 ( 
.A1(n_177),
.A2(n_152),
.B(n_32),
.Y(n_198)
);

AO21x1_ASAP7_75t_L g222 ( 
.A1(n_184),
.A2(n_196),
.B(n_199),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_158),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_186),
.B(n_193),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_167),
.B(n_129),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_198),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_188),
.Y(n_224)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_190),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_191),
.A2(n_194),
.B1(n_138),
.B2(n_124),
.Y(n_227)
);

BUFx5_ASAP7_75t_L g192 ( 
.A(n_154),
.Y(n_192)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_192),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_158),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_166),
.A2(n_134),
.B(n_131),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_156),
.Y(n_197)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_178),
.A2(n_127),
.B(n_131),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_156),
.Y(n_201)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_201),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_166),
.A2(n_127),
.B(n_133),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_202),
.B(n_138),
.Y(n_228)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_169),
.Y(n_203)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_203),
.Y(n_226)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_168),
.Y(n_204)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_204),
.A2(n_171),
.B1(n_157),
.B2(n_164),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_206),
.A2(n_213),
.B1(n_216),
.B2(n_217),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_201),
.Y(n_207)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_207),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_175),
.Y(n_208)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_208),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_188),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_212),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_180),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_179),
.A2(n_176),
.B1(n_162),
.B2(n_167),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_160),
.C(n_174),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_21),
.C(n_26),
.Y(n_244)
);

OA21x2_ASAP7_75t_L g215 ( 
.A1(n_202),
.A2(n_182),
.B(n_187),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_233),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_182),
.A2(n_172),
.B1(n_177),
.B2(n_170),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_203),
.A2(n_154),
.B1(n_141),
.B2(n_163),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_141),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_219),
.A2(n_195),
.B(n_151),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_183),
.A2(n_163),
.B1(n_124),
.B2(n_138),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_220),
.A2(n_230),
.B1(n_181),
.B2(n_193),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_225),
.B(n_232),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_227),
.A2(n_194),
.B1(n_189),
.B2(n_199),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_228),
.B(n_21),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_181),
.A2(n_38),
.B1(n_43),
.B2(n_37),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_229),
.A2(n_43),
.B1(n_38),
.B2(n_37),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_180),
.A2(n_124),
.B1(n_140),
.B2(n_47),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_190),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_192),
.Y(n_233)
);

XNOR2x1_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_185),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_235),
.A2(n_219),
.B1(n_221),
.B2(n_223),
.Y(n_263)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_237),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_238),
.A2(n_43),
.B1(n_37),
.B2(n_38),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_225),
.A2(n_189),
.B1(n_184),
.B2(n_196),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_239),
.A2(n_247),
.B1(n_224),
.B2(n_259),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_218),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_243),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_195),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_241),
.A2(n_220),
.B(n_230),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_242),
.A2(n_219),
.B(n_208),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_210),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_248),
.C(n_249),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_211),
.B(n_140),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_250),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_226),
.A2(n_140),
.B1(n_151),
.B2(n_2),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_211),
.B(n_151),
.C(n_62),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_214),
.B(n_61),
.C(n_53),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_53),
.C(n_91),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_39),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_253),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_222),
.B(n_39),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_213),
.B(n_215),
.Y(n_255)
);

BUFx12_ASAP7_75t_L g277 ( 
.A(n_255),
.Y(n_277)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_256),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_21),
.Y(n_257)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_257),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_210),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_205),
.Y(n_274)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_260),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_262),
.B(n_263),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_245),
.A2(n_207),
.B(n_221),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_264),
.A2(n_274),
.B(n_279),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_217),
.Y(n_266)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_266),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_267),
.A2(n_272),
.B1(n_282),
.B2(n_251),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_236),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_268),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_235),
.A2(n_206),
.B1(n_216),
.B2(n_224),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_237),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_278),
.A2(n_241),
.B1(n_244),
.B2(n_4),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_239),
.B(n_0),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_255),
.A2(n_1),
.B(n_2),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_281),
.A2(n_241),
.B(n_3),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_252),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_265),
.A2(n_238),
.B1(n_253),
.B2(n_247),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_283),
.A2(n_286),
.B1(n_279),
.B2(n_266),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_246),
.C(n_250),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_290),
.C(n_299),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_285),
.B(n_295),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_270),
.A2(n_234),
.B1(n_249),
.B2(n_248),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_287),
.A2(n_301),
.B1(n_271),
.B2(n_276),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_261),
.B(n_234),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_292),
.C(n_293),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_272),
.C(n_263),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_262),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_260),
.Y(n_293)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_294),
.Y(n_309)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_275),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_282),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_273),
.B(n_32),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_269),
.B(n_32),
.C(n_26),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_280),
.C(n_268),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_279),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_302),
.B(n_313),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_287),
.B(n_267),
.Y(n_304)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_304),
.Y(n_322)
);

BUFx24_ASAP7_75t_SL g306 ( 
.A(n_297),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_306),
.B(n_310),
.Y(n_331)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_307),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_284),
.B(n_264),
.Y(n_310)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_311),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_301),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_312),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_291),
.A2(n_277),
.B1(n_5),
.B2(n_6),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_314),
.A2(n_317),
.B1(n_312),
.B2(n_313),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_289),
.B(n_277),
.C(n_39),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_315),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_290),
.B(n_277),
.C(n_28),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_300),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_288),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_309),
.A2(n_285),
.B1(n_296),
.B2(n_292),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_318),
.B(n_8),
.Y(n_335)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_320),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_315),
.A2(n_316),
.B1(n_305),
.B2(n_308),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_321),
.A2(n_327),
.B1(n_11),
.B2(n_12),
.Y(n_340)
);

A2O1A1Ixp33_ASAP7_75t_L g323 ( 
.A1(n_305),
.A2(n_296),
.B(n_293),
.C(n_299),
.Y(n_323)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_323),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_330),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_303),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_28),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_322),
.B(n_7),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_334),
.B(n_13),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_335),
.A2(n_340),
.B1(n_324),
.B2(n_331),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_326),
.B(n_28),
.C(n_34),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_336),
.B(n_338),
.Y(n_344)
);

AOI21xp33_ASAP7_75t_L g337 ( 
.A1(n_319),
.A2(n_11),
.B(n_12),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_337),
.A2(n_15),
.B(n_16),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_326),
.B(n_34),
.C(n_12),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_325),
.B(n_34),
.C(n_15),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_341),
.B(n_15),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_342),
.B(n_345),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_339),
.A2(n_328),
.B(n_329),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_343),
.A2(n_346),
.B(n_348),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_338),
.Y(n_345)
);

AO21x1_ASAP7_75t_L g350 ( 
.A1(n_347),
.A2(n_349),
.B(n_336),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_333),
.A2(n_328),
.B1(n_324),
.B2(n_318),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_350),
.B(n_353),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_345),
.B(n_330),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_351),
.A2(n_352),
.B(n_344),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_348),
.B(n_332),
.Y(n_352)
);

OAI21x1_ASAP7_75t_L g358 ( 
.A1(n_355),
.A2(n_356),
.B(n_357),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_354),
.A2(n_341),
.B(n_332),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g359 ( 
.A(n_358),
.B(n_323),
.Y(n_359)
);

NAND3xp33_ASAP7_75t_L g360 ( 
.A(n_359),
.B(n_17),
.C(n_18),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_360),
.B(n_17),
.C(n_19),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_361),
.B(n_17),
.C(n_34),
.Y(n_362)
);

BUFx24_ASAP7_75t_SL g363 ( 
.A(n_362),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_363),
.B(n_34),
.Y(n_364)
);


endmodule