module fake_jpeg_4300_n_300 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx4_ASAP7_75t_SL g31 ( 
.A(n_22),
.Y(n_31)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_32),
.B(n_33),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_37),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx2_ASAP7_75t_R g37 ( 
.A(n_22),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_56),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_20),
.B1(n_17),
.B2(n_19),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_47),
.A2(n_33),
.B(n_28),
.C(n_18),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_15),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_49),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g49 ( 
.A(n_37),
.B(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_50),
.B(n_16),
.Y(n_72)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_19),
.B1(n_24),
.B2(n_20),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_53),
.A2(n_57),
.B1(n_58),
.B2(n_16),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_15),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_33),
.Y(n_70)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_37),
.A2(n_19),
.B1(n_24),
.B2(n_20),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_31),
.A2(n_16),
.B1(n_21),
.B2(n_23),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_39),
.Y(n_78)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_32),
.B(n_23),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_21),
.B(n_23),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_SL g92 ( 
.A1(n_65),
.A2(n_25),
.B(n_28),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_68),
.Y(n_101)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_69),
.A2(n_75),
.B1(n_81),
.B2(n_84),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_70),
.B(n_73),
.Y(n_103)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_74),
.Y(n_107)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_49),
.A2(n_39),
.B1(n_35),
.B2(n_41),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_60),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_76),
.Y(n_93)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_27),
.Y(n_79)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_43),
.B(n_18),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_80),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_27),
.Y(n_82)
);

NAND3xp33_ASAP7_75t_SL g108 ( 
.A(n_82),
.B(n_85),
.C(n_26),
.Y(n_108)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_43),
.B(n_27),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_75),
.A2(n_49),
.B(n_50),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_86),
.A2(n_92),
.B(n_102),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_74),
.C(n_75),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_85),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_65),
.A2(n_49),
.B1(n_38),
.B2(n_44),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_91),
.A2(n_65),
.B1(n_44),
.B2(n_78),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_47),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_98),
.Y(n_111)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_97),
.Y(n_125)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_76),
.Y(n_98)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_100),
.Y(n_130)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_77),
.B(n_45),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_51),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_73),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_93),
.Y(n_112)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_107),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_118),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_81),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_110),
.B(n_117),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_112),
.B(n_129),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_120),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_107),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_116),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_90),
.B(n_103),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_90),
.B(n_92),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_98),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_101),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_122),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_108),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_123),
.A2(n_88),
.B(n_94),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_80),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_124),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_79),
.Y(n_127)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_72),
.Y(n_128)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_82),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_102),
.A2(n_44),
.B1(n_46),
.B2(n_71),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_133),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_83),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_132),
.B(n_97),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_140),
.Y(n_163)
);

NOR2x1_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_102),
.Y(n_135)
);

FAx1_ASAP7_75t_SL g166 ( 
.A(n_135),
.B(n_143),
.CI(n_112),
.CON(n_166),
.SN(n_166)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_136),
.A2(n_138),
.B(n_128),
.Y(n_164)
);

AND2x2_ASAP7_75t_SL g138 ( 
.A(n_114),
.B(n_102),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_118),
.A2(n_89),
.B1(n_86),
.B2(n_94),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_139),
.A2(n_141),
.B1(n_99),
.B2(n_100),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_130),
.A2(n_86),
.B1(n_111),
.B2(n_102),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_91),
.C(n_105),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_151),
.C(n_152),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_116),
.A2(n_71),
.B1(n_84),
.B2(n_55),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_147),
.A2(n_55),
.B1(n_46),
.B2(n_56),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_105),
.C(n_64),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_45),
.C(n_99),
.Y(n_152)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_156),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_113),
.B(n_100),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_109),
.C(n_121),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_119),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_160),
.B(n_175),
.C(n_176),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_127),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_162),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_139),
.Y(n_162)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_164),
.A2(n_181),
.B(n_56),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_129),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_165),
.B(n_178),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_183),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_142),
.A2(n_136),
.B(n_157),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_168),
.Y(n_193)
);

BUFx12_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_110),
.Y(n_169)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_169),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_96),
.Y(n_170)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_144),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_179),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_152),
.A2(n_117),
.B(n_124),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_174),
.B(n_177),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_123),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_96),
.Y(n_177)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

OAI321xp33_ASAP7_75t_L g180 ( 
.A1(n_135),
.A2(n_95),
.A3(n_126),
.B1(n_132),
.B2(n_83),
.C(n_125),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_180),
.B(n_182),
.Y(n_205)
);

A2O1A1O1Ixp25_ASAP7_75t_L g181 ( 
.A1(n_143),
.A2(n_95),
.B(n_51),
.C(n_59),
.D(n_52),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_150),
.B(n_97),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_146),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_184),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_191),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_176),
.A2(n_141),
.B1(n_154),
.B2(n_137),
.Y(n_187)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_187),
.Y(n_226)
);

XNOR2x1_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_151),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_200),
.Y(n_221)
);

OA21x2_ASAP7_75t_L g191 ( 
.A1(n_166),
.A2(n_181),
.B(n_165),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_172),
.A2(n_137),
.B1(n_148),
.B2(n_150),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_194),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_171),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_196),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_159),
.A2(n_148),
.B1(n_155),
.B2(n_175),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_197),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_159),
.A2(n_155),
.B1(n_145),
.B2(n_38),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_199),
.A2(n_204),
.B(n_208),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_184),
.A2(n_38),
.B1(n_61),
.B2(n_46),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_201),
.B(n_68),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_161),
.A2(n_42),
.B1(n_55),
.B2(n_25),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_168),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_26),
.Y(n_217)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_209),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_207),
.B(n_160),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_221),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_R g213 ( 
.A(n_189),
.B(n_168),
.Y(n_213)
);

FAx1_ASAP7_75t_SL g244 ( 
.A(n_213),
.B(n_223),
.CI(n_40),
.CON(n_244),
.SN(n_244)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_188),
.B(n_198),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_185),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_35),
.C(n_39),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_218),
.C(n_227),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_217),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_197),
.C(n_203),
.Y(n_218)
);

FAx1_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_68),
.CI(n_30),
.CON(n_219),
.SN(n_219)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_219),
.A2(n_228),
.B(n_201),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_66),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_204),
.Y(n_233)
);

NAND3xp33_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_30),
.C(n_29),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_199),
.B(n_26),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_1),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_187),
.B(n_66),
.C(n_41),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_190),
.B(n_30),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_212),
.A2(n_190),
.B1(n_192),
.B2(n_194),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_230),
.A2(n_236),
.B1(n_239),
.B2(n_223),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_228),
.B(n_195),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_231),
.B(n_219),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_193),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_233),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_234),
.A2(n_227),
.B(n_224),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_210),
.A2(n_202),
.B1(n_191),
.B2(n_21),
.Y(n_236)
);

INVx11_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_244),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_226),
.A2(n_191),
.B1(n_30),
.B2(n_40),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_1),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_241),
.C(n_246),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_41),
.C(n_40),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_3),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_2),
.C(n_3),
.Y(n_246)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_247),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_248),
.Y(n_263)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

A2O1A1Ixp33_ASAP7_75t_L g252 ( 
.A1(n_233),
.A2(n_219),
.B(n_5),
.C(n_6),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_252),
.A2(n_240),
.B1(n_10),
.B2(n_12),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_243),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_253),
.B(n_259),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_4),
.Y(n_254)
);

AOI21xp33_ASAP7_75t_L g268 ( 
.A1(n_254),
.A2(n_261),
.B(n_257),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_4),
.C(n_5),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_237),
.C(n_229),
.Y(n_265)
);

OAI321xp33_ASAP7_75t_L g259 ( 
.A1(n_244),
.A2(n_4),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C(n_9),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_241),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_260),
.B(n_12),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_6),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_265),
.A2(n_255),
.B(n_252),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_237),
.C(n_232),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_266),
.A2(n_268),
.B(n_273),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_248),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_238),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_247),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_7),
.Y(n_272)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_272),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_7),
.C(n_10),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_12),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_281),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_255),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_277),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_278),
.A2(n_284),
.B(n_280),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_282),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_14),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_265),
.A2(n_13),
.B(n_14),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_283),
.B(n_13),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_13),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_284),
.Y(n_286)
);

AOI322xp5_ASAP7_75t_L g285 ( 
.A1(n_275),
.A2(n_262),
.A3(n_263),
.B1(n_267),
.B2(n_266),
.C1(n_269),
.C2(n_273),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_289),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_287),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_279),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_292),
.B(n_294),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_290),
.B(n_286),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_295),
.B(n_296),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_286),
.Y(n_296)
);

OAI21x1_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_293),
.B(n_296),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_297),
.Y(n_300)
);


endmodule