module fake_jpeg_4660_n_140 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_140);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx10_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_0),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_35),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_31),
.A2(n_16),
.B1(n_15),
.B2(n_17),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_44),
.B1(n_25),
.B2(n_24),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_29),
.A2(n_15),
.B1(n_16),
.B2(n_26),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_19),
.C(n_20),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_28),
.A2(n_21),
.B1(n_25),
.B2(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_47),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_18),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_49),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_40),
.B(n_21),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_33),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_52),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_14),
.Y(n_52)
);

FAx1_ASAP7_75t_SL g53 ( 
.A(n_40),
.B(n_35),
.CI(n_32),
.CON(n_53),
.SN(n_53)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_53),
.B(n_55),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_43),
.A2(n_23),
.B1(n_18),
.B2(n_27),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_61),
.B1(n_64),
.B2(n_0),
.Y(n_75)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_27),
.B(n_23),
.Y(n_56)
);

OR2x4_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_65),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_22),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_62),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_14),
.Y(n_58)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_9),
.B1(n_7),
.B2(n_4),
.Y(n_80)
);

O2A1O1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_45),
.A2(n_30),
.B(n_13),
.C(n_34),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_38),
.B1(n_1),
.B2(n_2),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_37),
.A2(n_20),
.B1(n_13),
.B2(n_34),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_37),
.A2(n_12),
.B1(n_11),
.B2(n_9),
.Y(n_64)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_38),
.B(n_34),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_67),
.A2(n_80),
.B1(n_61),
.B2(n_57),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_73),
.Y(n_89)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_77),
.Y(n_98)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_71),
.A2(n_46),
.B1(n_47),
.B2(n_62),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_96),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_86),
.B(n_91),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_51),
.C(n_56),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_79),
.C(n_74),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_51),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_67),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_78),
.B(n_53),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_53),
.Y(n_92)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_55),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_97),
.B(n_68),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_60),
.Y(n_95)
);

OAI21xp33_ASAP7_75t_SL g104 ( 
.A1(n_95),
.A2(n_94),
.B(n_97),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_38),
.B1(n_3),
.B2(n_4),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_38),
.Y(n_97)
);

AO21x1_ASAP7_75t_L g114 ( 
.A1(n_99),
.A2(n_109),
.B(n_96),
.Y(n_114)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_103),
.A2(n_104),
.B(n_108),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_72),
.Y(n_105)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_69),
.C(n_38),
.Y(n_108)
);

NAND2xp67_ASAP7_75t_SL g109 ( 
.A(n_95),
.B(n_80),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_109),
.A2(n_84),
.B1(n_95),
.B2(n_85),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_100),
.A2(n_107),
.B1(n_102),
.B2(n_99),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

AOI21x1_ASAP7_75t_L g120 ( 
.A1(n_114),
.A2(n_90),
.B(n_98),
.Y(n_120)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_117),
.B(n_88),
.C(n_103),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_101),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_119),
.C(n_123),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_120),
.A2(n_114),
.B(n_110),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_82),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_115),
.C(n_116),
.Y(n_130)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_126),
.Y(n_129)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_128),
.B(n_77),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_131),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_116),
.C(n_81),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_132),
.A2(n_2),
.B(n_4),
.Y(n_134)
);

NAND3xp33_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_128),
.C(n_3),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_133),
.B(n_134),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_135),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_5),
.C(n_6),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_6),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_137),
.Y(n_140)
);


endmodule