module fake_jpeg_14632_n_330 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_41),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_30),
.B1(n_26),
.B2(n_25),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_47),
.A2(n_50),
.B1(n_56),
.B2(n_32),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_20),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_48),
.B(n_32),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_43),
.A2(n_26),
.B1(n_31),
.B2(n_27),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_49),
.A2(n_51),
.B1(n_64),
.B2(n_19),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_34),
.A2(n_26),
.B1(n_25),
.B2(n_18),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_35),
.A2(n_31),
.B1(n_22),
.B2(n_28),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_19),
.B1(n_28),
.B2(n_27),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_52),
.A2(n_63),
.B1(n_20),
.B2(n_19),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_59),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_18),
.B1(n_25),
.B2(n_16),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_39),
.A2(n_24),
.B1(n_16),
.B2(n_21),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_39),
.A2(n_22),
.B1(n_28),
.B2(n_27),
.Y(n_64)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_70),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_22),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_68),
.B(n_74),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_63),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_90),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_72),
.A2(n_0),
.B(n_1),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_73),
.A2(n_89),
.B1(n_71),
.B2(n_76),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_57),
.B(n_20),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_24),
.Y(n_75)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

AO22x2_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_41),
.B1(n_25),
.B2(n_18),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_76),
.A2(n_79),
.B1(n_66),
.B2(n_16),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_51),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_78),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_29),
.Y(n_78)
);

OAI32xp33_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_49),
.A3(n_47),
.B1(n_50),
.B2(n_59),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_29),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_L g116 ( 
.A1(n_80),
.A2(n_92),
.B(n_93),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_81),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_24),
.Y(n_82)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_44),
.A2(n_18),
.B1(n_21),
.B2(n_32),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_83),
.A2(n_54),
.B1(n_17),
.B2(n_29),
.Y(n_119)
);

INVx13_ASAP7_75t_SL g85 ( 
.A(n_53),
.Y(n_85)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_46),
.A2(n_55),
.B1(n_60),
.B2(n_44),
.Y(n_89)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_29),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_61),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_94),
.A2(n_79),
.B1(n_76),
.B2(n_73),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_21),
.B(n_65),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_96),
.A2(n_79),
.B(n_76),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_98),
.A2(n_105),
.B1(n_107),
.B2(n_118),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_62),
.C(n_61),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_80),
.C(n_93),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_76),
.A2(n_66),
.B1(n_62),
.B2(n_54),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_102),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.Y(n_137)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_103),
.B(n_106),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_69),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_72),
.A2(n_54),
.B1(n_45),
.B2(n_29),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_68),
.B(n_45),
.Y(n_112)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_74),
.B(n_45),
.Y(n_113)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_17),
.Y(n_115)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

INVxp33_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_SL g131 ( 
.A1(n_117),
.A2(n_76),
.B(n_86),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_78),
.A2(n_54),
.B1(n_1),
.B2(n_2),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_119),
.A2(n_88),
.B1(n_81),
.B2(n_29),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_122),
.A2(n_137),
.B1(n_144),
.B2(n_102),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_123),
.A2(n_131),
.B(n_135),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_101),
.C(n_116),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_75),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_126),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_110),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_82),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_129),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_83),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_91),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_132),
.B(n_134),
.Y(n_173)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_100),
.B(n_76),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_111),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_89),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_139),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_96),
.B(n_84),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_96),
.B(n_84),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_94),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_141),
.A2(n_103),
.B1(n_119),
.B2(n_95),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_104),
.Y(n_142)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_143),
.B(n_111),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_97),
.A2(n_15),
.B1(n_1),
.B2(n_2),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_146),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_146),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_153),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_149),
.A2(n_99),
.B1(n_135),
.B2(n_114),
.Y(n_194)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_101),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_151),
.A2(n_159),
.B(n_169),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_145),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_122),
.A2(n_98),
.B1(n_97),
.B2(n_94),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_154),
.A2(n_156),
.B1(n_163),
.B2(n_164),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_109),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_155),
.B(n_138),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_121),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_165),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_168),
.C(n_172),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_140),
.A2(n_105),
.B(n_100),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_141),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_147),
.A2(n_98),
.B1(n_107),
.B2(n_105),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_147),
.A2(n_107),
.B1(n_116),
.B2(n_95),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_124),
.B(n_115),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_123),
.A2(n_113),
.B(n_109),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_125),
.B(n_118),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_126),
.Y(n_174)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_163),
.A2(n_123),
.B1(n_134),
.B2(n_131),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_176),
.A2(n_187),
.B1(n_194),
.B2(n_199),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_155),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_178),
.B(n_182),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_128),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_200),
.C(n_160),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_195),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_169),
.A2(n_136),
.B(n_127),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_181),
.A2(n_185),
.B(n_180),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_162),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_159),
.A2(n_136),
.B(n_127),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_162),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_186),
.B(n_188),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_164),
.A2(n_144),
.B1(n_118),
.B2(n_145),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_173),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_152),
.B(n_130),
.Y(n_189)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_130),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_191),
.B(n_196),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_193),
.B(n_167),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_173),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_99),
.Y(n_196)
);

INVxp33_ASAP7_75t_L g197 ( 
.A(n_157),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_197),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_171),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_171),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_149),
.A2(n_114),
.B1(n_120),
.B2(n_121),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_121),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_217),
.C(n_193),
.Y(n_234)
);

AO22x2_ASAP7_75t_L g204 ( 
.A1(n_178),
.A2(n_170),
.B1(n_154),
.B2(n_161),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_204),
.A2(n_205),
.B1(n_209),
.B2(n_212),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_199),
.A2(n_170),
.B1(n_156),
.B2(n_167),
.Y(n_205)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_206),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_208),
.B(n_222),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_184),
.A2(n_151),
.B1(n_166),
.B2(n_114),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_151),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_214),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_194),
.A2(n_120),
.B1(n_103),
.B2(n_133),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_133),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_179),
.B(n_142),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_220),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_142),
.C(n_88),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_184),
.A2(n_142),
.B1(n_88),
.B2(n_3),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_219),
.A2(n_221),
.B1(n_175),
.B2(n_189),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_177),
.B(n_17),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_188),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_175),
.B(n_15),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_223),
.B(n_0),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_190),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_190),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_226),
.Y(n_262)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_210),
.Y(n_227)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_183),
.Y(n_228)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_228),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_206),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_229),
.A2(n_237),
.B(n_241),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_213),
.B(n_174),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_230),
.B(n_243),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_235),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_233),
.B(n_240),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_239),
.C(n_244),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_225),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_218),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_177),
.C(n_185),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_207),
.B(n_182),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_181),
.C(n_195),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_204),
.A2(n_186),
.B(n_176),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_245),
.A2(n_219),
.B(n_220),
.Y(n_253)
);

NOR3xp33_ASAP7_75t_SL g247 ( 
.A(n_241),
.B(n_204),
.C(n_222),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_236),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_R g248 ( 
.A(n_229),
.B(n_204),
.Y(n_248)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_248),
.Y(n_272)
);

XNOR2x1_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_211),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_258),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_245),
.A2(n_209),
.B1(n_201),
.B2(n_202),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_252),
.A2(n_253),
.B1(n_259),
.B2(n_0),
.Y(n_275)
);

A2O1A1O1Ixp25_ASAP7_75t_L g255 ( 
.A1(n_246),
.A2(n_208),
.B(n_205),
.C(n_202),
.D(n_203),
.Y(n_255)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_255),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_217),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_237),
.A2(n_187),
.B1(n_198),
.B2(n_212),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_221),
.C(n_29),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_263),
.C(n_264),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_17),
.C(n_2),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_17),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_244),
.C(n_231),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_269),
.C(n_280),
.Y(n_287)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_268),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_231),
.C(n_242),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_257),
.Y(n_270)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_270),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_262),
.A2(n_235),
.B1(n_243),
.B2(n_232),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_271),
.A2(n_274),
.B1(n_5),
.B2(n_6),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_248),
.A2(n_227),
.B1(n_236),
.B2(n_246),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_253),
.Y(n_284)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_250),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_279),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_265),
.B(n_260),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_278),
.B(n_281),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_252),
.B(n_259),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_263),
.C(n_261),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_17),
.C(n_4),
.Y(n_281)
);

AOI21x1_ASAP7_75t_L g282 ( 
.A1(n_274),
.A2(n_247),
.B(n_250),
.Y(n_282)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_282),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_284),
.B(n_288),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_264),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_291),
.C(n_293),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_276),
.A2(n_249),
.B(n_255),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_289),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_3),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_5),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_5),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_5),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_266),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_271),
.Y(n_299)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_299),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_266),
.Y(n_301)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_301),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_6),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_281),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_304),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_290),
.B(n_291),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_284),
.A2(n_273),
.B1(n_7),
.B2(n_8),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_9),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_283),
.A2(n_273),
.B(n_7),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_287),
.A2(n_285),
.B1(n_7),
.B2(n_8),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_287),
.C(n_8),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_312),
.C(n_296),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_309),
.A2(n_313),
.B(n_9),
.Y(n_321)
);

AOI21x1_ASAP7_75t_SL g310 ( 
.A1(n_300),
.A2(n_6),
.B(n_8),
.Y(n_310)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_310),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_9),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_298),
.A2(n_9),
.B(n_10),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_316),
.B(n_10),
.Y(n_323)
);

NOR2x1_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_297),
.Y(n_317)
);

OAI321xp33_ASAP7_75t_L g325 ( 
.A1(n_317),
.A2(n_320),
.A3(n_311),
.B1(n_309),
.B2(n_314),
.C(n_12),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_319),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_308),
.Y(n_319)
);

AO21x1_ASAP7_75t_L g324 ( 
.A1(n_321),
.A2(n_322),
.B(n_323),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_305),
.C(n_11),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_325),
.A2(n_317),
.B1(n_12),
.B2(n_13),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_324),
.B1(n_12),
.B2(n_11),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_328),
.A2(n_326),
.B(n_11),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_11),
.Y(n_330)
);


endmodule