module fake_jpeg_11931_n_476 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_476);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_476;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_48),
.Y(n_133)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_50),
.Y(n_123)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_51),
.Y(n_141)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_30),
.B(n_16),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_55),
.B(n_66),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g148 ( 
.A(n_57),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_59),
.Y(n_139)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_26),
.B(n_16),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_72),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_28),
.B(n_16),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_63),
.B(n_75),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_26),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_68),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_39),
.Y(n_69)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_19),
.Y(n_71)
);

BUFx4f_ASAP7_75t_SL g109 ( 
.A(n_71),
.Y(n_109)
);

NAND2x1_ASAP7_75t_SL g72 ( 
.A(n_28),
.B(n_15),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_73),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_74),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_33),
.B(n_35),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_76),
.Y(n_149)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_77),
.Y(n_140)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_79),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_80),
.Y(n_145)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_81),
.Y(n_147)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_87),
.Y(n_138)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_88),
.B(n_0),
.Y(n_144)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_89),
.B(n_0),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_17),
.B(n_14),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_92),
.Y(n_101)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_91),
.B(n_18),
.Y(n_136)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_51),
.B(n_38),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_95),
.B(n_126),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_69),
.A2(n_41),
.B1(n_27),
.B2(n_44),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_98),
.A2(n_106),
.B1(n_107),
.B2(n_110),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_75),
.A2(n_44),
.B1(n_35),
.B2(n_41),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_99),
.A2(n_105),
.B1(n_127),
.B2(n_13),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_86),
.A2(n_85),
.B1(n_55),
.B2(n_80),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_78),
.A2(n_41),
.B1(n_44),
.B2(n_38),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_47),
.A2(n_17),
.B1(n_34),
.B2(n_31),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_87),
.A2(n_38),
.B1(n_42),
.B2(n_46),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_L g111 ( 
.A1(n_54),
.A2(n_46),
.B1(n_42),
.B2(n_36),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_111),
.A2(n_112),
.B1(n_114),
.B2(n_116),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_70),
.A2(n_38),
.B1(n_36),
.B2(n_29),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_61),
.A2(n_38),
.B1(n_34),
.B2(n_31),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_76),
.A2(n_33),
.B1(n_24),
.B2(n_21),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_63),
.B(n_72),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_121),
.B(n_136),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_61),
.A2(n_24),
.B1(n_21),
.B2(n_20),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_64),
.C(n_58),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_74),
.A2(n_20),
.B1(n_18),
.B2(n_14),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_56),
.B(n_0),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_142),
.B(n_71),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_144),
.B(n_10),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_141),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_150),
.B(n_152),
.Y(n_232)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_151),
.Y(n_208)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_115),
.Y(n_153)
);

INVx3_ASAP7_75t_SL g237 ( 
.A(n_153),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_101),
.B(n_0),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_154),
.B(n_160),
.Y(n_231)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_97),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_155),
.Y(n_218)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_104),
.Y(n_156)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_156),
.Y(n_206)
);

NOR2x1_ASAP7_75t_L g215 ( 
.A(n_157),
.B(n_178),
.Y(n_215)
);

INVx3_ASAP7_75t_SL g159 ( 
.A(n_115),
.Y(n_159)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_159),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_100),
.B(n_1),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_95),
.B(n_1),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_161),
.B(n_175),
.Y(n_246)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_163),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_164),
.Y(n_229)
);

BUFx12_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_165),
.Y(n_253)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_166),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_96),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_167),
.Y(n_228)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_168),
.Y(n_223)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_104),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_169),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_95),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_170),
.B(n_183),
.Y(n_207)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_118),
.Y(n_171)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_171),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_99),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_172)
);

OAI22x1_ASAP7_75t_L g224 ( 
.A1(n_172),
.A2(n_173),
.B1(n_185),
.B2(n_197),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_105),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_94),
.B(n_5),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_93),
.B(n_7),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_193),
.C(n_195),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_96),
.Y(n_177)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_177),
.Y(n_245)
);

A2O1A1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_122),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_108),
.Y(n_179)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_179),
.Y(n_238)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_118),
.Y(n_180)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_180),
.Y(n_247)
);

BUFx8_ASAP7_75t_L g181 ( 
.A(n_109),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_181),
.Y(n_250)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_182),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_133),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_116),
.A2(n_125),
.B1(n_106),
.B2(n_98),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_184),
.A2(n_201),
.B1(n_129),
.B2(n_120),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_127),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_132),
.Y(n_186)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_186),
.Y(n_242)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_135),
.Y(n_187)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_187),
.Y(n_243)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_149),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_188),
.B(n_189),
.Y(n_252)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_139),
.Y(n_189)
);

INVx11_ASAP7_75t_L g190 ( 
.A(n_109),
.Y(n_190)
);

INVx3_ASAP7_75t_SL g240 ( 
.A(n_190),
.Y(n_240)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_139),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_192),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_123),
.B(n_8),
.C(n_9),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_140),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_194),
.B(n_198),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_130),
.B(n_8),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_138),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_196),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_128),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_137),
.B(n_10),
.Y(n_199)
);

MAJx2_ASAP7_75t_L g234 ( 
.A(n_199),
.B(n_198),
.C(n_193),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_147),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_202),
.Y(n_225)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_143),
.Y(n_202)
);

A2O1A1Ixp33_ASAP7_75t_L g203 ( 
.A1(n_114),
.A2(n_124),
.B(n_111),
.C(n_109),
.Y(n_203)
);

FAx1_ASAP7_75t_SL g230 ( 
.A(n_203),
.B(n_190),
.CI(n_161),
.CON(n_230),
.SN(n_230)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_120),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_148),
.Y(n_226)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_128),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_205),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_211),
.A2(n_212),
.B1(n_216),
.B2(n_220),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_174),
.A2(n_145),
.B1(n_117),
.B2(n_119),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_158),
.A2(n_129),
.B1(n_148),
.B2(n_112),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_213),
.A2(n_162),
.B(n_151),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_157),
.A2(n_119),
.B1(n_113),
.B2(n_146),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_162),
.A2(n_113),
.B1(n_146),
.B2(n_110),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_203),
.A2(n_148),
.B1(n_162),
.B2(n_160),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_221),
.A2(n_180),
.B1(n_192),
.B2(n_189),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_226),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_175),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_227),
.B(n_235),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_230),
.B(n_214),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_234),
.B(n_214),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_154),
.B(n_198),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_176),
.B(n_199),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_239),
.B(n_241),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_195),
.B(n_196),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_166),
.A2(n_159),
.B1(n_205),
.B2(n_171),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_256),
.B(n_275),
.Y(n_319)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_206),
.Y(n_257)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_257),
.Y(n_324)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_217),
.Y(n_258)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_258),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_211),
.A2(n_178),
.B1(n_153),
.B2(n_164),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_259),
.A2(n_266),
.B1(n_271),
.B2(n_291),
.Y(n_321)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_206),
.Y(n_260)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_260),
.Y(n_307)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_217),
.Y(n_262)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_262),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_215),
.A2(n_181),
.B(n_165),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_264),
.A2(n_273),
.B(n_250),
.Y(n_304)
);

XNOR2x1_ASAP7_75t_L g305 ( 
.A(n_265),
.B(n_281),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_212),
.A2(n_188),
.B1(n_182),
.B2(n_167),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_215),
.A2(n_177),
.B1(n_156),
.B2(n_169),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_267),
.A2(n_288),
.B1(n_240),
.B2(n_237),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_219),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_268),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_240),
.A2(n_165),
.B1(n_181),
.B2(n_213),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_269),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_228),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_270),
.B(n_276),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_215),
.A2(n_230),
.B1(n_220),
.B2(n_216),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_245),
.Y(n_272)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_272),
.Y(n_310)
);

O2A1O1Ixp33_ASAP7_75t_L g275 ( 
.A1(n_230),
.A2(n_207),
.B(n_232),
.C(n_208),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_252),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_208),
.Y(n_277)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_277),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_252),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_280),
.Y(n_303)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_242),
.Y(n_279)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_279),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_244),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_231),
.B(n_209),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_295),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_252),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_283),
.B(n_285),
.Y(n_306)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_248),
.Y(n_284)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_284),
.Y(n_335)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_232),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_225),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_286),
.B(n_294),
.Y(n_325)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_248),
.Y(n_287)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_287),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_231),
.A2(n_246),
.B1(n_224),
.B2(n_234),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_246),
.B(n_238),
.C(n_210),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_292),
.C(n_251),
.Y(n_301)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_242),
.Y(n_290)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_290),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_224),
.A2(n_236),
.B1(n_218),
.B2(n_238),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_223),
.B(n_210),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_243),
.Y(n_293)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_293),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_251),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_236),
.A2(n_218),
.B1(n_223),
.B2(n_237),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_243),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_296),
.B(n_297),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_253),
.B(n_233),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_267),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_300),
.B(n_322),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_301),
.B(n_272),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_304),
.A2(n_265),
.B(n_263),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_261),
.A2(n_240),
.B1(n_237),
.B2(n_250),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_311),
.A2(n_261),
.B1(n_268),
.B2(n_229),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_281),
.B(n_253),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_312),
.B(n_271),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_289),
.B(n_292),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_314),
.B(n_323),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_316),
.A2(n_328),
.B1(n_254),
.B2(n_276),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_264),
.A2(n_233),
.B(n_222),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_317),
.A2(n_304),
.B(n_331),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_295),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_318),
.B(n_333),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_294),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_282),
.B(n_274),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_288),
.B(n_222),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_327),
.B(n_293),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_273),
.A2(n_229),
.B1(n_219),
.B2(n_247),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_256),
.B(n_247),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_331),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_284),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_255),
.B(n_245),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g343 ( 
.A(n_334),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_325),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_336),
.B(n_346),
.Y(n_382)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_299),
.Y(n_337)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_337),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_338),
.B(n_356),
.C(n_313),
.Y(n_386)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_324),
.Y(n_339)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_339),
.Y(n_377)
);

INVx5_ASAP7_75t_L g340 ( 
.A(n_324),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_340),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_342),
.A2(n_347),
.B(n_348),
.Y(n_368)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_344),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_300),
.A2(n_275),
.B1(n_277),
.B2(n_258),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_317),
.Y(n_349)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_349),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_315),
.A2(n_270),
.B(n_280),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_350),
.A2(n_302),
.B(n_307),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_321),
.A2(n_262),
.B1(n_296),
.B2(n_279),
.Y(n_351)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_351),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_329),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_352),
.Y(n_387)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_353),
.Y(n_376)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_299),
.Y(n_354)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_354),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_316),
.A2(n_290),
.B1(n_260),
.B2(n_257),
.Y(n_355)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_355),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_308),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_357),
.B(n_359),
.Y(n_385)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_309),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_321),
.A2(n_229),
.B1(n_287),
.B2(n_318),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_360),
.A2(n_362),
.B1(n_363),
.B2(n_364),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_327),
.A2(n_298),
.B1(n_328),
.B2(n_319),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_298),
.A2(n_323),
.B1(n_306),
.B2(n_315),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_305),
.A2(n_301),
.B1(n_314),
.B2(n_319),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_303),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_365),
.Y(n_372)
);

BUFx4f_ASAP7_75t_L g366 ( 
.A(n_333),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_366),
.Y(n_378)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_309),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_367),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_338),
.B(n_312),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_370),
.B(n_392),
.Y(n_405)
);

NOR2xp67_ASAP7_75t_SL g373 ( 
.A(n_346),
.B(n_331),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_373),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_345),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_380),
.B(n_336),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_349),
.A2(n_348),
.B1(n_353),
.B2(n_358),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_381),
.A2(n_391),
.B1(n_362),
.B2(n_344),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_358),
.A2(n_319),
.B(n_305),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_384),
.A2(n_390),
.B(n_367),
.Y(n_407)
);

MAJx2_ASAP7_75t_L g411 ( 
.A(n_386),
.B(n_330),
.C(n_307),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_364),
.A2(n_313),
.B1(n_320),
.B2(n_332),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_356),
.B(n_332),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_394),
.A2(n_393),
.B1(n_388),
.B2(n_371),
.Y(n_426)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_385),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_395),
.B(n_400),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_370),
.B(n_341),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_396),
.B(n_408),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_392),
.B(n_341),
.C(n_347),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_397),
.B(n_398),
.C(n_404),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_386),
.B(n_361),
.C(n_352),
.Y(n_398)
);

CKINVDCx14_ASAP7_75t_R g422 ( 
.A(n_399),
.Y(n_422)
);

AOI21xp33_ASAP7_75t_L g400 ( 
.A1(n_387),
.A2(n_343),
.B(n_350),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_387),
.B(n_337),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_401),
.B(n_402),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_372),
.A2(n_369),
.B1(n_374),
.B2(n_393),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_382),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_403),
.B(n_406),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_391),
.B(n_384),
.C(n_369),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_382),
.Y(n_406)
);

NAND2xp33_ASAP7_75t_SL g416 ( 
.A(n_407),
.B(n_368),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g408 ( 
.A(n_381),
.B(n_355),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_371),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_409),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_374),
.A2(n_359),
.B1(n_354),
.B2(n_320),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_410),
.A2(n_388),
.B1(n_383),
.B2(n_378),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_411),
.B(n_375),
.C(n_376),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_376),
.B(n_373),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_412),
.B(n_413),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_379),
.B(n_310),
.Y(n_413)
);

AOI21xp33_ASAP7_75t_L g414 ( 
.A1(n_368),
.A2(n_302),
.B(n_330),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_414),
.A2(n_366),
.B(n_326),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_416),
.A2(n_407),
.B(n_415),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_423),
.B(n_411),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_405),
.B(n_375),
.C(n_390),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_424),
.B(n_428),
.Y(n_440)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_426),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_427),
.A2(n_429),
.B1(n_430),
.B2(n_394),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_405),
.B(n_383),
.C(n_310),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_404),
.A2(n_377),
.B1(n_389),
.B2(n_339),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_415),
.A2(n_377),
.B1(n_389),
.B2(n_340),
.Y(n_430)
);

OR2x2_ASAP7_75t_L g439 ( 
.A(n_432),
.B(n_433),
.Y(n_439)
);

FAx1_ASAP7_75t_SL g433 ( 
.A(n_397),
.B(n_366),
.CI(n_326),
.CON(n_433),
.SN(n_433)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_435),
.B(n_438),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_431),
.B(n_398),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_436),
.B(n_446),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_431),
.B(n_401),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_437),
.B(n_441),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_424),
.B(n_396),
.Y(n_438)
);

OAI21x1_ASAP7_75t_SL g454 ( 
.A1(n_442),
.A2(n_432),
.B(n_433),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_421),
.B(n_412),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_443),
.B(n_417),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_421),
.B(n_408),
.C(n_410),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_444),
.B(n_445),
.C(n_418),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_428),
.B(n_409),
.C(n_335),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_416),
.A2(n_422),
.B(n_423),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_447),
.B(n_454),
.Y(n_457)
);

AOI211xp5_ASAP7_75t_L g448 ( 
.A1(n_434),
.A2(n_425),
.B(n_420),
.C(n_422),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_448),
.A2(n_439),
.B1(n_419),
.B2(n_442),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_435),
.A2(n_426),
.B1(n_420),
.B2(n_425),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_449),
.B(n_452),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_438),
.B(n_417),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_455),
.B(n_440),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_444),
.B(n_429),
.C(n_418),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_456),
.B(n_445),
.C(n_443),
.Y(n_458)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_458),
.Y(n_464)
);

NOR2xp67_ASAP7_75t_L g459 ( 
.A(n_451),
.B(n_441),
.Y(n_459)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_459),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_461),
.A2(n_462),
.B(n_463),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_453),
.B(n_447),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_458),
.A2(n_439),
.B(n_456),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_466),
.B(n_457),
.Y(n_468)
);

OAI21x1_ASAP7_75t_L g470 ( 
.A1(n_468),
.A2(n_469),
.B(n_465),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_467),
.A2(n_460),
.B1(n_419),
.B2(n_457),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_L g472 ( 
.A1(n_470),
.A2(n_471),
.B1(n_427),
.B2(n_430),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_468),
.A2(n_464),
.B(n_461),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_472),
.A2(n_433),
.B(n_450),
.Y(n_473)
);

BUFx24_ASAP7_75t_SL g474 ( 
.A(n_473),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_474),
.B(n_450),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_475),
.B(n_455),
.Y(n_476)
);


endmodule