module fake_ariane_1654_n_1750 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1750);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1750;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_45),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_78),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_135),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_109),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_0),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_121),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_54),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_108),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_143),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_39),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_44),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_106),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_44),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_62),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_76),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_13),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_79),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_65),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_21),
.Y(n_173)
);

BUFx10_ASAP7_75t_L g174 ( 
.A(n_4),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_148),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_91),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_32),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_0),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_59),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_63),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_26),
.Y(n_181)
);

BUFx8_ASAP7_75t_SL g182 ( 
.A(n_111),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_151),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_25),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_7),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_56),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_125),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_71),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_10),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_104),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_129),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_112),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_140),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_81),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_149),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_128),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_25),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_6),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_42),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_80),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_97),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_147),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_114),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_42),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_146),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_13),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_6),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_35),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_17),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_101),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_33),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_83),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_34),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_37),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_27),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_34),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_95),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_72),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_87),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_40),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_138),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_142),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_58),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_116),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_119),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_2),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_14),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_7),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_11),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_17),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_74),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_139),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_127),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_24),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_16),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_33),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_31),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_45),
.Y(n_238)
);

BUFx10_ASAP7_75t_L g239 ( 
.A(n_132),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_154),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_19),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_96),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_105),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_19),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_120),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_11),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_16),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_77),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_70),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_66),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_86),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_14),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_69),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_40),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_27),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_51),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_53),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_133),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_75),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_123),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_23),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_35),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_137),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_21),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_103),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_67),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_39),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_153),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_107),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_1),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_113),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_88),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_68),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_136),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_23),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_73),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_15),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_94),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_46),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_38),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_32),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_15),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_82),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_93),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_134),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_122),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_115),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_43),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_84),
.Y(n_289)
);

BUFx5_ASAP7_75t_L g290 ( 
.A(n_30),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_89),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_48),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_37),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_28),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_30),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_31),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_92),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_49),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_117),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_46),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_12),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_9),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_36),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_64),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_38),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_130),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_18),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_290),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_290),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_182),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_290),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_157),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_292),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_292),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_196),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_290),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_238),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_155),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_290),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_290),
.Y(n_320)
);

NOR2xp67_ASAP7_75t_L g321 ( 
.A(n_305),
.B(n_1),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_290),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_L g323 ( 
.A(n_305),
.B(n_2),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_265),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_283),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_290),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_212),
.B(n_3),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_290),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_156),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_292),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_212),
.B(n_3),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_299),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_156),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_306),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_164),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_229),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_161),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_161),
.Y(n_338)
);

INVxp33_ASAP7_75t_L g339 ( 
.A(n_159),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_166),
.B(n_4),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_166),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_171),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g343 ( 
.A(n_292),
.Y(n_343)
);

NOR2xp67_ASAP7_75t_L g344 ( 
.A(n_189),
.B(n_5),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_171),
.B(n_5),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_170),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_292),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g348 ( 
.A(n_189),
.B(n_8),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_159),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_288),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_158),
.B(n_8),
.Y(n_351)
);

NOR2xp67_ASAP7_75t_L g352 ( 
.A(n_235),
.B(n_9),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_239),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_188),
.B(n_10),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_173),
.Y(n_355)
);

OR2x2_ASAP7_75t_L g356 ( 
.A(n_235),
.B(n_12),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_239),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_188),
.Y(n_358)
);

INVxp33_ASAP7_75t_L g359 ( 
.A(n_165),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_186),
.Y(n_360)
);

INVxp67_ASAP7_75t_SL g361 ( 
.A(n_165),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_190),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_177),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_190),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_191),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_178),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_181),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_191),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_218),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_218),
.B(n_18),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_184),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_185),
.Y(n_372)
);

NOR2xp67_ASAP7_75t_L g373 ( 
.A(n_237),
.B(n_20),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_222),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_222),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_198),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_199),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_239),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_186),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_195),
.B(n_224),
.Y(n_380)
);

INVxp33_ASAP7_75t_SL g381 ( 
.A(n_204),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_209),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_224),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_308),
.Y(n_384)
);

AND2x2_ASAP7_75t_SL g385 ( 
.A(n_327),
.B(n_210),
.Y(n_385)
);

INVx4_ASAP7_75t_L g386 ( 
.A(n_379),
.Y(n_386)
);

CKINVDCx8_ASAP7_75t_R g387 ( 
.A(n_310),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_308),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_318),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_309),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_309),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_311),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_313),
.B(n_225),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_335),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_329),
.B(n_237),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_346),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_311),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_330),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_312),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_316),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_316),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_314),
.B(n_225),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_319),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_319),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_329),
.B(n_280),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_330),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_330),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_380),
.B(n_210),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_320),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_320),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_322),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_322),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_326),
.Y(n_413)
);

INVx4_ASAP7_75t_L g414 ( 
.A(n_379),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_326),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_333),
.B(n_280),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_328),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_328),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_379),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_379),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_343),
.B(n_248),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_379),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_333),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_379),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_337),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_347),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_337),
.Y(n_427)
);

OAI21x1_ASAP7_75t_L g428 ( 
.A1(n_338),
.A2(n_257),
.B(n_248),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_338),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_341),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_341),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_342),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_342),
.B(n_257),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_358),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_358),
.B(n_362),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_380),
.B(n_266),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_362),
.B(n_181),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_364),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_364),
.B(n_266),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_355),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_365),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_365),
.Y(n_442)
);

INVx6_ASAP7_75t_L g443 ( 
.A(n_360),
.Y(n_443)
);

NOR3xp33_ASAP7_75t_L g444 ( 
.A(n_331),
.B(n_351),
.C(n_345),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_368),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_368),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_369),
.Y(n_447)
);

BUFx8_ASAP7_75t_L g448 ( 
.A(n_360),
.Y(n_448)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_360),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_369),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_374),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_374),
.Y(n_452)
);

BUFx6f_ASAP7_75t_SL g453 ( 
.A(n_385),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_394),
.B(n_366),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_388),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_394),
.B(n_372),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_423),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_423),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g459 ( 
.A(n_448),
.Y(n_459)
);

NAND2xp33_ASAP7_75t_L g460 ( 
.A(n_444),
.B(n_376),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_426),
.B(n_357),
.Y(n_461)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_435),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_426),
.B(n_357),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_425),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_425),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_399),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_435),
.B(n_339),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_385),
.B(n_375),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_425),
.Y(n_469)
);

BUFx6f_ASAP7_75t_SL g470 ( 
.A(n_385),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_449),
.B(n_381),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_425),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_388),
.Y(n_473)
);

AOI22xp33_ASAP7_75t_L g474 ( 
.A1(n_385),
.A2(n_354),
.B1(n_370),
.B2(n_340),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_436),
.B(n_435),
.Y(n_475)
);

NAND2xp33_ASAP7_75t_L g476 ( 
.A(n_444),
.B(n_425),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_425),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_443),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_443),
.Y(n_479)
);

AOI22xp33_ASAP7_75t_L g480 ( 
.A1(n_436),
.A2(n_321),
.B1(n_323),
.B2(n_359),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_388),
.Y(n_481)
);

INVxp33_ASAP7_75t_L g482 ( 
.A(n_389),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_425),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_394),
.B(n_382),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_386),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_425),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_387),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_388),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_391),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_391),
.Y(n_490)
);

OAI22xp33_ASAP7_75t_SL g491 ( 
.A1(n_408),
.A2(n_356),
.B1(n_348),
.B2(n_349),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_441),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_408),
.A2(n_323),
.B1(n_321),
.B2(n_167),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_435),
.B(n_363),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_422),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_448),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_441),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_391),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_386),
.Y(n_499)
);

OR2x6_ASAP7_75t_L g500 ( 
.A(n_396),
.B(n_348),
.Y(n_500)
);

OR2x6_ASAP7_75t_L g501 ( 
.A(n_396),
.B(n_356),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_441),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_442),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_435),
.B(n_375),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_449),
.B(n_371),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_435),
.B(n_383),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_442),
.Y(n_507)
);

INVx5_ASAP7_75t_L g508 ( 
.A(n_425),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_449),
.B(n_383),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_442),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_445),
.Y(n_511)
);

NAND2xp33_ASAP7_75t_L g512 ( 
.A(n_434),
.B(n_272),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_391),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_449),
.B(n_377),
.Y(n_514)
);

INVx6_ASAP7_75t_L g515 ( 
.A(n_449),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_397),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_434),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_386),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_434),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_397),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_386),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_449),
.B(n_317),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_440),
.B(n_315),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_440),
.B(n_325),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_387),
.B(n_332),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_434),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_434),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_429),
.B(n_361),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_397),
.Y(n_529)
);

OAI22xp33_ASAP7_75t_L g530 ( 
.A1(n_389),
.A2(n_246),
.B1(n_255),
.B2(n_262),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_437),
.B(n_367),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_386),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_397),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_415),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_387),
.B(n_334),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_434),
.Y(n_536)
);

NOR2x1p5_ASAP7_75t_L g537 ( 
.A(n_433),
.B(n_206),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_415),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_399),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_434),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_434),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_415),
.Y(n_542)
);

AO22x2_ASAP7_75t_L g543 ( 
.A1(n_437),
.A2(n_202),
.B1(n_286),
.B2(n_294),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_443),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_443),
.B(n_353),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_437),
.B(n_344),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_415),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_418),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_445),
.Y(n_549)
);

OAI22xp33_ASAP7_75t_L g550 ( 
.A1(n_433),
.A2(n_344),
.B1(n_373),
.B2(n_352),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_445),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_447),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_447),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_429),
.B(n_378),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_429),
.B(n_179),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_429),
.B(n_213),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_447),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_448),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_427),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_427),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_443),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_430),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_422),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_434),
.Y(n_564)
);

OAI22xp33_ASAP7_75t_L g565 ( 
.A1(n_439),
.A2(n_373),
.B1(n_352),
.B2(n_261),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_429),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_443),
.B(n_393),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_430),
.B(n_250),
.Y(n_568)
);

OR2x6_ASAP7_75t_L g569 ( 
.A(n_405),
.B(n_206),
.Y(n_569)
);

INVxp33_ASAP7_75t_SL g570 ( 
.A(n_405),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_418),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_386),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_431),
.B(n_272),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_418),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_414),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_418),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_431),
.B(n_273),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_413),
.Y(n_578)
);

OR2x6_ASAP7_75t_L g579 ( 
.A(n_405),
.B(n_207),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_432),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_422),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_414),
.Y(n_582)
);

INVx4_ASAP7_75t_L g583 ( 
.A(n_443),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_437),
.A2(n_226),
.B1(n_256),
.B2(n_234),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_414),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_432),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_413),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_414),
.Y(n_588)
);

AND3x2_ASAP7_75t_L g589 ( 
.A(n_416),
.B(n_208),
.C(n_207),
.Y(n_589)
);

AND2x6_ASAP7_75t_L g590 ( 
.A(n_437),
.B(n_273),
.Y(n_590)
);

NAND2xp33_ASAP7_75t_L g591 ( 
.A(n_390),
.B(n_274),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_452),
.B(n_274),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_413),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_422),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_452),
.B(n_202),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_437),
.B(n_214),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_432),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_448),
.B(n_393),
.Y(n_598)
);

INVx4_ASAP7_75t_L g599 ( 
.A(n_390),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_413),
.Y(n_600)
);

AO22x2_ASAP7_75t_L g601 ( 
.A1(n_453),
.A2(n_256),
.B1(n_208),
.B2(n_211),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_455),
.Y(n_602)
);

INVx5_ASAP7_75t_L g603 ( 
.A(n_515),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_487),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_566),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_462),
.B(n_448),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_539),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_460),
.A2(n_402),
.B1(n_421),
.B2(n_395),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_566),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_457),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_475),
.B(n_448),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_462),
.B(n_439),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_458),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_570),
.B(n_402),
.Y(n_614)
);

NAND2xp33_ASAP7_75t_L g615 ( 
.A(n_590),
.B(n_384),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_453),
.A2(n_395),
.B1(n_450),
.B2(n_446),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_462),
.B(n_421),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_L g618 ( 
.A1(n_474),
.A2(n_451),
.B1(n_450),
.B2(n_446),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_455),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_539),
.B(n_416),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_570),
.B(n_413),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_453),
.A2(n_395),
.B1(n_450),
.B2(n_446),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_531),
.B(n_404),
.Y(n_623)
);

OR2x2_ASAP7_75t_L g624 ( 
.A(n_466),
.B(n_416),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_492),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_478),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_497),
.Y(n_627)
);

OR2x6_ASAP7_75t_L g628 ( 
.A(n_500),
.B(n_395),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_460),
.B(n_404),
.Y(n_629)
);

BUFx2_ASAP7_75t_L g630 ( 
.A(n_500),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_531),
.B(n_432),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_487),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_531),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_578),
.Y(n_634)
);

NOR3xp33_ASAP7_75t_L g635 ( 
.A(n_454),
.B(n_197),
.C(n_211),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_470),
.A2(n_395),
.B1(n_450),
.B2(n_446),
.Y(n_636)
);

BUFx4f_ASAP7_75t_L g637 ( 
.A(n_500),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_467),
.B(n_384),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_467),
.B(n_384),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_502),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_473),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_461),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_463),
.B(n_392),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_503),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_471),
.B(n_392),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_505),
.B(n_392),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_514),
.B(n_400),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_528),
.B(n_480),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_546),
.B(n_400),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_500),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_507),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_546),
.B(n_400),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_468),
.B(n_401),
.Y(n_653)
);

INVxp67_ASAP7_75t_SL g654 ( 
.A(n_459),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_546),
.B(n_401),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_473),
.Y(n_656)
);

NOR2xp67_ASAP7_75t_L g657 ( 
.A(n_522),
.B(n_438),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_568),
.B(n_401),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_481),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_501),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_510),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_504),
.B(n_409),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_511),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_470),
.A2(n_395),
.B1(n_438),
.B2(n_451),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_506),
.B(n_409),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_491),
.B(n_482),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_559),
.B(n_409),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_549),
.Y(n_668)
);

O2A1O1Ixp5_ASAP7_75t_L g669 ( 
.A1(n_556),
.A2(n_417),
.B(n_411),
.C(n_412),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_501),
.B(n_324),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_560),
.B(n_411),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_578),
.B(n_411),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_481),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_562),
.B(n_412),
.Y(n_674)
);

NAND2xp33_ASAP7_75t_L g675 ( 
.A(n_590),
.B(n_412),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_494),
.B(n_417),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_587),
.B(n_417),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_501),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_551),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_567),
.B(n_438),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_501),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_600),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_587),
.B(n_390),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_590),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_470),
.A2(n_543),
.B1(n_590),
.B2(n_584),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_552),
.Y(n_686)
);

HB1xp67_ASAP7_75t_L g687 ( 
.A(n_569),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_555),
.B(n_438),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_545),
.B(n_451),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_590),
.B(n_451),
.Y(n_690)
);

AOI22x1_ASAP7_75t_L g691 ( 
.A1(n_593),
.A2(n_414),
.B1(n_403),
.B2(n_390),
.Y(n_691)
);

NAND3xp33_ASAP7_75t_L g692 ( 
.A(n_476),
.B(n_216),
.C(n_215),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_590),
.B(n_390),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_488),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_596),
.B(n_414),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_569),
.B(n_390),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_569),
.B(n_336),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_593),
.B(n_390),
.Y(n_698)
);

INVx1_ASAP7_75t_SL g699 ( 
.A(n_523),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_600),
.B(n_390),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_456),
.B(n_220),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_478),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_488),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_569),
.B(n_350),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_537),
.B(n_390),
.Y(n_705)
);

O2A1O1Ixp5_ASAP7_75t_L g706 ( 
.A1(n_599),
.A2(n_419),
.B(n_424),
.C(n_420),
.Y(n_706)
);

AOI22xp5_ASAP7_75t_L g707 ( 
.A1(n_476),
.A2(n_286),
.B1(n_260),
.B2(n_194),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_553),
.A2(n_230),
.B1(n_267),
.B2(n_277),
.Y(n_708)
);

NAND3xp33_ASAP7_75t_L g709 ( 
.A(n_484),
.B(n_524),
.C(n_554),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_565),
.B(n_228),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_557),
.B(n_403),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_489),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_479),
.Y(n_713)
);

INVx1_ASAP7_75t_SL g714 ( 
.A(n_525),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_485),
.A2(n_410),
.B(n_403),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_550),
.B(n_403),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_493),
.B(n_236),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_580),
.B(n_403),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_579),
.A2(n_168),
.B1(n_253),
.B2(n_251),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_580),
.B(n_403),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_489),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_490),
.Y(n_722)
);

NOR3xp33_ASAP7_75t_L g723 ( 
.A(n_535),
.B(n_226),
.C(n_227),
.Y(n_723)
);

AO221x1_ASAP7_75t_L g724 ( 
.A1(n_530),
.A2(n_543),
.B1(n_234),
.B2(n_254),
.C(n_295),
.Y(n_724)
);

INVxp67_ASAP7_75t_L g725 ( 
.A(n_579),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_490),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_586),
.B(n_403),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_459),
.B(n_241),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_586),
.Y(n_729)
);

O2A1O1Ixp33_ASAP7_75t_L g730 ( 
.A1(n_597),
.A2(n_295),
.B(n_293),
.C(n_281),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_597),
.B(n_403),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_509),
.B(n_403),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_579),
.B(n_410),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_498),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_579),
.B(n_410),
.Y(n_735)
);

OR2x6_ASAP7_75t_L g736 ( 
.A(n_496),
.B(n_227),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_498),
.B(n_410),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_513),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_513),
.B(n_410),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_516),
.B(n_410),
.Y(n_740)
);

INVx4_ASAP7_75t_L g741 ( 
.A(n_479),
.Y(n_741)
);

OR2x6_ASAP7_75t_L g742 ( 
.A(n_496),
.B(n_252),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_SL g743 ( 
.A1(n_558),
.A2(n_282),
.B1(n_279),
.B2(n_270),
.Y(n_743)
);

OR2x6_ASAP7_75t_L g744 ( 
.A(n_558),
.B(n_252),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_516),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_485),
.B(n_410),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_485),
.B(n_499),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_543),
.A2(n_542),
.B1(n_576),
.B2(n_547),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_520),
.B(n_410),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_520),
.Y(n_750)
);

NAND3xp33_ASAP7_75t_L g751 ( 
.A(n_591),
.B(n_296),
.C(n_298),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_589),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_543),
.A2(n_244),
.B1(n_300),
.B2(n_247),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_599),
.B(n_410),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_599),
.B(n_428),
.Y(n_755)
);

O2A1O1Ixp5_ASAP7_75t_L g756 ( 
.A1(n_529),
.A2(n_419),
.B(n_424),
.C(n_420),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_529),
.A2(n_428),
.B1(n_254),
.B2(n_264),
.Y(n_757)
);

AND2x4_ASAP7_75t_L g758 ( 
.A(n_598),
.B(n_264),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_573),
.B(n_174),
.Y(n_759)
);

INVxp67_ASAP7_75t_R g760 ( 
.A(n_533),
.Y(n_760)
);

OAI22xp33_ASAP7_75t_L g761 ( 
.A1(n_577),
.A2(n_592),
.B1(n_595),
.B2(n_275),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_533),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_534),
.Y(n_763)
);

NOR2xp67_ASAP7_75t_SL g764 ( 
.A(n_499),
.B(n_275),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_499),
.B(n_301),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_518),
.B(n_428),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_518),
.B(n_302),
.Y(n_767)
);

INVx5_ASAP7_75t_L g768 ( 
.A(n_515),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_534),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_538),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_538),
.B(n_174),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_542),
.B(n_419),
.Y(n_772)
);

AO21x1_ASAP7_75t_L g773 ( 
.A1(n_629),
.A2(n_465),
.B(n_464),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_633),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_629),
.A2(n_518),
.B1(n_588),
.B2(n_585),
.Y(n_775)
);

INVxp67_ASAP7_75t_L g776 ( 
.A(n_607),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_602),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_614),
.B(n_547),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_602),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_633),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_614),
.B(n_548),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_604),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_642),
.B(n_521),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_621),
.B(n_643),
.Y(n_784)
);

AOI21x1_ASAP7_75t_L g785 ( 
.A1(n_766),
.A2(n_465),
.B(n_464),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_621),
.B(n_548),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_645),
.A2(n_571),
.B(n_574),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_605),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_699),
.B(n_521),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_771),
.B(n_571),
.Y(n_790)
);

BUFx4f_ASAP7_75t_L g791 ( 
.A(n_628),
.Y(n_791)
);

AO21x1_ASAP7_75t_L g792 ( 
.A1(n_611),
.A2(n_689),
.B(n_647),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_637),
.B(n_521),
.Y(n_793)
);

INVxp67_ASAP7_75t_L g794 ( 
.A(n_624),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_619),
.Y(n_795)
);

OAI21xp5_ASAP7_75t_L g796 ( 
.A1(n_706),
.A2(n_574),
.B(n_576),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_626),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_632),
.B(n_532),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_637),
.B(n_532),
.Y(n_799)
);

BUFx4f_ASAP7_75t_L g800 ( 
.A(n_628),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_766),
.A2(n_526),
.B(n_483),
.Y(n_801)
);

AO21x1_ASAP7_75t_L g802 ( 
.A1(n_647),
.A2(n_540),
.B(n_483),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_755),
.A2(n_653),
.B(n_646),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_755),
.A2(n_526),
.B(n_517),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_626),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_609),
.Y(n_806)
);

INVx2_ASAP7_75t_SL g807 ( 
.A(n_632),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_653),
.A2(n_720),
.B(n_718),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_714),
.B(n_532),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_727),
.A2(n_486),
.B(n_536),
.Y(n_810)
);

NOR3xp33_ASAP7_75t_L g811 ( 
.A(n_709),
.B(n_281),
.C(n_294),
.Y(n_811)
);

A2O1A1Ixp33_ASAP7_75t_L g812 ( 
.A1(n_676),
.A2(n_519),
.B(n_472),
.C(n_477),
.Y(n_812)
);

A2O1A1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_676),
.A2(n_519),
.B(n_472),
.C(n_477),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_626),
.Y(n_814)
);

BUFx2_ASAP7_75t_L g815 ( 
.A(n_628),
.Y(n_815)
);

BUFx12f_ASAP7_75t_L g816 ( 
.A(n_660),
.Y(n_816)
);

NOR2xp67_ASAP7_75t_L g817 ( 
.A(n_678),
.B(n_419),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_620),
.B(n_572),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_623),
.B(n_572),
.Y(n_819)
);

AO21x2_ASAP7_75t_L g820 ( 
.A1(n_657),
.A2(n_564),
.B(n_527),
.Y(n_820)
);

INVx2_ASAP7_75t_SL g821 ( 
.A(n_670),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_610),
.Y(n_822)
);

OAI21xp33_ASAP7_75t_SL g823 ( 
.A1(n_658),
.A2(n_541),
.B(n_564),
.Y(n_823)
);

A2O1A1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_696),
.A2(n_527),
.B(n_486),
.C(n_469),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_731),
.A2(n_541),
.B(n_536),
.Y(n_825)
);

NAND2x1_ASAP7_75t_L g826 ( 
.A(n_634),
.B(n_682),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_613),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_681),
.Y(n_828)
);

BUFx3_ASAP7_75t_L g829 ( 
.A(n_697),
.Y(n_829)
);

BUFx2_ASAP7_75t_L g830 ( 
.A(n_630),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_725),
.B(n_544),
.Y(n_831)
);

BUFx3_ASAP7_75t_L g832 ( 
.A(n_650),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_684),
.B(n_572),
.Y(n_833)
);

OA22x2_ASAP7_75t_L g834 ( 
.A1(n_724),
.A2(n_307),
.B1(n_303),
.B2(n_293),
.Y(n_834)
);

AOI22xp5_ASAP7_75t_L g835 ( 
.A1(n_696),
.A2(n_575),
.B1(n_588),
.B2(n_585),
.Y(n_835)
);

INVx2_ASAP7_75t_SL g836 ( 
.A(n_704),
.Y(n_836)
);

OR2x6_ASAP7_75t_L g837 ( 
.A(n_687),
.B(n_544),
.Y(n_837)
);

INVx4_ASAP7_75t_L g838 ( 
.A(n_603),
.Y(n_838)
);

OAI22xp5_ASAP7_75t_L g839 ( 
.A1(n_638),
.A2(n_575),
.B1(n_588),
.B2(n_585),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_733),
.Y(n_840)
);

AO21x2_ASAP7_75t_L g841 ( 
.A1(n_680),
.A2(n_469),
.B(n_517),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_641),
.Y(n_842)
);

INVx5_ASAP7_75t_L g843 ( 
.A(n_603),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_684),
.B(n_575),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_737),
.A2(n_540),
.B(n_582),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_739),
.A2(n_582),
.B(n_591),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_603),
.B(n_582),
.Y(n_847)
);

AOI21x1_ASAP7_75t_L g848 ( 
.A1(n_764),
.A2(n_420),
.B(n_424),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_740),
.A2(n_544),
.B(n_583),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_749),
.A2(n_561),
.B(n_583),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_625),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_608),
.B(n_515),
.Y(n_852)
);

BUFx8_ASAP7_75t_SL g853 ( 
.A(n_759),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_639),
.B(n_515),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_648),
.B(n_561),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_627),
.B(n_561),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_656),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_626),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_640),
.B(n_583),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_656),
.Y(n_860)
);

OAI21xp5_ASAP7_75t_L g861 ( 
.A1(n_756),
.A2(n_512),
.B(n_508),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_644),
.B(n_508),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_666),
.B(n_174),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_754),
.A2(n_594),
.B(n_581),
.Y(n_864)
);

INVx1_ASAP7_75t_SL g865 ( 
.A(n_752),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_754),
.A2(n_594),
.B(n_581),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_651),
.B(n_508),
.Y(n_867)
);

NOR3xp33_ASAP7_75t_L g868 ( 
.A(n_701),
.B(n_512),
.C(n_419),
.Y(n_868)
);

AOI21x1_ASAP7_75t_L g869 ( 
.A1(n_672),
.A2(n_420),
.B(n_424),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_715),
.A2(n_746),
.B(n_732),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_661),
.B(n_508),
.Y(n_871)
);

NOR2x1_ASAP7_75t_L g872 ( 
.A(n_736),
.B(n_242),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_663),
.B(n_508),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_668),
.Y(n_874)
);

AO21x1_ASAP7_75t_L g875 ( 
.A1(n_618),
.A2(n_242),
.B(n_422),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_746),
.A2(n_594),
.B(n_581),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_743),
.B(n_495),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_601),
.B(n_398),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_683),
.A2(n_594),
.B(n_581),
.Y(n_879)
);

INVx4_ASAP7_75t_L g880 ( 
.A(n_603),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_683),
.A2(n_594),
.B(n_581),
.Y(n_881)
);

O2A1O1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_612),
.A2(n_398),
.B(n_406),
.C(n_407),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_679),
.B(n_686),
.Y(n_883)
);

NAND2x1p5_ASAP7_75t_L g884 ( 
.A(n_768),
.B(n_398),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_659),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_698),
.A2(n_563),
.B(n_495),
.Y(n_886)
);

O2A1O1Ixp33_ASAP7_75t_SL g887 ( 
.A1(n_698),
.A2(n_407),
.B(n_406),
.C(n_398),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_765),
.B(n_495),
.Y(n_888)
);

AO21x1_ASAP7_75t_L g889 ( 
.A1(n_716),
.A2(n_422),
.B(n_495),
.Y(n_889)
);

O2A1O1Ixp5_ASAP7_75t_SL g890 ( 
.A1(n_753),
.A2(n_407),
.B(n_406),
.C(n_398),
.Y(n_890)
);

OAI21xp33_ASAP7_75t_SL g891 ( 
.A1(n_685),
.A2(n_406),
.B(n_407),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_700),
.A2(n_563),
.B(n_495),
.Y(n_892)
);

AND2x2_ASAP7_75t_SL g893 ( 
.A(n_685),
.B(n_563),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_702),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_736),
.A2(n_742),
.B1(n_744),
.B2(n_615),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_601),
.B(n_406),
.Y(n_896)
);

NOR2xp67_ASAP7_75t_L g897 ( 
.A(n_719),
.B(n_407),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_765),
.B(n_563),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_717),
.B(n_563),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_768),
.B(n_761),
.Y(n_900)
);

NOR2xp67_ASAP7_75t_L g901 ( 
.A(n_705),
.B(n_160),
.Y(n_901)
);

NOR3xp33_ASAP7_75t_L g902 ( 
.A(n_708),
.B(n_172),
.C(n_304),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_729),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_702),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_758),
.B(n_422),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_736),
.B(n_162),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_758),
.B(n_422),
.Y(n_907)
);

NOR2xp67_ASAP7_75t_L g908 ( 
.A(n_692),
.B(n_163),
.Y(n_908)
);

OAI21xp5_ASAP7_75t_L g909 ( 
.A1(n_747),
.A2(n_175),
.B(n_297),
.Y(n_909)
);

INVx11_ASAP7_75t_L g910 ( 
.A(n_723),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_700),
.A2(n_422),
.B(n_169),
.Y(n_911)
);

OAI21xp5_ASAP7_75t_L g912 ( 
.A1(n_747),
.A2(n_291),
.B(n_289),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_711),
.A2(n_287),
.B(n_285),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_672),
.A2(n_284),
.B(n_278),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_631),
.B(n_649),
.Y(n_915)
);

AOI22x1_ASAP7_75t_L g916 ( 
.A1(n_634),
.A2(n_682),
.B1(n_734),
.B2(n_762),
.Y(n_916)
);

AO21x1_ASAP7_75t_L g917 ( 
.A1(n_688),
.A2(n_144),
.B(n_152),
.Y(n_917)
);

OAI21xp5_ASAP7_75t_L g918 ( 
.A1(n_677),
.A2(n_276),
.B(n_271),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_677),
.A2(n_269),
.B(n_268),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_652),
.B(n_655),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_617),
.B(n_263),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_659),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_662),
.A2(n_259),
.B(n_258),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_665),
.A2(n_249),
.B(n_245),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_742),
.B(n_744),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_742),
.B(n_243),
.Y(n_926)
);

O2A1O1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_667),
.A2(n_20),
.B(n_22),
.C(n_24),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_671),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_735),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_768),
.B(n_616),
.Y(n_930)
);

O2A1O1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_674),
.A2(n_22),
.B(n_26),
.C(n_28),
.Y(n_931)
);

INVx2_ASAP7_75t_SL g932 ( 
.A(n_601),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_772),
.A2(n_240),
.B(n_233),
.Y(n_933)
);

CKINVDCx6p67_ASAP7_75t_R g934 ( 
.A(n_744),
.Y(n_934)
);

O2A1O1Ixp5_ASAP7_75t_L g935 ( 
.A1(n_767),
.A2(n_29),
.B(n_36),
.C(n_41),
.Y(n_935)
);

INVx1_ASAP7_75t_SL g936 ( 
.A(n_710),
.Y(n_936)
);

NAND2x1p5_ASAP7_75t_L g937 ( 
.A(n_768),
.B(n_124),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_616),
.B(n_232),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_675),
.A2(n_231),
.B(n_223),
.Y(n_939)
);

O2A1O1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_730),
.A2(n_29),
.B(n_41),
.C(n_43),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_693),
.A2(n_221),
.B(n_219),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_622),
.B(n_217),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_728),
.B(n_205),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_690),
.A2(n_203),
.B(n_201),
.Y(n_944)
);

AOI21x1_ASAP7_75t_L g945 ( 
.A1(n_673),
.A2(n_200),
.B(n_193),
.Y(n_945)
);

NOR3xp33_ASAP7_75t_L g946 ( 
.A(n_635),
.B(n_192),
.C(n_187),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_695),
.A2(n_770),
.B(n_769),
.Y(n_947)
);

HB1xp67_ASAP7_75t_L g948 ( 
.A(n_664),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_694),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_669),
.A2(n_183),
.B(n_180),
.Y(n_950)
);

OAI21xp5_ASAP7_75t_L g951 ( 
.A1(n_757),
.A2(n_176),
.B(n_98),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_694),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_695),
.B(n_47),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_703),
.A2(n_47),
.B(n_48),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_703),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_712),
.A2(n_49),
.B(n_50),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_622),
.B(n_50),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_712),
.A2(n_51),
.B(n_52),
.Y(n_958)
);

A2O1A1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_953),
.A2(n_707),
.B(n_757),
.C(n_748),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_784),
.A2(n_654),
.B(n_606),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_888),
.A2(n_741),
.B(n_769),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_794),
.B(n_760),
.Y(n_962)
);

O2A1O1Ixp5_ASAP7_75t_L g963 ( 
.A1(n_792),
.A2(n_741),
.B(n_763),
.C(n_726),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_895),
.B(n_636),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_776),
.B(n_636),
.Y(n_965)
);

INVx3_ASAP7_75t_L g966 ( 
.A(n_838),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_898),
.A2(n_770),
.B(n_763),
.Y(n_967)
);

AOI21x1_ASAP7_75t_L g968 ( 
.A1(n_803),
.A2(n_726),
.B(n_750),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_775),
.A2(n_722),
.B(n_750),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_934),
.B(n_722),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_777),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_786),
.A2(n_721),
.B(n_745),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_779),
.Y(n_973)
);

NAND2x2_ASAP7_75t_L g974 ( 
.A(n_807),
.B(n_52),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_782),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_928),
.B(n_748),
.Y(n_976)
);

AOI21xp33_ASAP7_75t_L g977 ( 
.A1(n_951),
.A2(n_745),
.B(n_738),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_778),
.A2(n_781),
.B(n_803),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_789),
.A2(n_751),
.B(n_738),
.C(n_713),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_822),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_791),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_816),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_809),
.B(n_702),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_893),
.A2(n_713),
.B1(n_702),
.B2(n_691),
.Y(n_984)
);

O2A1O1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_940),
.A2(n_713),
.B(n_57),
.C(n_60),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_783),
.B(n_713),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_890),
.A2(n_870),
.B(n_808),
.Y(n_987)
);

OAI21xp33_ASAP7_75t_SL g988 ( 
.A1(n_883),
.A2(n_835),
.B(n_920),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_821),
.B(n_55),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_827),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_SL g991 ( 
.A1(n_798),
.A2(n_61),
.B(n_85),
.C(n_90),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_818),
.B(n_99),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_903),
.A2(n_100),
.B1(n_102),
.B2(n_110),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_795),
.Y(n_994)
);

NOR3xp33_ASAP7_75t_SL g995 ( 
.A(n_927),
.B(n_931),
.C(n_924),
.Y(n_995)
);

AND3x1_ASAP7_75t_SL g996 ( 
.A(n_851),
.B(n_118),
.C(n_126),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_788),
.Y(n_997)
);

OAI21xp5_ASAP7_75t_L g998 ( 
.A1(n_870),
.A2(n_131),
.B(n_141),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_948),
.B(n_145),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_925),
.B(n_150),
.Y(n_1000)
);

BUFx4f_ASAP7_75t_L g1001 ( 
.A(n_774),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_843),
.B(n_791),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_829),
.B(n_830),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_832),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_806),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_874),
.B(n_906),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_815),
.B(n_774),
.Y(n_1007)
);

OAI21x1_ASAP7_75t_L g1008 ( 
.A1(n_801),
.A2(n_804),
.B(n_785),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_853),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_843),
.B(n_800),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_940),
.A2(n_902),
.B(n_931),
.C(n_927),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_949),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_840),
.B(n_915),
.Y(n_1013)
);

O2A1O1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_909),
.A2(n_912),
.B(n_811),
.C(n_813),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_955),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_843),
.B(n_800),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_774),
.B(n_780),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_780),
.B(n_936),
.Y(n_1018)
);

INVx4_ASAP7_75t_L g1019 ( 
.A(n_843),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_957),
.A2(n_819),
.B1(n_852),
.B2(n_854),
.Y(n_1020)
);

AOI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_836),
.A2(n_828),
.B1(n_877),
.B2(n_926),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_876),
.A2(n_808),
.B(n_849),
.Y(n_1022)
);

AOI22xp33_ASAP7_75t_L g1023 ( 
.A1(n_932),
.A2(n_834),
.B1(n_863),
.B2(n_878),
.Y(n_1023)
);

BUFx8_ASAP7_75t_L g1024 ( 
.A(n_780),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_842),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_910),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_876),
.A2(n_849),
.B(n_850),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_823),
.A2(n_943),
.B(n_899),
.C(n_923),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_865),
.B(n_896),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_793),
.B(n_799),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_838),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_923),
.A2(n_924),
.B(n_918),
.C(n_872),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_831),
.A2(n_900),
.B1(n_930),
.B2(n_837),
.Y(n_1033)
);

NOR2xp67_ASAP7_75t_SL g1034 ( 
.A(n_880),
.B(n_805),
.Y(n_1034)
);

INVxp67_ASAP7_75t_SL g1035 ( 
.A(n_905),
.Y(n_1035)
);

BUFx4f_ASAP7_75t_L g1036 ( 
.A(n_837),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_790),
.A2(n_859),
.B1(n_856),
.B2(n_839),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_929),
.B(n_831),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_837),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_921),
.B(n_938),
.Y(n_1040)
);

BUFx2_ASAP7_75t_SL g1041 ( 
.A(n_817),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_857),
.B(n_860),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_812),
.A2(n_846),
.B(n_845),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_885),
.B(n_922),
.Y(n_1044)
);

INVx3_ASAP7_75t_L g1045 ( 
.A(n_880),
.Y(n_1045)
);

NAND3xp33_ASAP7_75t_L g1046 ( 
.A(n_946),
.B(n_935),
.C(n_954),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_850),
.A2(n_825),
.B(n_810),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_942),
.B(n_797),
.Y(n_1048)
);

BUFx3_ASAP7_75t_L g1049 ( 
.A(n_805),
.Y(n_1049)
);

INVx2_ASAP7_75t_SL g1050 ( 
.A(n_805),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_810),
.A2(n_825),
.B(n_866),
.Y(n_1051)
);

BUFx8_ASAP7_75t_L g1052 ( 
.A(n_814),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_R g1053 ( 
.A(n_797),
.B(n_858),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_814),
.B(n_858),
.Y(n_1054)
);

INVx6_ASAP7_75t_L g1055 ( 
.A(n_814),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_864),
.A2(n_866),
.B(n_845),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_894),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_824),
.A2(n_958),
.B(n_956),
.C(n_954),
.Y(n_1058)
);

OA22x2_ASAP7_75t_L g1059 ( 
.A1(n_907),
.A2(n_950),
.B1(n_952),
.B2(n_873),
.Y(n_1059)
);

NOR2xp67_ASAP7_75t_L g1060 ( 
.A(n_894),
.B(n_904),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_956),
.A2(n_958),
.B1(n_834),
.B2(n_867),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_904),
.B(n_787),
.Y(n_1062)
);

AOI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_891),
.A2(n_897),
.B1(n_844),
.B2(n_833),
.Y(n_1063)
);

OAI21xp33_ASAP7_75t_L g1064 ( 
.A1(n_914),
.A2(n_919),
.B(n_862),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_882),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_787),
.B(n_947),
.Y(n_1066)
);

OAI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_846),
.A2(n_801),
.B(n_804),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_871),
.A2(n_855),
.B1(n_939),
.B2(n_916),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_947),
.B(n_773),
.Y(n_1069)
);

O2A1O1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_933),
.A2(n_887),
.B(n_913),
.C(n_802),
.Y(n_1070)
);

INVxp67_ASAP7_75t_L g1071 ( 
.A(n_908),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_868),
.B(n_884),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_864),
.A2(n_886),
.B(n_892),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_826),
.Y(n_1074)
);

BUFx2_ASAP7_75t_L g1075 ( 
.A(n_884),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_L g1076 ( 
.A1(n_901),
.A2(n_841),
.B1(n_820),
.B2(n_933),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_879),
.A2(n_886),
.B(n_892),
.Y(n_1077)
);

O2A1O1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_913),
.A2(n_944),
.B(n_847),
.C(n_911),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_841),
.B(n_820),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_945),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_879),
.A2(n_881),
.B(n_796),
.Y(n_1081)
);

AOI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_939),
.A2(n_917),
.B1(n_889),
.B2(n_937),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_937),
.Y(n_1083)
);

CKINVDCx10_ASAP7_75t_R g1084 ( 
.A(n_944),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_861),
.B(n_875),
.Y(n_1085)
);

O2A1O1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_911),
.A2(n_941),
.B(n_881),
.C(n_869),
.Y(n_1086)
);

AOI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_941),
.A2(n_604),
.B1(n_487),
.B2(n_539),
.Y(n_1087)
);

BUFx12f_ASAP7_75t_L g1088 ( 
.A(n_848),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_784),
.A2(n_898),
.B(n_888),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_782),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_SL g1091 ( 
.A1(n_782),
.A2(n_324),
.B1(n_350),
.B2(n_336),
.Y(n_1091)
);

HB1xp67_ASAP7_75t_L g1092 ( 
.A(n_776),
.Y(n_1092)
);

BUFx3_ASAP7_75t_L g1093 ( 
.A(n_782),
.Y(n_1093)
);

BUFx8_ASAP7_75t_SL g1094 ( 
.A(n_782),
.Y(n_1094)
);

INVx5_ASAP7_75t_L g1095 ( 
.A(n_843),
.Y(n_1095)
);

AOI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_953),
.A2(n_604),
.B1(n_487),
.B2(n_539),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_776),
.B(n_539),
.Y(n_1097)
);

O2A1O1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_784),
.A2(n_460),
.B(n_642),
.C(n_614),
.Y(n_1098)
);

OAI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_784),
.A2(n_953),
.B1(n_928),
.B2(n_629),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_801),
.A2(n_804),
.B(n_785),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_776),
.B(n_539),
.Y(n_1101)
);

O2A1O1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_784),
.A2(n_460),
.B(n_642),
.C(n_614),
.Y(n_1102)
);

INVx1_ASAP7_75t_SL g1103 ( 
.A(n_1004),
.Y(n_1103)
);

AND2x4_ASAP7_75t_L g1104 ( 
.A(n_981),
.B(n_1007),
.Y(n_1104)
);

AO31x2_ASAP7_75t_L g1105 ( 
.A1(n_1079),
.A2(n_1069),
.A3(n_1068),
.B(n_1061),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_971),
.Y(n_1106)
);

INVxp67_ASAP7_75t_SL g1107 ( 
.A(n_1099),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1012),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1099),
.A2(n_1089),
.B(n_988),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1096),
.B(n_1097),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_1029),
.B(n_1101),
.Y(n_1111)
);

NOR3xp33_ASAP7_75t_L g1112 ( 
.A(n_1011),
.B(n_1102),
.C(n_1098),
.Y(n_1112)
);

NAND3xp33_ASAP7_75t_L g1113 ( 
.A(n_995),
.B(n_1028),
.C(n_1040),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_968),
.A2(n_1100),
.B(n_1008),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_1014),
.A2(n_959),
.B(n_985),
.C(n_999),
.Y(n_1115)
);

O2A1O1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_1032),
.A2(n_1092),
.B(n_998),
.C(n_1058),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1015),
.Y(n_1117)
);

INVxp67_ASAP7_75t_L g1118 ( 
.A(n_1003),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_978),
.A2(n_1027),
.B(n_1047),
.Y(n_1119)
);

NOR2xp67_ASAP7_75t_SL g1120 ( 
.A(n_1009),
.B(n_975),
.Y(n_1120)
);

AO21x1_ASAP7_75t_L g1121 ( 
.A1(n_998),
.A2(n_999),
.B(n_1020),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_1030),
.A2(n_1046),
.B(n_1048),
.C(n_960),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1022),
.A2(n_1037),
.B(n_1068),
.Y(n_1123)
);

AO32x2_ASAP7_75t_L g1124 ( 
.A1(n_1061),
.A2(n_1020),
.A3(n_1037),
.B1(n_984),
.B2(n_993),
.Y(n_1124)
);

NOR2xp67_ASAP7_75t_L g1125 ( 
.A(n_1026),
.B(n_1095),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_1006),
.B(n_1095),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1051),
.A2(n_1066),
.B(n_1056),
.Y(n_1127)
);

OAI21xp5_ASAP7_75t_SL g1128 ( 
.A1(n_1087),
.A2(n_1023),
.B(n_993),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_1094),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1077),
.A2(n_1073),
.B(n_1081),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_980),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_L g1132 ( 
.A1(n_1091),
.A2(n_964),
.B1(n_965),
.B2(n_976),
.Y(n_1132)
);

BUFx10_ASAP7_75t_L g1133 ( 
.A(n_982),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_977),
.A2(n_992),
.B(n_1043),
.Y(n_1134)
);

AO31x2_ASAP7_75t_L g1135 ( 
.A1(n_1079),
.A2(n_1080),
.A3(n_967),
.B(n_1062),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1021),
.A2(n_1033),
.B1(n_1036),
.B2(n_1065),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_973),
.Y(n_1137)
);

NOR2xp67_ASAP7_75t_L g1138 ( 
.A(n_1095),
.B(n_981),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_1095),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_977),
.A2(n_1043),
.B(n_987),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1042),
.Y(n_1141)
);

OAI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_963),
.A2(n_969),
.B(n_1070),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1013),
.B(n_962),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1067),
.A2(n_1086),
.B(n_961),
.Y(n_1144)
);

NAND2xp33_ASAP7_75t_SL g1145 ( 
.A(n_1053),
.B(n_1034),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1042),
.Y(n_1146)
);

INVx1_ASAP7_75t_SL g1147 ( 
.A(n_1090),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_990),
.Y(n_1148)
);

NAND3xp33_ASAP7_75t_L g1149 ( 
.A(n_1063),
.B(n_1071),
.C(n_1076),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_1067),
.A2(n_972),
.B(n_1078),
.Y(n_1150)
);

CKINVDCx11_ASAP7_75t_R g1151 ( 
.A(n_1093),
.Y(n_1151)
);

AOI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_970),
.A2(n_1036),
.B1(n_1039),
.B2(n_1007),
.Y(n_1152)
);

INVx4_ASAP7_75t_L g1153 ( 
.A(n_1001),
.Y(n_1153)
);

INVx3_ASAP7_75t_SL g1154 ( 
.A(n_1017),
.Y(n_1154)
);

A2O1A1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_1064),
.A2(n_1082),
.B(n_979),
.C(n_1085),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1059),
.A2(n_984),
.B(n_1083),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_1018),
.B(n_1001),
.Y(n_1157)
);

INVx2_ASAP7_75t_SL g1158 ( 
.A(n_1024),
.Y(n_1158)
);

INVx1_ASAP7_75t_SL g1159 ( 
.A(n_1017),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_986),
.A2(n_983),
.B(n_991),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_1024),
.Y(n_1161)
);

INVx1_ASAP7_75t_SL g1162 ( 
.A(n_1055),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1035),
.A2(n_1072),
.B(n_1074),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_SL g1164 ( 
.A(n_1052),
.B(n_1019),
.Y(n_1164)
);

A2O1A1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_997),
.A2(n_1005),
.B(n_1000),
.C(n_1038),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_989),
.B(n_1049),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1054),
.A2(n_1060),
.B(n_1045),
.Y(n_1167)
);

OAI22xp33_ASAP7_75t_L g1168 ( 
.A1(n_974),
.A2(n_1075),
.B1(n_1057),
.B2(n_1016),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_966),
.A2(n_1045),
.B(n_1031),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1025),
.Y(n_1170)
);

AO32x2_ASAP7_75t_L g1171 ( 
.A1(n_1050),
.A2(n_1019),
.A3(n_996),
.B1(n_1084),
.B2(n_1088),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_994),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_SL g1173 ( 
.A1(n_1055),
.A2(n_1041),
.B1(n_1057),
.B2(n_1031),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_1052),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1055),
.B(n_1057),
.Y(n_1175)
);

INVxp67_ASAP7_75t_SL g1176 ( 
.A(n_1044),
.Y(n_1176)
);

AOI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1002),
.A2(n_539),
.B1(n_1096),
.B2(n_604),
.Y(n_1177)
);

AO31x2_ASAP7_75t_L g1178 ( 
.A1(n_1010),
.A2(n_889),
.A3(n_1079),
.B(n_792),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_966),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_1094),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_968),
.A2(n_1100),
.B(n_1008),
.Y(n_1181)
);

NAND3xp33_ASAP7_75t_L g1182 ( 
.A(n_1099),
.B(n_1011),
.C(n_460),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1099),
.A2(n_642),
.B(n_784),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_980),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1096),
.B(n_642),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_981),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1096),
.B(n_642),
.Y(n_1187)
);

OAI22x1_ASAP7_75t_L g1188 ( 
.A1(n_1096),
.A2(n_1021),
.B1(n_1087),
.B2(n_539),
.Y(n_1188)
);

INVx4_ASAP7_75t_L g1189 ( 
.A(n_1095),
.Y(n_1189)
);

OAI22x1_ASAP7_75t_L g1190 ( 
.A1(n_1096),
.A2(n_1021),
.B1(n_1087),
.B2(n_539),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1099),
.A2(n_784),
.B(n_1089),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1099),
.A2(n_784),
.B(n_1089),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_1004),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1029),
.B(n_620),
.Y(n_1194)
);

AND2x4_ASAP7_75t_L g1195 ( 
.A(n_981),
.B(n_1007),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_980),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1012),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1099),
.A2(n_642),
.B(n_784),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_980),
.Y(n_1199)
);

INVx6_ASAP7_75t_SL g1200 ( 
.A(n_1017),
.Y(n_1200)
);

O2A1O1Ixp33_ASAP7_75t_SL g1201 ( 
.A1(n_1099),
.A2(n_784),
.B(n_1102),
.C(n_1098),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1099),
.A2(n_460),
.B(n_642),
.C(n_1098),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1096),
.B(n_642),
.Y(n_1203)
);

AND2x6_ASAP7_75t_L g1204 ( 
.A(n_981),
.B(n_895),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1012),
.Y(n_1205)
);

A2O1A1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1099),
.A2(n_1098),
.B(n_1102),
.C(n_1040),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1099),
.B(n_637),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1099),
.A2(n_784),
.B(n_1089),
.Y(n_1208)
);

OR2x6_ASAP7_75t_L g1209 ( 
.A(n_981),
.B(n_539),
.Y(n_1209)
);

NOR4xp25_ASAP7_75t_L g1210 ( 
.A(n_1011),
.B(n_1098),
.C(n_1102),
.D(n_940),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_971),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1096),
.B(n_642),
.Y(n_1212)
);

AOI221x1_ASAP7_75t_L g1213 ( 
.A1(n_1099),
.A2(n_998),
.B1(n_1028),
.B2(n_1061),
.C(n_953),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1099),
.A2(n_784),
.B(n_1089),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_968),
.A2(n_1100),
.B(n_1008),
.Y(n_1215)
);

OR2x2_ASAP7_75t_L g1216 ( 
.A(n_1029),
.B(n_607),
.Y(n_1216)
);

OA21x2_ASAP7_75t_L g1217 ( 
.A1(n_987),
.A2(n_1027),
.B(n_1022),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_968),
.A2(n_1100),
.B(n_1008),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_981),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1091),
.A2(n_893),
.B1(n_697),
.B2(n_324),
.Y(n_1220)
);

BUFx10_ASAP7_75t_L g1221 ( 
.A(n_975),
.Y(n_1221)
);

AOI221xp5_ASAP7_75t_SL g1222 ( 
.A1(n_1098),
.A2(n_460),
.B1(n_1102),
.B2(n_1011),
.C(n_474),
.Y(n_1222)
);

O2A1O1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1099),
.A2(n_460),
.B(n_642),
.C(n_1098),
.Y(n_1223)
);

INVx4_ASAP7_75t_L g1224 ( 
.A(n_1095),
.Y(n_1224)
);

INVx3_ASAP7_75t_L g1225 ( 
.A(n_1095),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1099),
.A2(n_1098),
.B(n_1102),
.C(n_1040),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1099),
.A2(n_784),
.B(n_1089),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1099),
.A2(n_784),
.B(n_1089),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_971),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1099),
.A2(n_784),
.B(n_1089),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_968),
.A2(n_1100),
.B(n_1008),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1096),
.B(n_642),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_968),
.A2(n_1100),
.B(n_1008),
.Y(n_1233)
);

INVx2_ASAP7_75t_SL g1234 ( 
.A(n_1024),
.Y(n_1234)
);

AOI31xp67_ASAP7_75t_L g1235 ( 
.A1(n_1059),
.A2(n_1082),
.A3(n_1066),
.B(n_1069),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_968),
.A2(n_1100),
.B(n_1008),
.Y(n_1236)
);

OAI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1099),
.A2(n_642),
.B(n_784),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1099),
.A2(n_784),
.B(n_1089),
.Y(n_1238)
);

NOR2x1_ASAP7_75t_R g1239 ( 
.A(n_1026),
.B(n_487),
.Y(n_1239)
);

O2A1O1Ixp5_ASAP7_75t_SL g1240 ( 
.A1(n_1080),
.A2(n_1061),
.B(n_987),
.C(n_998),
.Y(n_1240)
);

OR2x2_ASAP7_75t_L g1241 ( 
.A(n_1029),
.B(n_607),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_981),
.Y(n_1242)
);

AO32x2_ASAP7_75t_L g1243 ( 
.A1(n_1061),
.A2(n_1020),
.A3(n_932),
.B1(n_1099),
.B2(n_1068),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_971),
.Y(n_1244)
);

OA21x2_ASAP7_75t_L g1245 ( 
.A1(n_987),
.A2(n_1027),
.B(n_1022),
.Y(n_1245)
);

O2A1O1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1099),
.A2(n_460),
.B(n_642),
.C(n_1098),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1107),
.A2(n_1182),
.B1(n_1183),
.B2(n_1237),
.Y(n_1247)
);

INVx2_ASAP7_75t_SL g1248 ( 
.A(n_1174),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1220),
.A2(n_1132),
.B1(n_1190),
.B2(n_1188),
.Y(n_1249)
);

AOI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1128),
.A2(n_1136),
.B1(n_1110),
.B2(n_1204),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1109),
.A2(n_1123),
.B(n_1191),
.Y(n_1251)
);

CKINVDCx11_ASAP7_75t_R g1252 ( 
.A(n_1133),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_1154),
.Y(n_1253)
);

INVx6_ASAP7_75t_L g1254 ( 
.A(n_1221),
.Y(n_1254)
);

BUFx2_ASAP7_75t_SL g1255 ( 
.A(n_1125),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1113),
.A2(n_1149),
.B1(n_1194),
.B2(n_1207),
.Y(n_1256)
);

BUFx12f_ASAP7_75t_L g1257 ( 
.A(n_1161),
.Y(n_1257)
);

NAND2x1p5_ASAP7_75t_L g1258 ( 
.A(n_1189),
.B(n_1224),
.Y(n_1258)
);

BUFx2_ASAP7_75t_L g1259 ( 
.A(n_1193),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1198),
.A2(n_1212),
.B1(n_1203),
.B2(n_1232),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1204),
.A2(n_1121),
.B1(n_1111),
.B2(n_1244),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1204),
.A2(n_1172),
.B1(n_1211),
.B2(n_1229),
.Y(n_1262)
);

BUFx2_ASAP7_75t_SL g1263 ( 
.A(n_1158),
.Y(n_1263)
);

INVx8_ASAP7_75t_L g1264 ( 
.A(n_1209),
.Y(n_1264)
);

CKINVDCx20_ASAP7_75t_R g1265 ( 
.A(n_1129),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1148),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1204),
.A2(n_1137),
.B1(n_1185),
.B2(n_1187),
.Y(n_1267)
);

INVx3_ASAP7_75t_L g1268 ( 
.A(n_1224),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1184),
.Y(n_1269)
);

AO22x1_ASAP7_75t_L g1270 ( 
.A1(n_1104),
.A2(n_1195),
.B1(n_1234),
.B2(n_1242),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1170),
.Y(n_1271)
);

BUFx2_ASAP7_75t_SL g1272 ( 
.A(n_1153),
.Y(n_1272)
);

OAI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1213),
.A2(n_1177),
.B1(n_1209),
.B2(n_1216),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1196),
.Y(n_1274)
);

CKINVDCx20_ASAP7_75t_R g1275 ( 
.A(n_1180),
.Y(n_1275)
);

INVx6_ASAP7_75t_L g1276 ( 
.A(n_1221),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1241),
.A2(n_1141),
.B1(n_1146),
.B2(n_1112),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1199),
.Y(n_1278)
);

OAI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1118),
.A2(n_1143),
.B1(n_1147),
.B2(n_1103),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1141),
.A2(n_1146),
.B1(n_1176),
.B2(n_1166),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1108),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1206),
.A2(n_1226),
.B1(n_1115),
.B2(n_1238),
.Y(n_1282)
);

HB1xp67_ASAP7_75t_L g1283 ( 
.A(n_1117),
.Y(n_1283)
);

INVx1_ASAP7_75t_SL g1284 ( 
.A(n_1159),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1192),
.B(n_1208),
.Y(n_1285)
);

OAI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1164),
.A2(n_1152),
.B1(n_1153),
.B2(n_1168),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_SL g1287 ( 
.A1(n_1214),
.A2(n_1230),
.B1(n_1228),
.B2(n_1227),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1197),
.A2(n_1205),
.B1(n_1163),
.B2(n_1145),
.Y(n_1288)
);

AOI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1173),
.A2(n_1157),
.B1(n_1126),
.B2(n_1222),
.Y(n_1289)
);

INVx6_ASAP7_75t_L g1290 ( 
.A(n_1133),
.Y(n_1290)
);

CKINVDCx11_ASAP7_75t_R g1291 ( 
.A(n_1151),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_SL g1292 ( 
.A1(n_1124),
.A2(n_1171),
.B1(n_1134),
.B2(n_1140),
.Y(n_1292)
);

BUFx8_ASAP7_75t_L g1293 ( 
.A(n_1171),
.Y(n_1293)
);

OAI22x1_ASAP7_75t_SL g1294 ( 
.A1(n_1120),
.A2(n_1239),
.B1(n_1162),
.B2(n_1179),
.Y(n_1294)
);

CKINVDCx20_ASAP7_75t_R g1295 ( 
.A(n_1186),
.Y(n_1295)
);

OAI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1202),
.A2(n_1246),
.B(n_1223),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1135),
.Y(n_1297)
);

BUFx2_ASAP7_75t_SL g1298 ( 
.A(n_1138),
.Y(n_1298)
);

CKINVDCx11_ASAP7_75t_R g1299 ( 
.A(n_1186),
.Y(n_1299)
);

BUFx6f_ASAP7_75t_L g1300 ( 
.A(n_1219),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1210),
.B(n_1122),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_SL g1302 ( 
.A1(n_1124),
.A2(n_1156),
.B1(n_1243),
.B2(n_1195),
.Y(n_1302)
);

CKINVDCx20_ASAP7_75t_R g1303 ( 
.A(n_1219),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_SL g1304 ( 
.A(n_1104),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1243),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1200),
.A2(n_1242),
.B1(n_1219),
.B2(n_1160),
.Y(n_1306)
);

INVxp67_ASAP7_75t_SL g1307 ( 
.A(n_1217),
.Y(n_1307)
);

CKINVDCx16_ASAP7_75t_R g1308 ( 
.A(n_1242),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1116),
.A2(n_1155),
.B1(n_1165),
.B2(n_1124),
.Y(n_1309)
);

INVx4_ASAP7_75t_L g1310 ( 
.A(n_1139),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1175),
.A2(n_1142),
.B1(n_1167),
.B2(n_1225),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1243),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1144),
.A2(n_1127),
.B1(n_1169),
.B2(n_1201),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1119),
.A2(n_1130),
.B1(n_1217),
.B2(n_1245),
.Y(n_1314)
);

CKINVDCx16_ASAP7_75t_R g1315 ( 
.A(n_1139),
.Y(n_1315)
);

BUFx8_ASAP7_75t_L g1316 ( 
.A(n_1225),
.Y(n_1316)
);

INVx6_ASAP7_75t_L g1317 ( 
.A(n_1235),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_1178),
.Y(n_1318)
);

INVx6_ASAP7_75t_L g1319 ( 
.A(n_1240),
.Y(n_1319)
);

INVx4_ASAP7_75t_L g1320 ( 
.A(n_1245),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1105),
.Y(n_1321)
);

INVxp67_ASAP7_75t_SL g1322 ( 
.A(n_1150),
.Y(n_1322)
);

BUFx2_ASAP7_75t_L g1323 ( 
.A(n_1105),
.Y(n_1323)
);

CKINVDCx6p67_ASAP7_75t_R g1324 ( 
.A(n_1114),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1181),
.A2(n_1215),
.B1(n_1218),
.B2(n_1231),
.Y(n_1325)
);

INVxp67_ASAP7_75t_L g1326 ( 
.A(n_1233),
.Y(n_1326)
);

BUFx6f_ASAP7_75t_L g1327 ( 
.A(n_1236),
.Y(n_1327)
);

HB1xp67_ASAP7_75t_L g1328 ( 
.A(n_1105),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1131),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1131),
.Y(n_1330)
);

BUFx6f_ASAP7_75t_L g1331 ( 
.A(n_1154),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1220),
.A2(n_893),
.B1(n_601),
.B2(n_1132),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1107),
.A2(n_1099),
.B1(n_1182),
.B2(n_1183),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1111),
.B(n_1194),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_1129),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1220),
.A2(n_893),
.B1(n_601),
.B2(n_1132),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1131),
.Y(n_1337)
);

CKINVDCx11_ASAP7_75t_R g1338 ( 
.A(n_1133),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_SL g1339 ( 
.A1(n_1182),
.A2(n_893),
.B1(n_601),
.B2(n_932),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1131),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1107),
.A2(n_1099),
.B1(n_1182),
.B2(n_1183),
.Y(n_1341)
);

AOI21xp33_ASAP7_75t_L g1342 ( 
.A1(n_1113),
.A2(n_1011),
.B(n_1099),
.Y(n_1342)
);

NAND2x1p5_ASAP7_75t_L g1343 ( 
.A(n_1189),
.B(n_1036),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_SL g1344 ( 
.A1(n_1182),
.A2(n_893),
.B1(n_601),
.B2(n_932),
.Y(n_1344)
);

OAI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1128),
.A2(n_1096),
.B1(n_1110),
.B2(n_895),
.Y(n_1345)
);

BUFx6f_ASAP7_75t_L g1346 ( 
.A(n_1154),
.Y(n_1346)
);

CKINVDCx20_ASAP7_75t_R g1347 ( 
.A(n_1129),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1131),
.Y(n_1348)
);

NAND2x1p5_ASAP7_75t_L g1349 ( 
.A(n_1189),
.B(n_1036),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1106),
.Y(n_1350)
);

INVx2_ASAP7_75t_SL g1351 ( 
.A(n_1174),
.Y(n_1351)
);

CKINVDCx20_ASAP7_75t_R g1352 ( 
.A(n_1129),
.Y(n_1352)
);

BUFx12f_ASAP7_75t_L g1353 ( 
.A(n_1161),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1131),
.Y(n_1354)
);

INVx4_ASAP7_75t_L g1355 ( 
.A(n_1161),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1220),
.A2(n_893),
.B1(n_601),
.B2(n_1132),
.Y(n_1356)
);

AOI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1128),
.A2(n_1096),
.B1(n_539),
.B2(n_1188),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1220),
.A2(n_893),
.B1(n_601),
.B2(n_1132),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1106),
.Y(n_1359)
);

BUFx6f_ASAP7_75t_L g1360 ( 
.A(n_1154),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1281),
.Y(n_1361)
);

INVx3_ASAP7_75t_L g1362 ( 
.A(n_1320),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1305),
.B(n_1312),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1357),
.A2(n_1250),
.B1(n_1260),
.B2(n_1345),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1283),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1297),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1259),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1323),
.B(n_1260),
.Y(n_1368)
);

NOR2x1_ASAP7_75t_R g1369 ( 
.A(n_1291),
.B(n_1252),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1321),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1302),
.B(n_1292),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1321),
.Y(n_1372)
);

INVxp67_ASAP7_75t_L g1373 ( 
.A(n_1334),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1251),
.A2(n_1314),
.B(n_1325),
.Y(n_1374)
);

BUFx12f_ASAP7_75t_L g1375 ( 
.A(n_1338),
.Y(n_1375)
);

OAI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1342),
.A2(n_1282),
.B(n_1341),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1328),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1328),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1266),
.Y(n_1379)
);

AND2x4_ASAP7_75t_L g1380 ( 
.A(n_1320),
.B(n_1307),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1269),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1251),
.A2(n_1314),
.B(n_1325),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1274),
.Y(n_1383)
);

INVx1_ASAP7_75t_SL g1384 ( 
.A(n_1295),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1278),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1329),
.Y(n_1386)
);

BUFx2_ASAP7_75t_L g1387 ( 
.A(n_1324),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1330),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1302),
.B(n_1292),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1277),
.B(n_1301),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1337),
.Y(n_1391)
);

INVx3_ASAP7_75t_L g1392 ( 
.A(n_1327),
.Y(n_1392)
);

AOI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1313),
.A2(n_1285),
.B(n_1282),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1340),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1348),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1285),
.A2(n_1313),
.B(n_1296),
.Y(n_1396)
);

INVx3_ASAP7_75t_L g1397 ( 
.A(n_1317),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1326),
.Y(n_1398)
);

AO21x2_ASAP7_75t_L g1399 ( 
.A1(n_1309),
.A2(n_1307),
.B(n_1301),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1318),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1354),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1294),
.B(n_1355),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1309),
.B(n_1271),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1322),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1247),
.Y(n_1405)
);

INVx1_ASAP7_75t_SL g1406 ( 
.A(n_1303),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1322),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1333),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1296),
.B(n_1310),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1333),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1247),
.B(n_1267),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1341),
.A2(n_1288),
.B(n_1311),
.Y(n_1412)
);

CKINVDCx6p67_ASAP7_75t_R g1413 ( 
.A(n_1257),
.Y(n_1413)
);

BUFx4f_ASAP7_75t_L g1414 ( 
.A(n_1343),
.Y(n_1414)
);

OAI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1342),
.A2(n_1287),
.B(n_1289),
.Y(n_1415)
);

AOI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1249),
.A2(n_1332),
.B1(n_1358),
.B2(n_1356),
.Y(n_1416)
);

OAI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1287),
.A2(n_1273),
.B(n_1256),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1261),
.A2(n_1306),
.B(n_1258),
.Y(n_1418)
);

INVx2_ASAP7_75t_SL g1419 ( 
.A(n_1315),
.Y(n_1419)
);

AO21x2_ASAP7_75t_L g1420 ( 
.A1(n_1286),
.A2(n_1279),
.B(n_1359),
.Y(n_1420)
);

AO21x2_ASAP7_75t_L g1421 ( 
.A1(n_1350),
.A2(n_1319),
.B(n_1344),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1284),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1319),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1280),
.B(n_1284),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1264),
.B(n_1308),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1293),
.Y(n_1426)
);

INVx2_ASAP7_75t_SL g1427 ( 
.A(n_1316),
.Y(n_1427)
);

AO21x2_ASAP7_75t_L g1428 ( 
.A1(n_1339),
.A2(n_1344),
.B(n_1262),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1268),
.Y(n_1429)
);

AO21x2_ASAP7_75t_L g1430 ( 
.A1(n_1339),
.A2(n_1336),
.B(n_1270),
.Y(n_1430)
);

INVxp67_ASAP7_75t_L g1431 ( 
.A(n_1263),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1349),
.A2(n_1255),
.B(n_1316),
.Y(n_1432)
);

OA21x2_ASAP7_75t_L g1433 ( 
.A1(n_1248),
.A2(n_1351),
.B(n_1300),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1253),
.B(n_1360),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1298),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1399),
.B(n_1360),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1399),
.B(n_1360),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1399),
.B(n_1253),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1363),
.B(n_1253),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1365),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1363),
.B(n_1331),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1376),
.A2(n_1331),
.B(n_1346),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1368),
.B(n_1331),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1364),
.A2(n_1254),
.B1(n_1276),
.B2(n_1290),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1371),
.B(n_1346),
.Y(n_1445)
);

AND2x6_ASAP7_75t_L g1446 ( 
.A(n_1403),
.B(n_1346),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1431),
.B(n_1355),
.Y(n_1447)
);

INVx3_ASAP7_75t_L g1448 ( 
.A(n_1380),
.Y(n_1448)
);

NOR2x1_ASAP7_75t_SL g1449 ( 
.A(n_1368),
.B(n_1272),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1371),
.B(n_1254),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1387),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1415),
.A2(n_1304),
.B(n_1299),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1389),
.B(n_1276),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_SL g1454 ( 
.A1(n_1375),
.A2(n_1265),
.B1(n_1275),
.B2(n_1352),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1365),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1389),
.B(n_1290),
.Y(n_1456)
);

AOI221xp5_ASAP7_75t_L g1457 ( 
.A1(n_1390),
.A2(n_1335),
.B1(n_1347),
.B2(n_1353),
.C(n_1417),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1379),
.B(n_1381),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1401),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1422),
.B(n_1367),
.Y(n_1460)
);

AOI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1405),
.A2(n_1411),
.B(n_1396),
.Y(n_1461)
);

OAI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1412),
.A2(n_1408),
.B(n_1410),
.Y(n_1462)
);

O2A1O1Ixp33_ASAP7_75t_SL g1463 ( 
.A1(n_1408),
.A2(n_1410),
.B(n_1427),
.C(n_1419),
.Y(n_1463)
);

OA21x2_ASAP7_75t_L g1464 ( 
.A1(n_1374),
.A2(n_1382),
.B(n_1396),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1370),
.B(n_1372),
.Y(n_1465)
);

OAI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1416),
.A2(n_1373),
.B1(n_1409),
.B2(n_1419),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1412),
.A2(n_1382),
.B(n_1374),
.Y(n_1467)
);

OAI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1393),
.A2(n_1409),
.B(n_1423),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1379),
.B(n_1381),
.Y(n_1469)
);

OAI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1393),
.A2(n_1409),
.B(n_1418),
.Y(n_1470)
);

OAI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1409),
.A2(n_1418),
.B(n_1432),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_SL g1472 ( 
.A(n_1369),
.B(n_1375),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1383),
.Y(n_1473)
);

OA21x2_ASAP7_75t_L g1474 ( 
.A1(n_1404),
.A2(n_1407),
.B(n_1378),
.Y(n_1474)
);

BUFx2_ASAP7_75t_L g1475 ( 
.A(n_1387),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1384),
.B(n_1406),
.Y(n_1476)
);

O2A1O1Ixp33_ASAP7_75t_SL g1477 ( 
.A1(n_1427),
.A2(n_1402),
.B(n_1435),
.C(n_1429),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1383),
.B(n_1385),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1370),
.B(n_1372),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1428),
.A2(n_1430),
.B1(n_1416),
.B2(n_1400),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1386),
.B(n_1391),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1380),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1388),
.B(n_1391),
.Y(n_1483)
);

AOI221xp5_ASAP7_75t_L g1484 ( 
.A1(n_1388),
.A2(n_1395),
.B1(n_1394),
.B2(n_1377),
.C(n_1361),
.Y(n_1484)
);

OAI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1362),
.A2(n_1392),
.B(n_1397),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1482),
.B(n_1448),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1459),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1480),
.A2(n_1428),
.B1(n_1430),
.B2(n_1421),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1482),
.B(n_1380),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1448),
.B(n_1398),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1474),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1474),
.Y(n_1492)
);

CKINVDCx20_ASAP7_75t_R g1493 ( 
.A(n_1454),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1461),
.B(n_1394),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1474),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1460),
.B(n_1395),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1464),
.B(n_1458),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1464),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1458),
.B(n_1469),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1473),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1457),
.A2(n_1424),
.B1(n_1414),
.B2(n_1426),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1462),
.B(n_1366),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1478),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1465),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1440),
.B(n_1433),
.Y(n_1505)
);

NOR2xp67_ASAP7_75t_L g1506 ( 
.A(n_1467),
.B(n_1470),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1481),
.B(n_1483),
.Y(n_1507)
);

INVx3_ASAP7_75t_L g1508 ( 
.A(n_1485),
.Y(n_1508)
);

INVx3_ASAP7_75t_L g1509 ( 
.A(n_1485),
.Y(n_1509)
);

INVxp67_ASAP7_75t_SL g1510 ( 
.A(n_1465),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1504),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1494),
.B(n_1455),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1494),
.B(n_1436),
.Y(n_1513)
);

AOI21xp33_ASAP7_75t_L g1514 ( 
.A1(n_1501),
.A2(n_1437),
.B(n_1438),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1497),
.B(n_1439),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1510),
.B(n_1479),
.Y(n_1516)
);

NAND3xp33_ASAP7_75t_L g1517 ( 
.A(n_1506),
.B(n_1437),
.C(n_1438),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1497),
.B(n_1439),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1497),
.B(n_1499),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_1493),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1491),
.Y(n_1521)
);

NAND2x1_ASAP7_75t_L g1522 ( 
.A(n_1508),
.B(n_1446),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1504),
.Y(n_1523)
);

AO21x2_ASAP7_75t_L g1524 ( 
.A1(n_1492),
.A2(n_1468),
.B(n_1471),
.Y(n_1524)
);

NOR3xp33_ASAP7_75t_L g1525 ( 
.A(n_1501),
.B(n_1444),
.C(n_1442),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1487),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1508),
.B(n_1446),
.Y(n_1527)
);

AND2x4_ASAP7_75t_L g1528 ( 
.A(n_1508),
.B(n_1446),
.Y(n_1528)
);

OAI21xp33_ASAP7_75t_L g1529 ( 
.A1(n_1488),
.A2(n_1466),
.B(n_1472),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1499),
.B(n_1441),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1491),
.Y(n_1531)
);

BUFx3_ASAP7_75t_L g1532 ( 
.A(n_1508),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1487),
.Y(n_1533)
);

NAND2x1_ASAP7_75t_L g1534 ( 
.A(n_1508),
.B(n_1446),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1499),
.B(n_1443),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1491),
.Y(n_1536)
);

NAND2x1p5_ASAP7_75t_L g1537 ( 
.A(n_1506),
.B(n_1433),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1507),
.B(n_1449),
.Y(n_1538)
);

BUFx3_ASAP7_75t_L g1539 ( 
.A(n_1509),
.Y(n_1539)
);

INVx1_ASAP7_75t_SL g1540 ( 
.A(n_1505),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1492),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1507),
.B(n_1486),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_L g1543 ( 
.A(n_1496),
.B(n_1451),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1488),
.A2(n_1420),
.B1(n_1445),
.B2(n_1421),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1507),
.B(n_1451),
.Y(n_1545)
);

NAND3xp33_ASAP7_75t_L g1546 ( 
.A(n_1506),
.B(n_1463),
.C(n_1484),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1487),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1511),
.B(n_1510),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1526),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1526),
.Y(n_1550)
);

AND2x4_ASAP7_75t_L g1551 ( 
.A(n_1527),
.B(n_1509),
.Y(n_1551)
);

INVx3_ASAP7_75t_L g1552 ( 
.A(n_1522),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1512),
.B(n_1500),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1519),
.B(n_1486),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1541),
.Y(n_1555)
);

NOR3xp33_ASAP7_75t_SL g1556 ( 
.A(n_1520),
.B(n_1447),
.C(n_1476),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1533),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1519),
.B(n_1486),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1521),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1519),
.B(n_1486),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1527),
.B(n_1509),
.Y(n_1561)
);

INVx2_ASAP7_75t_SL g1562 ( 
.A(n_1522),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1521),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1542),
.B(n_1489),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1542),
.B(n_1489),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1542),
.B(n_1489),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1533),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1515),
.B(n_1489),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1529),
.A2(n_1445),
.B1(n_1452),
.B2(n_1420),
.Y(n_1569)
);

NAND2x1_ASAP7_75t_L g1570 ( 
.A(n_1527),
.B(n_1509),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1511),
.B(n_1505),
.Y(n_1571)
);

INVx3_ASAP7_75t_L g1572 ( 
.A(n_1522),
.Y(n_1572)
);

OAI21x1_ASAP7_75t_L g1573 ( 
.A1(n_1534),
.A2(n_1509),
.B(n_1498),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1512),
.B(n_1523),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1521),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1547),
.Y(n_1576)
);

HB1xp67_ASAP7_75t_L g1577 ( 
.A(n_1541),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1518),
.B(n_1490),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1518),
.B(n_1503),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1574),
.B(n_1543),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1574),
.B(n_1523),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1552),
.B(n_1369),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1564),
.B(n_1538),
.Y(n_1583)
);

OAI21xp33_ASAP7_75t_L g1584 ( 
.A1(n_1556),
.A2(n_1546),
.B(n_1529),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1549),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1549),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1549),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1550),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1553),
.B(n_1543),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1564),
.B(n_1538),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1564),
.B(n_1565),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1553),
.B(n_1513),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1565),
.B(n_1538),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1559),
.Y(n_1594)
);

O2A1O1Ixp33_ASAP7_75t_SL g1595 ( 
.A1(n_1562),
.A2(n_1493),
.B(n_1546),
.C(n_1534),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1548),
.B(n_1513),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1565),
.B(n_1566),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1550),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1566),
.B(n_1545),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1569),
.A2(n_1544),
.B1(n_1514),
.B2(n_1524),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1555),
.Y(n_1601)
);

OAI21xp5_ASAP7_75t_SL g1602 ( 
.A1(n_1569),
.A2(n_1525),
.B(n_1517),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1556),
.B(n_1545),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1568),
.B(n_1530),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1568),
.B(n_1530),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1562),
.B(n_1528),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1555),
.B(n_1540),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1577),
.B(n_1540),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1577),
.B(n_1535),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1548),
.B(n_1516),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1550),
.Y(n_1611)
);

XNOR2xp5_ASAP7_75t_L g1612 ( 
.A(n_1562),
.B(n_1450),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1548),
.B(n_1516),
.Y(n_1613)
);

AND2x4_ASAP7_75t_L g1614 ( 
.A(n_1562),
.B(n_1528),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1557),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1579),
.B(n_1535),
.Y(n_1616)
);

INVx1_ASAP7_75t_SL g1617 ( 
.A(n_1571),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1559),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1557),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1557),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1584),
.B(n_1579),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1580),
.B(n_1589),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1602),
.B(n_1579),
.Y(n_1623)
);

NOR2x1_ASAP7_75t_L g1624 ( 
.A(n_1582),
.B(n_1552),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1596),
.B(n_1571),
.Y(n_1625)
);

NOR3xp33_ASAP7_75t_L g1626 ( 
.A(n_1603),
.B(n_1525),
.C(n_1517),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1617),
.B(n_1579),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1604),
.B(n_1568),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1596),
.B(n_1571),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_SL g1630 ( 
.A(n_1612),
.B(n_1552),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1604),
.B(n_1558),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1609),
.B(n_1496),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1601),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1612),
.B(n_1413),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1585),
.Y(n_1635)
);

NOR4xp25_ASAP7_75t_L g1636 ( 
.A(n_1600),
.B(n_1595),
.C(n_1607),
.D(n_1608),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1585),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1592),
.B(n_1496),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1586),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1586),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1610),
.B(n_1516),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1587),
.Y(n_1642)
);

NOR2xp67_ASAP7_75t_L g1643 ( 
.A(n_1606),
.B(n_1552),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1610),
.B(n_1567),
.Y(n_1644)
);

NAND4xp75_ASAP7_75t_SL g1645 ( 
.A(n_1591),
.B(n_1558),
.C(n_1560),
.D(n_1554),
.Y(n_1645)
);

INVx3_ASAP7_75t_L g1646 ( 
.A(n_1606),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1613),
.B(n_1567),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1605),
.B(n_1578),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1587),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1594),
.Y(n_1650)
);

INVx2_ASAP7_75t_SL g1651 ( 
.A(n_1606),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1605),
.B(n_1578),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1613),
.B(n_1578),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1588),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1591),
.B(n_1597),
.Y(n_1655)
);

NAND2x1p5_ASAP7_75t_L g1656 ( 
.A(n_1646),
.B(n_1534),
.Y(n_1656)
);

NAND3xp33_ASAP7_75t_L g1657 ( 
.A(n_1626),
.B(n_1598),
.C(n_1588),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1646),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1635),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1622),
.B(n_1599),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1637),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_SL g1662 ( 
.A(n_1636),
.B(n_1626),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1646),
.Y(n_1663)
);

OAI22xp33_ASAP7_75t_L g1664 ( 
.A1(n_1623),
.A2(n_1514),
.B1(n_1537),
.B2(n_1502),
.Y(n_1664)
);

AOI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1630),
.A2(n_1621),
.B1(n_1524),
.B2(n_1544),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1634),
.B(n_1413),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1651),
.Y(n_1667)
);

INVx2_ASAP7_75t_SL g1668 ( 
.A(n_1651),
.Y(n_1668)
);

AOI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1630),
.A2(n_1524),
.B1(n_1537),
.B2(n_1450),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1639),
.Y(n_1670)
);

NOR2x1_ASAP7_75t_L g1671 ( 
.A(n_1634),
.B(n_1552),
.Y(n_1671)
);

OAI22xp33_ASAP7_75t_L g1672 ( 
.A1(n_1627),
.A2(n_1537),
.B1(n_1502),
.B2(n_1453),
.Y(n_1672)
);

A2O1A1Ixp33_ASAP7_75t_L g1673 ( 
.A1(n_1643),
.A2(n_1495),
.B(n_1492),
.C(n_1552),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1655),
.B(n_1597),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1633),
.B(n_1581),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1628),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1640),
.Y(n_1677)
);

O2A1O1Ixp33_ASAP7_75t_L g1678 ( 
.A1(n_1650),
.A2(n_1594),
.B(n_1618),
.C(n_1581),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1642),
.Y(n_1679)
);

NAND3xp33_ASAP7_75t_L g1680 ( 
.A(n_1649),
.B(n_1611),
.C(n_1598),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1662),
.B(n_1660),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1659),
.Y(n_1682)
);

AOI21xp33_ASAP7_75t_L g1683 ( 
.A1(n_1662),
.A2(n_1650),
.B(n_1654),
.Y(n_1683)
);

O2A1O1Ixp5_ASAP7_75t_L g1684 ( 
.A1(n_1664),
.A2(n_1653),
.B(n_1644),
.C(n_1647),
.Y(n_1684)
);

AOI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1665),
.A2(n_1524),
.B1(n_1537),
.B2(n_1453),
.Y(n_1685)
);

A2O1A1Ixp33_ASAP7_75t_L g1686 ( 
.A1(n_1669),
.A2(n_1678),
.B(n_1657),
.C(n_1675),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1661),
.Y(n_1687)
);

NOR2x1_ASAP7_75t_L g1688 ( 
.A(n_1666),
.B(n_1645),
.Y(n_1688)
);

INVx1_ASAP7_75t_SL g1689 ( 
.A(n_1667),
.Y(n_1689)
);

AOI211xp5_ASAP7_75t_L g1690 ( 
.A1(n_1664),
.A2(n_1625),
.B(n_1629),
.C(n_1641),
.Y(n_1690)
);

OAI221xp5_ASAP7_75t_L g1691 ( 
.A1(n_1673),
.A2(n_1624),
.B1(n_1618),
.B2(n_1536),
.C(n_1521),
.Y(n_1691)
);

AOI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1675),
.A2(n_1524),
.B1(n_1456),
.B2(n_1495),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1668),
.B(n_1628),
.Y(n_1693)
);

OAI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1672),
.A2(n_1495),
.B1(n_1572),
.B2(n_1652),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1674),
.B(n_1631),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_SL g1696 ( 
.A1(n_1680),
.A2(n_1575),
.B1(n_1563),
.B2(n_1559),
.Y(n_1696)
);

OAI22xp33_ASAP7_75t_L g1697 ( 
.A1(n_1672),
.A2(n_1572),
.B1(n_1648),
.B2(n_1638),
.Y(n_1697)
);

A2O1A1Ixp33_ASAP7_75t_L g1698 ( 
.A1(n_1673),
.A2(n_1572),
.B(n_1573),
.C(n_1532),
.Y(n_1698)
);

INVxp67_ASAP7_75t_SL g1699 ( 
.A(n_1666),
.Y(n_1699)
);

XNOR2xp5_ASAP7_75t_L g1700 ( 
.A(n_1681),
.B(n_1699),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1695),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1682),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1687),
.Y(n_1703)
);

AOI211xp5_ASAP7_75t_L g1704 ( 
.A1(n_1686),
.A2(n_1663),
.B(n_1658),
.C(n_1679),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1693),
.Y(n_1705)
);

INVx1_ASAP7_75t_SL g1706 ( 
.A(n_1689),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1684),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1683),
.Y(n_1708)
);

NOR4xp25_ASAP7_75t_L g1709 ( 
.A(n_1691),
.B(n_1677),
.C(n_1670),
.D(n_1676),
.Y(n_1709)
);

NAND3xp33_ASAP7_75t_SL g1710 ( 
.A(n_1709),
.B(n_1690),
.C(n_1696),
.Y(n_1710)
);

NOR2xp67_ASAP7_75t_L g1711 ( 
.A(n_1700),
.B(n_1572),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1700),
.B(n_1688),
.Y(n_1712)
);

A2O1A1Ixp33_ASAP7_75t_L g1713 ( 
.A1(n_1707),
.A2(n_1708),
.B(n_1685),
.C(n_1704),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1706),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1701),
.B(n_1631),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_SL g1716 ( 
.A(n_1705),
.B(n_1671),
.Y(n_1716)
);

NOR4xp25_ASAP7_75t_L g1717 ( 
.A(n_1707),
.B(n_1698),
.C(n_1697),
.D(n_1694),
.Y(n_1717)
);

NOR2x1_ASAP7_75t_L g1718 ( 
.A(n_1702),
.B(n_1645),
.Y(n_1718)
);

OAI21xp5_ASAP7_75t_L g1719 ( 
.A1(n_1710),
.A2(n_1696),
.B(n_1703),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_R g1720 ( 
.A(n_1714),
.B(n_1702),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1715),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1713),
.A2(n_1656),
.B1(n_1692),
.B2(n_1606),
.Y(n_1722)
);

OAI211xp5_ASAP7_75t_L g1723 ( 
.A1(n_1717),
.A2(n_1572),
.B(n_1570),
.C(n_1620),
.Y(n_1723)
);

NAND4xp25_ASAP7_75t_L g1724 ( 
.A(n_1719),
.B(n_1712),
.C(n_1718),
.D(n_1711),
.Y(n_1724)
);

AOI211xp5_ASAP7_75t_L g1725 ( 
.A1(n_1723),
.A2(n_1716),
.B(n_1614),
.C(n_1572),
.Y(n_1725)
);

O2A1O1Ixp33_ASAP7_75t_L g1726 ( 
.A1(n_1722),
.A2(n_1656),
.B(n_1611),
.C(n_1620),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1721),
.B(n_1614),
.Y(n_1727)
);

AOI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1720),
.A2(n_1614),
.B1(n_1619),
.B2(n_1615),
.Y(n_1728)
);

AOI221xp5_ASAP7_75t_L g1729 ( 
.A1(n_1719),
.A2(n_1615),
.B1(n_1619),
.B2(n_1559),
.C(n_1575),
.Y(n_1729)
);

NAND4xp75_ASAP7_75t_L g1730 ( 
.A(n_1727),
.B(n_1434),
.C(n_1456),
.D(n_1590),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1728),
.Y(n_1731)
);

NAND2x1p5_ASAP7_75t_L g1732 ( 
.A(n_1724),
.B(n_1475),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1729),
.B(n_1632),
.Y(n_1733)
);

AOI22xp5_ASAP7_75t_L g1734 ( 
.A1(n_1725),
.A2(n_1551),
.B1(n_1561),
.B2(n_1575),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1733),
.B(n_1616),
.Y(n_1735)
);

OAI321xp33_ASAP7_75t_L g1736 ( 
.A1(n_1732),
.A2(n_1731),
.A3(n_1726),
.B1(n_1734),
.B2(n_1730),
.C(n_1475),
.Y(n_1736)
);

NAND3x1_ASAP7_75t_L g1737 ( 
.A(n_1731),
.B(n_1593),
.C(n_1590),
.Y(n_1737)
);

OAI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1737),
.A2(n_1570),
.B1(n_1551),
.B2(n_1561),
.Y(n_1738)
);

AO22x2_ASAP7_75t_SL g1739 ( 
.A1(n_1738),
.A2(n_1736),
.B1(n_1735),
.B2(n_1583),
.Y(n_1739)
);

INVxp67_ASAP7_75t_L g1740 ( 
.A(n_1739),
.Y(n_1740)
);

O2A1O1Ixp33_ASAP7_75t_SL g1741 ( 
.A1(n_1739),
.A2(n_1570),
.B(n_1567),
.C(n_1576),
.Y(n_1741)
);

BUFx2_ASAP7_75t_L g1742 ( 
.A(n_1740),
.Y(n_1742)
);

NAND2x1_ASAP7_75t_L g1743 ( 
.A(n_1741),
.B(n_1599),
.Y(n_1743)
);

OAI21xp5_ASAP7_75t_L g1744 ( 
.A1(n_1742),
.A2(n_1563),
.B(n_1575),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1743),
.A2(n_1563),
.B1(n_1531),
.B2(n_1536),
.Y(n_1745)
);

XOR2xp5_ASAP7_75t_L g1746 ( 
.A(n_1744),
.B(n_1425),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1746),
.B(n_1745),
.Y(n_1747)
);

BUFx3_ASAP7_75t_L g1748 ( 
.A(n_1747),
.Y(n_1748)
);

OAI221xp5_ASAP7_75t_R g1749 ( 
.A1(n_1748),
.A2(n_1593),
.B1(n_1583),
.B2(n_1539),
.C(n_1532),
.Y(n_1749)
);

AOI211xp5_ASAP7_75t_L g1750 ( 
.A1(n_1749),
.A2(n_1463),
.B(n_1477),
.C(n_1425),
.Y(n_1750)
);


endmodule