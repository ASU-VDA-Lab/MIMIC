module fake_jpeg_3709_n_557 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_557);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_557;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_17),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx8_ASAP7_75t_SL g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx11_ASAP7_75t_SL g43 ( 
.A(n_2),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_57),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_59),
.Y(n_136)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_60),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_26),
.B(n_18),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_62),
.B(n_66),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_63),
.Y(n_139)
);

INVx11_ASAP7_75t_SL g64 ( 
.A(n_43),
.Y(n_64)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_64),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_38),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_69),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_26),
.B(n_16),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_67),
.Y(n_132)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_68),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_36),
.B(n_18),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_70),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g160 ( 
.A(n_74),
.Y(n_160)
);

BUFx10_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

BUFx10_ASAP7_75t_L g168 ( 
.A(n_75),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_36),
.B(n_0),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_77),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_0),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_78),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_79),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_82),
.Y(n_165)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_83),
.Y(n_133)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_30),
.B(n_45),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_84),
.B(n_91),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_85),
.Y(n_157)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_88),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_42),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_89),
.B(n_93),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_19),
.Y(n_90)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_90),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_41),
.B(n_1),
.Y(n_91)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

BUFx10_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_41),
.B(n_44),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_21),
.B(n_1),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_94),
.B(n_40),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_97),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_20),
.Y(n_98)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_98),
.Y(n_162)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_99),
.B(n_47),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_100),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_35),
.Y(n_101)
);

NAND2xp33_ASAP7_75t_SL g166 ( 
.A(n_101),
.B(n_105),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_28),
.Y(n_102)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_102),
.Y(n_164)
);

BUFx16f_ASAP7_75t_L g103 ( 
.A(n_35),
.Y(n_103)
);

BUFx10_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

BUFx10_ASAP7_75t_L g147 ( 
.A(n_104),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_20),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_57),
.B(n_37),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_113),
.B(n_117),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_21),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_93),
.A2(n_47),
.B1(n_22),
.B2(n_24),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_119),
.A2(n_121),
.B1(n_126),
.B2(n_128),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_58),
.B1(n_53),
.B2(n_80),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_81),
.A2(n_45),
.B1(n_22),
.B2(n_49),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_87),
.A2(n_45),
.B1(n_22),
.B2(n_49),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_91),
.A2(n_55),
.B1(n_79),
.B2(n_59),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_129),
.A2(n_135),
.B1(n_137),
.B2(n_150),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_24),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_130),
.B(n_143),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_84),
.A2(n_47),
.B1(n_22),
.B2(n_45),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_61),
.A2(n_40),
.B1(n_32),
.B2(n_33),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_148),
.B(n_103),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_63),
.A2(n_37),
.B1(n_32),
.B2(n_33),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_92),
.A2(n_46),
.B1(n_51),
.B2(n_49),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_151),
.A2(n_159),
.B1(n_157),
.B2(n_165),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_67),
.B(n_27),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_154),
.B(n_68),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_64),
.A2(n_51),
.B1(n_48),
.B2(n_46),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_82),
.A2(n_51),
.B1(n_48),
.B2(n_46),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_161),
.A2(n_29),
.B1(n_31),
.B2(n_48),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_84),
.B(n_27),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g219 ( 
.A(n_167),
.B(n_52),
.Y(n_219)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_169),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_83),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_170),
.B(n_172),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_127),
.B(n_73),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_173),
.Y(n_280)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_106),
.Y(n_174)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_174),
.Y(n_244)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_124),
.Y(n_175)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_175),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_149),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_177),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_127),
.A2(n_88),
.B1(n_70),
.B2(n_71),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_178),
.A2(n_168),
.B(n_112),
.Y(n_254)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_179),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_137),
.A2(n_105),
.B1(n_100),
.B2(n_98),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_181),
.A2(n_183),
.B1(n_8),
.B2(n_9),
.Y(n_282)
);

NAND2x1p5_ASAP7_75t_L g182 ( 
.A(n_148),
.B(n_103),
.Y(n_182)
);

OAI21xp33_ASAP7_75t_L g264 ( 
.A1(n_182),
.A2(n_195),
.B(n_204),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_85),
.B1(n_90),
.B2(n_95),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_133),
.Y(n_184)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_184),
.Y(n_248)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_108),
.Y(n_185)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_185),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_111),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_186),
.Y(n_257)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_141),
.Y(n_187)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_187),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_152),
.B(n_86),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_188),
.B(n_190),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_189),
.A2(n_201),
.B1(n_222),
.B2(n_138),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_110),
.B(n_31),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_156),
.Y(n_191)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_191),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_192),
.B(n_210),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_115),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_193),
.B(n_216),
.Y(n_238)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_134),
.Y(n_194)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_194),
.Y(n_252)
);

OR2x4_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_75),
.Y(n_195)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_145),
.Y(n_197)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_197),
.Y(n_256)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_146),
.Y(n_198)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_198),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_116),
.B(n_31),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_199),
.B(n_205),
.Y(n_246)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_162),
.Y(n_200)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_200),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_L g201 ( 
.A1(n_126),
.A2(n_74),
.B1(n_72),
.B2(n_29),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_160),
.Y(n_202)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_202),
.Y(n_284)
);

BUFx2_ASAP7_75t_SL g203 ( 
.A(n_118),
.Y(n_203)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_203),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_163),
.B(n_96),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_114),
.B(n_29),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_160),
.Y(n_206)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_206),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_161),
.B(n_1),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_207),
.B(n_221),
.Y(n_276)
);

NAND3xp33_ASAP7_75t_L g261 ( 
.A(n_208),
.B(n_219),
.C(n_220),
.Y(n_261)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_144),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_118),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_164),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_211),
.B(n_218),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_111),
.Y(n_212)
);

INVx8_ASAP7_75t_L g263 ( 
.A(n_212),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_132),
.B(n_75),
.Y(n_213)
);

AND2x2_ASAP7_75t_SL g239 ( 
.A(n_213),
.B(n_139),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_132),
.B(n_140),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_214),
.B(n_217),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_128),
.B(n_75),
.C(n_104),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_215),
.B(n_7),
.C(n_8),
.Y(n_272)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_107),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_107),
.B(n_140),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_122),
.B(n_2),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_115),
.B(n_52),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_109),
.B(n_2),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_159),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_109),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_223),
.B(n_227),
.Y(n_266)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_123),
.Y(n_224)
);

INVx8_ASAP7_75t_L g267 ( 
.A(n_224),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_225),
.A2(n_136),
.B1(n_125),
.B2(n_168),
.Y(n_251)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_165),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_226),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_122),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_120),
.B(n_3),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_228),
.B(n_15),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_120),
.B(n_3),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_229),
.B(n_6),
.Y(n_270)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_158),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_230),
.B(n_7),
.Y(n_277)
);

OAI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_176),
.A2(n_151),
.B1(n_123),
.B2(n_155),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_231),
.A2(n_235),
.B1(n_250),
.B2(n_282),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_233),
.B(n_272),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_176),
.A2(n_158),
.B1(n_138),
.B2(n_155),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_239),
.Y(n_333)
);

A2O1A1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_172),
.A2(n_115),
.B(n_147),
.C(n_168),
.Y(n_241)
);

A2O1A1Ixp33_ASAP7_75t_L g332 ( 
.A1(n_241),
.A2(n_13),
.B(n_261),
.C(n_254),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_170),
.B(n_147),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_243),
.B(n_258),
.C(n_273),
.Y(n_302)
);

NOR2x1p5_ASAP7_75t_L g245 ( 
.A(n_195),
.B(n_147),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_245),
.B(n_186),
.Y(n_325)
);

OAI22xp33_ASAP7_75t_L g250 ( 
.A1(n_207),
.A2(n_139),
.B1(n_136),
.B2(n_125),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_251),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_254),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_199),
.B(n_112),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_180),
.A2(n_112),
.B1(n_5),
.B2(n_6),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_259),
.A2(n_260),
.B1(n_285),
.B2(n_202),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_201),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_204),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_274),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_270),
.B(n_210),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_188),
.B(n_7),
.C(n_8),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_204),
.Y(n_274)
);

INVxp33_ASAP7_75t_L g308 ( 
.A(n_277),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_281),
.B(n_169),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_189),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_246),
.B(n_219),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_286),
.B(n_313),
.C(n_326),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_233),
.A2(n_178),
.B1(n_228),
.B2(n_221),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_287),
.A2(n_300),
.B1(n_241),
.B2(n_242),
.Y(n_345)
);

INVx5_ASAP7_75t_L g288 ( 
.A(n_263),
.Y(n_288)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_288),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_245),
.A2(n_220),
.B(n_205),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_289),
.B(n_314),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_291),
.B(n_307),
.Y(n_350)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_247),
.Y(n_292)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_292),
.Y(n_351)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_247),
.Y(n_293)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_293),
.Y(n_355)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_252),
.Y(n_294)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_294),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_296),
.A2(n_269),
.B1(n_248),
.B2(n_283),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_267),
.Y(n_297)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_297),
.Y(n_341)
);

NOR3xp33_ASAP7_75t_SL g298 ( 
.A(n_246),
.B(n_196),
.C(n_190),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_298),
.B(n_322),
.Y(n_352)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_252),
.Y(n_299)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_299),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_276),
.A2(n_171),
.B1(n_230),
.B2(n_223),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_279),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_301),
.B(n_303),
.Y(n_338)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_279),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_280),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_305),
.B(n_306),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_237),
.Y(n_307)
);

OAI32xp33_ASAP7_75t_L g310 ( 
.A1(n_232),
.A2(n_215),
.A3(n_194),
.B1(n_192),
.B2(n_182),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_310),
.B(n_312),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_237),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_311),
.B(n_317),
.Y(n_379)
);

INVx2_ASAP7_75t_SL g312 ( 
.A(n_284),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_258),
.B(n_232),
.C(n_243),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_245),
.A2(n_182),
.B(n_192),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_235),
.A2(n_209),
.B1(n_197),
.B2(n_198),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_315),
.A2(n_316),
.B1(n_329),
.B2(n_285),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_276),
.A2(n_200),
.B1(n_184),
.B2(n_175),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_266),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_240),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_318),
.B(n_319),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_236),
.B(n_216),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_264),
.A2(n_179),
.B(n_213),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_320),
.A2(n_325),
.B(n_332),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_281),
.B(n_191),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_321),
.B(n_323),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_262),
.B(n_226),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_236),
.B(n_213),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_240),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_324),
.B(n_330),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_242),
.B(n_212),
.C(n_224),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_255),
.B(n_11),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_328),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_259),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_273),
.B(n_13),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_277),
.B(n_13),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_331),
.B(n_334),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_238),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_242),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_335),
.B(n_239),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_336),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_309),
.A2(n_260),
.B1(n_239),
.B2(n_250),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_343),
.A2(n_349),
.B1(n_371),
.B2(n_377),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_288),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_344),
.B(n_346),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_345),
.B(n_364),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_290),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_305),
.Y(n_347)
);

CKINVDCx14_ASAP7_75t_R g389 ( 
.A(n_347),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_313),
.B(n_244),
.C(n_249),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_348),
.B(n_368),
.C(n_369),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_309),
.A2(n_327),
.B1(n_304),
.B2(n_325),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_295),
.A2(n_317),
.B1(n_335),
.B2(n_297),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_354),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_306),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_360),
.B(n_366),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_295),
.A2(n_267),
.B1(n_272),
.B2(n_283),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_363),
.A2(n_331),
.B1(n_294),
.B2(n_299),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_312),
.Y(n_366)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_367),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_302),
.B(n_275),
.C(n_248),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_302),
.B(n_278),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_312),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_370),
.B(n_311),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_327),
.A2(n_234),
.B1(n_263),
.B2(n_257),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_286),
.B(n_265),
.C(n_256),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_372),
.B(n_375),
.C(n_376),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_319),
.B(n_256),
.Y(n_373)
);

XNOR2x2_ASAP7_75t_L g405 ( 
.A(n_373),
.B(n_374),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_291),
.B(n_271),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_323),
.B(n_271),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_310),
.B(n_278),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_327),
.A2(n_257),
.B1(n_265),
.B2(n_253),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_346),
.B(n_334),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_380),
.B(n_391),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_369),
.B(n_289),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_387),
.B(n_388),
.C(n_393),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_339),
.B(n_320),
.C(n_333),
.Y(n_388)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_338),
.Y(n_390)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_390),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_338),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_338),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_392),
.B(n_400),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_339),
.B(n_333),
.C(n_314),
.Y(n_393)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_394),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_349),
.A2(n_287),
.B1(n_296),
.B2(n_325),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_395),
.A2(n_396),
.B1(n_404),
.B2(n_409),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_337),
.A2(n_332),
.B1(n_300),
.B2(n_308),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_378),
.B(n_321),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_397),
.B(n_407),
.C(n_408),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_337),
.A2(n_307),
.B(n_326),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_399),
.A2(n_403),
.B(n_355),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_360),
.B(n_330),
.Y(n_400)
);

INVx5_ASAP7_75t_L g401 ( 
.A(n_341),
.Y(n_401)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_401),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_379),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_402),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_359),
.A2(n_292),
.B(n_293),
.Y(n_403)
);

INVx4_ASAP7_75t_L g406 ( 
.A(n_344),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_406),
.B(n_347),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_368),
.B(n_301),
.C(n_303),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_348),
.B(n_316),
.C(n_318),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_343),
.A2(n_315),
.B1(n_329),
.B2(n_324),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_351),
.Y(n_410)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_410),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_362),
.Y(n_411)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_411),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_378),
.B(n_298),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_412),
.B(n_387),
.Y(n_420)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_351),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_415),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_352),
.B(n_253),
.Y(n_416)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_416),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_418),
.B(n_389),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_420),
.B(n_422),
.Y(n_465)
);

FAx1_ASAP7_75t_SL g421 ( 
.A(n_412),
.B(n_359),
.CI(n_353),
.CON(n_421),
.SN(n_421)
);

FAx1_ASAP7_75t_SL g458 ( 
.A(n_421),
.B(n_385),
.CI(n_429),
.CON(n_458),
.SN(n_458)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_384),
.B(n_376),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_398),
.A2(n_358),
.B1(n_357),
.B2(n_345),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_424),
.A2(n_431),
.B1(n_433),
.B2(n_436),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_384),
.B(n_353),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_427),
.B(n_430),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_SL g430 ( 
.A(n_397),
.B(n_375),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_386),
.A2(n_342),
.B1(n_357),
.B2(n_350),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_396),
.A2(n_371),
.B1(n_342),
.B2(n_377),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_413),
.A2(n_367),
.B1(n_370),
.B2(n_366),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_434),
.A2(n_437),
.B1(n_444),
.B2(n_417),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_386),
.A2(n_373),
.B1(n_374),
.B2(n_372),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_395),
.A2(n_356),
.B1(n_365),
.B2(n_361),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g439 ( 
.A(n_393),
.B(n_356),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_439),
.B(n_446),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_442),
.A2(n_403),
.B(n_382),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_388),
.B(n_355),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_443),
.B(n_439),
.C(n_447),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_399),
.A2(n_365),
.B1(n_361),
.B2(n_340),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_382),
.Y(n_445)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_445),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_407),
.B(n_340),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_385),
.B(n_381),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_447),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_432),
.A2(n_437),
.B1(n_442),
.B2(n_431),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_449),
.A2(n_469),
.B1(n_470),
.B2(n_454),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_451),
.A2(n_456),
.B(n_469),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_441),
.B(n_414),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_452),
.B(n_467),
.Y(n_498)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_455),
.Y(n_485)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_418),
.Y(n_456)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_456),
.Y(n_486)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_426),
.Y(n_457)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_457),
.Y(n_488)
);

MAJx2_ASAP7_75t_L g479 ( 
.A(n_458),
.B(n_423),
.C(n_429),
.Y(n_479)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_428),
.Y(n_459)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_459),
.Y(n_491)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_419),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_460),
.B(n_467),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_461),
.B(n_423),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_438),
.B(n_427),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_462),
.B(n_450),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_422),
.B(n_408),
.C(n_394),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_463),
.B(n_464),
.C(n_430),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_443),
.B(n_394),
.C(n_382),
.Y(n_464)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_435),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_466),
.B(n_472),
.Y(n_489)
);

INVxp33_ASAP7_75t_L g467 ( 
.A(n_440),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_425),
.A2(n_413),
.B1(n_383),
.B2(n_404),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_436),
.A2(n_383),
.B1(n_409),
.B2(n_406),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_448),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_471),
.Y(n_483)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_417),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_434),
.A2(n_405),
.B(n_415),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_473),
.A2(n_421),
.B(n_401),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_474),
.A2(n_444),
.B1(n_446),
.B2(n_405),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_476),
.A2(n_449),
.B1(n_399),
.B2(n_436),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_473),
.A2(n_421),
.B(n_420),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_SL g513 ( 
.A1(n_477),
.A2(n_482),
.B(n_495),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_478),
.B(n_480),
.Y(n_502)
);

FAx1_ASAP7_75t_SL g501 ( 
.A(n_479),
.B(n_458),
.CI(n_475),
.CON(n_501),
.SN(n_501)
);

BUFx24_ASAP7_75t_SL g481 ( 
.A(n_458),
.Y(n_481)
);

BUFx24_ASAP7_75t_SL g500 ( 
.A(n_481),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_463),
.B(n_465),
.C(n_464),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_484),
.B(n_487),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_465),
.B(n_475),
.C(n_453),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_490),
.A2(n_460),
.B(n_457),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_492),
.B(n_493),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_453),
.B(n_461),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_449),
.A2(n_470),
.B1(n_468),
.B2(n_451),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_494),
.B(n_490),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_496),
.B(n_498),
.Y(n_503)
);

BUFx12_ASAP7_75t_L g497 ( 
.A(n_455),
.Y(n_497)
);

INVx11_ASAP7_75t_L g515 ( 
.A(n_497),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_501),
.B(n_506),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_504),
.B(n_513),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_505),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_484),
.B(n_480),
.C(n_478),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_489),
.B(n_485),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_507),
.B(n_511),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_482),
.A2(n_476),
.B(n_477),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_508),
.B(n_514),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_493),
.B(n_491),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_509),
.B(n_499),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_487),
.B(n_479),
.C(n_494),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_486),
.B(n_495),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_512),
.B(n_516),
.Y(n_522)
);

FAx1_ASAP7_75t_SL g514 ( 
.A(n_497),
.B(n_488),
.CI(n_483),
.CON(n_514),
.SN(n_514)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_512),
.B(n_483),
.Y(n_519)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_519),
.Y(n_534)
);

FAx1_ASAP7_75t_L g520 ( 
.A(n_513),
.B(n_497),
.CI(n_508),
.CON(n_520),
.SN(n_520)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_520),
.B(n_514),
.Y(n_537)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_504),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_523),
.B(n_524),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_506),
.B(n_502),
.C(n_510),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_525),
.B(n_527),
.C(n_522),
.Y(n_538)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_503),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g535 ( 
.A(n_526),
.B(n_529),
.Y(n_535)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_516),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_510),
.B(n_502),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_530),
.A2(n_500),
.B(n_515),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_521),
.B(n_511),
.Y(n_531)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_531),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_532),
.B(n_533),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_SL g533 ( 
.A1(n_517),
.A2(n_501),
.B(n_515),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_528),
.A2(n_501),
.B(n_514),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_536),
.B(n_537),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_SL g544 ( 
.A(n_538),
.B(n_540),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_525),
.B(n_527),
.C(n_518),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_535),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_543),
.B(n_545),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_531),
.B(n_518),
.Y(n_545)
);

CKINVDCx16_ASAP7_75t_R g547 ( 
.A(n_546),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_547),
.B(n_544),
.Y(n_552)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_541),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g551 ( 
.A(n_548),
.B(n_550),
.Y(n_551)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_542),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_552),
.B(n_549),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_553),
.A2(n_554),
.B1(n_546),
.B2(n_537),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_551),
.B(n_549),
.C(n_539),
.Y(n_554)
);

CKINVDCx14_ASAP7_75t_R g556 ( 
.A(n_555),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_556),
.B(n_534),
.Y(n_557)
);


endmodule