module fake_aes_2318_n_36 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_36);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_36;
wire n_20;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_30;
wire n_13;
wire n_33;
wire n_26;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
INVx1_ASAP7_75t_L g11 ( .A(n_6), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_9), .Y(n_12) );
OA21x2_ASAP7_75t_L g13 ( .A1(n_3), .A2(n_0), .B(n_8), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_5), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_0), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_2), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_7), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_16), .Y(n_18) );
AND2x4_ASAP7_75t_L g19 ( .A(n_15), .B(n_1), .Y(n_19) );
INVx1_ASAP7_75t_SL g20 ( .A(n_12), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_11), .Y(n_21) );
INVx1_ASAP7_75t_SL g22 ( .A(n_12), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_20), .B(n_13), .Y(n_23) );
INVx4_ASAP7_75t_L g24 ( .A(n_19), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_18), .Y(n_25) );
O2A1O1Ixp5_ASAP7_75t_L g26 ( .A1(n_21), .A2(n_14), .B(n_17), .C(n_13), .Y(n_26) );
AND2x4_ASAP7_75t_L g27 ( .A(n_24), .B(n_19), .Y(n_27) );
AND2x2_ASAP7_75t_L g28 ( .A(n_25), .B(n_20), .Y(n_28) );
OR2x2_ASAP7_75t_L g29 ( .A(n_24), .B(n_22), .Y(n_29) );
AND2x2_ASAP7_75t_L g30 ( .A(n_28), .B(n_23), .Y(n_30) );
OAI21xp5_ASAP7_75t_SL g31 ( .A1(n_30), .A2(n_29), .B(n_27), .Y(n_31) );
NAND2xp5_ASAP7_75t_L g32 ( .A(n_31), .B(n_30), .Y(n_32) );
AO22x1_ASAP7_75t_SL g33 ( .A1(n_31), .A2(n_1), .B1(n_2), .B2(n_4), .Y(n_33) );
CKINVDCx16_ASAP7_75t_R g34 ( .A(n_32), .Y(n_34) );
HB1xp67_ASAP7_75t_L g35 ( .A(n_34), .Y(n_35) );
AOI22xp33_ASAP7_75t_L g36 ( .A1(n_35), .A2(n_33), .B1(n_26), .B2(n_10), .Y(n_36) );
endmodule