module fake_jpeg_31643_n_26 (n_3, n_2, n_1, n_0, n_4, n_5, n_26);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_26;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx8_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_4),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_1),
.B(n_4),
.Y(n_9)
);

INVx6_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

INVx13_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_13),
.Y(n_20)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_14),
.A2(n_15),
.B1(n_16),
.B2(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_8),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_15),
.B(n_6),
.C(n_9),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_17),
.A2(n_18),
.B(n_19),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_SL g18 ( 
.A(n_12),
.B(n_7),
.C(n_11),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_17),
.B(n_7),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_23),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_20),
.A2(n_13),
.B1(n_14),
.B2(n_11),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_5),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_25),
.Y(n_26)
);


endmodule