module fake_netlist_5_2496_n_7499 (n_924, n_1263, n_977, n_1378, n_611, n_1126, n_1423, n_1729, n_1166, n_469, n_1508, n_82, n_785, n_549, n_532, n_1161, n_1677, n_1150, n_226, n_1488, n_667, n_790, n_1055, n_1501, n_111, n_880, n_544, n_1007, n_155, n_552, n_1528, n_1370, n_1292, n_1198, n_1360, n_1099, n_956, n_564, n_423, n_21, n_105, n_1021, n_4, n_551, n_1323, n_1466, n_688, n_1695, n_1353, n_800, n_1347, n_1535, n_1666, n_671, n_819, n_1451, n_1022, n_915, n_1545, n_864, n_173, n_859, n_951, n_1264, n_447, n_247, n_1494, n_292, n_625, n_854, n_1462, n_1580, n_674, n_417, n_516, n_933, n_1152, n_497, n_1607, n_1563, n_606, n_275, n_26, n_877, n_2, n_1696, n_755, n_1118, n_6, n_1686, n_947, n_1285, n_373, n_307, n_1359, n_530, n_87, n_150, n_1107, n_1728, n_556, n_1230, n_668, n_375, n_301, n_929, n_1124, n_902, n_1576, n_191, n_1104, n_1294, n_659, n_51, n_1705, n_1257, n_171, n_1182, n_579, n_1698, n_1261, n_938, n_1098, n_320, n_1154, n_1242, n_1135, n_24, n_406, n_519, n_1016, n_1243, n_546, n_101, n_1280, n_281, n_240, n_291, n_231, n_257, n_731, n_371, n_1483, n_1314, n_1512, n_709, n_1490, n_317, n_1236, n_1633, n_569, n_227, n_920, n_1289, n_1517, n_94, n_335, n_1669, n_370, n_976, n_343, n_1449, n_308, n_1566, n_297, n_156, n_1078, n_1670, n_775, n_219, n_157, n_600, n_1484, n_1374, n_1328, n_223, n_264, n_1598, n_1723, n_955, n_163, n_339, n_1146, n_882, n_183, n_243, n_1036, n_1097, n_347, n_59, n_550, n_696, n_897, n_215, n_350, n_196, n_798, n_646, n_1428, n_436, n_1394, n_1414, n_1216, n_290, n_580, n_1040, n_578, n_926, n_344, n_1218, n_422, n_475, n_777, n_1070, n_1547, n_1030, n_72, n_415, n_1071, n_485, n_1165, n_1267, n_1561, n_496, n_1391, n_958, n_1034, n_670, n_1513, n_1600, n_48, n_521, n_663, n_845, n_673, n_837, n_1239, n_528, n_680, n_1473, n_1587, n_395, n_164, n_553, n_901, n_813, n_1521, n_1284, n_1590, n_214, n_1672, n_675, n_888, n_1167, n_1626, n_637, n_1384, n_1556, n_184, n_446, n_1064, n_144, n_858, n_114, n_96, n_923, n_691, n_1151, n_881, n_1405, n_1706, n_468, n_213, n_129, n_342, n_464, n_363, n_1582, n_197, n_1069, n_1075, n_1450, n_1322, n_1471, n_1459, n_460, n_889, n_973, n_1700, n_477, n_571, n_1585, n_461, n_1599, n_1211, n_1197, n_1523, n_907, n_1447, n_1377, n_190, n_989, n_1039, n_34, n_228, n_283, n_1403, n_488, n_736, n_892, n_1000, n_1202, n_1278, n_1002, n_1463, n_1581, n_49, n_310, n_54, n_593, n_12, n_748, n_586, n_1058, n_1667, n_838, n_332, n_1053, n_1224, n_349, n_1248, n_230, n_1331, n_953, n_279, n_1014, n_1241, n_70, n_289, n_963, n_1052, n_954, n_627, n_1385, n_440, n_793, n_478, n_476, n_1527, n_534, n_884, n_345, n_944, n_1623, n_91, n_1565, n_182, n_143, n_647, n_237, n_407, n_1072, n_832, n_857, n_207, n_561, n_1319, n_1712, n_1387, n_1532, n_18, n_1027, n_971, n_1156, n_117, n_326, n_794, n_404, n_686, n_847, n_1393, n_596, n_1368, n_558, n_702, n_1276, n_822, n_1412, n_1709, n_728, n_266, n_1162, n_272, n_1538, n_1199, n_352, n_53, n_1038, n_520, n_1369, n_409, n_1660, n_887, n_154, n_71, n_300, n_809, n_870, n_931, n_599, n_1711, n_1662, n_1481, n_434, n_1544, n_868, n_639, n_914, n_411, n_414, n_1629, n_1293, n_965, n_935, n_121, n_1175, n_817, n_360, n_36, n_1479, n_64, n_759, n_28, n_806, n_1477, n_324, n_1635, n_1571, n_187, n_1189, n_103, n_97, n_11, n_7, n_1259, n_1690, n_706, n_746, n_1649, n_747, n_52, n_784, n_110, n_1733, n_1244, n_431, n_1194, n_615, n_851, n_843, n_523, n_913, n_1537, n_705, n_865, n_61, n_678, n_697, n_127, n_1222, n_75, n_1679, n_776, n_1415, n_367, n_452, n_525, n_1260, n_1647, n_1464, n_649, n_547, n_43, n_1444, n_1191, n_1674, n_116, n_1710, n_284, n_1128, n_139, n_1734, n_744, n_590, n_629, n_1308, n_254, n_1680, n_1233, n_23, n_1615, n_1529, n_526, n_293, n_372, n_677, n_244, n_47, n_1333, n_1121, n_314, n_368, n_433, n_604, n_8, n_949, n_100, n_1443, n_1008, n_946, n_1539, n_1001, n_1503, n_498, n_1468, n_1559, n_689, n_738, n_1624, n_640, n_1510, n_252, n_624, n_1380, n_1617, n_295, n_133, n_1010, n_1231, n_739, n_1279, n_1406, n_1195, n_610, n_936, n_568, n_1500, n_39, n_1090, n_757, n_633, n_439, n_106, n_259, n_448, n_758, n_999, n_93, n_1656, n_1158, n_1509, n_563, n_1145, n_878, n_524, n_204, n_394, n_1678, n_1049, n_1153, n_741, n_1639, n_1306, n_1068, n_122, n_331, n_10, n_906, n_1163, n_1207, n_919, n_908, n_90, n_724, n_658, n_1362, n_1586, n_456, n_959, n_535, n_152, n_940, n_1445, n_9, n_1492, n_592, n_1169, n_45, n_1596, n_1692, n_1017, n_123, n_978, n_1434, n_1054, n_1474, n_1665, n_1269, n_1095, n_1614, n_267, n_514, n_457, n_1079, n_1045, n_1208, n_603, n_1431, n_484, n_1593, n_1033, n_442, n_131, n_636, n_660, n_1640, n_1732, n_1009, n_1148, n_109, n_742, n_750, n_995, n_454, n_1609, n_374, n_185, n_396, n_1383, n_1073, n_255, n_662, n_459, n_218, n_962, n_1215, n_1171, n_1578, n_723, n_1065, n_1592, n_1336, n_1721, n_1574, n_473, n_1309, n_1426, n_1043, n_355, n_486, n_1548, n_614, n_337, n_1421, n_88, n_1286, n_1177, n_1355, n_168, n_974, n_727, n_1159, n_957, n_773, n_208, n_142, n_743, n_299, n_303, n_296, n_613, n_1119, n_1240, n_65, n_829, n_1612, n_1416, n_1724, n_361, n_700, n_1237, n_573, n_69, n_1420, n_1132, n_388, n_1366, n_1300, n_1127, n_761, n_1568, n_1006, n_329, n_274, n_1270, n_1664, n_1486, n_582, n_1332, n_1390, n_73, n_19, n_309, n_30, n_512, n_1591, n_84, n_130, n_322, n_1682, n_1249, n_652, n_1111, n_1365, n_25, n_1349, n_1093, n_288, n_1031, n_263, n_609, n_1041, n_1265, n_44, n_224, n_1562, n_383, n_834, n_112, n_765, n_893, n_1015, n_1140, n_891, n_1651, n_239, n_630, n_55, n_504, n_511, n_874, n_358, n_1101, n_77, n_102, n_1106, n_1456, n_1304, n_1324, n_987, n_261, n_174, n_1455, n_767, n_993, n_1407, n_1551, n_545, n_441, n_860, n_450, n_429, n_948, n_1217, n_628, n_365, n_729, n_1131, n_1084, n_970, n_911, n_1430, n_83, n_513, n_1094, n_1354, n_560, n_1534, n_340, n_1351, n_1044, n_1205, n_346, n_1209, n_1552, n_495, n_602, n_574, n_1435, n_879, n_16, n_58, n_623, n_405, n_824, n_359, n_1645, n_490, n_1327, n_996, n_921, n_1684, n_233, n_1717, n_572, n_366, n_815, n_128, n_120, n_327, n_135, n_1381, n_1611, n_1037, n_1080, n_1274, n_1316, n_1708, n_426, n_1438, n_1082, n_589, n_716, n_1630, n_562, n_1436, n_62, n_1691, n_952, n_1229, n_391, n_701, n_1437, n_1023, n_645, n_539, n_803, n_1092, n_238, n_531, n_890, n_764, n_1056, n_1424, n_162, n_960, n_222, n_1290, n_1123, n_1467, n_1047, n_634, n_199, n_32, n_1252, n_348, n_1382, n_1029, n_925, n_1206, n_424, n_1311, n_1519, n_256, n_950, n_1553, n_380, n_419, n_1346, n_444, n_1299, n_1060, n_1141, n_316, n_389, n_418, n_248, n_136, n_86, n_146, n_912, n_315, n_968, n_451, n_619, n_408, n_1386, n_1699, n_376, n_967, n_1442, n_74, n_1139, n_515, n_57, n_351, n_885, n_397, n_1432, n_1357, n_483, n_683, n_1632, n_1057, n_1051, n_1085, n_1066, n_721, n_1157, n_841, n_1050, n_22, n_802, n_46, n_1608, n_983, n_38, n_280, n_1305, n_873, n_378, n_1112, n_762, n_1283, n_1644, n_17, n_690, n_33, n_583, n_302, n_1343, n_1203, n_1631, n_821, n_321, n_1179, n_621, n_753, n_455, n_1048, n_1719, n_1288, n_212, n_385, n_507, n_1560, n_1605, n_330, n_1228, n_972, n_692, n_820, n_1200, n_1301, n_1363, n_1668, n_1185, n_991, n_828, n_779, n_576, n_1143, n_1579, n_1329, n_1312, n_1439, n_804, n_537, n_1688, n_945, n_492, n_153, n_1504, n_943, n_341, n_250, n_992, n_543, n_260, n_842, n_650, n_984, n_694, n_286, n_1643, n_883, n_470, n_325, n_449, n_1594, n_132, n_1214, n_1342, n_1400, n_900, n_856, n_918, n_942, n_189, n_1147, n_1557, n_1610, n_13, n_1077, n_1422, n_540, n_618, n_896, n_323, n_195, n_356, n_894, n_1636, n_1730, n_831, n_964, n_1373, n_1350, n_1511, n_1470, n_1096, n_234, n_1575, n_1697, n_1735, n_833, n_5, n_1646, n_225, n_1307, n_988, n_814, n_192, n_1549, n_1201, n_1114, n_655, n_1616, n_1446, n_669, n_472, n_1458, n_1176, n_1472, n_387, n_1149, n_398, n_1671, n_635, n_763, n_1020, n_1062, n_211, n_1219, n_3, n_1204, n_178, n_1035, n_287, n_555, n_783, n_1188, n_1722, n_661, n_41, n_849, n_15, n_336, n_584, n_681, n_1638, n_50, n_430, n_510, n_216, n_311, n_830, n_1296, n_1413, n_801, n_241, n_875, n_357, n_1110, n_1655, n_445, n_749, n_1134, n_1358, n_717, n_165, n_939, n_482, n_1088, n_588, n_1173, n_789, n_1232, n_1603, n_734, n_638, n_866, n_107, n_969, n_1401, n_1019, n_1105, n_249, n_304, n_1338, n_577, n_1522, n_1687, n_1637, n_1419, n_338, n_149, n_1653, n_693, n_1506, n_14, n_836, n_990, n_1389, n_975, n_1256, n_1702, n_567, n_1465, n_778, n_1122, n_151, n_306, n_458, n_770, n_1375, n_1102, n_711, n_1499, n_85, n_1187, n_1441, n_1392, n_1597, n_1164, n_1659, n_489, n_1174, n_1371, n_617, n_1303, n_1572, n_876, n_1516, n_1190, n_1736, n_1685, n_118, n_601, n_917, n_1714, n_966, n_253, n_1116, n_1661, n_1212, n_1541, n_172, n_206, n_217, n_726, n_982, n_1573, n_1453, n_1731, n_818, n_861, n_1713, n_1183, n_1658, n_899, n_1253, n_210, n_1737, n_774, n_1628, n_1335, n_1514, n_1059, n_1345, n_176, n_1133, n_557, n_1410, n_1005, n_607, n_1003, n_679, n_710, n_527, n_1168, n_707, n_937, n_1427, n_393, n_108, n_487, n_1584, n_665, n_1726, n_66, n_1440, n_177, n_421, n_1356, n_910, n_1657, n_768, n_1475, n_1302, n_1725, n_205, n_1136, n_1313, n_1491, n_754, n_1496, n_179, n_1125, n_125, n_410, n_708, n_529, n_735, n_232, n_1109, n_126, n_895, n_1310, n_202, n_427, n_1399, n_1543, n_791, n_732, n_1533, n_193, n_808, n_797, n_1025, n_500, n_1067, n_1720, n_148, n_435, n_159, n_766, n_1457, n_541, n_538, n_1117, n_799, n_687, n_715, n_1480, n_1482, n_1213, n_1266, n_536, n_872, n_594, n_200, n_1291, n_1297, n_1155, n_1418, n_89, n_1524, n_1689, n_1485, n_115, n_1011, n_1184, n_985, n_869, n_810, n_416, n_827, n_401, n_1703, n_1352, n_626, n_1650, n_1144, n_1137, n_1570, n_1170, n_305, n_137, n_676, n_294, n_318, n_653, n_642, n_1602, n_194, n_855, n_1178, n_1461, n_850, n_684, n_124, n_268, n_664, n_503, n_235, n_1372, n_605, n_1273, n_353, n_620, n_643, n_916, n_1081, n_493, n_1235, n_703, n_698, n_980, n_1115, n_1282, n_1318, n_780, n_998, n_1454, n_467, n_1227, n_1531, n_840, n_1334, n_501, n_823, n_245, n_725, n_1388, n_1417, n_1295, n_672, n_581, n_382, n_554, n_1625, n_898, n_1013, n_1452, n_718, n_265, n_1120, n_719, n_443, n_198, n_714, n_1683, n_909, n_1497, n_1530, n_997, n_932, n_612, n_1409, n_788, n_1326, n_119, n_1268, n_559, n_825, n_508, n_506, n_1320, n_1663, n_737, n_1718, n_986, n_509, n_1317, n_147, n_1518, n_1715, n_1281, n_67, n_1192, n_1024, n_1063, n_209, n_1564, n_1613, n_733, n_1489, n_1376, n_941, n_981, n_1569, n_68, n_867, n_186, n_134, n_587, n_63, n_792, n_756, n_1429, n_399, n_1238, n_548, n_812, n_298, n_518, n_505, n_282, n_752, n_905, n_1476, n_1108, n_782, n_1100, n_1395, n_862, n_1425, n_760, n_1620, n_381, n_220, n_390, n_1330, n_31, n_481, n_1675, n_1727, n_1554, n_769, n_42, n_1046, n_271, n_934, n_1618, n_826, n_886, n_1221, n_654, n_1172, n_167, n_379, n_428, n_1341, n_570, n_1641, n_1361, n_1707, n_853, n_377, n_751, n_786, n_1083, n_1142, n_1129, n_392, n_158, n_704, n_787, n_138, n_961, n_771, n_276, n_95, n_1716, n_1225, n_1520, n_169, n_522, n_1287, n_1262, n_400, n_930, n_181, n_1411, n_221, n_622, n_1577, n_1087, n_386, n_994, n_1701, n_848, n_1550, n_1498, n_1223, n_1272, n_104, n_682, n_1567, n_56, n_141, n_1247, n_922, n_816, n_1648, n_591, n_145, n_1536, n_1344, n_313, n_631, n_479, n_1246, n_1339, n_1478, n_432, n_839, n_1210, n_1364, n_328, n_140, n_1250, n_369, n_871, n_598, n_685, n_928, n_608, n_1367, n_78, n_1460, n_772, n_1555, n_499, n_1589, n_517, n_98, n_402, n_413, n_1086, n_796, n_1619, n_236, n_1502, n_1469, n_1012, n_1, n_1396, n_1348, n_903, n_1525, n_740, n_203, n_384, n_1404, n_80, n_35, n_1315, n_277, n_1061, n_92, n_333, n_1298, n_1652, n_462, n_1193, n_1676, n_1255, n_258, n_1113, n_29, n_79, n_1226, n_722, n_1277, n_188, n_844, n_201, n_471, n_852, n_1487, n_40, n_1028, n_1601, n_781, n_474, n_542, n_463, n_1546, n_595, n_502, n_466, n_420, n_1337, n_1495, n_632, n_699, n_979, n_1515, n_1627, n_1245, n_846, n_1673, n_465, n_76, n_362, n_1321, n_170, n_27, n_161, n_273, n_585, n_270, n_616, n_81, n_745, n_1654, n_1103, n_648, n_1379, n_312, n_1076, n_1091, n_1408, n_494, n_641, n_730, n_1325, n_1595, n_354, n_575, n_480, n_425, n_795, n_695, n_180, n_656, n_1606, n_1220, n_37, n_1694, n_1540, n_229, n_437, n_1642, n_60, n_403, n_453, n_1130, n_720, n_0, n_1526, n_863, n_805, n_1604, n_1275, n_113, n_712, n_246, n_1583, n_1042, n_1402, n_269, n_285, n_412, n_1493, n_657, n_644, n_1160, n_1397, n_491, n_1258, n_1074, n_1621, n_251, n_160, n_566, n_565, n_1448, n_1507, n_1398, n_597, n_1181, n_1505, n_1634, n_1196, n_651, n_1340, n_334, n_811, n_1558, n_807, n_835, n_175, n_666, n_262, n_1433, n_1704, n_99, n_1254, n_1026, n_1234, n_319, n_364, n_1138, n_927, n_20, n_1089, n_1004, n_1186, n_1032, n_242, n_1681, n_1018, n_1693, n_438, n_713, n_904, n_1588, n_1622, n_166, n_1180, n_1271, n_533, n_1542, n_1251, n_278, n_7499);

input n_924;
input n_1263;
input n_977;
input n_1378;
input n_611;
input n_1126;
input n_1423;
input n_1729;
input n_1166;
input n_469;
input n_1508;
input n_82;
input n_785;
input n_549;
input n_532;
input n_1161;
input n_1677;
input n_1150;
input n_226;
input n_1488;
input n_667;
input n_790;
input n_1055;
input n_1501;
input n_111;
input n_880;
input n_544;
input n_1007;
input n_155;
input n_552;
input n_1528;
input n_1370;
input n_1292;
input n_1198;
input n_1360;
input n_1099;
input n_956;
input n_564;
input n_423;
input n_21;
input n_105;
input n_1021;
input n_4;
input n_551;
input n_1323;
input n_1466;
input n_688;
input n_1695;
input n_1353;
input n_800;
input n_1347;
input n_1535;
input n_1666;
input n_671;
input n_819;
input n_1451;
input n_1022;
input n_915;
input n_1545;
input n_864;
input n_173;
input n_859;
input n_951;
input n_1264;
input n_447;
input n_247;
input n_1494;
input n_292;
input n_625;
input n_854;
input n_1462;
input n_1580;
input n_674;
input n_417;
input n_516;
input n_933;
input n_1152;
input n_497;
input n_1607;
input n_1563;
input n_606;
input n_275;
input n_26;
input n_877;
input n_2;
input n_1696;
input n_755;
input n_1118;
input n_6;
input n_1686;
input n_947;
input n_1285;
input n_373;
input n_307;
input n_1359;
input n_530;
input n_87;
input n_150;
input n_1107;
input n_1728;
input n_556;
input n_1230;
input n_668;
input n_375;
input n_301;
input n_929;
input n_1124;
input n_902;
input n_1576;
input n_191;
input n_1104;
input n_1294;
input n_659;
input n_51;
input n_1705;
input n_1257;
input n_171;
input n_1182;
input n_579;
input n_1698;
input n_1261;
input n_938;
input n_1098;
input n_320;
input n_1154;
input n_1242;
input n_1135;
input n_24;
input n_406;
input n_519;
input n_1016;
input n_1243;
input n_546;
input n_101;
input n_1280;
input n_281;
input n_240;
input n_291;
input n_231;
input n_257;
input n_731;
input n_371;
input n_1483;
input n_1314;
input n_1512;
input n_709;
input n_1490;
input n_317;
input n_1236;
input n_1633;
input n_569;
input n_227;
input n_920;
input n_1289;
input n_1517;
input n_94;
input n_335;
input n_1669;
input n_370;
input n_976;
input n_343;
input n_1449;
input n_308;
input n_1566;
input n_297;
input n_156;
input n_1078;
input n_1670;
input n_775;
input n_219;
input n_157;
input n_600;
input n_1484;
input n_1374;
input n_1328;
input n_223;
input n_264;
input n_1598;
input n_1723;
input n_955;
input n_163;
input n_339;
input n_1146;
input n_882;
input n_183;
input n_243;
input n_1036;
input n_1097;
input n_347;
input n_59;
input n_550;
input n_696;
input n_897;
input n_215;
input n_350;
input n_196;
input n_798;
input n_646;
input n_1428;
input n_436;
input n_1394;
input n_1414;
input n_1216;
input n_290;
input n_580;
input n_1040;
input n_578;
input n_926;
input n_344;
input n_1218;
input n_422;
input n_475;
input n_777;
input n_1070;
input n_1547;
input n_1030;
input n_72;
input n_415;
input n_1071;
input n_485;
input n_1165;
input n_1267;
input n_1561;
input n_496;
input n_1391;
input n_958;
input n_1034;
input n_670;
input n_1513;
input n_1600;
input n_48;
input n_521;
input n_663;
input n_845;
input n_673;
input n_837;
input n_1239;
input n_528;
input n_680;
input n_1473;
input n_1587;
input n_395;
input n_164;
input n_553;
input n_901;
input n_813;
input n_1521;
input n_1284;
input n_1590;
input n_214;
input n_1672;
input n_675;
input n_888;
input n_1167;
input n_1626;
input n_637;
input n_1384;
input n_1556;
input n_184;
input n_446;
input n_1064;
input n_144;
input n_858;
input n_114;
input n_96;
input n_923;
input n_691;
input n_1151;
input n_881;
input n_1405;
input n_1706;
input n_468;
input n_213;
input n_129;
input n_342;
input n_464;
input n_363;
input n_1582;
input n_197;
input n_1069;
input n_1075;
input n_1450;
input n_1322;
input n_1471;
input n_1459;
input n_460;
input n_889;
input n_973;
input n_1700;
input n_477;
input n_571;
input n_1585;
input n_461;
input n_1599;
input n_1211;
input n_1197;
input n_1523;
input n_907;
input n_1447;
input n_1377;
input n_190;
input n_989;
input n_1039;
input n_34;
input n_228;
input n_283;
input n_1403;
input n_488;
input n_736;
input n_892;
input n_1000;
input n_1202;
input n_1278;
input n_1002;
input n_1463;
input n_1581;
input n_49;
input n_310;
input n_54;
input n_593;
input n_12;
input n_748;
input n_586;
input n_1058;
input n_1667;
input n_838;
input n_332;
input n_1053;
input n_1224;
input n_349;
input n_1248;
input n_230;
input n_1331;
input n_953;
input n_279;
input n_1014;
input n_1241;
input n_70;
input n_289;
input n_963;
input n_1052;
input n_954;
input n_627;
input n_1385;
input n_440;
input n_793;
input n_478;
input n_476;
input n_1527;
input n_534;
input n_884;
input n_345;
input n_944;
input n_1623;
input n_91;
input n_1565;
input n_182;
input n_143;
input n_647;
input n_237;
input n_407;
input n_1072;
input n_832;
input n_857;
input n_207;
input n_561;
input n_1319;
input n_1712;
input n_1387;
input n_1532;
input n_18;
input n_1027;
input n_971;
input n_1156;
input n_117;
input n_326;
input n_794;
input n_404;
input n_686;
input n_847;
input n_1393;
input n_596;
input n_1368;
input n_558;
input n_702;
input n_1276;
input n_822;
input n_1412;
input n_1709;
input n_728;
input n_266;
input n_1162;
input n_272;
input n_1538;
input n_1199;
input n_352;
input n_53;
input n_1038;
input n_520;
input n_1369;
input n_409;
input n_1660;
input n_887;
input n_154;
input n_71;
input n_300;
input n_809;
input n_870;
input n_931;
input n_599;
input n_1711;
input n_1662;
input n_1481;
input n_434;
input n_1544;
input n_868;
input n_639;
input n_914;
input n_411;
input n_414;
input n_1629;
input n_1293;
input n_965;
input n_935;
input n_121;
input n_1175;
input n_817;
input n_360;
input n_36;
input n_1479;
input n_64;
input n_759;
input n_28;
input n_806;
input n_1477;
input n_324;
input n_1635;
input n_1571;
input n_187;
input n_1189;
input n_103;
input n_97;
input n_11;
input n_7;
input n_1259;
input n_1690;
input n_706;
input n_746;
input n_1649;
input n_747;
input n_52;
input n_784;
input n_110;
input n_1733;
input n_1244;
input n_431;
input n_1194;
input n_615;
input n_851;
input n_843;
input n_523;
input n_913;
input n_1537;
input n_705;
input n_865;
input n_61;
input n_678;
input n_697;
input n_127;
input n_1222;
input n_75;
input n_1679;
input n_776;
input n_1415;
input n_367;
input n_452;
input n_525;
input n_1260;
input n_1647;
input n_1464;
input n_649;
input n_547;
input n_43;
input n_1444;
input n_1191;
input n_1674;
input n_116;
input n_1710;
input n_284;
input n_1128;
input n_139;
input n_1734;
input n_744;
input n_590;
input n_629;
input n_1308;
input n_254;
input n_1680;
input n_1233;
input n_23;
input n_1615;
input n_1529;
input n_526;
input n_293;
input n_372;
input n_677;
input n_244;
input n_47;
input n_1333;
input n_1121;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_949;
input n_100;
input n_1443;
input n_1008;
input n_946;
input n_1539;
input n_1001;
input n_1503;
input n_498;
input n_1468;
input n_1559;
input n_689;
input n_738;
input n_1624;
input n_640;
input n_1510;
input n_252;
input n_624;
input n_1380;
input n_1617;
input n_295;
input n_133;
input n_1010;
input n_1231;
input n_739;
input n_1279;
input n_1406;
input n_1195;
input n_610;
input n_936;
input n_568;
input n_1500;
input n_39;
input n_1090;
input n_757;
input n_633;
input n_439;
input n_106;
input n_259;
input n_448;
input n_758;
input n_999;
input n_93;
input n_1656;
input n_1158;
input n_1509;
input n_563;
input n_1145;
input n_878;
input n_524;
input n_204;
input n_394;
input n_1678;
input n_1049;
input n_1153;
input n_741;
input n_1639;
input n_1306;
input n_1068;
input n_122;
input n_331;
input n_10;
input n_906;
input n_1163;
input n_1207;
input n_919;
input n_908;
input n_90;
input n_724;
input n_658;
input n_1362;
input n_1586;
input n_456;
input n_959;
input n_535;
input n_152;
input n_940;
input n_1445;
input n_9;
input n_1492;
input n_592;
input n_1169;
input n_45;
input n_1596;
input n_1692;
input n_1017;
input n_123;
input n_978;
input n_1434;
input n_1054;
input n_1474;
input n_1665;
input n_1269;
input n_1095;
input n_1614;
input n_267;
input n_514;
input n_457;
input n_1079;
input n_1045;
input n_1208;
input n_603;
input n_1431;
input n_484;
input n_1593;
input n_1033;
input n_442;
input n_131;
input n_636;
input n_660;
input n_1640;
input n_1732;
input n_1009;
input n_1148;
input n_109;
input n_742;
input n_750;
input n_995;
input n_454;
input n_1609;
input n_374;
input n_185;
input n_396;
input n_1383;
input n_1073;
input n_255;
input n_662;
input n_459;
input n_218;
input n_962;
input n_1215;
input n_1171;
input n_1578;
input n_723;
input n_1065;
input n_1592;
input n_1336;
input n_1721;
input n_1574;
input n_473;
input n_1309;
input n_1426;
input n_1043;
input n_355;
input n_486;
input n_1548;
input n_614;
input n_337;
input n_1421;
input n_88;
input n_1286;
input n_1177;
input n_1355;
input n_168;
input n_974;
input n_727;
input n_1159;
input n_957;
input n_773;
input n_208;
input n_142;
input n_743;
input n_299;
input n_303;
input n_296;
input n_613;
input n_1119;
input n_1240;
input n_65;
input n_829;
input n_1612;
input n_1416;
input n_1724;
input n_361;
input n_700;
input n_1237;
input n_573;
input n_69;
input n_1420;
input n_1132;
input n_388;
input n_1366;
input n_1300;
input n_1127;
input n_761;
input n_1568;
input n_1006;
input n_329;
input n_274;
input n_1270;
input n_1664;
input n_1486;
input n_582;
input n_1332;
input n_1390;
input n_73;
input n_19;
input n_309;
input n_30;
input n_512;
input n_1591;
input n_84;
input n_130;
input n_322;
input n_1682;
input n_1249;
input n_652;
input n_1111;
input n_1365;
input n_25;
input n_1349;
input n_1093;
input n_288;
input n_1031;
input n_263;
input n_609;
input n_1041;
input n_1265;
input n_44;
input n_224;
input n_1562;
input n_383;
input n_834;
input n_112;
input n_765;
input n_893;
input n_1015;
input n_1140;
input n_891;
input n_1651;
input n_239;
input n_630;
input n_55;
input n_504;
input n_511;
input n_874;
input n_358;
input n_1101;
input n_77;
input n_102;
input n_1106;
input n_1456;
input n_1304;
input n_1324;
input n_987;
input n_261;
input n_174;
input n_1455;
input n_767;
input n_993;
input n_1407;
input n_1551;
input n_545;
input n_441;
input n_860;
input n_450;
input n_429;
input n_948;
input n_1217;
input n_628;
input n_365;
input n_729;
input n_1131;
input n_1084;
input n_970;
input n_911;
input n_1430;
input n_83;
input n_513;
input n_1094;
input n_1354;
input n_560;
input n_1534;
input n_340;
input n_1351;
input n_1044;
input n_1205;
input n_346;
input n_1209;
input n_1552;
input n_495;
input n_602;
input n_574;
input n_1435;
input n_879;
input n_16;
input n_58;
input n_623;
input n_405;
input n_824;
input n_359;
input n_1645;
input n_490;
input n_1327;
input n_996;
input n_921;
input n_1684;
input n_233;
input n_1717;
input n_572;
input n_366;
input n_815;
input n_128;
input n_120;
input n_327;
input n_135;
input n_1381;
input n_1611;
input n_1037;
input n_1080;
input n_1274;
input n_1316;
input n_1708;
input n_426;
input n_1438;
input n_1082;
input n_589;
input n_716;
input n_1630;
input n_562;
input n_1436;
input n_62;
input n_1691;
input n_952;
input n_1229;
input n_391;
input n_701;
input n_1437;
input n_1023;
input n_645;
input n_539;
input n_803;
input n_1092;
input n_238;
input n_531;
input n_890;
input n_764;
input n_1056;
input n_1424;
input n_162;
input n_960;
input n_222;
input n_1290;
input n_1123;
input n_1467;
input n_1047;
input n_634;
input n_199;
input n_32;
input n_1252;
input n_348;
input n_1382;
input n_1029;
input n_925;
input n_1206;
input n_424;
input n_1311;
input n_1519;
input n_256;
input n_950;
input n_1553;
input n_380;
input n_419;
input n_1346;
input n_444;
input n_1299;
input n_1060;
input n_1141;
input n_316;
input n_389;
input n_418;
input n_248;
input n_136;
input n_86;
input n_146;
input n_912;
input n_315;
input n_968;
input n_451;
input n_619;
input n_408;
input n_1386;
input n_1699;
input n_376;
input n_967;
input n_1442;
input n_74;
input n_1139;
input n_515;
input n_57;
input n_351;
input n_885;
input n_397;
input n_1432;
input n_1357;
input n_483;
input n_683;
input n_1632;
input n_1057;
input n_1051;
input n_1085;
input n_1066;
input n_721;
input n_1157;
input n_841;
input n_1050;
input n_22;
input n_802;
input n_46;
input n_1608;
input n_983;
input n_38;
input n_280;
input n_1305;
input n_873;
input n_378;
input n_1112;
input n_762;
input n_1283;
input n_1644;
input n_17;
input n_690;
input n_33;
input n_583;
input n_302;
input n_1343;
input n_1203;
input n_1631;
input n_821;
input n_321;
input n_1179;
input n_621;
input n_753;
input n_455;
input n_1048;
input n_1719;
input n_1288;
input n_212;
input n_385;
input n_507;
input n_1560;
input n_1605;
input n_330;
input n_1228;
input n_972;
input n_692;
input n_820;
input n_1200;
input n_1301;
input n_1363;
input n_1668;
input n_1185;
input n_991;
input n_828;
input n_779;
input n_576;
input n_1143;
input n_1579;
input n_1329;
input n_1312;
input n_1439;
input n_804;
input n_537;
input n_1688;
input n_945;
input n_492;
input n_153;
input n_1504;
input n_943;
input n_341;
input n_250;
input n_992;
input n_543;
input n_260;
input n_842;
input n_650;
input n_984;
input n_694;
input n_286;
input n_1643;
input n_883;
input n_470;
input n_325;
input n_449;
input n_1594;
input n_132;
input n_1214;
input n_1342;
input n_1400;
input n_900;
input n_856;
input n_918;
input n_942;
input n_189;
input n_1147;
input n_1557;
input n_1610;
input n_13;
input n_1077;
input n_1422;
input n_540;
input n_618;
input n_896;
input n_323;
input n_195;
input n_356;
input n_894;
input n_1636;
input n_1730;
input n_831;
input n_964;
input n_1373;
input n_1350;
input n_1511;
input n_1470;
input n_1096;
input n_234;
input n_1575;
input n_1697;
input n_1735;
input n_833;
input n_5;
input n_1646;
input n_225;
input n_1307;
input n_988;
input n_814;
input n_192;
input n_1549;
input n_1201;
input n_1114;
input n_655;
input n_1616;
input n_1446;
input n_669;
input n_472;
input n_1458;
input n_1176;
input n_1472;
input n_387;
input n_1149;
input n_398;
input n_1671;
input n_635;
input n_763;
input n_1020;
input n_1062;
input n_211;
input n_1219;
input n_3;
input n_1204;
input n_178;
input n_1035;
input n_287;
input n_555;
input n_783;
input n_1188;
input n_1722;
input n_661;
input n_41;
input n_849;
input n_15;
input n_336;
input n_584;
input n_681;
input n_1638;
input n_50;
input n_430;
input n_510;
input n_216;
input n_311;
input n_830;
input n_1296;
input n_1413;
input n_801;
input n_241;
input n_875;
input n_357;
input n_1110;
input n_1655;
input n_445;
input n_749;
input n_1134;
input n_1358;
input n_717;
input n_165;
input n_939;
input n_482;
input n_1088;
input n_588;
input n_1173;
input n_789;
input n_1232;
input n_1603;
input n_734;
input n_638;
input n_866;
input n_107;
input n_969;
input n_1401;
input n_1019;
input n_1105;
input n_249;
input n_304;
input n_1338;
input n_577;
input n_1522;
input n_1687;
input n_1637;
input n_1419;
input n_338;
input n_149;
input n_1653;
input n_693;
input n_1506;
input n_14;
input n_836;
input n_990;
input n_1389;
input n_975;
input n_1256;
input n_1702;
input n_567;
input n_1465;
input n_778;
input n_1122;
input n_151;
input n_306;
input n_458;
input n_770;
input n_1375;
input n_1102;
input n_711;
input n_1499;
input n_85;
input n_1187;
input n_1441;
input n_1392;
input n_1597;
input n_1164;
input n_1659;
input n_489;
input n_1174;
input n_1371;
input n_617;
input n_1303;
input n_1572;
input n_876;
input n_1516;
input n_1190;
input n_1736;
input n_1685;
input n_118;
input n_601;
input n_917;
input n_1714;
input n_966;
input n_253;
input n_1116;
input n_1661;
input n_1212;
input n_1541;
input n_172;
input n_206;
input n_217;
input n_726;
input n_982;
input n_1573;
input n_1453;
input n_1731;
input n_818;
input n_861;
input n_1713;
input n_1183;
input n_1658;
input n_899;
input n_1253;
input n_210;
input n_1737;
input n_774;
input n_1628;
input n_1335;
input n_1514;
input n_1059;
input n_1345;
input n_176;
input n_1133;
input n_557;
input n_1410;
input n_1005;
input n_607;
input n_1003;
input n_679;
input n_710;
input n_527;
input n_1168;
input n_707;
input n_937;
input n_1427;
input n_393;
input n_108;
input n_487;
input n_1584;
input n_665;
input n_1726;
input n_66;
input n_1440;
input n_177;
input n_421;
input n_1356;
input n_910;
input n_1657;
input n_768;
input n_1475;
input n_1302;
input n_1725;
input n_205;
input n_1136;
input n_1313;
input n_1491;
input n_754;
input n_1496;
input n_179;
input n_1125;
input n_125;
input n_410;
input n_708;
input n_529;
input n_735;
input n_232;
input n_1109;
input n_126;
input n_895;
input n_1310;
input n_202;
input n_427;
input n_1399;
input n_1543;
input n_791;
input n_732;
input n_1533;
input n_193;
input n_808;
input n_797;
input n_1025;
input n_500;
input n_1067;
input n_1720;
input n_148;
input n_435;
input n_159;
input n_766;
input n_1457;
input n_541;
input n_538;
input n_1117;
input n_799;
input n_687;
input n_715;
input n_1480;
input n_1482;
input n_1213;
input n_1266;
input n_536;
input n_872;
input n_594;
input n_200;
input n_1291;
input n_1297;
input n_1155;
input n_1418;
input n_89;
input n_1524;
input n_1689;
input n_1485;
input n_115;
input n_1011;
input n_1184;
input n_985;
input n_869;
input n_810;
input n_416;
input n_827;
input n_401;
input n_1703;
input n_1352;
input n_626;
input n_1650;
input n_1144;
input n_1137;
input n_1570;
input n_1170;
input n_305;
input n_137;
input n_676;
input n_294;
input n_318;
input n_653;
input n_642;
input n_1602;
input n_194;
input n_855;
input n_1178;
input n_1461;
input n_850;
input n_684;
input n_124;
input n_268;
input n_664;
input n_503;
input n_235;
input n_1372;
input n_605;
input n_1273;
input n_353;
input n_620;
input n_643;
input n_916;
input n_1081;
input n_493;
input n_1235;
input n_703;
input n_698;
input n_980;
input n_1115;
input n_1282;
input n_1318;
input n_780;
input n_998;
input n_1454;
input n_467;
input n_1227;
input n_1531;
input n_840;
input n_1334;
input n_501;
input n_823;
input n_245;
input n_725;
input n_1388;
input n_1417;
input n_1295;
input n_672;
input n_581;
input n_382;
input n_554;
input n_1625;
input n_898;
input n_1013;
input n_1452;
input n_718;
input n_265;
input n_1120;
input n_719;
input n_443;
input n_198;
input n_714;
input n_1683;
input n_909;
input n_1497;
input n_1530;
input n_997;
input n_932;
input n_612;
input n_1409;
input n_788;
input n_1326;
input n_119;
input n_1268;
input n_559;
input n_825;
input n_508;
input n_506;
input n_1320;
input n_1663;
input n_737;
input n_1718;
input n_986;
input n_509;
input n_1317;
input n_147;
input n_1518;
input n_1715;
input n_1281;
input n_67;
input n_1192;
input n_1024;
input n_1063;
input n_209;
input n_1564;
input n_1613;
input n_733;
input n_1489;
input n_1376;
input n_941;
input n_981;
input n_1569;
input n_68;
input n_867;
input n_186;
input n_134;
input n_587;
input n_63;
input n_792;
input n_756;
input n_1429;
input n_399;
input n_1238;
input n_548;
input n_812;
input n_298;
input n_518;
input n_505;
input n_282;
input n_752;
input n_905;
input n_1476;
input n_1108;
input n_782;
input n_1100;
input n_1395;
input n_862;
input n_1425;
input n_760;
input n_1620;
input n_381;
input n_220;
input n_390;
input n_1330;
input n_31;
input n_481;
input n_1675;
input n_1727;
input n_1554;
input n_769;
input n_42;
input n_1046;
input n_271;
input n_934;
input n_1618;
input n_826;
input n_886;
input n_1221;
input n_654;
input n_1172;
input n_167;
input n_379;
input n_428;
input n_1341;
input n_570;
input n_1641;
input n_1361;
input n_1707;
input n_853;
input n_377;
input n_751;
input n_786;
input n_1083;
input n_1142;
input n_1129;
input n_392;
input n_158;
input n_704;
input n_787;
input n_138;
input n_961;
input n_771;
input n_276;
input n_95;
input n_1716;
input n_1225;
input n_1520;
input n_169;
input n_522;
input n_1287;
input n_1262;
input n_400;
input n_930;
input n_181;
input n_1411;
input n_221;
input n_622;
input n_1577;
input n_1087;
input n_386;
input n_994;
input n_1701;
input n_848;
input n_1550;
input n_1498;
input n_1223;
input n_1272;
input n_104;
input n_682;
input n_1567;
input n_56;
input n_141;
input n_1247;
input n_922;
input n_816;
input n_1648;
input n_591;
input n_145;
input n_1536;
input n_1344;
input n_313;
input n_631;
input n_479;
input n_1246;
input n_1339;
input n_1478;
input n_432;
input n_839;
input n_1210;
input n_1364;
input n_328;
input n_140;
input n_1250;
input n_369;
input n_871;
input n_598;
input n_685;
input n_928;
input n_608;
input n_1367;
input n_78;
input n_1460;
input n_772;
input n_1555;
input n_499;
input n_1589;
input n_517;
input n_98;
input n_402;
input n_413;
input n_1086;
input n_796;
input n_1619;
input n_236;
input n_1502;
input n_1469;
input n_1012;
input n_1;
input n_1396;
input n_1348;
input n_903;
input n_1525;
input n_740;
input n_203;
input n_384;
input n_1404;
input n_80;
input n_35;
input n_1315;
input n_277;
input n_1061;
input n_92;
input n_333;
input n_1298;
input n_1652;
input n_462;
input n_1193;
input n_1676;
input n_1255;
input n_258;
input n_1113;
input n_29;
input n_79;
input n_1226;
input n_722;
input n_1277;
input n_188;
input n_844;
input n_201;
input n_471;
input n_852;
input n_1487;
input n_40;
input n_1028;
input n_1601;
input n_781;
input n_474;
input n_542;
input n_463;
input n_1546;
input n_595;
input n_502;
input n_466;
input n_420;
input n_1337;
input n_1495;
input n_632;
input n_699;
input n_979;
input n_1515;
input n_1627;
input n_1245;
input n_846;
input n_1673;
input n_465;
input n_76;
input n_362;
input n_1321;
input n_170;
input n_27;
input n_161;
input n_273;
input n_585;
input n_270;
input n_616;
input n_81;
input n_745;
input n_1654;
input n_1103;
input n_648;
input n_1379;
input n_312;
input n_1076;
input n_1091;
input n_1408;
input n_494;
input n_641;
input n_730;
input n_1325;
input n_1595;
input n_354;
input n_575;
input n_480;
input n_425;
input n_795;
input n_695;
input n_180;
input n_656;
input n_1606;
input n_1220;
input n_37;
input n_1694;
input n_1540;
input n_229;
input n_437;
input n_1642;
input n_60;
input n_403;
input n_453;
input n_1130;
input n_720;
input n_0;
input n_1526;
input n_863;
input n_805;
input n_1604;
input n_1275;
input n_113;
input n_712;
input n_246;
input n_1583;
input n_1042;
input n_1402;
input n_269;
input n_285;
input n_412;
input n_1493;
input n_657;
input n_644;
input n_1160;
input n_1397;
input n_491;
input n_1258;
input n_1074;
input n_1621;
input n_251;
input n_160;
input n_566;
input n_565;
input n_1448;
input n_1507;
input n_1398;
input n_597;
input n_1181;
input n_1505;
input n_1634;
input n_1196;
input n_651;
input n_1340;
input n_334;
input n_811;
input n_1558;
input n_807;
input n_835;
input n_175;
input n_666;
input n_262;
input n_1433;
input n_1704;
input n_99;
input n_1254;
input n_1026;
input n_1234;
input n_319;
input n_364;
input n_1138;
input n_927;
input n_20;
input n_1089;
input n_1004;
input n_1186;
input n_1032;
input n_242;
input n_1681;
input n_1018;
input n_1693;
input n_438;
input n_713;
input n_904;
input n_1588;
input n_1622;
input n_166;
input n_1180;
input n_1271;
input n_533;
input n_1542;
input n_1251;
input n_278;

output n_7499;

wire n_6643;
wire n_6122;
wire n_2253;
wire n_2417;
wire n_2756;
wire n_4706;
wire n_5567;
wire n_2380;
wire n_3241;
wire n_3006;
wire n_6579;
wire n_7164;
wire n_5287;
wire n_6546;
wire n_2327;
wire n_2899;
wire n_5484;
wire n_3619;
wire n_3541;
wire n_3622;
wire n_5978;
wire n_2395;
wire n_5161;
wire n_5776;
wire n_6551;
wire n_5512;
wire n_5207;
wire n_2347;
wire n_6786;
wire n_7206;
wire n_7303;
wire n_4963;
wire n_4240;
wire n_4508;
wire n_2021;
wire n_2391;
wire n_5035;
wire n_5282;
wire n_1960;
wire n_2843;
wire n_3615;
wire n_2059;
wire n_7461;
wire n_2487;
wire n_6649;
wire n_7154;
wire n_3202;
wire n_4977;
wire n_3813;
wire n_6810;
wire n_6276;
wire n_6072;
wire n_3341;
wire n_3587;
wire n_4128;
wire n_3445;
wire n_2001;
wire n_4145;
wire n_3785;
wire n_5033;
wire n_4211;
wire n_7024;
wire n_3448;
wire n_7205;
wire n_6742;
wire n_3019;
wire n_2096;
wire n_6694;
wire n_3776;
wire n_2530;
wire n_4517;
wire n_2483;
wire n_7486;
wire n_4425;
wire n_4950;
wire n_4988;
wire n_1860;
wire n_4615;
wire n_2076;
wire n_6090;
wire n_6580;
wire n_7010;
wire n_5480;
wire n_6549;
wire n_6913;
wire n_2147;
wire n_3010;
wire n_7315;
wire n_7004;
wire n_2770;
wire n_4131;
wire n_5402;
wire n_2584;
wire n_5851;
wire n_3188;
wire n_5509;
wire n_3403;
wire n_3624;
wire n_3461;
wire n_3082;
wire n_2189;
wire n_3796;
wire n_5154;
wire n_3283;
wire n_7468;
wire n_5469;
wire n_2323;
wire n_6431;
wire n_5744;
wire n_2597;
wire n_3340;
wire n_3277;
wire n_5453;
wire n_2052;
wire n_4499;
wire n_4927;
wire n_5202;
wire n_5648;
wire n_6931;
wire n_6618;
wire n_6408;
wire n_3214;
wire n_2091;
wire n_4311;
wire n_3631;
wire n_3806;
wire n_4691;
wire n_5922;
wire n_6698;
wire n_4678;
wire n_2032;
wire n_2587;
wire n_5848;
wire n_5406;
wire n_6085;
wire n_3947;
wire n_3490;
wire n_7421;
wire n_7306;
wire n_6214;
wire n_7493;
wire n_1948;
wire n_3868;
wire n_3183;
wire n_3437;
wire n_3353;
wire n_4203;
wire n_3687;
wire n_5241;
wire n_6939;
wire n_2384;
wire n_3156;
wire n_3376;
wire n_5037;
wire n_4468;
wire n_5661;
wire n_6991;
wire n_3653;
wire n_5562;
wire n_3702;
wire n_4976;
wire n_6586;
wire n_2202;
wire n_2648;
wire n_5008;
wire n_2159;
wire n_2976;
wire n_3876;
wire n_2353;
wire n_2439;
wire n_4811;
wire n_5398;
wire n_6096;
wire n_2276;
wire n_6707;
wire n_5852;
wire n_2089;
wire n_3420;
wire n_6920;
wire n_6868;
wire n_5144;
wire n_3361;
wire n_4758;
wire n_7402;
wire n_4255;
wire n_1796;
wire n_5577;
wire n_4484;
wire n_3668;
wire n_7152;
wire n_6512;
wire n_4237;
wire n_2934;
wire n_1880;
wire n_3550;
wire n_5689;
wire n_5894;
wire n_2079;
wire n_2238;
wire n_7463;
wire n_3418;
wire n_4901;
wire n_6725;
wire n_2859;
wire n_3395;
wire n_7083;
wire n_4917;
wire n_7086;
wire n_7349;
wire n_6464;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_5825;
wire n_2968;
wire n_7316;
wire n_6820;
wire n_2684;
wire n_3593;
wire n_5343;
wire n_4421;
wire n_6098;
wire n_7019;
wire n_6686;
wire n_4836;
wire n_5062;
wire n_4020;
wire n_2730;
wire n_2251;
wire n_3915;
wire n_4469;
wire n_4414;
wire n_6561;
wire n_6584;
wire n_7452;
wire n_5184;
wire n_4532;
wire n_3339;
wire n_3735;
wire n_3349;
wire n_7323;
wire n_2248;
wire n_7195;
wire n_6701;
wire n_7478;
wire n_3007;
wire n_6769;
wire n_6592;
wire n_5686;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_5463;
wire n_2100;
wire n_5236;
wire n_3487;
wire n_3310;
wire n_6062;
wire n_6191;
wire n_2258;
wire n_3983;
wire n_4405;
wire n_5433;
wire n_1926;
wire n_4195;
wire n_4969;
wire n_4504;
wire n_5909;
wire n_2776;
wire n_4408;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_4531;
wire n_6043;
wire n_2987;
wire n_6271;
wire n_7171;
wire n_4567;
wire n_4164;
wire n_5315;
wire n_4234;
wire n_4130;
wire n_3611;
wire n_2862;
wire n_5348;
wire n_2175;
wire n_5055;
wire n_6793;
wire n_2324;
wire n_2606;
wire n_3187;
wire n_2828;
wire n_7127;
wire n_5397;
wire n_4471;
wire n_6550;
wire n_5031;
wire n_3392;
wire n_3975;
wire n_3430;
wire n_4444;
wire n_5709;
wire n_3208;
wire n_6021;
wire n_3331;
wire n_4983;
wire n_2379;
wire n_5695;
wire n_2911;
wire n_2154;
wire n_4916;
wire n_5860;
wire n_6926;
wire n_3649;
wire n_4302;
wire n_6928;
wire n_2514;
wire n_5862;
wire n_6304;
wire n_5189;
wire n_6956;
wire n_5381;
wire n_4786;
wire n_3257;
wire n_7026;
wire n_4160;
wire n_6782;
wire n_2293;
wire n_5854;
wire n_5516;
wire n_4051;
wire n_2028;
wire n_3009;
wire n_7002;
wire n_3981;
wire n_7141;
wire n_5936;
wire n_6126;
wire n_1841;
wire n_6027;
wire n_6598;
wire n_2581;
wire n_3224;
wire n_4647;
wire n_3752;
wire n_6342;
wire n_6638;
wire n_1891;
wire n_7308;
wire n_5254;
wire n_3526;
wire n_6900;
wire n_2546;
wire n_3790;
wire n_7264;
wire n_3491;
wire n_7457;
wire n_4613;
wire n_4649;
wire n_1888;
wire n_6269;
wire n_5615;
wire n_1963;
wire n_4795;
wire n_2226;
wire n_2891;
wire n_5902;
wire n_4028;
wire n_5479;
wire n_3819;
wire n_6013;
wire n_7357;
wire n_2449;
wire n_5083;
wire n_6927;
wire n_6503;
wire n_5888;
wire n_4186;
wire n_2297;
wire n_7310;
wire n_4731;
wire n_1759;
wire n_2177;
wire n_3747;
wire n_5698;
wire n_5592;
wire n_2227;
wire n_4618;
wire n_2190;
wire n_3346;
wire n_4742;
wire n_6256;
wire n_2876;
wire n_4099;
wire n_7406;
wire n_3484;
wire n_3620;
wire n_1746;
wire n_2479;
wire n_5870;
wire n_4295;
wire n_5303;
wire n_7076;
wire n_4694;
wire n_4533;
wire n_3038;
wire n_5081;
wire n_5124;
wire n_3068;
wire n_2871;
wire n_5807;
wire n_5863;
wire n_5943;
wire n_4244;
wire n_4603;
wire n_2943;
wire n_4254;
wire n_3143;
wire n_3168;
wire n_6982;
wire n_4697;
wire n_7286;
wire n_7137;
wire n_2607;
wire n_3994;
wire n_4190;
wire n_4810;
wire n_6727;
wire n_3317;
wire n_7229;
wire n_4391;
wire n_5954;
wire n_3263;
wire n_2582;
wire n_4157;
wire n_4283;
wire n_4681;
wire n_4638;
wire n_3455;
wire n_6097;
wire n_5047;
wire n_3452;
wire n_5346;
wire n_1994;
wire n_5517;
wire n_7125;
wire n_6677;
wire n_4707;
wire n_2577;
wire n_4527;
wire n_5109;
wire n_6624;
wire n_7121;
wire n_2796;
wire n_6466;
wire n_2342;
wire n_4156;
wire n_1851;
wire n_4848;
wire n_2937;
wire n_6008;
wire n_3095;
wire n_2805;
wire n_5624;
wire n_4918;
wire n_5714;
wire n_5806;
wire n_3856;
wire n_2914;
wire n_4898;
wire n_1964;
wire n_2869;
wire n_6221;
wire n_7160;
wire n_4002;
wire n_6805;
wire n_6185;
wire n_5010;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_2925;
wire n_3773;
wire n_3918;
wire n_2398;
wire n_6568;
wire n_2857;
wire n_5358;
wire n_4528;
wire n_3932;
wire n_4619;
wire n_4673;
wire n_6004;
wire n_6351;
wire n_3516;
wire n_4822;
wire n_2155;
wire n_2516;
wire n_3797;
wire n_6901;
wire n_2947;
wire n_5580;
wire n_4299;
wire n_5937;
wire n_4801;
wire n_7183;
wire n_6411;
wire n_3515;
wire n_2886;
wire n_2093;
wire n_2473;
wire n_3287;
wire n_3378;
wire n_5435;
wire n_6873;
wire n_4279;
wire n_4769;
wire n_4632;
wire n_5373;
wire n_5745;
wire n_7139;
wire n_4294;
wire n_5279;
wire n_4125;
wire n_4232;
wire n_4949;
wire n_2941;
wire n_6594;
wire n_2457;
wire n_5493;
wire n_4790;
wire n_2536;
wire n_6387;
wire n_7223;
wire n_1758;
wire n_2952;
wire n_4847;
wire n_6179;
wire n_7338;
wire n_5321;
wire n_3058;
wire n_5096;
wire n_4365;
wire n_1878;
wire n_6019;
wire n_6222;
wire n_7165;
wire n_3505;
wire n_6223;
wire n_4610;
wire n_6435;
wire n_3730;
wire n_4489;
wire n_7235;
wire n_5210;
wire n_6976;
wire n_4967;
wire n_6486;
wire n_5657;
wire n_6889;
wire n_6083;
wire n_4992;
wire n_6844;
wire n_3001;
wire n_7404;
wire n_3945;
wire n_4542;
wire n_2261;
wire n_2729;
wire n_6295;
wire n_3597;
wire n_2897;
wire n_2077;
wire n_4198;
wire n_2909;
wire n_5857;
wire n_4534;
wire n_4500;
wire n_7437;
wire n_5014;
wire n_6241;
wire n_3185;
wire n_6087;
wire n_3523;
wire n_1785;
wire n_2829;
wire n_4597;
wire n_6846;
wire n_4329;
wire n_4087;
wire n_3811;
wire n_3200;
wire n_5756;
wire n_2231;
wire n_6041;
wire n_2017;
wire n_2604;
wire n_6994;
wire n_4257;
wire n_3453;
wire n_7449;
wire n_7329;
wire n_2390;
wire n_5708;
wire n_3213;
wire n_6790;
wire n_3077;
wire n_7194;
wire n_6273;
wire n_3474;
wire n_3984;
wire n_6807;
wire n_5927;
wire n_2151;
wire n_2106;
wire n_2716;
wire n_4665;
wire n_1913;
wire n_1823;
wire n_3679;
wire n_3422;
wire n_3888;
wire n_5638;
wire n_7115;
wire n_4189;
wire n_5670;
wire n_1875;
wire n_2803;
wire n_3707;
wire n_1846;
wire n_5584;
wire n_3429;
wire n_1903;
wire n_3849;
wire n_3946;
wire n_5965;
wire n_3229;
wire n_4463;
wire n_1805;
wire n_4687;
wire n_5751;
wire n_5664;
wire n_4670;
wire n_4084;
wire n_4703;
wire n_5641;
wire n_4037;
wire n_6218;
wire n_7281;
wire n_2922;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_2727;
wire n_3421;
wire n_2240;
wire n_2436;
wire n_6824;
wire n_6189;
wire n_3618;
wire n_2593;
wire n_5262;
wire n_6993;
wire n_3683;
wire n_6037;
wire n_7245;
wire n_3642;
wire n_3286;
wire n_3808;
wire n_5963;
wire n_5980;
wire n_4763;
wire n_3590;
wire n_5310;
wire n_4594;
wire n_6153;
wire n_3424;
wire n_5970;
wire n_6418;
wire n_6564;
wire n_2301;
wire n_3583;
wire n_3560;
wire n_4076;
wire n_4714;
wire n_3215;
wire n_2419;
wire n_5146;
wire n_4776;
wire n_2122;
wire n_2512;
wire n_4102;
wire n_2786;
wire n_7192;
wire n_3171;
wire n_6671;
wire n_6591;
wire n_6266;
wire n_7161;
wire n_7153;
wire n_5213;
wire n_3020;
wire n_3677;
wire n_3462;
wire n_5441;
wire n_6517;
wire n_3468;
wire n_2910;
wire n_1893;
wire n_7350;
wire n_5690;
wire n_2163;
wire n_6967;
wire n_5885;
wire n_2254;
wire n_6433;
wire n_3546;
wire n_6893;
wire n_2647;
wire n_4443;
wire n_5461;
wire n_4507;
wire n_7178;
wire n_7480;
wire n_2443;
wire n_1811;
wire n_2624;
wire n_3012;
wire n_4575;
wire n_3244;
wire n_6501;
wire n_6028;
wire n_3130;
wire n_3822;
wire n_3569;
wire n_5629;
wire n_4452;
wire n_4348;
wire n_5634;
wire n_5430;
wire n_5362;
wire n_6709;
wire n_4355;
wire n_3494;
wire n_6798;
wire n_5702;
wire n_5050;
wire n_5063;
wire n_5229;
wire n_3771;
wire n_2125;
wire n_5199;
wire n_3110;
wire n_3073;
wire n_4572;
wire n_5527;
wire n_6986;
wire n_5609;
wire n_5416;
wire n_4026;
wire n_2265;
wire n_4104;
wire n_4512;
wire n_3554;
wire n_4377;
wire n_5266;
wire n_7471;
wire n_3178;
wire n_5355;
wire n_2334;
wire n_6745;
wire n_4521;
wire n_4488;
wire n_5977;
wire n_6811;
wire n_2289;
wire n_3051;
wire n_2783;
wire n_6209;
wire n_2263;
wire n_6875;
wire n_3750;
wire n_2341;
wire n_3632;
wire n_4588;
wire n_2733;
wire n_2785;
wire n_2415;
wire n_3299;
wire n_6853;
wire n_4519;
wire n_5551;
wire n_3715;
wire n_7340;
wire n_6699;
wire n_6073;
wire n_5767;
wire n_6324;
wire n_3040;
wire n_1938;
wire n_5640;
wire n_2499;
wire n_3568;
wire n_5655;
wire n_5475;
wire n_3737;
wire n_6138;
wire n_1967;
wire n_3255;
wire n_5692;
wire n_4856;
wire n_7494;
wire n_2997;
wire n_5921;
wire n_4400;
wire n_5168;
wire n_3326;
wire n_6477;
wire n_3734;
wire n_4778;
wire n_2429;
wire n_6159;
wire n_6283;
wire n_7396;
wire n_5322;
wire n_7116;
wire n_1793;
wire n_4352;
wire n_4441;
wire n_6943;
wire n_4761;
wire n_6827;
wire n_6173;
wire n_1804;
wire n_4347;
wire n_4095;
wire n_3196;
wire n_4593;
wire n_6312;
wire n_2533;
wire n_2364;
wire n_3492;
wire n_2780;
wire n_4727;
wire n_4568;
wire n_5371;
wire n_2291;
wire n_4043;
wire n_3601;
wire n_6997;
wire n_5418;
wire n_1865;
wire n_2973;
wire n_2094;
wire n_2393;
wire n_5316;
wire n_3831;
wire n_3801;
wire n_6300;
wire n_2043;
wire n_2751;
wire n_6131;
wire n_4893;
wire n_5032;
wire n_1934;
wire n_6537;
wire n_5933;
wire n_4948;
wire n_4000;
wire n_3240;
wire n_2025;
wire n_4406;
wire n_2758;
wire n_7023;
wire n_1807;
wire n_2618;
wire n_7428;
wire n_5112;
wire n_5386;
wire n_2559;
wire n_6783;
wire n_4748;
wire n_7465;
wire n_2295;
wire n_3931;
wire n_4010;
wire n_2840;
wire n_5017;
wire n_1814;
wire n_2822;
wire n_4710;
wire n_4607;
wire n_5123;
wire n_4117;
wire n_3636;
wire n_2441;
wire n_1802;
wire n_3083;
wire n_4487;
wire n_5001;
wire n_7149;
wire n_2795;
wire n_6459;
wire n_2981;
wire n_2282;
wire n_2800;
wire n_4817;
wire n_3380;
wire n_5644;
wire n_2098;
wire n_3460;
wire n_3409;
wire n_3538;
wire n_6869;
wire n_2068;
wire n_4849;
wire n_4867;
wire n_5424;
wire n_3198;
wire n_2641;
wire n_1895;
wire n_4728;
wire n_7117;
wire n_4247;
wire n_4933;
wire n_6977;
wire n_4018;
wire n_3900;
wire n_4902;
wire n_4518;
wire n_4409;
wire n_4411;
wire n_6313;
wire n_3872;
wire n_4336;
wire n_6569;
wire n_2270;
wire n_4777;
wire n_2653;
wire n_2496;
wire n_1908;
wire n_2259;
wire n_6555;
wire n_3877;
wire n_6639;
wire n_2995;
wire n_5496;
wire n_2494;
wire n_3547;
wire n_3977;
wire n_4052;
wire n_5864;
wire n_6536;
wire n_3459;
wire n_4398;
wire n_3155;
wire n_6490;
wire n_2633;
wire n_6961;
wire n_4954;
wire n_2435;
wire n_2097;
wire n_5460;
wire n_4304;
wire n_6761;
wire n_3911;
wire n_5333;
wire n_6294;
wire n_6767;
wire n_4431;
wire n_7427;
wire n_4192;
wire n_6802;
wire n_5570;
wire n_3736;
wire n_6326;
wire n_4805;
wire n_4885;
wire n_5983;
wire n_5804;
wire n_6376;
wire n_3565;
wire n_6167;
wire n_4701;
wire n_2575;
wire n_5910;
wire n_7411;
wire n_7101;
wire n_5040;
wire n_6730;
wire n_6948;
wire n_6582;
wire n_1904;
wire n_6996;
wire n_1899;
wire n_6974;
wire n_6765;
wire n_6921;
wire n_2067;
wire n_2219;
wire n_3533;
wire n_2877;
wire n_2148;
wire n_4631;
wire n_3035;
wire n_5194;
wire n_6898;
wire n_6710;
wire n_5717;
wire n_7162;
wire n_5464;
wire n_6565;
wire n_5886;
wire n_7080;
wire n_3639;
wire n_7302;
wire n_6533;
wire n_2501;
wire n_3079;
wire n_4965;
wire n_6960;
wire n_6426;
wire n_6634;
wire n_7180;
wire n_1915;
wire n_5610;
wire n_5239;
wire n_6836;
wire n_2605;
wire n_4747;
wire n_5197;
wire n_1979;
wire n_6972;
wire n_2924;
wire n_7111;
wire n_4111;
wire n_2484;
wire n_5785;
wire n_4587;
wire n_3731;
wire n_2946;
wire n_6344;
wire n_5305;
wire n_6093;
wire n_4538;
wire n_5994;
wire n_6010;
wire n_7247;
wire n_6833;
wire n_2754;
wire n_1742;
wire n_5376;
wire n_2489;
wire n_7481;
wire n_5204;
wire n_7292;
wire n_2012;
wire n_4094;
wire n_3503;
wire n_7150;
wire n_2866;
wire n_3561;
wire n_2917;
wire n_2425;
wire n_3536;
wire n_3661;
wire n_4150;
wire n_4878;
wire n_6265;
wire n_6821;
wire n_3934;
wire n_4985;
wire n_6373;
wire n_6988;
wire n_5788;
wire n_3922;
wire n_3846;
wire n_5897;
wire n_6887;
wire n_2103;
wire n_2160;
wire n_2498;
wire n_2697;
wire n_3074;
wire n_1999;
wire n_6676;
wire n_2372;
wire n_3673;
wire n_6347;
wire n_6492;
wire n_7016;
wire n_3768;
wire n_2861;
wire n_2630;
wire n_3943;
wire n_2430;
wire n_2433;
wire n_3293;
wire n_5795;
wire n_7072;
wire n_5508;
wire n_5582;
wire n_4022;
wire n_7374;
wire n_7440;
wire n_4852;
wire n_2528;
wire n_4869;
wire n_4700;
wire n_7201;
wire n_4035;
wire n_2316;
wire n_1898;
wire n_3294;
wire n_4426;
wire n_3415;
wire n_2284;
wire n_5746;
wire n_2817;
wire n_3139;
wire n_5292;
wire n_2598;
wire n_6648;
wire n_4601;
wire n_2687;
wire n_1890;
wire n_4220;
wire n_1944;
wire n_5630;
wire n_3431;
wire n_3169;
wire n_3151;
wire n_2078;
wire n_3284;
wire n_3070;
wire n_4066;
wire n_2884;
wire n_4515;
wire n_4351;
wire n_5264;
wire n_3126;
wire n_7413;
wire n_4403;
wire n_1981;
wire n_4509;
wire n_4858;
wire n_3700;
wire n_5504;
wire n_7005;
wire n_4223;
wire n_7353;
wire n_6219;
wire n_1889;
wire n_6965;
wire n_5025;
wire n_2966;
wire n_2326;
wire n_6720;
wire n_2188;
wire n_6032;
wire n_7174;
wire n_6205;
wire n_6362;
wire n_6402;
wire n_4644;
wire n_7166;
wire n_4456;
wire n_5060;
wire n_5334;
wire n_2448;
wire n_4346;
wire n_3170;
wire n_5775;
wire n_3311;
wire n_2748;
wire n_3272;
wire n_7282;
wire n_6491;
wire n_2898;
wire n_2717;
wire n_7151;
wire n_6229;
wire n_1861;
wire n_5731;
wire n_5581;
wire n_3628;
wire n_3691;
wire n_6668;
wire n_7446;
wire n_4235;
wire n_1867;
wire n_1945;
wire n_3018;
wire n_7053;
wire n_5831;
wire n_2573;
wire n_7473;
wire n_4435;
wire n_2939;
wire n_6835;
wire n_6419;
wire n_6039;
wire n_3807;
wire n_5884;
wire n_2447;
wire n_4764;
wire n_5653;
wire n_6258;
wire n_7070;
wire n_5394;
wire n_6755;
wire n_2774;
wire n_7276;
wire n_7351;
wire n_4655;
wire n_3161;
wire n_4581;
wire n_6084;
wire n_4827;
wire n_7412;
wire n_7157;
wire n_6436;
wire n_2488;
wire n_6472;
wire n_3477;
wire n_5421;
wire n_2476;
wire n_7211;
wire n_4399;
wire n_6531;
wire n_2781;
wire n_5309;
wire n_2778;
wire n_4782;
wire n_4363;
wire n_2887;
wire n_4864;
wire n_2691;
wire n_7368;
wire n_3054;
wire n_4335;
wire n_6567;
wire n_5889;
wire n_6771;
wire n_2526;
wire n_6389;
wire n_2703;
wire n_2167;
wire n_5764;
wire n_5428;
wire n_6910;
wire n_6442;
wire n_3391;
wire n_6102;
wire n_4259;
wire n_5541;
wire n_2709;
wire n_6441;
wire n_5543;
wire n_5678;
wire n_5935;
wire n_4865;
wire n_4056;
wire n_4564;
wire n_3840;
wire n_5085;
wire n_3518;
wire n_2956;
wire n_3733;
wire n_5950;
wire n_2173;
wire n_1842;
wire n_3738;
wire n_5995;
wire n_6162;
wire n_5116;
wire n_3464;
wire n_2018;
wire n_4526;
wire n_6331;
wire n_6006;
wire n_3245;
wire n_4417;
wire n_6109;
wire n_6278;
wire n_6787;
wire n_6872;
wire n_4899;
wire n_6208;
wire n_2119;
wire n_2157;
wire n_2552;
wire n_6632;
wire n_5411;
wire n_2453;
wire n_4798;
wire n_7027;
wire n_3509;
wire n_3352;
wire n_5671;
wire n_3076;
wire n_6990;
wire n_3535;
wire n_2182;
wire n_6349;
wire n_3251;
wire n_2931;
wire n_6830;
wire n_5185;
wire n_6359;
wire n_3118;
wire n_3511;
wire n_3443;
wire n_2146;
wire n_7498;
wire n_3644;
wire n_5076;
wire n_3336;
wire n_3935;
wire n_7377;
wire n_3521;
wire n_5379;
wire n_3562;
wire n_3948;
wire n_4750;
wire n_6301;
wire n_2918;
wire n_3232;
wire n_5945;
wire n_2112;
wire n_1739;
wire n_2958;
wire n_6744;
wire n_4981;
wire n_3114;
wire n_3125;
wire n_2394;
wire n_3612;
wire n_2954;
wire n_4835;
wire n_5811;
wire n_4430;
wire n_6439;
wire n_7381;
wire n_5565;
wire n_4081;
wire n_3132;
wire n_4407;
wire n_7291;
wire n_3951;
wire n_4894;
wire n_5780;
wire n_5643;
wire n_3238;
wire n_3210;
wire n_5846;
wire n_2036;
wire n_7430;
wire n_3267;
wire n_4995;
wire n_5524;
wire n_3964;
wire n_3772;
wire n_1956;
wire n_2279;
wire n_3373;
wire n_4446;
wire n_6104;
wire n_3884;
wire n_6475;
wire n_6465;
wire n_3726;
wire n_6496;
wire n_2525;
wire n_2892;
wire n_2907;
wire n_6998;
wire n_6145;
wire n_3577;
wire n_2820;
wire n_7305;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1741;
wire n_4057;
wire n_4332;
wire n_4314;
wire n_3347;
wire n_3216;
wire n_3809;
wire n_2113;
wire n_7075;
wire n_4288;
wire n_6076;
wire n_3567;
wire n_6194;
wire n_5066;
wire n_3939;
wire n_6092;
wire n_7275;
wire n_5401;
wire n_6357;
wire n_5843;
wire n_4241;
wire n_3321;
wire n_3212;
wire n_3152;
wire n_2256;
wire n_7489;
wire n_5106;
wire n_5468;
wire n_2920;
wire n_4265;
wire n_6335;
wire n_5883;
wire n_6985;
wire n_5319;
wire n_2247;
wire n_7451;
wire n_6238;
wire n_3705;
wire n_6548;
wire n_2802;
wire n_4705;
wire n_3159;
wire n_5455;
wire n_2268;
wire n_3778;
wire n_5706;
wire n_5337;
wire n_6366;
wire n_3304;
wire n_3912;
wire n_7236;
wire n_2739;
wire n_2771;
wire n_4604;
wire n_7269;
wire n_5223;
wire n_5962;
wire n_3795;
wire n_5020;
wire n_6602;
wire n_4419;
wire n_4477;
wire n_6620;
wire n_3179;
wire n_6502;
wire n_3256;
wire n_7326;
wire n_7060;
wire n_2386;
wire n_3086;
wire n_6885;
wire n_2369;
wire n_2927;
wire n_4217;
wire n_4395;
wire n_2821;
wire n_5074;
wire n_2568;
wire n_5364;
wire n_6529;
wire n_1738;
wire n_3728;
wire n_3064;
wire n_3088;
wire n_5895;
wire n_4639;
wire n_6951;
wire n_3713;
wire n_3663;
wire n_5649;
wire n_5046;
wire n_5166;
wire n_7169;
wire n_6423;
wire n_3246;
wire n_2495;
wire n_1789;
wire n_7140;
wire n_7233;
wire n_5088;
wire n_2302;
wire n_6558;
wire n_5457;
wire n_7352;
wire n_7134;
wire n_5532;
wire n_2069;
wire n_6950;
wire n_7246;
wire n_6525;
wire n_3434;
wire n_1806;
wire n_6631;
wire n_6892;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_2024;
wire n_4780;
wire n_7056;
wire n_4243;
wire n_4982;
wire n_3695;
wire n_4330;
wire n_6683;
wire n_2482;
wire n_2677;
wire n_6292;
wire n_5544;
wire n_3832;
wire n_3987;
wire n_7339;
wire n_5987;
wire n_6180;
wire n_5352;
wire n_5824;
wire n_4991;
wire n_5538;
wire n_6658;
wire n_6264;
wire n_6925;
wire n_5919;
wire n_2329;
wire n_2142;
wire n_6176;
wire n_5410;
wire n_3332;
wire n_7146;
wire n_3048;
wire n_3937;
wire n_6124;
wire n_2203;
wire n_4525;
wire n_3782;
wire n_7482;
wire n_6864;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_4208;
wire n_7090;
wire n_3786;
wire n_7158;
wire n_2888;
wire n_7156;
wire n_5742;
wire n_3638;
wire n_5992;
wire n_6494;
wire n_5503;
wire n_4177;
wire n_6199;
wire n_3763;
wire n_2669;
wire n_1778;
wire n_2306;
wire n_5958;
wire n_6614;
wire n_3022;
wire n_4264;
wire n_3087;
wire n_3489;
wire n_2566;
wire n_7360;
wire n_7301;
wire n_5129;
wire n_2149;
wire n_7375;
wire n_7102;
wire n_5500;
wire n_3060;
wire n_4276;
wire n_7366;
wire n_5219;
wire n_5605;
wire n_3013;
wire n_1984;
wire n_5170;
wire n_5654;
wire n_2408;
wire n_7025;
wire n_5320;
wire n_1877;
wire n_3049;
wire n_6947;
wire n_5107;
wire n_5999;
wire n_4485;
wire n_7309;
wire n_4626;
wire n_6863;
wire n_6637;
wire n_6100;
wire n_6735;
wire n_2659;
wire n_4975;
wire n_6358;
wire n_1852;
wire n_5602;
wire n_3089;
wire n_6050;
wire n_2470;
wire n_7244;
wire n_5405;
wire n_3985;
wire n_5253;
wire n_4760;
wire n_4652;
wire n_4624;
wire n_2551;
wire n_2682;
wire n_5903;
wire n_6371;
wire n_7043;
wire n_3440;
wire n_6171;
wire n_6510;
wire n_1748;
wire n_4569;
wire n_6468;
wire n_2699;
wire n_4897;
wire n_2769;
wire n_3542;
wire n_3436;
wire n_5491;
wire n_2615;
wire n_3940;
wire n_5842;
wire n_6352;
wire n_2985;
wire n_5722;
wire n_5636;
wire n_5065;
wire n_2753;
wire n_7287;
wire n_7032;
wire n_3637;
wire n_2842;
wire n_4523;
wire n_1836;
wire n_2868;
wire n_5492;
wire n_3141;
wire n_5084;
wire n_6850;
wire n_5667;
wire n_3164;
wire n_3570;
wire n_5260;
wire n_7119;
wire n_4919;
wire n_4025;
wire n_2712;
wire n_5328;
wire n_3936;
wire n_6354;
wire n_5918;
wire n_4503;
wire n_3507;
wire n_6959;
wire n_3821;
wire n_6909;
wire n_2700;
wire n_6332;
wire n_3367;
wire n_4464;
wire n_7006;
wire n_5877;
wire n_3096;
wire n_6306;
wire n_3496;
wire n_4114;
wire n_2544;
wire n_6434;
wire n_2356;
wire n_6751;
wire n_7068;
wire n_4556;
wire n_6322;
wire n_5454;
wire n_2620;
wire n_6667;
wire n_6530;
wire n_4089;
wire n_7376;
wire n_6156;
wire n_5913;
wire n_7268;
wire n_7044;
wire n_5621;
wire n_2919;
wire n_4327;
wire n_4218;
wire n_6429;
wire n_2150;
wire n_3146;
wire n_5165;
wire n_2241;
wire n_7239;
wire n_2757;
wire n_5573;
wire n_6405;
wire n_6613;
wire n_4353;
wire n_2042;
wire n_6248;
wire n_1754;
wire n_2921;
wire n_2720;
wire n_1854;
wire n_4990;
wire n_6088;
wire n_5529;
wire n_6894;
wire n_1856;
wire n_7267;
wire n_4959;
wire n_4161;
wire n_5800;
wire n_3992;
wire n_2616;
wire n_1906;
wire n_4103;
wire n_4466;
wire n_2262;
wire n_6204;
wire n_2462;
wire n_3625;
wire n_7387;
wire n_7431;
wire n_2798;
wire n_2945;
wire n_2331;
wire n_2837;
wire n_4844;
wire n_6296;
wire n_2979;
wire n_5257;
wire n_6290;
wire n_6288;
wire n_3655;
wire n_4688;
wire n_4765;
wire n_2548;
wire n_5645;
wire n_5180;
wire n_2108;
wire n_3640;
wire n_5779;
wire n_4388;
wire n_4206;
wire n_6140;
wire n_1779;
wire n_7441;
wire n_4738;
wire n_6211;
wire n_3909;
wire n_6307;
wire n_6164;
wire n_3207;
wire n_3944;
wire n_7394;
wire n_4434;
wire n_4837;
wire n_7022;
wire n_3042;
wire n_1942;
wire n_6860;
wire n_2510;
wire n_4219;
wire n_3659;
wire n_2804;
wire n_2120;
wire n_5012;
wire n_1876;
wire n_4620;
wire n_5697;
wire n_7188;
wire n_1810;
wire n_2813;
wire n_4438;
wire n_2009;
wire n_7087;
wire n_2222;
wire n_3510;
wire n_6147;
wire n_3218;
wire n_2667;
wire n_6515;
wire n_6011;
wire n_6645;
wire n_3150;
wire n_6984;
wire n_4325;
wire n_2413;
wire n_7193;
wire n_3775;
wire n_4133;
wire n_6897;
wire n_7256;
wire n_4184;
wire n_5203;
wire n_2518;
wire n_2629;
wire n_4481;
wire n_3416;
wire n_6460;
wire n_4379;
wire n_7128;
wire n_2181;
wire n_1829;
wire n_6183;
wire n_5882;
wire n_4030;
wire n_7436;
wire n_4490;
wire n_3138;
wire n_7380;
wire n_7012;
wire n_4397;
wire n_2928;
wire n_7335;
wire n_7103;
wire n_4820;
wire n_6246;
wire n_3770;
wire n_5094;
wire n_6383;
wire n_4938;
wire n_7020;
wire n_4179;
wire n_3469;
wire n_5336;
wire n_2723;
wire n_5672;
wire n_3220;
wire n_4641;
wire n_2539;
wire n_5548;
wire n_5601;
wire n_7248;
wire n_3855;
wire n_2054;
wire n_5339;
wire n_4931;
wire n_1765;
wire n_6099;
wire n_3158;
wire n_5693;
wire n_1744;
wire n_2623;
wire n_3113;
wire n_6904;
wire n_2718;
wire n_3760;
wire n_4078;
wire n_1760;
wire n_2856;
wire n_1832;
wire n_4146;
wire n_4360;
wire n_3666;
wire n_3828;
wire n_3288;
wire n_5514;
wire n_4404;
wire n_5091;
wire n_1874;
wire n_4787;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_3667;
wire n_6626;
wire n_6563;
wire n_5486;
wire n_6611;
wire n_3703;
wire n_4903;
wire n_3558;
wire n_2545;
wire n_2787;
wire n_5599;
wire n_6116;
wire n_7186;
wire n_4356;
wire n_6819;
wire n_2061;
wire n_4432;
wire n_5251;
wire n_2378;
wire n_1740;
wire n_6473;
wire n_4291;
wire n_5403;
wire n_4386;
wire n_4149;
wire n_6310;
wire n_2982;
wire n_2481;
wire n_7429;
wire n_3545;
wire n_6688;
wire n_2507;
wire n_4019;
wire n_2900;
wire n_2339;
wire n_7148;
wire n_5782;
wire n_6714;
wire n_4637;
wire n_7017;
wire n_7250;
wire n_7462;
wire n_4935;
wire n_6365;
wire n_4785;
wire n_3426;
wire n_3454;
wire n_3820;
wire n_5608;
wire n_3741;
wire n_3410;
wire n_7401;
wire n_6828;
wire n_2029;
wire n_5298;
wire n_6355;
wire n_5596;
wire n_1887;
wire n_4413;
wire n_6777;
wire n_5728;
wire n_2346;
wire n_3990;
wire n_4493;
wire n_3475;
wire n_6420;
wire n_6945;
wire n_2882;
wire n_7356;
wire n_2338;
wire n_5726;
wire n_7288;
wire n_7124;
wire n_3672;
wire n_7294;
wire n_5290;
wire n_3197;
wire n_7018;
wire n_3109;
wire n_2721;
wire n_7321;
wire n_5095;
wire n_3002;
wire n_6754;
wire n_6583;
wire n_6622;
wire n_6936;
wire n_5324;
wire n_3897;
wire n_5928;
wire n_3845;
wire n_7108;
wire n_6882;
wire n_2081;
wire n_4570;
wire n_7386;
wire n_2156;
wire n_5101;
wire n_4296;
wire n_1820;
wire n_5019;
wire n_5911;
wire n_7362;
wire n_7417;
wire n_2418;
wire n_7187;
wire n_5589;
wire n_5841;
wire n_2179;
wire n_2521;
wire n_3458;
wire n_5712;
wire n_3330;
wire n_4606;
wire n_6166;
wire n_4774;
wire n_2477;
wire n_6966;
wire n_3887;
wire n_6781;
wire n_7255;
wire n_4093;
wire n_7120;
wire n_7218;
wire n_4672;
wire n_7147;
wire n_3519;
wire n_7221;
wire n_4174;
wire n_3374;
wire n_3045;
wire n_2367;
wire n_1870;
wire n_4766;
wire n_5633;
wire n_2896;
wire n_4074;
wire n_4600;
wire n_6980;
wire n_1927;
wire n_5583;
wire n_4460;
wire n_3645;
wire n_3223;
wire n_3929;
wire n_6110;
wire n_6064;
wire n_6237;
wire n_7196;
wire n_2255;
wire n_2272;
wire n_6341;
wire n_1965;
wire n_1902;
wire n_6590;
wire n_1941;
wire n_5501;
wire n_3938;
wire n_5377;
wire n_2878;
wire n_6697;
wire n_5652;
wire n_6453;
wire n_6135;
wire n_3498;
wire n_2015;
wire n_1982;
wire n_4110;
wire n_7081;
wire n_3189;
wire n_2066;
wire n_6449;
wire n_3154;
wire n_6141;
wire n_2905;
wire n_3965;
wire n_3566;
wire n_2220;
wire n_4349;
wire n_3788;
wire n_4313;
wire n_2410;
wire n_6983;
wire n_1935;
wire n_6036;
wire n_3366;
wire n_2696;
wire n_4863;
wire n_7222;
wire n_3242;
wire n_6071;
wire n_3525;
wire n_3486;
wire n_6808;
wire n_2405;
wire n_6724;
wire n_3995;
wire n_2953;
wire n_2088;
wire n_4036;
wire n_6571;
wire n_5100;
wire n_7470;
wire n_1795;
wire n_5849;
wire n_6251;
wire n_7400;
wire n_2578;
wire n_3483;
wire n_6635;
wire n_1821;
wire n_3894;
wire n_3478;
wire n_4015;
wire n_3890;
wire n_2740;
wire n_5367;
wire n_2656;
wire n_3524;
wire n_5616;
wire n_5034;
wire n_6733;
wire n_7071;
wire n_5988;
wire n_6467;
wire n_6035;
wire n_3549;
wire n_6522;
wire n_7109;
wire n_2092;
wire n_5959;
wire n_2075;
wire n_3658;
wire n_6732;
wire n_1776;
wire n_4807;
wire n_6562;
wire n_6150;
wire n_2281;
wire n_2131;
wire n_3026;
wire n_1757;
wire n_1919;
wire n_4230;
wire n_3419;
wire n_2053;
wire n_1958;
wire n_5917;
wire n_5754;
wire n_6016;
wire n_3784;
wire n_2969;
wire n_3941;
wire n_2864;
wire n_3195;
wire n_3190;
wire n_7212;
wire n_3678;
wire n_2664;
wire n_3456;
wire n_5628;
wire n_1808;
wire n_6726;
wire n_2266;
wire n_2650;
wire n_4428;
wire n_5003;
wire n_5252;
wire n_7009;
wire n_6554;
wire n_6689;
wire n_2731;
wire n_6143;
wire n_5614;
wire n_5134;
wire n_3953;
wire n_3166;
wire n_4122;
wire n_3976;
wire n_7355;
wire n_3979;
wire n_7365;
wire n_4582;
wire n_2998;
wire n_6277;
wire n_4684;
wire n_7395;
wire n_5981;
wire n_6095;
wire n_6247;
wire n_4840;
wire n_3162;
wire n_2760;
wire n_6880;
wire n_3377;
wire n_3749;
wire n_5720;
wire n_3962;
wire n_1826;
wire n_2304;
wire n_5325;
wire n_5696;
wire n_2637;
wire n_5375;
wire n_4384;
wire n_6499;
wire n_6837;
wire n_4423;
wire n_4096;
wire n_7393;
wire n_2881;
wire n_6616;
wire n_3282;
wire n_1763;
wire n_3231;
wire n_1966;
wire n_6946;
wire n_4996;
wire n_2475;
wire n_4598;
wire n_5064;
wire n_5759;
wire n_4478;
wire n_5753;
wire n_2646;
wire n_5536;
wire n_7484;
wire n_5173;
wire n_6305;
wire n_6317;
wire n_3920;
wire n_4890;
wire n_5691;
wire n_5794;
wire n_5027;
wire n_5647;
wire n_7231;
wire n_3203;
wire n_3866;
wire n_2903;
wire n_3921;
wire n_7272;
wire n_4106;
wire n_3717;
wire n_5738;
wire n_2743;
wire n_2675;
wire n_3052;
wire n_5215;
wire n_7324;
wire n_6693;
wire n_3743;
wire n_6734;
wire n_7135;
wire n_7014;
wire n_1932;
wire n_4721;
wire n_5597;
wire n_5635;
wire n_6382;
wire n_7328;
wire n_1983;
wire n_6404;
wire n_5975;
wire n_4029;
wire n_3870;
wire n_6379;
wire n_7066;
wire n_4496;
wire n_3529;
wire n_7358;
wire n_1977;
wire n_2153;
wire n_6235;
wire n_4338;
wire n_7277;
wire n_6504;
wire n_3094;
wire n_2310;
wire n_3952;
wire n_7265;
wire n_2287;
wire n_2860;
wire n_2056;
wire n_6789;
wire n_7184;
wire n_6440;
wire n_6417;
wire n_2318;
wire n_2502;
wire n_2504;
wire n_4495;
wire n_4762;
wire n_7491;
wire n_5942;
wire n_2974;
wire n_2901;
wire n_1940;
wire n_2793;
wire n_3442;
wire n_7219;
wire n_7479;
wire n_3998;
wire n_2285;
wire n_3147;
wire n_4141;
wire n_7270;
wire n_5940;
wire n_7390;
wire n_5121;
wire n_1824;
wire n_3386;
wire n_1917;
wire n_4107;
wire n_4667;
wire n_2325;
wire n_5555;
wire n_6914;
wire n_2446;
wire n_3488;
wire n_7182;
wire n_4547;
wire n_2893;
wire n_2588;
wire n_2962;
wire n_4004;
wire n_5784;
wire n_6272;
wire n_6484;
wire n_6236;
wire n_5576;
wire n_4668;
wire n_4953;
wire n_5466;
wire n_6958;
wire n_6840;
wire n_3898;
wire n_6871;
wire n_1786;
wire n_5284;
wire n_4997;
wire n_5308;
wire n_4274;
wire n_2627;
wire n_6768;
wire n_4759;
wire n_4467;
wire n_2377;
wire n_2080;
wire n_2340;
wire n_3552;
wire n_6717;
wire n_3684;
wire n_4735;
wire n_3137;
wire n_7048;
wire n_5578;
wire n_2361;
wire n_4113;
wire n_1998;
wire n_4686;
wire n_5530;
wire n_3759;
wire n_6196;
wire n_7416;
wire n_4321;
wire n_4342;
wire n_2034;
wire n_5741;
wire n_5991;
wire n_3933;
wire n_7330;
wire n_3206;
wire n_5506;
wire n_3966;
wire n_5243;
wire n_5449;
wire n_5221;
wire n_6992;
wire n_4183;
wire n_4068;
wire n_4872;
wire n_6000;
wire n_4233;
wire n_7283;
wire n_3192;
wire n_7099;
wire n_3764;
wire n_4709;
wire n_5038;
wire n_5311;
wire n_6448;
wire n_2649;
wire n_6655;
wire n_7304;
wire n_5792;
wire n_6657;
wire n_1929;
wire n_5575;
wire n_2807;
wire n_2542;
wire n_2313;
wire n_3324;
wire n_3914;
wire n_4625;
wire n_2558;
wire n_2063;
wire n_3803;
wire n_3742;
wire n_7474;
wire n_2252;
wire n_6113;
wire n_4819;
wire n_6242;
wire n_7088;
wire n_6519;
wire n_2576;
wire n_4900;
wire n_6842;
wire n_3390;
wire n_6206;
wire n_6414;
wire n_3746;
wire n_2373;
wire n_3817;
wire n_2745;
wire n_6801;
wire n_2493;
wire n_4930;
wire n_5276;
wire n_6308;
wire n_7398;
wire n_6906;
wire n_5078;
wire n_4537;
wire n_7230;
wire n_2885;
wire n_6629;
wire n_5011;
wire n_3318;
wire n_4070;
wire n_6968;
wire n_4282;
wire n_6615;
wire n_3485;
wire n_4180;
wire n_7378;
wire n_3839;
wire n_5205;
wire n_3333;
wire n_5651;
wire n_2845;
wire n_6144;
wire n_4143;
wire n_4659;
wire n_6188;
wire n_2602;
wire n_5819;
wire n_4579;
wire n_4616;
wire n_3014;
wire n_2547;
wire n_5998;
wire n_6398;
wire n_5023;
wire n_1812;
wire n_4105;
wire n_5721;
wire n_5673;
wire n_2532;
wire n_3791;
wire n_2665;
wire n_5351;
wire n_3905;
wire n_3368;
wire n_3530;
wire n_1930;
wire n_1955;
wire n_3329;
wire n_2765;
wire n_6415;
wire n_2994;
wire n_6857;
wire n_2401;
wire n_3135;
wire n_5476;
wire n_2003;
wire n_5856;
wire n_5446;
wire n_4895;
wire n_6722;
wire n_3573;
wire n_3148;
wire n_6428;
wire n_5944;
wire n_2264;
wire n_3534;
wire n_6413;
wire n_4275;
wire n_3970;
wire n_6361;
wire n_3438;
wire n_6231;
wire n_4098;
wire n_5684;
wire n_5861;
wire n_5976;
wire n_4789;
wire n_1972;
wire n_2806;
wire n_5312;
wire n_2184;
wire n_5850;
wire n_3217;
wire n_3425;
wire n_3404;
wire n_5111;
wire n_5890;
wire n_4055;
wire n_2926;
wire n_3540;
wire n_3670;
wire n_3973;
wire n_7167;
wire n_2023;
wire n_3249;
wire n_2351;
wire n_5113;
wire n_4442;
wire n_4698;
wire n_6712;
wire n_5687;
wire n_4779;
wire n_2286;
wire n_4966;
wire n_2065;
wire n_4017;
wire n_5839;
wire n_3397;
wire n_3740;
wire n_6953;
wire n_4418;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_2977;
wire n_6303;
wire n_6474;
wire n_6182;
wire n_3723;
wire n_5674;
wire n_3600;
wire n_6573;
wire n_4134;
wire n_6053;
wire n_7234;
wire n_2836;
wire n_5682;
wire n_6392;
wire n_2130;
wire n_5167;
wire n_3239;
wire n_5117;
wire n_2773;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_4913;
wire n_5612;
wire n_6125;
wire n_6599;
wire n_6685;
wire n_1791;
wire n_2850;
wire n_1747;
wire n_4251;
wire n_1817;
wire n_3982;
wire n_2654;
wire n_4621;
wire n_6560;
wire n_3176;
wire n_4559;
wire n_2186;
wire n_4368;
wire n_6253;
wire n_4740;
wire n_7382;
wire n_5301;
wire n_5007;
wire n_3581;
wire n_2562;
wire n_4077;
wire n_4642;
wire n_5898;
wire n_2221;
wire n_3576;
wire n_7298;
wire n_1792;
wire n_1868;
wire n_4049;
wire n_6641;
wire n_3862;
wire n_5214;
wire n_5563;
wire n_5487;
wire n_6593;
wire n_3495;
wire n_3879;
wire n_2348;
wire n_6673;
wire n_7172;
wire n_7074;
wire n_5497;
wire n_4724;
wire n_5832;
wire n_7190;
wire n_7112;
wire n_1772;
wire n_5526;
wire n_2818;
wire n_3646;
wire n_6367;
wire n_2129;
wire n_3345;
wire n_4546;
wire n_6195;
wire n_3584;
wire n_6356;
wire n_3756;
wire n_2889;
wire n_7001;
wire n_5593;
wire n_5021;
wire n_6514;
wire n_2772;
wire n_7369;
wire n_5444;
wire n_1924;
wire n_4382;
wire n_3999;
wire n_2844;
wire n_2138;
wire n_5211;
wire n_5230;
wire n_6559;
wire n_7359;
wire n_2260;
wire n_5389;
wire n_1813;
wire n_7144;
wire n_4833;
wire n_6841;
wire n_3056;
wire n_2345;
wire n_5110;
wire n_6653;
wire n_3295;
wire n_2382;
wire n_4719;
wire n_4178;
wire n_3062;
wire n_2317;
wire n_7450;
wire n_5425;
wire n_3289;
wire n_1973;
wire n_5737;
wire n_2579;
wire n_6825;
wire n_6923;
wire n_1770;
wire n_4228;
wire n_4401;
wire n_1756;
wire n_6112;
wire n_2788;
wire n_6547;
wire n_2984;
wire n_6198;
wire n_7439;
wire n_3364;
wire n_5560;
wire n_6399;
wire n_1873;
wire n_3201;
wire n_6275;
wire n_5666;
wire n_6575;
wire n_3472;
wire n_6151;
wire n_2874;
wire n_5179;
wire n_7227;
wire n_7040;
wire n_4605;
wire n_4877;
wire n_3235;
wire n_7325;
wire n_4968;
wire n_6469;
wire n_6756;
wire n_5030;
wire n_3949;
wire n_5961;
wire n_3543;
wire n_7191;
wire n_7459;
wire n_7096;
wire n_3050;
wire n_3903;
wire n_4834;
wire n_5272;
wire n_2183;
wire n_3314;
wire n_4158;
wire n_2742;
wire n_6826;
wire n_2360;
wire n_6015;
wire n_3254;
wire n_5361;
wire n_5683;
wire n_4171;
wire n_5847;
wire n_4045;
wire n_6678;
wire n_4562;
wire n_5068;
wire n_3634;
wire n_5740;
wire n_2834;
wire n_2531;
wire n_5015;
wire n_2702;
wire n_5729;
wire n_7485;
wire n_6748;
wire n_2030;
wire n_3115;
wire n_4749;
wire n_4390;
wire n_5302;
wire n_4979;
wire n_1794;
wire n_6752;
wire n_2234;
wire n_4804;
wire n_5545;
wire n_6553;
wire n_2209;
wire n_6500;
wire n_4270;
wire n_2797;
wire n_7051;
wire n_5152;
wire n_2321;
wire n_3680;
wire n_6628;
wire n_6297;
wire n_5905;
wire n_3497;
wire n_6975;
wire n_5409;
wire n_6329;
wire n_2940;
wire n_5688;
wire n_2612;
wire n_5128;
wire n_4566;
wire n_2841;
wire n_6293;
wire n_3322;
wire n_4576;
wire n_2427;
wire n_2505;
wire n_4061;
wire n_3250;
wire n_2070;
wire n_6905;
wire n_7425;
wire n_2594;
wire n_5798;
wire n_6381;
wire n_6521;
wire n_1914;
wire n_2335;
wire n_2904;
wire n_5307;
wire n_4767;
wire n_4328;
wire n_3004;
wire n_5986;
wire n_3112;
wire n_2349;
wire n_6581;
wire n_3874;
wire n_6215;
wire n_7095;
wire n_5415;
wire n_4676;
wire n_5770;
wire n_7064;
wire n_5892;
wire n_4544;
wire n_2170;
wire n_6577;
wire n_6899;
wire n_5676;
wire n_7307;
wire n_6545;
wire n_5802;
wire n_3175;
wire n_3522;
wire n_4429;
wire n_4591;
wire n_6370;
wire n_3266;
wire n_7210;
wire n_4646;
wire n_5769;
wire n_6065;
wire n_7039;
wire n_6987;
wire n_4725;
wire n_4563;
wire n_2210;
wire n_4169;
wire n_5331;
wire n_6190;
wire n_6859;
wire n_3247;
wire n_3091;
wire n_3066;
wire n_6309;
wire n_6623;
wire n_2426;
wire n_6527;
wire n_7443;
wire n_5341;
wire n_4320;
wire n_5930;
wire n_5814;
wire n_4881;
wire n_5979;
wire n_5271;
wire n_5089;
wire n_7015;
wire n_5263;
wire n_3613;
wire n_3444;
wire n_6929;
wire n_4012;
wire n_5518;
wire n_4636;
wire n_5637;
wire n_4584;
wire n_5622;
wire n_3910;
wire n_4711;
wire n_3319;
wire n_7348;
wire n_5240;
wire n_3335;
wire n_5813;
wire n_3413;
wire n_5495;
wire n_1969;
wire n_4680;
wire n_2044;
wire n_5546;
wire n_2689;
wire n_3259;
wire n_7143;
wire n_5482;
wire n_7312;
wire n_4191;
wire n_5224;
wire n_4293;
wire n_2010;
wire n_7155;
wire n_3688;
wire n_6865;
wire n_3016;
wire n_5393;
wire n_2599;
wire n_6535;
wire n_7213;
wire n_3338;
wire n_3414;
wire n_1827;
wire n_4671;
wire n_4209;
wire n_5966;
wire n_7456;
wire n_5041;
wire n_7420;
wire n_1751;
wire n_5431;
wire n_3261;
wire n_2200;
wire n_6482;
wire n_5026;
wire n_3863;
wire n_3027;
wire n_2746;
wire n_5059;
wire n_5505;
wire n_3127;
wire n_1780;
wire n_3732;
wire n_6605;
wire n_4250;
wire n_5329;
wire n_3596;
wire n_4699;
wire n_7007;
wire n_3906;
wire n_4127;
wire n_3297;
wire n_2683;
wire n_2388;
wire n_4292;
wire n_3641;
wire n_4577;
wire n_4854;
wire n_6018;
wire n_5908;
wire n_4202;
wire n_7168;
wire n_5212;
wire n_5000;
wire n_2853;
wire n_5939;
wire n_7177;
wire n_3766;
wire n_2880;
wire n_7379;
wire n_3350;
wire n_2389;
wire n_4165;
wire n_4866;
wire n_7444;
wire n_5931;
wire n_7435;
wire n_4038;
wire n_4109;
wire n_5297;
wire n_7030;
wire n_5420;
wire n_6311;
wire n_4412;
wire n_3407;
wire n_3599;
wire n_6424;
wire n_6654;
wire n_6816;
wire n_6220;
wire n_3621;
wire n_5234;
wire n_6740;
wire n_7122;
wire n_5835;
wire n_7049;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_6029;
wire n_6879;
wire n_2538;
wire n_2105;
wire n_5259;
wire n_3163;
wire n_5440;
wire n_5679;
wire n_3710;
wire n_5938;
wire n_6702;
wire n_4155;
wire n_2031;
wire n_3891;
wire n_5891;
wire n_4144;
wire n_5724;
wire n_5774;
wire n_2165;
wire n_6452;
wire n_3379;
wire n_4374;
wire n_6791;
wire n_3532;
wire n_5131;
wire n_7280;
wire n_1818;
wire n_2127;
wire n_6915;
wire n_7110;
wire n_6856;
wire n_3531;
wire n_2963;
wire n_3834;
wire n_7232;
wire n_4548;
wire n_7345;
wire n_5923;
wire n_5790;
wire n_3258;
wire n_4989;
wire n_4622;
wire n_4315;
wire n_2959;
wire n_2047;
wire n_6364;
wire n_6451;
wire n_6552;
wire n_1845;
wire n_2193;
wire n_2478;
wire n_5140;
wire n_6328;
wire n_4816;
wire n_6363;
wire n_2983;
wire n_7159;
wire n_3810;
wire n_2715;
wire n_6132;
wire n_6578;
wire n_6406;
wire n_5598;
wire n_2085;
wire n_5306;
wire n_6978;
wire n_4483;
wire n_5342;
wire n_2782;
wire n_2672;
wire n_2651;
wire n_4358;
wire n_7477;
wire n_5147;
wire n_3656;
wire n_6918;
wire n_2071;
wire n_2561;
wire n_2643;
wire n_4793;
wire n_7363;
wire n_6612;
wire n_5677;
wire n_4168;
wire n_3446;
wire n_5997;
wire n_5511;
wire n_5680;
wire n_3028;
wire n_4806;
wire n_4350;
wire n_7295;
wire n_5533;
wire n_5838;
wire n_6058;
wire n_5280;
wire n_6375;
wire n_6479;
wire n_6866;
wire n_5235;
wire n_3836;
wire n_3963;
wire n_1872;
wire n_3389;
wire n_6170;
wire n_1931;
wire n_4187;
wire n_4166;
wire n_6447;
wire n_6263;
wire n_7093;
wire n_5206;
wire n_3222;
wire n_7466;
wire n_1801;
wire n_5419;
wire n_6130;
wire n_2970;
wire n_2235;
wire n_4937;
wire n_3980;
wire n_2791;
wire n_5103;
wire n_3755;
wire n_5803;
wire n_4258;
wire n_6014;
wire n_4498;
wire n_6935;
wire n_2174;
wire n_2714;
wire n_5285;
wire n_3563;
wire n_2506;
wire n_4064;
wire n_4936;
wire n_5387;
wire n_1863;
wire n_3841;
wire n_2118;
wire n_4770;
wire n_5985;
wire n_2944;
wire n_2407;
wire n_4907;
wire n_5058;
wire n_6907;
wire n_6158;
wire n_6541;
wire n_3262;
wire n_6119;
wire n_5018;
wire n_4006;
wire n_5896;
wire n_4861;
wire n_3690;
wire n_2358;
wire n_5192;
wire n_5141;
wire n_3716;
wire n_5133;
wire n_2833;
wire n_4712;
wire n_6226;
wire n_3191;
wire n_3837;
wire n_3193;
wire n_1971;
wire n_3252;
wire n_7145;
wire n_2275;
wire n_2855;
wire n_3273;
wire n_3544;
wire n_4310;
wire n_6338;
wire n_1950;
wire n_2370;
wire n_5159;
wire n_3954;
wire n_3025;
wire n_4674;
wire n_4908;
wire n_7467;
wire n_5097;
wire n_2750;
wire n_5730;
wire n_3899;
wire n_4159;
wire n_3714;
wire n_3071;
wire n_3739;
wire n_5816;
wire n_4069;
wire n_2784;
wire n_3718;
wire n_3092;
wire n_3470;
wire n_4862;
wire n_7241;
wire n_2557;
wire n_5300;
wire n_4850;
wire n_6625;
wire n_3781;
wire n_4912;
wire n_4813;
wire n_7464;
wire n_2590;
wire n_6302;
wire n_2330;
wire n_5748;
wire n_2942;
wire n_6759;
wire n_5525;
wire n_3106;
wire n_1882;
wire n_3328;
wire n_6706;
wire n_3889;
wire n_6139;
wire n_4256;
wire n_7434;
wire n_6999;
wire n_7054;
wire n_4224;
wire n_6403;
wire n_3508;
wire n_6483;
wire n_4024;
wire n_2267;
wire n_2218;
wire n_6228;
wire n_5650;
wire n_2636;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_5400;
wire n_2759;
wire n_4415;
wire n_5552;
wire n_7299;
wire n_4702;
wire n_6888;
wire n_4252;
wire n_4457;
wire n_6063;
wire n_6800;
wire n_5139;
wire n_2319;
wire n_6922;
wire n_3481;
wire n_5481;
wire n_6890;
wire n_2808;
wire n_6070;
wire n_2676;
wire n_2679;
wire n_6651;
wire n_5821;
wire n_7091;
wire n_4491;
wire n_7273;
wire n_6647;
wire n_7296;
wire n_2930;
wire n_5733;
wire n_1838;
wire n_3514;
wire n_2777;
wire n_2434;
wire n_4132;
wire n_2660;
wire n_5871;
wire n_2611;
wire n_4261;
wire n_6184;
wire n_4886;
wire n_4090;
wire n_2529;
wire n_2698;
wire n_5043;
wire n_5707;
wire n_4001;
wire n_3047;
wire n_2454;
wire n_4371;
wire n_5836;
wire n_5281;
wire n_6716;
wire n_6422;
wire n_4473;
wire n_3120;
wire n_4007;
wire n_1743;
wire n_4268;
wire n_5048;
wire n_5521;
wire n_5028;
wire n_4480;
wire n_2350;
wire n_3895;
wire n_7475;
wire n_4194;
wire n_5585;
wire n_6397;
wire n_4824;
wire n_1892;
wire n_4120;
wire n_4427;
wire n_3745;
wire n_2990;
wire n_1766;
wire n_7033;
wire n_6121;
wire n_3119;
wire n_4142;
wire n_4082;
wire n_5561;
wire n_3479;
wire n_4085;
wire n_4073;
wire n_4260;
wire n_4163;
wire n_4439;
wire n_2064;
wire n_6981;
wire n_3867;
wire n_4372;
wire n_3500;
wire n_6954;
wire n_3279;
wire n_2621;
wire n_5799;
wire n_5073;
wire n_5024;
wire n_5875;
wire n_4262;
wire n_2671;
wire n_6646;
wire n_1798;
wire n_1790;
wire n_4720;
wire n_7131;
wire n_6903;
wire n_4685;
wire n_6101;
wire n_5968;
wire n_2563;
wire n_2387;
wire n_4334;
wire n_6941;
wire n_1830;
wire n_2073;
wire n_4511;
wire n_5812;
wire n_6148;
wire n_5515;
wire n_6106;
wire n_6604;
wire n_4014;
wire n_7418;
wire n_5250;
wire n_3144;
wire n_4757;
wire n_2913;
wire n_2336;
wire n_5607;
wire n_4175;
wire n_2005;
wire n_1916;
wire n_4648;
wire n_5006;
wire n_6566;
wire n_5734;
wire n_6081;
wire n_4892;
wire n_7204;
wire n_3823;
wire n_1866;
wire n_4173;
wire n_4970;
wire n_3816;
wire n_5404;
wire n_4108;
wire n_4486;
wire n_6047;
wire n_2960;
wire n_5438;
wire n_4627;
wire n_7354;
wire n_7448;
wire n_6244;
wire n_2290;
wire n_6861;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_2040;
wire n_3199;
wire n_3843;
wire n_2145;
wire n_5725;
wire n_3030;
wire n_2580;
wire n_3685;
wire n_4249;
wire n_5163;
wire n_2039;
wire n_5768;
wire n_4961;
wire n_3753;
wire n_2035;
wire n_4718;
wire n_3555;
wire n_3579;
wire n_5190;
wire n_7422;
wire n_2509;
wire n_3236;
wire n_4317;
wire n_4855;
wire n_3969;
wire n_2459;
wire n_4154;
wire n_6588;
wire n_3396;
wire n_7050;
wire n_4023;
wire n_4420;
wire n_5685;
wire n_1923;
wire n_5773;
wire n_7136;
wire n_7318;
wire n_6055;
wire n_5138;
wire n_5374;
wire n_6108;
wire n_2116;
wire n_6165;
wire n_1828;
wire n_6621;
wire n_2320;
wire n_7175;
wire n_5349;
wire n_2038;
wire n_2137;
wire n_4973;
wire n_4640;
wire n_2583;
wire n_6323;
wire n_4396;
wire n_5127;
wire n_6587;
wire n_4367;
wire n_6480;
wire n_2087;
wire n_6731;
wire n_5485;
wire n_5766;
wire n_5216;
wire n_6597;
wire n_1989;
wire n_3818;
wire n_2523;
wire n_6933;
wire n_4387;
wire n_4951;
wire n_4453;
wire n_4170;
wire n_6881;
wire n_7289;
wire n_5805;
wire n_3719;
wire n_1959;
wire n_3681;
wire n_2737;
wire n_2399;
wire n_4308;
wire n_2812;
wire n_2355;
wire n_2133;
wire n_6216;
wire n_3830;
wire n_2585;
wire n_6817;
wire n_7170;
wire n_7314;
wire n_2725;
wire n_6949;
wire n_6509;
wire n_5175;
wire n_3883;
wire n_7260;
wire n_4152;
wire n_2565;
wire n_7263;
wire n_5948;
wire n_4392;
wire n_4660;
wire n_3149;
wire n_5611;
wire n_6911;
wire n_3268;
wire n_4281;
wire n_4661;
wire n_4200;
wire n_3614;
wire n_2111;
wire n_3301;
wire n_5900;
wire n_3466;
wire n_4962;
wire n_6327;
wire n_2595;
wire n_6607;
wire n_3411;
wire n_4958;
wire n_4271;
wire n_7209;
wire n_5171;
wire n_3586;
wire n_6401;
wire n_5554;
wire n_6227;
wire n_7240;
wire n_4071;
wire n_4921;
wire n_1980;
wire n_5427;
wire n_5639;
wire n_3065;
wire n_4361;
wire n_5417;
wire n_4614;
wire n_2681;
wire n_3103;
wire n_4945;
wire n_2424;
wire n_4922;
wire n_4732;
wire n_7278;
wire n_2775;
wire n_6416;
wire n_4693;
wire n_5488;
wire n_4326;
wire n_6695;
wire n_3557;
wire n_2230;
wire n_5447;
wire n_5383;
wire n_4744;
wire n_6127;
wire n_2851;
wire n_4305;
wire n_5781;
wire n_6600;
wire n_2490;
wire n_7410;
wire n_4213;
wire n_2849;
wire n_7097;
wire n_3692;
wire n_2204;
wire n_6421;
wire n_5747;
wire n_7414;
wire n_7495;
wire n_5969;
wire n_4929;
wire n_1961;
wire n_4964;
wire n_6079;
wire n_4802;
wire n_6192;
wire n_6458;
wire n_4139;
wire n_3029;
wire n_6746;
wire n_2508;
wire n_4031;
wire n_6719;
wire n_2416;
wire n_5437;
wire n_5826;
wire n_3881;
wire n_2461;
wire n_6506;
wire n_2243;
wire n_4583;
wire n_6287;
wire n_6662;
wire n_4210;
wire n_5245;
wire n_7189;
wire n_4666;
wire n_2929;
wire n_3751;
wire n_2555;
wire n_2662;
wire n_2368;
wire n_6851;
wire n_6687;
wire n_2890;
wire n_6884;
wire n_2554;
wire n_3698;
wire n_3927;
wire n_1840;
wire n_4540;
wire n_3961;
wire n_6780;
wire n_6513;
wire n_4891;
wire n_6619;
wire n_5603;
wire n_6804;
wire n_3559;
wire n_2661;
wire n_2572;
wire n_5716;
wire n_3993;
wire n_4940;
wire n_6516;
wire n_5208;
wire n_7490;
wire n_3588;
wire n_6924;
wire n_2308;
wire n_4590;
wire n_7492;
wire n_5606;
wire n_4830;
wire n_5231;
wire n_5237;
wire n_4664;
wire n_3860;
wire n_5456;
wire n_3160;
wire n_7073;
wire n_2191;
wire n_5093;
wire n_2428;
wire n_6040;
wire n_3847;
wire n_4946;
wire n_4906;
wire n_5727;
wire n_2158;
wire n_3290;
wire n_4663;
wire n_5390;
wire n_7114;
wire n_5347;
wire n_2824;
wire n_3033;
wire n_3298;
wire n_6788;
wire n_2440;
wire n_4883;
wire n_2923;
wire n_4162;
wire n_3665;
wire n_5115;
wire n_3264;
wire n_6393;
wire n_2333;
wire n_2916;
wire n_6249;
wire n_4297;
wire n_5833;
wire n_6849;
wire n_3800;
wire n_2403;
wire n_5407;
wire n_4608;
wire n_5232;
wire n_2792;
wire n_2870;
wire n_7271;
wire n_3991;
wire n_3134;
wire n_6572;
wire n_4172;
wire n_4791;
wire n_6739;
wire n_4536;
wire n_5149;
wire n_5967;
wire n_2463;
wire n_5151;
wire n_7003;
wire n_4773;
wire n_5345;
wire n_5357;
wire n_4497;
wire n_6666;
wire n_2472;
wire n_4611;
wire n_6812;
wire n_4755;
wire n_5982;
wire n_1768;
wire n_2294;
wire n_4960;
wire n_2993;
wire n_3864;
wire n_4658;
wire n_5135;
wire n_2732;
wire n_2948;
wire n_2309;
wire n_7419;
wire n_5827;
wire n_5494;
wire n_4362;
wire n_4306;
wire n_6200;
wire n_2123;
wire n_3209;
wire n_3504;
wire n_2037;
wire n_2685;
wire n_1953;
wire n_4422;
wire n_6123;
wire n_6934;
wire n_2589;
wire n_7094;
wire n_3482;
wire n_6082;
wire n_2233;
wire n_4555;
wire n_2827;
wire n_5136;
wire n_5228;
wire n_7129;
wire n_3956;
wire n_5758;
wire n_5323;
wire n_3572;
wire n_4215;
wire n_6952;
wire n_4280;
wire n_7062;
wire n_3375;
wire n_4047;
wire n_5471;
wire n_5434;
wire n_2082;
wire n_5941;
wire n_7045;
wire n_5879;
wire n_3167;
wire n_5558;
wire n_5350;
wire n_3423;
wire n_2362;
wire n_2609;
wire n_5338;
wire n_7238;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_7126;
wire n_5669;
wire n_3854;
wire n_2468;
wire n_3078;
wire n_6979;
wire n_6203;
wire n_7405;
wire n_3253;
wire n_7207;
wire n_4027;
wire n_2280;
wire n_7454;
wire n_4599;
wire n_5830;
wire n_6796;
wire n_3363;
wire n_4812;
wire n_5760;
wire n_6368;
wire n_3689;
wire n_6556;
wire n_2020;
wire n_4628;
wire n_5668;
wire n_1881;
wire n_2749;
wire n_3451;
wire n_4873;
wire n_5878;
wire n_5588;
wire n_4657;
wire n_2971;
wire n_2311;
wire n_5765;
wire n_3950;
wire n_4458;
wire n_6596;
wire n_4121;
wire n_5090;
wire n_6870;
wire n_4476;
wire n_5613;
wire n_2298;
wire n_4756;
wire n_3869;
wire n_4307;
wire n_5104;
wire n_5042;
wire n_4860;
wire n_4359;
wire n_7251;
wire n_2303;
wire n_2810;
wire n_2747;
wire n_6080;
wire n_7059;
wire n_7035;
wire n_1848;
wire n_5571;
wire n_2126;
wire n_4573;
wire n_5289;
wire n_4118;
wire n_6713;
wire n_5513;
wire n_6747;
wire n_6281;
wire n_4803;
wire n_5972;
wire n_4079;
wire n_4091;
wire n_5916;
wire n_5984;
wire n_7029;
wire n_7317;
wire n_2002;
wire n_5145;
wire n_3712;
wire n_2371;
wire n_6094;
wire n_2935;
wire n_6444;
wire n_5132;
wire n_5191;
wire n_6333;
wire n_6262;
wire n_3085;
wire n_5869;
wire n_5925;
wire n_6240;
wire n_5359;
wire n_6412;
wire n_2574;
wire n_5293;
wire n_7220;
wire n_4316;
wire n_3697;
wire n_7438;
wire n_2638;
wire n_4044;
wire n_4062;
wire n_6684;
wire n_4524;
wire n_4843;
wire n_3971;
wire n_7065;
wire n_5510;
wire n_6046;
wire n_2016;
wire n_6973;
wire n_2949;
wire n_2711;
wire n_5363;
wire n_7285;
wire n_5200;
wire n_5659;
wire n_5618;
wire n_6325;
wire n_2867;
wire n_1894;
wire n_2794;
wire n_3145;
wire n_3124;
wire n_6737;
wire n_6454;
wire n_4253;
wire n_5356;
wire n_6721;
wire n_5369;
wire n_2608;
wire n_5258;
wire n_2657;
wire n_5255;
wire n_2852;
wire n_2392;
wire n_7008;
wire n_3517;
wire n_3100;
wire n_2522;
wire n_6111;
wire n_1834;
wire n_3758;
wire n_3356;
wire n_2835;
wire n_6260;
wire n_1968;
wire n_3269;
wire n_5080;
wire n_6665;
wire n_7055;
wire n_3506;
wire n_3605;
wire n_2409;
wire n_5858;
wire n_5817;
wire n_6690;
wire n_3402;
wire n_5723;
wire n_5295;
wire n_6137;
wire n_4679;
wire n_4115;
wire n_6201;
wire n_7113;
wire n_4998;
wire n_2988;
wire n_1970;
wire n_2766;
wire n_5627;
wire n_2201;
wire n_2117;
wire n_4167;
wire n_7242;
wire n_1993;
wire n_5155;
wire n_3835;
wire n_6461;
wire n_2205;
wire n_1777;
wire n_1957;
wire n_3967;
wire n_5016;
wire n_1912;
wire n_6212;
wire n_3401;
wire n_6908;
wire n_3226;
wire n_6570;
wire n_6498;
wire n_3902;
wire n_4730;
wire n_7228;
wire n_6692;
wire n_6074;
wire n_2779;
wire n_6380;
wire n_3654;
wire n_2164;
wire n_5996;
wire n_2115;
wire n_2232;
wire n_5327;
wire n_6045;
wire n_1774;
wire n_4713;
wire n_5137;
wire n_6505;
wire n_2811;
wire n_3348;
wire n_7415;
wire n_5796;
wire n_6320;
wire n_6489;
wire n_6068;
wire n_3358;
wire n_5791;
wire n_2121;
wire n_1803;
wire n_4204;
wire n_5098;
wire n_6877;
wire n_2224;
wire n_1991;
wire n_6772;
wire n_6823;
wire n_6806;
wire n_7426;
wire n_5906;
wire n_4743;
wire n_3805;
wire n_3825;
wire n_6831;
wire n_3657;
wire n_4924;
wire n_3928;
wire n_4859;
wire n_7217;
wire n_2692;
wire n_2008;
wire n_6284;
wire n_7058;
wire n_4654;
wire n_6157;
wire n_5423;
wire n_7497;
wire n_6785;
wire n_6374;
wire n_6930;
wire n_4733;
wire n_3792;
wire n_6017;
wire n_4272;
wire n_3974;
wire n_3871;
wire n_1753;
wire n_2283;
wire n_3278;
wire n_4269;
wire n_4695;
wire n_1855;
wire n_6838;
wire n_5736;
wire n_6937;
wire n_6443;
wire n_3312;
wire n_6105;
wire n_2197;
wire n_2199;
wire n_5069;
wire n_7442;
wire n_5700;
wire n_6543;
wire n_3285;
wire n_3968;
wire n_5099;
wire n_2228;
wire n_4704;
wire n_4551;
wire n_5052;
wire n_6091;
wire n_2421;
wire n_2902;
wire n_4957;
wire n_6674;
wire n_2480;
wire n_6034;
wire n_2363;
wire n_4072;
wire n_5579;
wire n_7085;
wire n_4781;
wire n_3606;
wire n_6652;
wire n_7098;
wire n_5004;
wire n_2550;
wire n_6762;
wire n_7341;
wire n_4424;
wire n_7391;
wire n_3055;
wire n_3711;
wire n_3315;
wire n_5837;
wire n_3172;
wire n_3292;
wire n_4436;
wire n_6895;
wire n_3878;
wire n_4450;
wire n_5642;
wire n_3553;
wire n_7224;
wire n_5880;
wire n_6169;
wire n_4746;
wire n_5713;
wire n_6005;
wire n_3131;
wire n_5118;
wire n_5105;
wire n_3850;
wire n_4459;
wire n_2996;
wire n_5793;
wire n_5591;
wire n_4050;
wire n_7496;
wire n_2315;
wire n_3228;
wire n_2102;
wire n_5623;
wire n_5681;
wire n_4853;
wire n_7399;
wire n_2422;
wire n_6213;
wire n_2239;
wire n_6118;
wire n_5256;
wire n_2950;
wire n_5220;
wire n_5732;
wire n_3852;
wire n_5178;
wire n_4520;
wire n_6814;
wire n_7342;
wire n_2057;
wire n_4008;
wire n_5507;
wire n_7214;
wire n_7472;
wire n_5077;
wire n_5872;
wire n_3858;
wire n_7408;
wire n_1901;
wire n_6115;
wire n_4502;
wire n_6858;
wire n_3032;
wire n_4851;
wire n_5735;
wire n_7254;
wire n_6944;
wire n_7384;
wire n_3072;
wire n_3081;
wire n_3313;
wire n_2710;
wire n_1745;
wire n_3924;
wire n_4571;
wire n_2006;
wire n_6430;
wire n_6193;
wire n_5314;
wire n_6462;
wire n_2343;
wire n_3439;
wire n_5049;
wire n_6757;
wire n_6822;
wire n_2535;
wire n_4205;
wire n_5953;
wire n_2726;
wire n_5277;
wire n_4723;
wire n_5176;
wire n_6779;
wire n_6518;
wire n_6797;
wire n_2799;
wire n_4454;
wire n_4229;
wire n_5952;
wire n_4739;
wire n_5820;
wire n_2376;
wire n_5483;
wire n_3017;
wire n_5718;
wire n_6916;
wire n_2456;
wire n_3904;
wire n_5150;
wire n_2678;
wire n_4838;
wire n_2872;
wire n_2451;
wire n_5075;
wire n_4879;
wire n_5051;
wire n_3926;
wire n_6152;
wire n_1962;
wire n_3996;
wire n_4221;
wire n_2854;
wire n_4181;
wire n_5777;
wire n_2764;
wire n_7046;
wire n_4225;
wire n_2567;
wire n_5142;
wire n_3102;
wire n_4153;
wire n_5156;
wire n_5926;
wire n_3627;
wire n_4300;
wire n_3551;
wire n_1769;
wire n_4783;
wire n_2964;
wire n_3769;
wire n_6589;
wire n_2673;
wire n_4530;
wire n_4267;
wire n_2292;
wire n_3865;
wire n_3859;
wire n_3722;
wire n_7173;
wire n_5951;
wire n_7092;
wire n_2442;
wire n_6197;
wire n_6971;
wire n_1943;
wire n_7460;
wire n_3117;
wire n_3428;
wire n_2961;
wire n_3351;
wire n_3527;
wire n_6154;
wire n_7344;
wire n_6020;
wire n_2883;
wire n_1752;
wire n_4182;
wire n_2912;
wire n_4825;
wire n_5701;
wire n_4440;
wire n_4549;
wire n_1910;
wire n_3955;
wire n_7079;
wire n_5120;
wire n_5470;
wire n_4565;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_4303;
wire n_4574;
wire n_5797;
wire n_6696;
wire n_4839;
wire n_5222;
wire n_5743;
wire n_4016;
wire n_6210;
wire n_5772;
wire n_3435;
wire n_3575;
wire n_6964;
wire n_5801;
wire n_6117;
wire n_4231;
wire n_6202;
wire n_7279;
wire n_3165;
wire n_4923;
wire n_3652;
wire n_4097;
wire n_6681;
wire n_4083;
wire n_1937;
wire n_5971;
wire n_4461;
wire n_3234;
wire n_5392;
wire n_2381;
wire n_6661;
wire n_3303;
wire n_6640;
wire n_3916;
wire n_2569;
wire n_3556;
wire n_7371;
wire n_6962;
wire n_4101;
wire n_6455;
wire n_2196;
wire n_3591;
wire n_4273;
wire n_3024;
wire n_5443;
wire n_3512;
wire n_5600;
wire n_4939;
wire n_5169;
wire n_6963;
wire n_6644;
wire n_4389;
wire n_6896;
wire n_3930;
wire n_4448;
wire n_6832;
wire n_2161;
wire n_6160;
wire n_2404;
wire n_2083;
wire n_6718;
wire n_2503;
wire n_6542;
wire n_1936;
wire n_6031;
wire n_5502;
wire n_2027;
wire n_5568;
wire n_2642;
wire n_2500;
wire n_1918;
wire n_5656;
wire n_6763;
wire n_4831;
wire n_2513;
wire n_5974;
wire n_3480;
wire n_2695;
wire n_3057;
wire n_3194;
wire n_6280;
wire n_2414;
wire n_6438;
wire n_3662;
wire n_6316;
wire n_7383;
wire n_4319;
wire n_5474;
wire n_2229;
wire n_5413;
wire n_4596;
wire n_6758;
wire n_2004;
wire n_5412;
wire n_3694;
wire n_2586;
wire n_6069;
wire n_5752;
wire n_6874;
wire n_4726;
wire n_1879;
wire n_4751;
wire n_4222;
wire n_2274;
wire n_2972;
wire n_3225;
wire n_6030;
wire n_6077;
wire n_4119;
wire n_3799;
wire n_4298;
wire n_5201;
wire n_6299;
wire n_4474;
wire n_6386;
wire n_5217;
wire n_5957;
wire n_2511;
wire n_3383;
wire n_3585;
wire n_2975;
wire n_5490;
wire n_5029;
wire n_2704;
wire n_4214;
wire n_5158;
wire n_4884;
wire n_6708;
wire n_7433;
wire n_4366;
wire n_4009;
wire n_7347;
wire n_4580;
wire n_6792;
wire n_6177;
wire n_5912;
wire n_4129;
wire n_4871;
wire n_2617;
wire n_4999;
wire n_6033;
wire n_1859;
wire n_5557;
wire n_7397;
wire n_7389;
wire n_5472;
wire n_2955;
wire n_4112;
wire n_6002;
wire n_4337;
wire n_5711;
wire n_4138;
wire n_5396;
wire n_5335;
wire n_2520;
wire n_6557;
wire n_7300;
wire n_2134;
wire n_5960;
wire n_4236;
wire n_2185;
wire n_3270;
wire n_2143;
wire n_5002;
wire n_3595;
wire n_5143;
wire n_4238;
wire n_6142;
wire n_6917;
wire n_2374;
wire n_5859;
wire n_1947;
wire n_2114;
wire n_3571;
wire n_2396;
wire n_1799;
wire n_4734;
wire n_1939;
wire n_2486;
wire n_6163;
wire n_4635;
wire n_3501;
wire n_7118;
wire n_1869;
wire n_4013;
wire n_3039;
wire n_2011;
wire n_6285;
wire n_6778;
wire n_6025;
wire n_7257;
wire n_4242;
wire n_6862;
wire n_6319;
wire n_7067;
wire n_4984;
wire n_3851;
wire n_2543;
wire n_3036;
wire n_1896;
wire n_3180;
wire n_5283;
wire n_5268;
wire n_6318;
wire n_4561;
wire n_2639;
wire n_6089;
wire n_3325;
wire n_3107;
wire n_4021;
wire n_3880;
wire n_5122;
wire n_6315;
wire n_3186;
wire n_4955;
wire n_5556;
wire n_5462;
wire n_4501;
wire n_3696;
wire n_3650;
wire n_5840;
wire n_2761;
wire n_6343;
wire n_3157;
wire n_2537;
wire n_2144;
wire n_6049;
wire n_6919;
wire n_7423;
wire n_2515;
wire n_2466;
wire n_2652;
wire n_6052;
wire n_2635;
wire n_5330;
wire n_4197;
wire n_4829;
wire n_7069;
wire n_6886;
wire n_1949;
wire n_2936;
wire n_1946;
wire n_6912;
wire n_5914;
wire n_4715;
wire n_5039;
wire n_2141;
wire n_6061;
wire n_4369;
wire n_5378;
wire n_4543;
wire n_2099;
wire n_4941;
wire n_7252;
wire n_5542;
wire n_1831;
wire n_4394;
wire n_7133;
wire n_1850;
wire n_6883;
wire n_5519;
wire n_1749;
wire n_3101;
wire n_3669;
wire n_6009;
wire n_7061;
wire n_5278;
wire n_2663;
wire n_5586;
wire n_2693;
wire n_3798;
wire n_4065;
wire n_6378;
wire n_5187;
wire n_4944;
wire n_5675;
wire n_2180;
wire n_2249;
wire n_4135;
wire n_2632;
wire n_6601;
wire n_5771;
wire n_7216;
wire n_6407;
wire n_1755;
wire n_6749;
wire n_6839;
wire n_2908;
wire n_3744;
wire n_4263;
wire n_1862;
wire n_2915;
wire n_2300;
wire n_3291;
wire n_6051;
wire n_4716;
wire n_4942;
wire n_6217;
wire n_6680;
wire n_5844;
wire n_2432;
wire n_6532;
wire n_3405;
wire n_4745;
wire n_6155;
wire n_6446;
wire n_6738;
wire n_6250;
wire n_7458;
wire n_2337;
wire n_3907;
wire n_6736;
wire n_5344;
wire n_6526;
wire n_4629;
wire n_6339;
wire n_2932;
wire n_2980;
wire n_5225;
wire n_6350;
wire n_7013;
wire n_3306;
wire n_1784;
wire n_5662;
wire n_4857;
wire n_3136;
wire n_4080;
wire n_4226;
wire n_4741;
wire n_2101;
wire n_1986;
wire n_4752;
wire n_5265;
wire n_1750;
wire n_3986;
wire n_4376;
wire n_5705;
wire n_4753;
wire n_4552;
wire n_3885;
wire n_6845;
wire n_7105;
wire n_2713;
wire n_5196;
wire n_5181;
wire n_2644;
wire n_2951;
wire n_3008;
wire n_3709;
wire n_6829;
wire n_5574;
wire n_5126;
wire n_6508;
wire n_2214;
wire n_2055;
wire n_3427;
wire n_4067;
wire n_5553;
wire n_4176;
wire n_4042;
wire n_4385;
wire n_3320;
wire n_7052;
wire n_5009;
wire n_7262;
wire n_2688;
wire n_5368;
wire n_5626;
wire n_6603;
wire n_6114;
wire n_6576;
wire n_3651;
wire n_4333;
wire n_7364;
wire n_3359;
wire n_7208;
wire n_6245;
wire n_2865;
wire n_2706;
wire n_5499;
wire n_6703;
wire n_3676;
wire n_4375;
wire n_4788;
wire n_4717;
wire n_4986;
wire n_5604;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_4815;
wire n_7202;
wire n_4246;
wire n_3580;
wire n_7011;
wire n_2139;
wire n_4609;
wire n_5291;
wire n_5876;
wire n_6970;
wire n_5114;
wire n_2674;
wire n_6409;
wire n_6704;
wire n_4088;
wire n_6876;
wire n_3682;
wire n_4357;
wire n_3371;
wire n_1809;
wire n_7028;
wire n_4462;
wire n_4472;
wire n_3433;
wire n_7320;
wire n_6255;
wire n_7313;
wire n_7343;
wire n_5288;
wire n_2305;
wire n_5540;
wire n_5699;
wire n_2450;
wire n_3447;
wire n_5810;
wire n_3305;
wire n_4148;
wire n_4151;
wire n_3528;
wire n_6938;
wire n_4373;
wire n_5762;
wire n_4934;
wire n_5218;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_7337;
wire n_6989;
wire n_4630;
wire n_5408;
wire n_4643;
wire n_4331;
wire n_6427;
wire n_3989;
wire n_4475;
wire n_4846;
wire n_3804;
wire n_4344;
wire n_1775;
wire n_3296;
wire n_2762;
wire n_7038;
wire n_4683;
wire n_5366;
wire n_1847;
wire n_2767;
wire n_6360;
wire n_2603;
wire n_3116;
wire n_1884;
wire n_3602;
wire n_2967;
wire n_6146;
wire n_6270;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_2195;
wire n_5477;
wire n_5451;
wire n_3923;
wire n_4696;
wire n_2626;
wire n_3441;
wire n_1978;
wire n_5086;
wire n_2801;
wire n_5901;
wire n_6353;
wire n_4011;
wire n_4905;
wire n_2763;
wire n_2825;
wire n_3643;
wire n_4876;
wire n_6345;
wire n_1997;
wire n_6691;
wire n_3748;
wire n_3142;
wire n_4278;
wire n_4623;
wire n_4910;
wire n_2690;
wire n_4410;
wire n_3370;
wire n_7392;
wire n_2215;
wire n_5053;
wire n_6239;
wire n_4553;
wire n_6803;
wire n_3978;
wire n_6340;
wire n_4809;
wire n_5226;
wire n_1925;
wire n_3660;
wire n_1815;
wire n_5867;
wire n_6048;
wire n_1788;
wire n_2491;
wire n_5079;
wire n_5590;
wire n_6773;
wire n_3833;
wire n_5632;
wire n_4841;
wire n_2022;
wire n_6336;
wire n_3814;
wire n_7041;
wire n_2592;
wire n_2838;
wire n_4842;
wire n_4911;
wire n_4340;
wire n_7370;
wire n_3513;
wire n_3133;
wire n_5660;
wire n_4645;
wire n_2992;
wire n_6174;
wire n_3725;
wire n_1833;
wire n_4920;
wire n_4972;
wire n_6023;
wire n_2517;
wire n_6776;
wire n_3128;
wire n_5426;
wire n_6463;
wire n_2631;
wire n_2178;
wire n_1767;
wire n_6372;
wire n_7176;
wire n_2469;
wire n_5625;
wire n_5778;
wire n_6396;
wire n_3355;
wire n_2007;
wire n_3917;
wire n_6669;
wire n_3942;
wire n_2736;
wire n_3765;
wire n_5531;
wire n_3000;
wire n_5429;
wire n_3108;
wire n_3111;
wire n_1837;
wire n_1839;
wire n_5818;
wire n_5646;
wire n_6940;
wire n_4557;
wire n_5248;
wire n_4451;
wire n_6394;
wire n_2875;
wire n_3844;
wire n_3280;
wire n_4054;
wire n_5448;
wire n_3471;
wire n_5432;
wire n_3205;
wire n_2046;
wire n_2848;
wire n_5160;
wire n_2741;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_6995;
wire n_7185;
wire n_3564;
wire n_3988;
wire n_6254;
wire n_6161;
wire n_3457;
wire n_4324;
wire n_4821;
wire n_1871;
wire n_5445;
wire n_3630;
wire n_3271;
wire n_7332;
wire n_6660;
wire n_4771;
wire n_5719;
wire n_7225;
wire n_6128;
wire n_4086;
wire n_2412;
wire n_7037;
wire n_4814;
wire n_1781;
wire n_2084;
wire n_3648;
wire n_5749;
wire n_3075;
wire n_3173;
wire n_5332;
wire n_5108;
wire n_7409;
wire n_4692;
wire n_3031;
wire n_7258;
wire n_7432;
wire n_3701;
wire n_1773;
wire n_3243;
wire n_6334;
wire n_3385;
wire n_2666;
wire n_6848;
wire n_2171;
wire n_4708;
wire n_6321;
wire n_2768;
wire n_2314;
wire n_6794;
wire n_4826;
wire n_3343;
wire n_2420;
wire n_7197;
wire n_5489;
wire n_6400;
wire n_3767;
wire n_2873;
wire n_2299;
wire n_2540;
wire n_4589;
wire n_5057;
wire n_4578;
wire n_6705;
wire n_2162;
wire n_2847;
wire n_2051;
wire n_3221;
wire n_5436;
wire n_5907;
wire n_2168;
wire n_2790;
wire n_5072;
wire n_3629;
wire n_3021;
wire n_6044;
wire n_2359;
wire n_3674;
wire n_5286;
wire n_3502;
wire n_3098;
wire n_6495;
wire n_5013;
wire n_2312;
wire n_7403;
wire n_6902;
wire n_6470;
wire n_3015;
wire n_1920;
wire n_5569;
wire n_5439;
wire n_5619;
wire n_4147;
wire n_2048;
wire n_6481;
wire n_3607;
wire n_4925;
wire n_1921;
wire n_6534;
wire n_4974;
wire n_1800;
wire n_4932;
wire n_4510;
wire n_2571;
wire n_6181;
wire n_3276;
wire n_6728;
wire n_3787;
wire n_5119;
wire n_2124;
wire n_5715;
wire n_6133;
wire n_6528;
wire n_7407;
wire n_3827;
wire n_3354;
wire n_2519;
wire n_2724;
wire n_4447;
wire n_6670;
wire n_6774;
wire n_4285;
wire n_5887;
wire n_4651;
wire n_6741;
wire n_7424;
wire n_6038;
wire n_4818;
wire n_4514;
wire n_4800;
wire n_3960;
wire n_3248;
wire n_2277;
wire n_6282;
wire n_2110;
wire n_4433;
wire n_2879;
wire n_2474;
wire n_2090;
wire n_3153;
wire n_6700;
wire n_7334;
wire n_2033;
wire n_4341;
wire n_4312;
wire n_3399;
wire n_2628;
wire n_5932;
wire n_6178;
wire n_2132;
wire n_6234;
wire n_6012;
wire n_2400;
wire n_4633;
wire n_3838;
wire n_1909;
wire n_4277;
wire n_4140;
wire n_3675;
wire n_5092;
wire n_3387;
wire n_5186;
wire n_7367;
wire n_4662;
wire n_3779;
wire n_2464;
wire n_6715;
wire n_5828;
wire n_2831;
wire n_7200;
wire n_4882;
wire n_4993;
wire n_2365;
wire n_4832;
wire n_4207;
wire n_4545;
wire n_3037;
wire n_6337;
wire n_4868;
wire n_1885;
wire n_2452;
wire n_6770;
wire n_6743;
wire n_3925;
wire n_2176;
wire n_1816;
wire n_5238;
wire n_4059;
wire n_2455;
wire n_4595;
wire n_1849;
wire n_6682;
wire n_5054;
wire n_5631;
wire n_2467;
wire n_6539;
wire n_7243;
wire n_7179;
wire n_2288;
wire n_4063;
wire n_5399;
wire n_6314;
wire n_6617;
wire n_3592;
wire n_5694;
wire n_4650;
wire n_4888;
wire n_7274;
wire n_5326;
wire n_3394;
wire n_4874;
wire n_3793;
wire n_4669;
wire n_4339;
wire n_6595;
wire n_4041;
wire n_5459;
wire n_2858;
wire n_4060;
wire n_2658;
wire n_2895;
wire n_2128;
wire n_5528;
wire n_3097;
wire n_5391;
wire n_4541;
wire n_3824;
wire n_5422;
wire n_6385;
wire n_6289;
wire n_3388;
wire n_5267;
wire n_4494;
wire n_3059;
wire n_5523;
wire n_3465;
wire n_4796;
wire n_7373;
wire n_3589;
wire n_2534;
wire n_6186;
wire n_4799;
wire n_5153;
wire n_6257;
wire n_3449;
wire n_2694;
wire n_2198;
wire n_2610;
wire n_2989;
wire n_6852;
wire n_2789;
wire n_6346;
wire n_4775;
wire n_2216;
wire n_5044;
wire n_5809;
wire n_1897;
wire n_5365;
wire n_2933;
wire n_5045;
wire n_4381;
wire n_4266;
wire n_3886;
wire n_5354;
wire n_4455;
wire n_6274;
wire n_7372;
wire n_2328;
wire n_4248;
wire n_5915;
wire n_6818;
wire n_5452;
wire n_7226;
wire n_4754;
wire n_7057;
wire n_4554;
wire n_5595;
wire n_6609;
wire n_4845;
wire n_6815;
wire n_6753;
wire n_3053;
wire n_3893;
wire n_2465;
wire n_3548;
wire n_4585;
wire n_3334;
wire n_4383;
wire n_2541;
wire n_6764;
wire n_5535;
wire n_3875;
wire n_5370;
wire n_6391;
wire n_4003;
wire n_5372;
wire n_5299;
wire n_2402;
wire n_5594;
wire n_4301;
wire n_4586;
wire n_1954;
wire n_4048;
wire n_6471;
wire n_1844;
wire n_3777;
wire n_6627;
wire n_5761;
wire n_4784;
wire n_7203;
wire n_2999;
wire n_5550;
wire n_5082;
wire n_4046;
wire n_1974;
wire n_2086;
wire n_3537;
wire n_5209;
wire n_7215;
wire n_3080;
wire n_6636;
wire n_4199;
wire n_2701;
wire n_5929;
wire n_3362;
wire n_5559;
wire n_3105;
wire n_5478;
wire n_7388;
wire n_6243;
wire n_6488;
wire n_4286;
wire n_5102;
wire n_2556;
wire n_2269;
wire n_3274;
wire n_3041;
wire n_6022;
wire n_6457;
wire n_4470;
wire n_2236;
wire n_2816;
wire n_1911;
wire n_3616;
wire n_4058;
wire n_2460;
wire n_3664;
wire n_4188;
wire n_3913;
wire n_6867;
wire n_3417;
wire n_5868;
wire n_6230;
wire n_4034;
wire n_6538;
wire n_6633;
wire n_6187;
wire n_3327;
wire n_6172;
wire n_5275;
wire n_4689;
wire n_5071;
wire n_3067;
wire n_7311;
wire n_2755;
wire n_5989;
wire n_3237;
wire n_6574;
wire n_1992;
wire n_6395;
wire n_4402;
wire n_4239;
wire n_6854;
wire n_3400;
wire n_6233;
wire n_4550;
wire n_6456;
wire n_3382;
wire n_7488;
wire n_3574;
wire n_5227;
wire n_2169;
wire n_7198;
wire n_4201;
wire n_6784;
wire n_6168;
wire n_3316;
wire n_6766;
wire n_5242;
wire n_3099;
wire n_3704;
wire n_2596;
wire n_3603;
wire n_4123;
wire n_6330;
wire n_2192;
wire n_5520;
wire n_3633;
wire n_4479;
wire n_7249;
wire n_2670;
wire n_5947;
wire n_7336;
wire n_4416;
wire n_3372;
wire n_7031;
wire n_4539;
wire n_2707;
wire n_6799;
wire n_5920;
wire n_6672;
wire n_2471;
wire n_6149;
wire n_7142;
wire n_3230;
wire n_5808;
wire n_3342;
wire n_6054;
wire n_7089;
wire n_4682;
wire n_5353;
wire n_3708;
wire n_5294;
wire n_6450;
wire n_3729;
wire n_4978;
wire n_4690;
wire n_4437;
wire n_5458;
wire n_3861;
wire n_5617;
wire n_4736;
wire n_7042;
wire n_3780;
wire n_1928;
wire n_5244;
wire n_6523;
wire n_5382;
wire n_6107;
wire n_3957;
wire n_6775;
wire n_5274;
wire n_3848;
wire n_4284;
wire n_2600;
wire n_3919;
wire n_6232;
wire n_6445;
wire n_7181;
wire n_6134;
wire n_5384;
wire n_3608;
wire n_6056;
wire n_6932;
wire n_7036;
wire n_4513;
wire n_3233;
wire n_3829;
wire n_3177;
wire n_4053;
wire n_2352;
wire n_5125;
wire n_4040;
wire n_2207;
wire n_5587;
wire n_2619;
wire n_6855;
wire n_2444;
wire n_5789;
wire n_3123;
wire n_5787;
wire n_6585;
wire n_6369;
wire n_5056;
wire n_5249;
wire n_3393;
wire n_7447;
wire n_5198;
wire n_5360;
wire n_7455;
wire n_5233;
wire n_4887;
wire n_5829;
wire n_4617;
wire n_5269;
wire n_3520;
wire n_2492;
wire n_6252;
wire n_5866;
wire n_6493;
wire n_4005;
wire n_4904;
wire n_5899;
wire n_4792;
wire n_7104;
wire n_3578;
wire n_3812;
wire n_1886;
wire n_4980;
wire n_6026;
wire n_4290;
wire n_5247;
wire n_5865;
wire n_3727;
wire n_5317;
wire n_6544;
wire n_3774;
wire n_3093;
wire n_1843;
wire n_3061;
wire n_7138;
wire n_7290;
wire n_2431;
wire n_6679;
wire n_4956;
wire n_5380;
wire n_2206;
wire n_5924;
wire n_3182;
wire n_5822;
wire n_2564;
wire n_6259;
wire n_4947;
wire n_7284;
wire n_4656;
wire n_3896;
wire n_3958;
wire n_6390;
wire n_3450;
wire n_4729;
wire n_5786;
wire n_4987;
wire n_5182;
wire n_4971;
wire n_2000;
wire n_2074;
wire n_3174;
wire n_2217;
wire n_6630;
wire n_3398;
wire n_2307;
wire n_5658;
wire n_3408;
wire n_2722;
wire n_5388;
wire n_2640;
wire n_4823;
wire n_4875;
wire n_3432;
wire n_6279;
wire n_1771;
wire n_3090;
wire n_3762;
wire n_2437;
wire n_6813;
wire n_5564;
wire n_2445;
wire n_1835;
wire n_1988;
wire n_7106;
wire n_6042;
wire n_1853;
wire n_6057;
wire n_1787;
wire n_4137;
wire n_6675;
wire n_2634;
wire n_4529;
wire n_4323;
wire n_3034;
wire n_2212;
wire n_6476;
wire n_3972;
wire n_6207;
wire n_5539;
wire n_6268;
wire n_6878;
wire n_6286;
wire n_3308;
wire n_6524;
wire n_5036;
wire n_5547;
wire n_4772;
wire n_3467;
wire n_6225;
wire n_4322;
wire n_7297;
wire n_6291;
wire n_2830;
wire n_5893;
wire n_4354;
wire n_4653;
wire n_2354;
wire n_2246;
wire n_7199;
wire n_5273;
wire n_4677;
wire n_3901;
wire n_5261;
wire n_6520;
wire n_3757;
wire n_3381;
wire n_5193;
wire n_2245;
wire n_1782;
wire n_4909;
wire n_2965;
wire n_3635;
wire n_6024;
wire n_5022;
wire n_5005;
wire n_2814;
wire n_3882;
wire n_3046;
wire n_7487;
wire n_2213;
wire n_6425;
wire n_5993;
wire n_3826;
wire n_3211;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_5703;
wire n_4634;
wire n_3337;
wire n_2527;
wire n_6432;
wire n_5534;
wire n_3204;
wire n_7259;
wire n_2136;
wire n_6540;
wire n_6955;
wire n_5174;
wire n_1822;
wire n_4952;
wire n_5157;
wire n_3005;
wire n_4380;
wire n_3129;
wire n_4126;
wire n_7237;
wire n_1783;
wire n_2601;
wire n_5087;
wire n_3043;
wire n_3802;
wire n_2375;
wire n_4506;
wire n_6388;
wire n_5904;
wire n_4880;
wire n_6760;
wire n_1907;
wire n_2686;
wire n_2344;
wire n_3892;
wire n_4896;
wire n_5620;
wire n_5061;
wire n_5572;
wire n_5750;
wire n_7063;
wire n_1985;
wire n_2107;
wire n_3219;
wire n_2906;
wire n_4943;
wire n_2187;
wire n_1762;
wire n_3023;
wire n_6795;
wire n_5881;
wire n_6664;
wire n_5815;
wire n_6261;
wire n_4193;
wire n_5873;
wire n_4075;
wire n_3104;
wire n_6487;
wire n_4737;
wire n_6729;
wire n_3647;
wire n_5755;
wire n_2819;
wire n_5949;
wire n_5195;
wire n_7483;
wire n_3609;
wire n_4136;
wire n_6608;
wire n_1952;
wire n_4393;
wire n_7385;
wire n_3720;
wire n_4535;
wire n_1922;
wire n_2560;
wire n_4522;
wire n_6663;
wire n_4794;
wire n_5955;
wire n_7476;
wire n_3959;
wire n_7327;
wire n_5763;
wire n_6656;
wire n_6843;
wire n_3140;
wire n_5246;
wire n_5964;
wire n_3724;
wire n_2104;
wire n_3011;
wire n_7266;
wire n_5164;
wire n_4196;
wire n_6969;
wire n_4592;
wire n_4675;
wire n_5340;
wire n_5665;
wire n_6485;
wire n_3069;
wire n_5498;
wire n_7100;
wire n_4370;
wire n_1900;
wire n_5783;
wire n_5183;
wire n_6075;
wire n_7082;
wire n_3084;
wire n_6120;
wire n_6659;
wire n_2735;
wire n_6750;
wire n_3412;
wire n_2497;
wire n_1995;
wire n_5549;
wire n_2411;
wire n_3761;
wire n_4889;
wire n_7132;
wire n_2014;
wire n_2986;
wire n_5442;
wire n_5739;
wire n_3184;
wire n_4828;
wire n_6003;
wire n_5385;
wire n_4558;
wire n_6478;
wire n_2172;
wire n_6066;
wire n_7034;
wire n_6086;
wire n_4722;
wire n_6650;
wire n_6224;
wire n_3626;
wire n_4768;
wire n_4100;
wire n_2250;
wire n_7084;
wire n_5845;
wire n_7293;
wire n_4092;
wire n_5990;
wire n_3908;
wire n_6175;
wire n_6060;
wire n_7253;
wire n_2423;
wire n_3671;
wire n_6891;
wire n_5663;
wire n_6410;
wire n_3344;
wire n_2194;
wire n_4465;
wire n_5973;
wire n_3302;
wire n_5537;
wire n_5304;
wire n_2680;
wire n_6059;
wire n_5130;
wire n_3122;
wire n_5162;
wire n_4808;
wire n_3842;
wire n_6103;
wire n_6809;
wire n_3265;
wire n_1857;
wire n_4482;
wire n_2041;
wire n_6267;
wire n_1797;
wire n_2957;
wire n_5855;
wire n_2357;
wire n_5757;
wire n_6437;
wire n_3309;
wire n_7331;
wire n_6610;
wire n_3260;
wire n_4926;
wire n_3357;
wire n_4116;
wire n_6957;
wire n_5704;
wire n_7163;
wire n_2570;
wire n_1858;
wire n_2815;
wire n_5473;
wire n_3754;
wire n_4612;
wire n_5946;
wire n_2744;
wire n_6711;
wire n_4287;
wire n_2397;
wire n_7445;
wire n_2208;
wire n_6847;
wire n_3063;
wire n_5177;
wire n_3617;
wire n_7123;
wire n_6384;
wire n_4516;
wire n_3794;
wire n_2809;
wire n_2050;
wire n_4505;
wire n_6298;
wire n_2591;
wire n_3384;
wire n_7361;
wire n_4602;
wire n_5172;
wire n_4449;
wire n_1864;
wire n_7322;
wire n_5710;
wire n_7453;
wire n_6067;
wire n_5070;
wire n_6377;
wire n_4445;
wire n_5566;
wire n_5414;
wire n_4870;
wire n_2438;
wire n_2832;
wire n_1975;
wire n_2296;
wire n_3181;
wire n_6348;
wire n_2278;
wire n_4915;
wire n_5296;
wire n_6129;
wire n_2135;
wire n_5450;
wire n_3493;
wire n_6834;
wire n_5313;
wire n_3323;
wire n_2734;
wire n_4914;
wire n_6136;
wire n_7261;
wire n_6723;
wire n_5834;
wire n_2823;
wire n_1761;
wire n_5874;
wire n_7021;
wire n_5270;
wire n_5956;
wire n_4345;
wire n_5188;
wire n_3281;
wire n_6078;
wire n_3307;
wire n_7000;
wire n_4318;
wire n_2485;
wire n_2655;
wire n_4185;
wire n_4797;
wire n_2366;
wire n_7130;
wire n_5823;
wire n_3997;
wire n_5465;
wire n_4032;
wire n_1764;
wire n_3582;
wire n_5853;
wire n_2826;
wire n_3539;
wire n_7077;
wire n_4343;
wire n_4212;
wire n_6642;
wire n_4124;
wire n_5467;
wire n_5522;
wire n_4492;
wire n_7346;
wire n_2708;
wire n_5148;
wire n_4994;
wire n_7333;
wire n_4245;
wire n_4364;
wire n_4928;
wire n_2225;
wire n_4378;
wire n_2383;
wire n_1996;
wire n_3406;
wire n_3604;
wire n_3853;
wire n_4216;
wire n_5934;
wire n_6942;
wire n_2019;
wire n_2166;
wire n_2938;
wire n_4309;
wire n_3594;
wire n_6511;
wire n_3721;
wire n_6507;
wire n_2026;
wire n_2109;
wire n_2013;
wire n_1990;
wire n_2614;
wire n_7319;
wire n_2991;
wire n_6497;
wire n_6001;
wire n_6007;
wire n_2242;
wire n_2752;
wire n_2894;
wire n_6606;
wire n_3473;
wire n_4560;
wire n_5318;
wire n_2839;
wire n_5395;
wire n_2237;
wire n_7078;
wire n_3463;
wire n_7047;
wire n_3699;
wire n_5067;
wire n_7107;
wire n_3360;
wire n_2524;
wire n_3873;
wire n_3693;
wire n_7469;
wire n_2728;
wire n_3857;

CKINVDCx5p33_ASAP7_75t_R g1738 ( 
.A(n_1600),
.Y(n_1738)
);

INVx3_ASAP7_75t_L g1739 ( 
.A(n_170),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_1145),
.Y(n_1740)
);

BUFx2_ASAP7_75t_L g1741 ( 
.A(n_1562),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_1426),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_318),
.Y(n_1743)
);

BUFx3_ASAP7_75t_L g1744 ( 
.A(n_514),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1001),
.Y(n_1745)
);

CKINVDCx5p33_ASAP7_75t_R g1746 ( 
.A(n_1450),
.Y(n_1746)
);

CKINVDCx5p33_ASAP7_75t_R g1747 ( 
.A(n_803),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1497),
.Y(n_1748)
);

CKINVDCx20_ASAP7_75t_R g1749 ( 
.A(n_794),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_1436),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_1469),
.Y(n_1751)
);

INVx1_ASAP7_75t_SL g1752 ( 
.A(n_372),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_405),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_1506),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_392),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_1647),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_1574),
.Y(n_1757)
);

CKINVDCx5p33_ASAP7_75t_R g1758 ( 
.A(n_1116),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1572),
.Y(n_1759)
);

CKINVDCx5p33_ASAP7_75t_R g1760 ( 
.A(n_961),
.Y(n_1760)
);

CKINVDCx5p33_ASAP7_75t_R g1761 ( 
.A(n_791),
.Y(n_1761)
);

CKINVDCx5p33_ASAP7_75t_R g1762 ( 
.A(n_460),
.Y(n_1762)
);

BUFx3_ASAP7_75t_L g1763 ( 
.A(n_1554),
.Y(n_1763)
);

BUFx10_ASAP7_75t_L g1764 ( 
.A(n_715),
.Y(n_1764)
);

CKINVDCx5p33_ASAP7_75t_R g1765 ( 
.A(n_649),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_532),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_86),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_1381),
.Y(n_1768)
);

CKINVDCx5p33_ASAP7_75t_R g1769 ( 
.A(n_500),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_1283),
.Y(n_1770)
);

CKINVDCx5p33_ASAP7_75t_R g1771 ( 
.A(n_42),
.Y(n_1771)
);

CKINVDCx5p33_ASAP7_75t_R g1772 ( 
.A(n_158),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_1557),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_842),
.Y(n_1774)
);

CKINVDCx5p33_ASAP7_75t_R g1775 ( 
.A(n_90),
.Y(n_1775)
);

CKINVDCx5p33_ASAP7_75t_R g1776 ( 
.A(n_1665),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_1292),
.Y(n_1777)
);

HB1xp67_ASAP7_75t_L g1778 ( 
.A(n_1659),
.Y(n_1778)
);

INVx2_ASAP7_75t_SL g1779 ( 
.A(n_343),
.Y(n_1779)
);

CKINVDCx5p33_ASAP7_75t_R g1780 ( 
.A(n_381),
.Y(n_1780)
);

CKINVDCx5p33_ASAP7_75t_R g1781 ( 
.A(n_891),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_605),
.Y(n_1782)
);

BUFx10_ASAP7_75t_L g1783 ( 
.A(n_246),
.Y(n_1783)
);

CKINVDCx5p33_ASAP7_75t_R g1784 ( 
.A(n_1455),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_87),
.Y(n_1785)
);

CKINVDCx20_ASAP7_75t_R g1786 ( 
.A(n_448),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1700),
.Y(n_1787)
);

CKINVDCx5p33_ASAP7_75t_R g1788 ( 
.A(n_1648),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1222),
.Y(n_1789)
);

CKINVDCx5p33_ASAP7_75t_R g1790 ( 
.A(n_1720),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_873),
.Y(n_1791)
);

CKINVDCx5p33_ASAP7_75t_R g1792 ( 
.A(n_703),
.Y(n_1792)
);

CKINVDCx20_ASAP7_75t_R g1793 ( 
.A(n_1379),
.Y(n_1793)
);

CKINVDCx20_ASAP7_75t_R g1794 ( 
.A(n_371),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1703),
.Y(n_1795)
);

CKINVDCx20_ASAP7_75t_R g1796 ( 
.A(n_1244),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_543),
.Y(n_1797)
);

CKINVDCx5p33_ASAP7_75t_R g1798 ( 
.A(n_1656),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1074),
.Y(n_1799)
);

CKINVDCx5p33_ASAP7_75t_R g1800 ( 
.A(n_1673),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_194),
.Y(n_1801)
);

BUFx2_ASAP7_75t_L g1802 ( 
.A(n_111),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1570),
.Y(n_1803)
);

CKINVDCx5p33_ASAP7_75t_R g1804 ( 
.A(n_1490),
.Y(n_1804)
);

CKINVDCx5p33_ASAP7_75t_R g1805 ( 
.A(n_1584),
.Y(n_1805)
);

CKINVDCx5p33_ASAP7_75t_R g1806 ( 
.A(n_239),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1735),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_1579),
.Y(n_1808)
);

CKINVDCx16_ASAP7_75t_R g1809 ( 
.A(n_1251),
.Y(n_1809)
);

CKINVDCx5p33_ASAP7_75t_R g1810 ( 
.A(n_16),
.Y(n_1810)
);

CKINVDCx5p33_ASAP7_75t_R g1811 ( 
.A(n_1097),
.Y(n_1811)
);

INVx1_ASAP7_75t_SL g1812 ( 
.A(n_437),
.Y(n_1812)
);

CKINVDCx5p33_ASAP7_75t_R g1813 ( 
.A(n_1530),
.Y(n_1813)
);

CKINVDCx5p33_ASAP7_75t_R g1814 ( 
.A(n_218),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_210),
.Y(n_1815)
);

CKINVDCx5p33_ASAP7_75t_R g1816 ( 
.A(n_1391),
.Y(n_1816)
);

HB1xp67_ASAP7_75t_L g1817 ( 
.A(n_809),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1411),
.Y(n_1818)
);

CKINVDCx5p33_ASAP7_75t_R g1819 ( 
.A(n_1717),
.Y(n_1819)
);

CKINVDCx5p33_ASAP7_75t_R g1820 ( 
.A(n_808),
.Y(n_1820)
);

CKINVDCx5p33_ASAP7_75t_R g1821 ( 
.A(n_448),
.Y(n_1821)
);

BUFx10_ASAP7_75t_L g1822 ( 
.A(n_1553),
.Y(n_1822)
);

CKINVDCx5p33_ASAP7_75t_R g1823 ( 
.A(n_162),
.Y(n_1823)
);

CKINVDCx5p33_ASAP7_75t_R g1824 ( 
.A(n_1581),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1689),
.Y(n_1825)
);

CKINVDCx5p33_ASAP7_75t_R g1826 ( 
.A(n_829),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1598),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_685),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_1466),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1472),
.Y(n_1830)
);

CKINVDCx5p33_ASAP7_75t_R g1831 ( 
.A(n_838),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1370),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_790),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1662),
.Y(n_1834)
);

BUFx3_ASAP7_75t_L g1835 ( 
.A(n_229),
.Y(n_1835)
);

BUFx2_ASAP7_75t_L g1836 ( 
.A(n_12),
.Y(n_1836)
);

CKINVDCx5p33_ASAP7_75t_R g1837 ( 
.A(n_576),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_546),
.Y(n_1838)
);

CKINVDCx5p33_ASAP7_75t_R g1839 ( 
.A(n_1030),
.Y(n_1839)
);

CKINVDCx5p33_ASAP7_75t_R g1840 ( 
.A(n_1577),
.Y(n_1840)
);

CKINVDCx5p33_ASAP7_75t_R g1841 ( 
.A(n_1537),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_530),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1107),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_1633),
.Y(n_1844)
);

CKINVDCx5p33_ASAP7_75t_R g1845 ( 
.A(n_34),
.Y(n_1845)
);

CKINVDCx5p33_ASAP7_75t_R g1846 ( 
.A(n_1565),
.Y(n_1846)
);

CKINVDCx5p33_ASAP7_75t_R g1847 ( 
.A(n_506),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1523),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_172),
.Y(n_1849)
);

CKINVDCx5p33_ASAP7_75t_R g1850 ( 
.A(n_402),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1223),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1048),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_370),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_1649),
.Y(n_1854)
);

CKINVDCx20_ASAP7_75t_R g1855 ( 
.A(n_121),
.Y(n_1855)
);

CKINVDCx5p33_ASAP7_75t_R g1856 ( 
.A(n_162),
.Y(n_1856)
);

CKINVDCx5p33_ASAP7_75t_R g1857 ( 
.A(n_1507),
.Y(n_1857)
);

CKINVDCx5p33_ASAP7_75t_R g1858 ( 
.A(n_1620),
.Y(n_1858)
);

CKINVDCx20_ASAP7_75t_R g1859 ( 
.A(n_256),
.Y(n_1859)
);

CKINVDCx5p33_ASAP7_75t_R g1860 ( 
.A(n_1164),
.Y(n_1860)
);

CKINVDCx5p33_ASAP7_75t_R g1861 ( 
.A(n_135),
.Y(n_1861)
);

CKINVDCx5p33_ASAP7_75t_R g1862 ( 
.A(n_819),
.Y(n_1862)
);

CKINVDCx20_ASAP7_75t_R g1863 ( 
.A(n_1611),
.Y(n_1863)
);

CKINVDCx5p33_ASAP7_75t_R g1864 ( 
.A(n_1037),
.Y(n_1864)
);

CKINVDCx5p33_ASAP7_75t_R g1865 ( 
.A(n_1249),
.Y(n_1865)
);

CKINVDCx5p33_ASAP7_75t_R g1866 ( 
.A(n_1629),
.Y(n_1866)
);

CKINVDCx5p33_ASAP7_75t_R g1867 ( 
.A(n_1483),
.Y(n_1867)
);

CKINVDCx5p33_ASAP7_75t_R g1868 ( 
.A(n_403),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_546),
.Y(n_1869)
);

CKINVDCx5p33_ASAP7_75t_R g1870 ( 
.A(n_873),
.Y(n_1870)
);

INVxp67_ASAP7_75t_L g1871 ( 
.A(n_1417),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1177),
.Y(n_1872)
);

BUFx3_ASAP7_75t_L g1873 ( 
.A(n_635),
.Y(n_1873)
);

CKINVDCx5p33_ASAP7_75t_R g1874 ( 
.A(n_1008),
.Y(n_1874)
);

CKINVDCx5p33_ASAP7_75t_R g1875 ( 
.A(n_371),
.Y(n_1875)
);

CKINVDCx5p33_ASAP7_75t_R g1876 ( 
.A(n_1007),
.Y(n_1876)
);

CKINVDCx5p33_ASAP7_75t_R g1877 ( 
.A(n_217),
.Y(n_1877)
);

CKINVDCx5p33_ASAP7_75t_R g1878 ( 
.A(n_1135),
.Y(n_1878)
);

INVxp67_ASAP7_75t_L g1879 ( 
.A(n_367),
.Y(n_1879)
);

CKINVDCx16_ASAP7_75t_R g1880 ( 
.A(n_105),
.Y(n_1880)
);

CKINVDCx5p33_ASAP7_75t_R g1881 ( 
.A(n_706),
.Y(n_1881)
);

CKINVDCx20_ASAP7_75t_R g1882 ( 
.A(n_508),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1371),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_520),
.Y(n_1884)
);

CKINVDCx16_ASAP7_75t_R g1885 ( 
.A(n_729),
.Y(n_1885)
);

CKINVDCx5p33_ASAP7_75t_R g1886 ( 
.A(n_1697),
.Y(n_1886)
);

CKINVDCx5p33_ASAP7_75t_R g1887 ( 
.A(n_231),
.Y(n_1887)
);

CKINVDCx5p33_ASAP7_75t_R g1888 ( 
.A(n_233),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_796),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1526),
.Y(n_1890)
);

BUFx6f_ASAP7_75t_L g1891 ( 
.A(n_1605),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_874),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1726),
.Y(n_1893)
);

BUFx3_ASAP7_75t_L g1894 ( 
.A(n_1639),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1671),
.Y(n_1895)
);

CKINVDCx5p33_ASAP7_75t_R g1896 ( 
.A(n_1019),
.Y(n_1896)
);

CKINVDCx5p33_ASAP7_75t_R g1897 ( 
.A(n_1339),
.Y(n_1897)
);

CKINVDCx5p33_ASAP7_75t_R g1898 ( 
.A(n_1560),
.Y(n_1898)
);

CKINVDCx5p33_ASAP7_75t_R g1899 ( 
.A(n_940),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_375),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_740),
.Y(n_1901)
);

CKINVDCx14_ASAP7_75t_R g1902 ( 
.A(n_1638),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_645),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1501),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1488),
.Y(n_1905)
);

INVx1_ASAP7_75t_SL g1906 ( 
.A(n_780),
.Y(n_1906)
);

CKINVDCx5p33_ASAP7_75t_R g1907 ( 
.A(n_708),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_1695),
.Y(n_1908)
);

CKINVDCx5p33_ASAP7_75t_R g1909 ( 
.A(n_1270),
.Y(n_1909)
);

CKINVDCx5p33_ASAP7_75t_R g1910 ( 
.A(n_555),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_572),
.Y(n_1911)
);

CKINVDCx5p33_ASAP7_75t_R g1912 ( 
.A(n_86),
.Y(n_1912)
);

CKINVDCx5p33_ASAP7_75t_R g1913 ( 
.A(n_1080),
.Y(n_1913)
);

CKINVDCx5p33_ASAP7_75t_R g1914 ( 
.A(n_1593),
.Y(n_1914)
);

CKINVDCx5p33_ASAP7_75t_R g1915 ( 
.A(n_1109),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_390),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1034),
.Y(n_1917)
);

CKINVDCx5p33_ASAP7_75t_R g1918 ( 
.A(n_1372),
.Y(n_1918)
);

CKINVDCx5p33_ASAP7_75t_R g1919 ( 
.A(n_1457),
.Y(n_1919)
);

INVx1_ASAP7_75t_SL g1920 ( 
.A(n_1666),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_1595),
.Y(n_1921)
);

CKINVDCx5p33_ASAP7_75t_R g1922 ( 
.A(n_616),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1038),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1388),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_835),
.Y(n_1925)
);

CKINVDCx5p33_ASAP7_75t_R g1926 ( 
.A(n_859),
.Y(n_1926)
);

BUFx2_ASAP7_75t_L g1927 ( 
.A(n_1065),
.Y(n_1927)
);

CKINVDCx5p33_ASAP7_75t_R g1928 ( 
.A(n_42),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1694),
.Y(n_1929)
);

CKINVDCx5p33_ASAP7_75t_R g1930 ( 
.A(n_1190),
.Y(n_1930)
);

CKINVDCx5p33_ASAP7_75t_R g1931 ( 
.A(n_1650),
.Y(n_1931)
);

CKINVDCx5p33_ASAP7_75t_R g1932 ( 
.A(n_674),
.Y(n_1932)
);

CKINVDCx5p33_ASAP7_75t_R g1933 ( 
.A(n_362),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_231),
.Y(n_1934)
);

INVx1_ASAP7_75t_SL g1935 ( 
.A(n_230),
.Y(n_1935)
);

CKINVDCx5p33_ASAP7_75t_R g1936 ( 
.A(n_1737),
.Y(n_1936)
);

CKINVDCx5p33_ASAP7_75t_R g1937 ( 
.A(n_1631),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1563),
.Y(n_1938)
);

CKINVDCx5p33_ASAP7_75t_R g1939 ( 
.A(n_1051),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1576),
.Y(n_1940)
);

CKINVDCx5p33_ASAP7_75t_R g1941 ( 
.A(n_737),
.Y(n_1941)
);

CKINVDCx5p33_ASAP7_75t_R g1942 ( 
.A(n_838),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1622),
.Y(n_1943)
);

CKINVDCx16_ASAP7_75t_R g1944 ( 
.A(n_428),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1653),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1533),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1503),
.Y(n_1947)
);

CKINVDCx5p33_ASAP7_75t_R g1948 ( 
.A(n_1669),
.Y(n_1948)
);

CKINVDCx5p33_ASAP7_75t_R g1949 ( 
.A(n_1589),
.Y(n_1949)
);

CKINVDCx5p33_ASAP7_75t_R g1950 ( 
.A(n_940),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1696),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1102),
.Y(n_1952)
);

BUFx3_ASAP7_75t_L g1953 ( 
.A(n_1569),
.Y(n_1953)
);

CKINVDCx20_ASAP7_75t_R g1954 ( 
.A(n_274),
.Y(n_1954)
);

CKINVDCx5p33_ASAP7_75t_R g1955 ( 
.A(n_1733),
.Y(n_1955)
);

CKINVDCx5p33_ASAP7_75t_R g1956 ( 
.A(n_91),
.Y(n_1956)
);

CKINVDCx5p33_ASAP7_75t_R g1957 ( 
.A(n_1539),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_758),
.Y(n_1958)
);

CKINVDCx20_ASAP7_75t_R g1959 ( 
.A(n_762),
.Y(n_1959)
);

CKINVDCx5p33_ASAP7_75t_R g1960 ( 
.A(n_443),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1618),
.Y(n_1961)
);

CKINVDCx5p33_ASAP7_75t_R g1962 ( 
.A(n_1044),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1176),
.Y(n_1963)
);

CKINVDCx5p33_ASAP7_75t_R g1964 ( 
.A(n_1247),
.Y(n_1964)
);

CKINVDCx20_ASAP7_75t_R g1965 ( 
.A(n_1435),
.Y(n_1965)
);

CKINVDCx20_ASAP7_75t_R g1966 ( 
.A(n_1556),
.Y(n_1966)
);

CKINVDCx5p33_ASAP7_75t_R g1967 ( 
.A(n_325),
.Y(n_1967)
);

BUFx3_ASAP7_75t_L g1968 ( 
.A(n_1607),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_1558),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_749),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_14),
.Y(n_1971)
);

CKINVDCx5p33_ASAP7_75t_R g1972 ( 
.A(n_125),
.Y(n_1972)
);

INVx2_ASAP7_75t_SL g1973 ( 
.A(n_1006),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_549),
.Y(n_1974)
);

CKINVDCx5p33_ASAP7_75t_R g1975 ( 
.A(n_533),
.Y(n_1975)
);

CKINVDCx5p33_ASAP7_75t_R g1976 ( 
.A(n_1133),
.Y(n_1976)
);

CKINVDCx20_ASAP7_75t_R g1977 ( 
.A(n_1479),
.Y(n_1977)
);

CKINVDCx20_ASAP7_75t_R g1978 ( 
.A(n_770),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1131),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_65),
.Y(n_1980)
);

BUFx6f_ASAP7_75t_L g1981 ( 
.A(n_1621),
.Y(n_1981)
);

CKINVDCx5p33_ASAP7_75t_R g1982 ( 
.A(n_1015),
.Y(n_1982)
);

CKINVDCx20_ASAP7_75t_R g1983 ( 
.A(n_1664),
.Y(n_1983)
);

BUFx3_ASAP7_75t_L g1984 ( 
.A(n_153),
.Y(n_1984)
);

CKINVDCx5p33_ASAP7_75t_R g1985 ( 
.A(n_1016),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1730),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_692),
.Y(n_1987)
);

CKINVDCx5p33_ASAP7_75t_R g1988 ( 
.A(n_781),
.Y(n_1988)
);

BUFx3_ASAP7_75t_L g1989 ( 
.A(n_1517),
.Y(n_1989)
);

CKINVDCx5p33_ASAP7_75t_R g1990 ( 
.A(n_1510),
.Y(n_1990)
);

CKINVDCx14_ASAP7_75t_R g1991 ( 
.A(n_1686),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1058),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_285),
.Y(n_1993)
);

CKINVDCx5p33_ASAP7_75t_R g1994 ( 
.A(n_1112),
.Y(n_1994)
);

CKINVDCx5p33_ASAP7_75t_R g1995 ( 
.A(n_715),
.Y(n_1995)
);

CKINVDCx5p33_ASAP7_75t_R g1996 ( 
.A(n_1679),
.Y(n_1996)
);

CKINVDCx5p33_ASAP7_75t_R g1997 ( 
.A(n_452),
.Y(n_1997)
);

BUFx5_ASAP7_75t_L g1998 ( 
.A(n_1464),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_433),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1615),
.Y(n_2000)
);

CKINVDCx5p33_ASAP7_75t_R g2001 ( 
.A(n_56),
.Y(n_2001)
);

CKINVDCx14_ASAP7_75t_R g2002 ( 
.A(n_1674),
.Y(n_2002)
);

CKINVDCx5p33_ASAP7_75t_R g2003 ( 
.A(n_62),
.Y(n_2003)
);

CKINVDCx5p33_ASAP7_75t_R g2004 ( 
.A(n_76),
.Y(n_2004)
);

CKINVDCx5p33_ASAP7_75t_R g2005 ( 
.A(n_503),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1452),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1502),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1603),
.Y(n_2008)
);

CKINVDCx5p33_ASAP7_75t_R g2009 ( 
.A(n_1393),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_287),
.Y(n_2010)
);

CKINVDCx5p33_ASAP7_75t_R g2011 ( 
.A(n_1604),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1364),
.Y(n_2012)
);

CKINVDCx5p33_ASAP7_75t_R g2013 ( 
.A(n_314),
.Y(n_2013)
);

CKINVDCx16_ASAP7_75t_R g2014 ( 
.A(n_989),
.Y(n_2014)
);

CKINVDCx20_ASAP7_75t_R g2015 ( 
.A(n_40),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1627),
.Y(n_2016)
);

CKINVDCx5p33_ASAP7_75t_R g2017 ( 
.A(n_1447),
.Y(n_2017)
);

CKINVDCx5p33_ASAP7_75t_R g2018 ( 
.A(n_79),
.Y(n_2018)
);

CKINVDCx5p33_ASAP7_75t_R g2019 ( 
.A(n_180),
.Y(n_2019)
);

CKINVDCx5p33_ASAP7_75t_R g2020 ( 
.A(n_1706),
.Y(n_2020)
);

CKINVDCx5p33_ASAP7_75t_R g2021 ( 
.A(n_1441),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1021),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1050),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1168),
.Y(n_2024)
);

CKINVDCx20_ASAP7_75t_R g2025 ( 
.A(n_294),
.Y(n_2025)
);

CKINVDCx5p33_ASAP7_75t_R g2026 ( 
.A(n_522),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1532),
.Y(n_2027)
);

CKINVDCx5p33_ASAP7_75t_R g2028 ( 
.A(n_1406),
.Y(n_2028)
);

INVx2_ASAP7_75t_SL g2029 ( 
.A(n_1016),
.Y(n_2029)
);

CKINVDCx5p33_ASAP7_75t_R g2030 ( 
.A(n_1654),
.Y(n_2030)
);

CKINVDCx5p33_ASAP7_75t_R g2031 ( 
.A(n_981),
.Y(n_2031)
);

CKINVDCx5p33_ASAP7_75t_R g2032 ( 
.A(n_1651),
.Y(n_2032)
);

CKINVDCx5p33_ASAP7_75t_R g2033 ( 
.A(n_232),
.Y(n_2033)
);

CKINVDCx5p33_ASAP7_75t_R g2034 ( 
.A(n_1522),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1481),
.Y(n_2035)
);

INVx1_ASAP7_75t_SL g2036 ( 
.A(n_359),
.Y(n_2036)
);

BUFx3_ASAP7_75t_L g2037 ( 
.A(n_1106),
.Y(n_2037)
);

BUFx3_ASAP7_75t_L g2038 ( 
.A(n_344),
.Y(n_2038)
);

CKINVDCx5p33_ASAP7_75t_R g2039 ( 
.A(n_1049),
.Y(n_2039)
);

CKINVDCx20_ASAP7_75t_R g2040 ( 
.A(n_1358),
.Y(n_2040)
);

BUFx6f_ASAP7_75t_L g2041 ( 
.A(n_92),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1529),
.Y(n_2042)
);

CKINVDCx5p33_ASAP7_75t_R g2043 ( 
.A(n_1036),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_140),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_792),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1192),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1054),
.Y(n_2047)
);

CKINVDCx5p33_ASAP7_75t_R g2048 ( 
.A(n_1003),
.Y(n_2048)
);

INVx1_ASAP7_75t_SL g2049 ( 
.A(n_258),
.Y(n_2049)
);

INVxp67_ASAP7_75t_SL g2050 ( 
.A(n_955),
.Y(n_2050)
);

CKINVDCx5p33_ASAP7_75t_R g2051 ( 
.A(n_1729),
.Y(n_2051)
);

CKINVDCx5p33_ASAP7_75t_R g2052 ( 
.A(n_976),
.Y(n_2052)
);

INVx1_ASAP7_75t_SL g2053 ( 
.A(n_658),
.Y(n_2053)
);

CKINVDCx5p33_ASAP7_75t_R g2054 ( 
.A(n_1601),
.Y(n_2054)
);

INVx2_ASAP7_75t_SL g2055 ( 
.A(n_1701),
.Y(n_2055)
);

CKINVDCx16_ASAP7_75t_R g2056 ( 
.A(n_1307),
.Y(n_2056)
);

CKINVDCx5p33_ASAP7_75t_R g2057 ( 
.A(n_76),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_805),
.Y(n_2058)
);

CKINVDCx5p33_ASAP7_75t_R g2059 ( 
.A(n_70),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1245),
.Y(n_2060)
);

CKINVDCx20_ASAP7_75t_R g2061 ( 
.A(n_689),
.Y(n_2061)
);

CKINVDCx5p33_ASAP7_75t_R g2062 ( 
.A(n_1478),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_666),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_521),
.Y(n_2064)
);

CKINVDCx5p33_ASAP7_75t_R g2065 ( 
.A(n_1670),
.Y(n_2065)
);

CKINVDCx5p33_ASAP7_75t_R g2066 ( 
.A(n_692),
.Y(n_2066)
);

CKINVDCx5p33_ASAP7_75t_R g2067 ( 
.A(n_62),
.Y(n_2067)
);

CKINVDCx5p33_ASAP7_75t_R g2068 ( 
.A(n_1429),
.Y(n_2068)
);

BUFx10_ASAP7_75t_L g2069 ( 
.A(n_772),
.Y(n_2069)
);

CKINVDCx5p33_ASAP7_75t_R g2070 ( 
.A(n_333),
.Y(n_2070)
);

CKINVDCx5p33_ASAP7_75t_R g2071 ( 
.A(n_1511),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_989),
.Y(n_2072)
);

CKINVDCx5p33_ASAP7_75t_R g2073 ( 
.A(n_712),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_885),
.Y(n_2074)
);

INVx1_ASAP7_75t_SL g2075 ( 
.A(n_1053),
.Y(n_2075)
);

INVx1_ASAP7_75t_SL g2076 ( 
.A(n_1645),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1405),
.Y(n_2077)
);

CKINVDCx5p33_ASAP7_75t_R g2078 ( 
.A(n_976),
.Y(n_2078)
);

CKINVDCx5p33_ASAP7_75t_R g2079 ( 
.A(n_260),
.Y(n_2079)
);

CKINVDCx5p33_ASAP7_75t_R g2080 ( 
.A(n_1567),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1486),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_680),
.Y(n_2082)
);

CKINVDCx5p33_ASAP7_75t_R g2083 ( 
.A(n_1493),
.Y(n_2083)
);

CKINVDCx5p33_ASAP7_75t_R g2084 ( 
.A(n_343),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_511),
.Y(n_2085)
);

CKINVDCx5p33_ASAP7_75t_R g2086 ( 
.A(n_601),
.Y(n_2086)
);

CKINVDCx5p33_ASAP7_75t_R g2087 ( 
.A(n_907),
.Y(n_2087)
);

CKINVDCx5p33_ASAP7_75t_R g2088 ( 
.A(n_58),
.Y(n_2088)
);

CKINVDCx20_ASAP7_75t_R g2089 ( 
.A(n_447),
.Y(n_2089)
);

CKINVDCx5p33_ASAP7_75t_R g2090 ( 
.A(n_954),
.Y(n_2090)
);

INVx1_ASAP7_75t_SL g2091 ( 
.A(n_1520),
.Y(n_2091)
);

CKINVDCx5p33_ASAP7_75t_R g2092 ( 
.A(n_986),
.Y(n_2092)
);

CKINVDCx5p33_ASAP7_75t_R g2093 ( 
.A(n_635),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1313),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_125),
.Y(n_2095)
);

CKINVDCx5p33_ASAP7_75t_R g2096 ( 
.A(n_1053),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1422),
.Y(n_2097)
);

CKINVDCx5p33_ASAP7_75t_R g2098 ( 
.A(n_1413),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_646),
.Y(n_2099)
);

CKINVDCx5p33_ASAP7_75t_R g2100 ( 
.A(n_712),
.Y(n_2100)
);

CKINVDCx5p33_ASAP7_75t_R g2101 ( 
.A(n_1081),
.Y(n_2101)
);

CKINVDCx5p33_ASAP7_75t_R g2102 ( 
.A(n_1420),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1043),
.Y(n_2103)
);

CKINVDCx5p33_ASAP7_75t_R g2104 ( 
.A(n_1683),
.Y(n_2104)
);

CKINVDCx5p33_ASAP7_75t_R g2105 ( 
.A(n_1734),
.Y(n_2105)
);

CKINVDCx5p33_ASAP7_75t_R g2106 ( 
.A(n_1202),
.Y(n_2106)
);

CKINVDCx5p33_ASAP7_75t_R g2107 ( 
.A(n_1715),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_991),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_896),
.Y(n_2109)
);

CKINVDCx5p33_ASAP7_75t_R g2110 ( 
.A(n_1203),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_17),
.Y(n_2111)
);

CKINVDCx5p33_ASAP7_75t_R g2112 ( 
.A(n_286),
.Y(n_2112)
);

CKINVDCx5p33_ASAP7_75t_R g2113 ( 
.A(n_996),
.Y(n_2113)
);

CKINVDCx5p33_ASAP7_75t_R g2114 ( 
.A(n_853),
.Y(n_2114)
);

BUFx6f_ASAP7_75t_L g2115 ( 
.A(n_799),
.Y(n_2115)
);

CKINVDCx5p33_ASAP7_75t_R g2116 ( 
.A(n_1090),
.Y(n_2116)
);

CKINVDCx5p33_ASAP7_75t_R g2117 ( 
.A(n_650),
.Y(n_2117)
);

CKINVDCx5p33_ASAP7_75t_R g2118 ( 
.A(n_1586),
.Y(n_2118)
);

CKINVDCx5p33_ASAP7_75t_R g2119 ( 
.A(n_466),
.Y(n_2119)
);

INVxp67_ASAP7_75t_L g2120 ( 
.A(n_1484),
.Y(n_2120)
);

CKINVDCx5p33_ASAP7_75t_R g2121 ( 
.A(n_1678),
.Y(n_2121)
);

CKINVDCx5p33_ASAP7_75t_R g2122 ( 
.A(n_472),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1262),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_154),
.Y(n_2124)
);

CKINVDCx5p33_ASAP7_75t_R g2125 ( 
.A(n_705),
.Y(n_2125)
);

CKINVDCx5p33_ASAP7_75t_R g2126 ( 
.A(n_456),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1519),
.Y(n_2127)
);

CKINVDCx5p33_ASAP7_75t_R g2128 ( 
.A(n_150),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1566),
.Y(n_2129)
);

CKINVDCx5p33_ASAP7_75t_R g2130 ( 
.A(n_1685),
.Y(n_2130)
);

CKINVDCx5p33_ASAP7_75t_R g2131 ( 
.A(n_777),
.Y(n_2131)
);

CKINVDCx16_ASAP7_75t_R g2132 ( 
.A(n_275),
.Y(n_2132)
);

BUFx3_ASAP7_75t_L g2133 ( 
.A(n_339),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_596),
.Y(n_2134)
);

CKINVDCx5p33_ASAP7_75t_R g2135 ( 
.A(n_1152),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_388),
.Y(n_2136)
);

CKINVDCx5p33_ASAP7_75t_R g2137 ( 
.A(n_856),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_1068),
.Y(n_2138)
);

CKINVDCx20_ASAP7_75t_R g2139 ( 
.A(n_678),
.Y(n_2139)
);

CKINVDCx5p33_ASAP7_75t_R g2140 ( 
.A(n_1591),
.Y(n_2140)
);

INVx2_ASAP7_75t_SL g2141 ( 
.A(n_1369),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_730),
.Y(n_2142)
);

CKINVDCx20_ASAP7_75t_R g2143 ( 
.A(n_824),
.Y(n_2143)
);

CKINVDCx5p33_ASAP7_75t_R g2144 ( 
.A(n_24),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_1334),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1368),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_467),
.Y(n_2147)
);

CKINVDCx5p33_ASAP7_75t_R g2148 ( 
.A(n_1728),
.Y(n_2148)
);

CKINVDCx16_ASAP7_75t_R g2149 ( 
.A(n_844),
.Y(n_2149)
);

CKINVDCx5p33_ASAP7_75t_R g2150 ( 
.A(n_361),
.Y(n_2150)
);

CKINVDCx5p33_ASAP7_75t_R g2151 ( 
.A(n_1637),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_1434),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_1230),
.Y(n_2153)
);

CKINVDCx5p33_ASAP7_75t_R g2154 ( 
.A(n_1026),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1658),
.Y(n_2155)
);

CKINVDCx5p33_ASAP7_75t_R g2156 ( 
.A(n_44),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_999),
.Y(n_2157)
);

INVx1_ASAP7_75t_SL g2158 ( 
.A(n_147),
.Y(n_2158)
);

CKINVDCx5p33_ASAP7_75t_R g2159 ( 
.A(n_181),
.Y(n_2159)
);

CKINVDCx20_ASAP7_75t_R g2160 ( 
.A(n_699),
.Y(n_2160)
);

CKINVDCx5p33_ASAP7_75t_R g2161 ( 
.A(n_1337),
.Y(n_2161)
);

INVx2_ASAP7_75t_SL g2162 ( 
.A(n_922),
.Y(n_2162)
);

CKINVDCx5p33_ASAP7_75t_R g2163 ( 
.A(n_1206),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_1636),
.Y(n_2164)
);

CKINVDCx5p33_ASAP7_75t_R g2165 ( 
.A(n_1505),
.Y(n_2165)
);

CKINVDCx5p33_ASAP7_75t_R g2166 ( 
.A(n_1704),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_169),
.Y(n_2167)
);

CKINVDCx5p33_ASAP7_75t_R g2168 ( 
.A(n_1626),
.Y(n_2168)
);

INVxp33_ASAP7_75t_SL g2169 ( 
.A(n_859),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1617),
.Y(n_2170)
);

CKINVDCx5p33_ASAP7_75t_R g2171 ( 
.A(n_803),
.Y(n_2171)
);

CKINVDCx5p33_ASAP7_75t_R g2172 ( 
.A(n_1267),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_808),
.Y(n_2173)
);

CKINVDCx5p33_ASAP7_75t_R g2174 ( 
.A(n_830),
.Y(n_2174)
);

CKINVDCx5p33_ASAP7_75t_R g2175 ( 
.A(n_146),
.Y(n_2175)
);

CKINVDCx5p33_ASAP7_75t_R g2176 ( 
.A(n_192),
.Y(n_2176)
);

CKINVDCx5p33_ASAP7_75t_R g2177 ( 
.A(n_870),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1561),
.Y(n_2178)
);

CKINVDCx5p33_ASAP7_75t_R g2179 ( 
.A(n_1232),
.Y(n_2179)
);

CKINVDCx5p33_ASAP7_75t_R g2180 ( 
.A(n_1415),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1518),
.Y(n_2181)
);

BUFx2_ASAP7_75t_SL g2182 ( 
.A(n_1398),
.Y(n_2182)
);

INVx1_ASAP7_75t_SL g2183 ( 
.A(n_428),
.Y(n_2183)
);

CKINVDCx5p33_ASAP7_75t_R g2184 ( 
.A(n_911),
.Y(n_2184)
);

CKINVDCx5p33_ASAP7_75t_R g2185 ( 
.A(n_1536),
.Y(n_2185)
);

CKINVDCx5p33_ASAP7_75t_R g2186 ( 
.A(n_791),
.Y(n_2186)
);

CKINVDCx5p33_ASAP7_75t_R g2187 ( 
.A(n_670),
.Y(n_2187)
);

CKINVDCx5p33_ASAP7_75t_R g2188 ( 
.A(n_666),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1465),
.Y(n_2189)
);

CKINVDCx16_ASAP7_75t_R g2190 ( 
.A(n_1046),
.Y(n_2190)
);

CKINVDCx16_ASAP7_75t_R g2191 ( 
.A(n_1180),
.Y(n_2191)
);

CKINVDCx5p33_ASAP7_75t_R g2192 ( 
.A(n_359),
.Y(n_2192)
);

CKINVDCx20_ASAP7_75t_R g2193 ( 
.A(n_1708),
.Y(n_2193)
);

BUFx8_ASAP7_75t_SL g2194 ( 
.A(n_1646),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_1357),
.Y(n_2195)
);

INVxp67_ASAP7_75t_L g2196 ( 
.A(n_865),
.Y(n_2196)
);

CKINVDCx5p33_ASAP7_75t_R g2197 ( 
.A(n_1236),
.Y(n_2197)
);

CKINVDCx5p33_ASAP7_75t_R g2198 ( 
.A(n_523),
.Y(n_2198)
);

HB1xp67_ASAP7_75t_L g2199 ( 
.A(n_1439),
.Y(n_2199)
);

CKINVDCx5p33_ASAP7_75t_R g2200 ( 
.A(n_149),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1540),
.Y(n_2201)
);

CKINVDCx5p33_ASAP7_75t_R g2202 ( 
.A(n_266),
.Y(n_2202)
);

CKINVDCx5p33_ASAP7_75t_R g2203 ( 
.A(n_1521),
.Y(n_2203)
);

CKINVDCx5p33_ASAP7_75t_R g2204 ( 
.A(n_584),
.Y(n_2204)
);

HB1xp67_ASAP7_75t_L g2205 ( 
.A(n_1559),
.Y(n_2205)
);

CKINVDCx5p33_ASAP7_75t_R g2206 ( 
.A(n_1241),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1635),
.Y(n_2207)
);

BUFx3_ASAP7_75t_L g2208 ( 
.A(n_1019),
.Y(n_2208)
);

CKINVDCx5p33_ASAP7_75t_R g2209 ( 
.A(n_1187),
.Y(n_2209)
);

CKINVDCx5p33_ASAP7_75t_R g2210 ( 
.A(n_1736),
.Y(n_2210)
);

CKINVDCx20_ASAP7_75t_R g2211 ( 
.A(n_1020),
.Y(n_2211)
);

CKINVDCx5p33_ASAP7_75t_R g2212 ( 
.A(n_931),
.Y(n_2212)
);

CKINVDCx5p33_ASAP7_75t_R g2213 ( 
.A(n_1419),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_1491),
.Y(n_2214)
);

CKINVDCx20_ASAP7_75t_R g2215 ( 
.A(n_1463),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1543),
.Y(n_2216)
);

CKINVDCx5p33_ASAP7_75t_R g2217 ( 
.A(n_647),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_824),
.Y(n_2218)
);

CKINVDCx5p33_ASAP7_75t_R g2219 ( 
.A(n_1018),
.Y(n_2219)
);

CKINVDCx5p33_ASAP7_75t_R g2220 ( 
.A(n_1545),
.Y(n_2220)
);

CKINVDCx5p33_ASAP7_75t_R g2221 ( 
.A(n_1527),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_964),
.Y(n_2222)
);

INVxp33_ASAP7_75t_SL g2223 ( 
.A(n_432),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_538),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1395),
.Y(n_2225)
);

CKINVDCx20_ASAP7_75t_R g2226 ( 
.A(n_408),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_117),
.Y(n_2227)
);

CKINVDCx5p33_ASAP7_75t_R g2228 ( 
.A(n_1642),
.Y(n_2228)
);

CKINVDCx5p33_ASAP7_75t_R g2229 ( 
.A(n_1059),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_556),
.Y(n_2230)
);

CKINVDCx5p33_ASAP7_75t_R g2231 ( 
.A(n_1573),
.Y(n_2231)
);

BUFx10_ASAP7_75t_L g2232 ( 
.A(n_507),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_478),
.Y(n_2233)
);

CKINVDCx5p33_ASAP7_75t_R g2234 ( 
.A(n_1361),
.Y(n_2234)
);

CKINVDCx5p33_ASAP7_75t_R g2235 ( 
.A(n_1013),
.Y(n_2235)
);

CKINVDCx5p33_ASAP7_75t_R g2236 ( 
.A(n_579),
.Y(n_2236)
);

CKINVDCx5p33_ASAP7_75t_R g2237 ( 
.A(n_1535),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_1655),
.Y(n_2238)
);

INVx1_ASAP7_75t_SL g2239 ( 
.A(n_118),
.Y(n_2239)
);

CKINVDCx5p33_ASAP7_75t_R g2240 ( 
.A(n_1316),
.Y(n_2240)
);

CKINVDCx5p33_ASAP7_75t_R g2241 ( 
.A(n_798),
.Y(n_2241)
);

CKINVDCx16_ASAP7_75t_R g2242 ( 
.A(n_754),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_340),
.Y(n_2243)
);

CKINVDCx20_ASAP7_75t_R g2244 ( 
.A(n_403),
.Y(n_2244)
);

BUFx6f_ASAP7_75t_L g2245 ( 
.A(n_527),
.Y(n_2245)
);

CKINVDCx5p33_ASAP7_75t_R g2246 ( 
.A(n_1123),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_1713),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_742),
.Y(n_2248)
);

CKINVDCx5p33_ASAP7_75t_R g2249 ( 
.A(n_984),
.Y(n_2249)
);

INVx2_ASAP7_75t_L g2250 ( 
.A(n_768),
.Y(n_2250)
);

INVx2_ASAP7_75t_L g2251 ( 
.A(n_1296),
.Y(n_2251)
);

INVx1_ASAP7_75t_SL g2252 ( 
.A(n_1710),
.Y(n_2252)
);

CKINVDCx5p33_ASAP7_75t_R g2253 ( 
.A(n_34),
.Y(n_2253)
);

CKINVDCx16_ASAP7_75t_R g2254 ( 
.A(n_1614),
.Y(n_2254)
);

CKINVDCx5p33_ASAP7_75t_R g2255 ( 
.A(n_136),
.Y(n_2255)
);

INVx2_ASAP7_75t_L g2256 ( 
.A(n_99),
.Y(n_2256)
);

CKINVDCx5p33_ASAP7_75t_R g2257 ( 
.A(n_1467),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_1599),
.Y(n_2258)
);

BUFx5_ASAP7_75t_L g2259 ( 
.A(n_237),
.Y(n_2259)
);

CKINVDCx5p33_ASAP7_75t_R g2260 ( 
.A(n_1693),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1071),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_1031),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_1014),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_560),
.Y(n_2264)
);

CKINVDCx5p33_ASAP7_75t_R g2265 ( 
.A(n_1017),
.Y(n_2265)
);

CKINVDCx5p33_ASAP7_75t_R g2266 ( 
.A(n_1677),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_1412),
.Y(n_2267)
);

CKINVDCx5p33_ASAP7_75t_R g2268 ( 
.A(n_1681),
.Y(n_2268)
);

BUFx3_ASAP7_75t_L g2269 ( 
.A(n_897),
.Y(n_2269)
);

CKINVDCx5p33_ASAP7_75t_R g2270 ( 
.A(n_980),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_536),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_995),
.Y(n_2272)
);

BUFx6f_ASAP7_75t_L g2273 ( 
.A(n_1538),
.Y(n_2273)
);

CKINVDCx5p33_ASAP7_75t_R g2274 ( 
.A(n_583),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_1205),
.Y(n_2275)
);

CKINVDCx5p33_ASAP7_75t_R g2276 ( 
.A(n_1397),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_575),
.Y(n_2277)
);

CKINVDCx5p33_ASAP7_75t_R g2278 ( 
.A(n_469),
.Y(n_2278)
);

CKINVDCx5p33_ASAP7_75t_R g2279 ( 
.A(n_972),
.Y(n_2279)
);

CKINVDCx20_ASAP7_75t_R g2280 ( 
.A(n_232),
.Y(n_2280)
);

INVx2_ASAP7_75t_L g2281 ( 
.A(n_1229),
.Y(n_2281)
);

CKINVDCx5p33_ASAP7_75t_R g2282 ( 
.A(n_804),
.Y(n_2282)
);

BUFx8_ASAP7_75t_SL g2283 ( 
.A(n_1375),
.Y(n_2283)
);

BUFx5_ASAP7_75t_L g2284 ( 
.A(n_1731),
.Y(n_2284)
);

CKINVDCx5p33_ASAP7_75t_R g2285 ( 
.A(n_271),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_1725),
.Y(n_2286)
);

CKINVDCx5p33_ASAP7_75t_R g2287 ( 
.A(n_202),
.Y(n_2287)
);

CKINVDCx5p33_ASAP7_75t_R g2288 ( 
.A(n_1516),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_1182),
.Y(n_2289)
);

CKINVDCx5p33_ASAP7_75t_R g2290 ( 
.A(n_558),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_743),
.Y(n_2291)
);

CKINVDCx5p33_ASAP7_75t_R g2292 ( 
.A(n_398),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_1682),
.Y(n_2293)
);

INVx2_ASAP7_75t_L g2294 ( 
.A(n_614),
.Y(n_2294)
);

HB1xp67_ASAP7_75t_L g2295 ( 
.A(n_889),
.Y(n_2295)
);

CKINVDCx5p33_ASAP7_75t_R g2296 ( 
.A(n_1632),
.Y(n_2296)
);

CKINVDCx5p33_ASAP7_75t_R g2297 ( 
.A(n_965),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_1320),
.Y(n_2298)
);

INVx4_ASAP7_75t_R g2299 ( 
.A(n_661),
.Y(n_2299)
);

CKINVDCx5p33_ASAP7_75t_R g2300 ( 
.A(n_562),
.Y(n_2300)
);

CKINVDCx5p33_ASAP7_75t_R g2301 ( 
.A(n_1336),
.Y(n_2301)
);

CKINVDCx5p33_ASAP7_75t_R g2302 ( 
.A(n_816),
.Y(n_2302)
);

INVx1_ASAP7_75t_SL g2303 ( 
.A(n_2),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_154),
.Y(n_2304)
);

CKINVDCx5p33_ASAP7_75t_R g2305 ( 
.A(n_850),
.Y(n_2305)
);

BUFx2_ASAP7_75t_L g2306 ( 
.A(n_197),
.Y(n_2306)
);

CKINVDCx5p33_ASAP7_75t_R g2307 ( 
.A(n_10),
.Y(n_2307)
);

INVx2_ASAP7_75t_SL g2308 ( 
.A(n_1547),
.Y(n_2308)
);

CKINVDCx5p33_ASAP7_75t_R g2309 ( 
.A(n_481),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_987),
.Y(n_2310)
);

CKINVDCx5p33_ASAP7_75t_R g2311 ( 
.A(n_1028),
.Y(n_2311)
);

CKINVDCx5p33_ASAP7_75t_R g2312 ( 
.A(n_1204),
.Y(n_2312)
);

CKINVDCx5p33_ASAP7_75t_R g2313 ( 
.A(n_1509),
.Y(n_2313)
);

CKINVDCx5p33_ASAP7_75t_R g2314 ( 
.A(n_1005),
.Y(n_2314)
);

BUFx3_ASAP7_75t_L g2315 ( 
.A(n_1054),
.Y(n_2315)
);

CKINVDCx5p33_ASAP7_75t_R g2316 ( 
.A(n_1237),
.Y(n_2316)
);

CKINVDCx5p33_ASAP7_75t_R g2317 ( 
.A(n_461),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_150),
.Y(n_2318)
);

CKINVDCx5p33_ASAP7_75t_R g2319 ( 
.A(n_1513),
.Y(n_2319)
);

CKINVDCx5p33_ASAP7_75t_R g2320 ( 
.A(n_515),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_720),
.Y(n_2321)
);

CKINVDCx5p33_ASAP7_75t_R g2322 ( 
.A(n_1476),
.Y(n_2322)
);

CKINVDCx5p33_ASAP7_75t_R g2323 ( 
.A(n_1078),
.Y(n_2323)
);

CKINVDCx5p33_ASAP7_75t_R g2324 ( 
.A(n_1327),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_1367),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_435),
.Y(n_2326)
);

CKINVDCx20_ASAP7_75t_R g2327 ( 
.A(n_110),
.Y(n_2327)
);

CKINVDCx5p33_ASAP7_75t_R g2328 ( 
.A(n_1134),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_492),
.Y(n_2329)
);

CKINVDCx5p33_ASAP7_75t_R g2330 ( 
.A(n_1477),
.Y(n_2330)
);

CKINVDCx5p33_ASAP7_75t_R g2331 ( 
.A(n_1719),
.Y(n_2331)
);

CKINVDCx5p33_ASAP7_75t_R g2332 ( 
.A(n_1057),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_85),
.Y(n_2333)
);

CKINVDCx5p33_ASAP7_75t_R g2334 ( 
.A(n_1471),
.Y(n_2334)
);

CKINVDCx5p33_ASAP7_75t_R g2335 ( 
.A(n_175),
.Y(n_2335)
);

CKINVDCx5p33_ASAP7_75t_R g2336 ( 
.A(n_947),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_471),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_1089),
.Y(n_2338)
);

CKINVDCx5p33_ASAP7_75t_R g2339 ( 
.A(n_1114),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_1238),
.Y(n_2340)
);

CKINVDCx5p33_ASAP7_75t_R g2341 ( 
.A(n_82),
.Y(n_2341)
);

CKINVDCx5p33_ASAP7_75t_R g2342 ( 
.A(n_69),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_409),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_983),
.Y(n_2344)
);

CKINVDCx5p33_ASAP7_75t_R g2345 ( 
.A(n_329),
.Y(n_2345)
);

CKINVDCx5p33_ASAP7_75t_R g2346 ( 
.A(n_1209),
.Y(n_2346)
);

INVx2_ASAP7_75t_SL g2347 ( 
.A(n_847),
.Y(n_2347)
);

CKINVDCx5p33_ASAP7_75t_R g2348 ( 
.A(n_1727),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_1243),
.Y(n_2349)
);

CKINVDCx5p33_ASAP7_75t_R g2350 ( 
.A(n_1608),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_107),
.Y(n_2351)
);

CKINVDCx5p33_ASAP7_75t_R g2352 ( 
.A(n_1255),
.Y(n_2352)
);

CKINVDCx20_ASAP7_75t_R g2353 ( 
.A(n_1691),
.Y(n_2353)
);

CKINVDCx5p33_ASAP7_75t_R g2354 ( 
.A(n_1260),
.Y(n_2354)
);

INVxp33_ASAP7_75t_SL g2355 ( 
.A(n_167),
.Y(n_2355)
);

CKINVDCx5p33_ASAP7_75t_R g2356 ( 
.A(n_1394),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_985),
.Y(n_2357)
);

CKINVDCx5p33_ASAP7_75t_R g2358 ( 
.A(n_1011),
.Y(n_2358)
);

CKINVDCx5p33_ASAP7_75t_R g2359 ( 
.A(n_10),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_787),
.Y(n_2360)
);

CKINVDCx5p33_ASAP7_75t_R g2361 ( 
.A(n_1475),
.Y(n_2361)
);

CKINVDCx5p33_ASAP7_75t_R g2362 ( 
.A(n_1039),
.Y(n_2362)
);

CKINVDCx5p33_ASAP7_75t_R g2363 ( 
.A(n_1154),
.Y(n_2363)
);

CKINVDCx5p33_ASAP7_75t_R g2364 ( 
.A(n_1542),
.Y(n_2364)
);

CKINVDCx5p33_ASAP7_75t_R g2365 ( 
.A(n_323),
.Y(n_2365)
);

CKINVDCx5p33_ASAP7_75t_R g2366 ( 
.A(n_218),
.Y(n_2366)
);

CKINVDCx20_ASAP7_75t_R g2367 ( 
.A(n_1195),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_440),
.Y(n_2368)
);

CKINVDCx5p33_ASAP7_75t_R g2369 ( 
.A(n_97),
.Y(n_2369)
);

CKINVDCx5p33_ASAP7_75t_R g2370 ( 
.A(n_43),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_1644),
.Y(n_2371)
);

BUFx10_ASAP7_75t_L g2372 ( 
.A(n_596),
.Y(n_2372)
);

BUFx3_ASAP7_75t_L g2373 ( 
.A(n_921),
.Y(n_2373)
);

INVx1_ASAP7_75t_SL g2374 ( 
.A(n_982),
.Y(n_2374)
);

CKINVDCx5p33_ASAP7_75t_R g2375 ( 
.A(n_374),
.Y(n_2375)
);

CKINVDCx5p33_ASAP7_75t_R g2376 ( 
.A(n_1287),
.Y(n_2376)
);

BUFx3_ASAP7_75t_L g2377 ( 
.A(n_1310),
.Y(n_2377)
);

CKINVDCx5p33_ASAP7_75t_R g2378 ( 
.A(n_1239),
.Y(n_2378)
);

CKINVDCx5p33_ASAP7_75t_R g2379 ( 
.A(n_954),
.Y(n_2379)
);

BUFx3_ASAP7_75t_L g2380 ( 
.A(n_354),
.Y(n_2380)
);

CKINVDCx16_ASAP7_75t_R g2381 ( 
.A(n_628),
.Y(n_2381)
);

CKINVDCx5p33_ASAP7_75t_R g2382 ( 
.A(n_1344),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_1606),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_1025),
.Y(n_2384)
);

CKINVDCx5p33_ASAP7_75t_R g2385 ( 
.A(n_1167),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_1625),
.Y(n_2386)
);

CKINVDCx5p33_ASAP7_75t_R g2387 ( 
.A(n_1281),
.Y(n_2387)
);

CKINVDCx5p33_ASAP7_75t_R g2388 ( 
.A(n_1056),
.Y(n_2388)
);

CKINVDCx5p33_ASAP7_75t_R g2389 ( 
.A(n_1498),
.Y(n_2389)
);

CKINVDCx20_ASAP7_75t_R g2390 ( 
.A(n_1200),
.Y(n_2390)
);

BUFx6f_ASAP7_75t_L g2391 ( 
.A(n_1451),
.Y(n_2391)
);

BUFx6f_ASAP7_75t_L g2392 ( 
.A(n_643),
.Y(n_2392)
);

CKINVDCx16_ASAP7_75t_R g2393 ( 
.A(n_1707),
.Y(n_2393)
);

INVx1_ASAP7_75t_SL g2394 ( 
.A(n_579),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_1174),
.Y(n_2395)
);

CKINVDCx5p33_ASAP7_75t_R g2396 ( 
.A(n_670),
.Y(n_2396)
);

CKINVDCx5p33_ASAP7_75t_R g2397 ( 
.A(n_1585),
.Y(n_2397)
);

INVxp67_ASAP7_75t_L g2398 ( 
.A(n_101),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_460),
.Y(n_2399)
);

CKINVDCx5p33_ASAP7_75t_R g2400 ( 
.A(n_272),
.Y(n_2400)
);

BUFx3_ASAP7_75t_L g2401 ( 
.A(n_44),
.Y(n_2401)
);

CKINVDCx5p33_ASAP7_75t_R g2402 ( 
.A(n_105),
.Y(n_2402)
);

CKINVDCx5p33_ASAP7_75t_R g2403 ( 
.A(n_93),
.Y(n_2403)
);

CKINVDCx5p33_ASAP7_75t_R g2404 ( 
.A(n_876),
.Y(n_2404)
);

CKINVDCx5p33_ASAP7_75t_R g2405 ( 
.A(n_1541),
.Y(n_2405)
);

CKINVDCx5p33_ASAP7_75t_R g2406 ( 
.A(n_1220),
.Y(n_2406)
);

CKINVDCx5p33_ASAP7_75t_R g2407 ( 
.A(n_1083),
.Y(n_2407)
);

CKINVDCx5p33_ASAP7_75t_R g2408 ( 
.A(n_358),
.Y(n_2408)
);

CKINVDCx5p33_ASAP7_75t_R g2409 ( 
.A(n_866),
.Y(n_2409)
);

CKINVDCx5p33_ASAP7_75t_R g2410 ( 
.A(n_627),
.Y(n_2410)
);

CKINVDCx5p33_ASAP7_75t_R g2411 ( 
.A(n_946),
.Y(n_2411)
);

CKINVDCx20_ASAP7_75t_R g2412 ( 
.A(n_1403),
.Y(n_2412)
);

BUFx2_ASAP7_75t_R g2413 ( 
.A(n_444),
.Y(n_2413)
);

CKINVDCx5p33_ASAP7_75t_R g2414 ( 
.A(n_793),
.Y(n_2414)
);

CKINVDCx5p33_ASAP7_75t_R g2415 ( 
.A(n_109),
.Y(n_2415)
);

INVx1_ASAP7_75t_SL g2416 ( 
.A(n_1032),
.Y(n_2416)
);

CKINVDCx5p33_ASAP7_75t_R g2417 ( 
.A(n_667),
.Y(n_2417)
);

CKINVDCx5p33_ASAP7_75t_R g2418 ( 
.A(n_681),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_664),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_612),
.Y(n_2420)
);

CKINVDCx5p33_ASAP7_75t_R g2421 ( 
.A(n_1146),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_721),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_66),
.Y(n_2423)
);

CKINVDCx5p33_ASAP7_75t_R g2424 ( 
.A(n_1128),
.Y(n_2424)
);

CKINVDCx14_ASAP7_75t_R g2425 ( 
.A(n_760),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_724),
.Y(n_2426)
);

CKINVDCx5p33_ASAP7_75t_R g2427 ( 
.A(n_926),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_773),
.Y(n_2428)
);

CKINVDCx5p33_ASAP7_75t_R g2429 ( 
.A(n_1549),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_1612),
.Y(n_2430)
);

INVx2_ASAP7_75t_L g2431 ( 
.A(n_992),
.Y(n_2431)
);

CKINVDCx5p33_ASAP7_75t_R g2432 ( 
.A(n_1534),
.Y(n_2432)
);

CKINVDCx5p33_ASAP7_75t_R g2433 ( 
.A(n_1047),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_1425),
.Y(n_2434)
);

CKINVDCx16_ASAP7_75t_R g2435 ( 
.A(n_288),
.Y(n_2435)
);

CKINVDCx5p33_ASAP7_75t_R g2436 ( 
.A(n_1548),
.Y(n_2436)
);

CKINVDCx5p33_ASAP7_75t_R g2437 ( 
.A(n_488),
.Y(n_2437)
);

INVx2_ASAP7_75t_SL g2438 ( 
.A(n_164),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_1551),
.Y(n_2439)
);

CKINVDCx5p33_ASAP7_75t_R g2440 ( 
.A(n_1034),
.Y(n_2440)
);

CKINVDCx5p33_ASAP7_75t_R g2441 ( 
.A(n_1594),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_1544),
.Y(n_2442)
);

INVx1_ASAP7_75t_SL g2443 ( 
.A(n_1583),
.Y(n_2443)
);

CKINVDCx5p33_ASAP7_75t_R g2444 ( 
.A(n_684),
.Y(n_2444)
);

CKINVDCx5p33_ASAP7_75t_R g2445 ( 
.A(n_697),
.Y(n_2445)
);

CKINVDCx16_ASAP7_75t_R g2446 ( 
.A(n_611),
.Y(n_2446)
);

INVx2_ASAP7_75t_SL g2447 ( 
.A(n_153),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_729),
.Y(n_2448)
);

CKINVDCx5p33_ASAP7_75t_R g2449 ( 
.A(n_1353),
.Y(n_2449)
);

CKINVDCx5p33_ASAP7_75t_R g2450 ( 
.A(n_1546),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_888),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_1711),
.Y(n_2452)
);

CKINVDCx5p33_ASAP7_75t_R g2453 ( 
.A(n_102),
.Y(n_2453)
);

CKINVDCx5p33_ASAP7_75t_R g2454 ( 
.A(n_1596),
.Y(n_2454)
);

INVxp67_ASAP7_75t_SL g2455 ( 
.A(n_468),
.Y(n_2455)
);

CKINVDCx5p33_ASAP7_75t_R g2456 ( 
.A(n_1515),
.Y(n_2456)
);

CKINVDCx5p33_ASAP7_75t_R g2457 ( 
.A(n_1722),
.Y(n_2457)
);

BUFx3_ASAP7_75t_L g2458 ( 
.A(n_990),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_1663),
.Y(n_2459)
);

CKINVDCx5p33_ASAP7_75t_R g2460 ( 
.A(n_829),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_494),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_1575),
.Y(n_2462)
);

INVx1_ASAP7_75t_SL g2463 ( 
.A(n_67),
.Y(n_2463)
);

CKINVDCx5p33_ASAP7_75t_R g2464 ( 
.A(n_796),
.Y(n_2464)
);

INVx2_ASAP7_75t_SL g2465 ( 
.A(n_948),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_1025),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_1219),
.Y(n_2467)
);

INVx1_ASAP7_75t_SL g2468 ( 
.A(n_322),
.Y(n_2468)
);

CKINVDCx5p33_ASAP7_75t_R g2469 ( 
.A(n_151),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_1193),
.Y(n_2470)
);

INVx2_ASAP7_75t_SL g2471 ( 
.A(n_1018),
.Y(n_2471)
);

CKINVDCx5p33_ASAP7_75t_R g2472 ( 
.A(n_1473),
.Y(n_2472)
);

CKINVDCx5p33_ASAP7_75t_R g2473 ( 
.A(n_693),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_746),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_679),
.Y(n_2475)
);

CKINVDCx5p33_ASAP7_75t_R g2476 ( 
.A(n_88),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_15),
.Y(n_2477)
);

CKINVDCx5p33_ASAP7_75t_R g2478 ( 
.A(n_988),
.Y(n_2478)
);

CKINVDCx5p33_ASAP7_75t_R g2479 ( 
.A(n_1592),
.Y(n_2479)
);

CKINVDCx5p33_ASAP7_75t_R g2480 ( 
.A(n_65),
.Y(n_2480)
);

CKINVDCx5p33_ASAP7_75t_R g2481 ( 
.A(n_507),
.Y(n_2481)
);

INVx2_ASAP7_75t_L g2482 ( 
.A(n_320),
.Y(n_2482)
);

CKINVDCx5p33_ASAP7_75t_R g2483 ( 
.A(n_677),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_1508),
.Y(n_2484)
);

INVx2_ASAP7_75t_SL g2485 ( 
.A(n_1279),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_928),
.Y(n_2486)
);

CKINVDCx5p33_ASAP7_75t_R g2487 ( 
.A(n_13),
.Y(n_2487)
);

CKINVDCx5p33_ASAP7_75t_R g2488 ( 
.A(n_1352),
.Y(n_2488)
);

CKINVDCx5p33_ASAP7_75t_R g2489 ( 
.A(n_1550),
.Y(n_2489)
);

INVx2_ASAP7_75t_L g2490 ( 
.A(n_849),
.Y(n_2490)
);

CKINVDCx5p33_ASAP7_75t_R g2491 ( 
.A(n_74),
.Y(n_2491)
);

CKINVDCx20_ASAP7_75t_R g2492 ( 
.A(n_783),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_997),
.Y(n_2493)
);

BUFx6f_ASAP7_75t_L g2494 ( 
.A(n_1474),
.Y(n_2494)
);

CKINVDCx20_ASAP7_75t_R g2495 ( 
.A(n_1623),
.Y(n_2495)
);

INVx1_ASAP7_75t_SL g2496 ( 
.A(n_1186),
.Y(n_2496)
);

INVx2_ASAP7_75t_SL g2497 ( 
.A(n_939),
.Y(n_2497)
);

CKINVDCx5p33_ASAP7_75t_R g2498 ( 
.A(n_907),
.Y(n_2498)
);

BUFx3_ASAP7_75t_L g2499 ( 
.A(n_243),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_700),
.Y(n_2500)
);

BUFx8_ASAP7_75t_SL g2501 ( 
.A(n_1482),
.Y(n_2501)
);

CKINVDCx5p33_ASAP7_75t_R g2502 ( 
.A(n_536),
.Y(n_2502)
);

CKINVDCx5p33_ASAP7_75t_R g2503 ( 
.A(n_1355),
.Y(n_2503)
);

INVx2_ASAP7_75t_SL g2504 ( 
.A(n_1184),
.Y(n_2504)
);

CKINVDCx5p33_ASAP7_75t_R g2505 ( 
.A(n_56),
.Y(n_2505)
);

CKINVDCx5p33_ASAP7_75t_R g2506 ( 
.A(n_1500),
.Y(n_2506)
);

CKINVDCx20_ASAP7_75t_R g2507 ( 
.A(n_1231),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_1189),
.Y(n_2508)
);

INVx2_ASAP7_75t_SL g2509 ( 
.A(n_862),
.Y(n_2509)
);

BUFx3_ASAP7_75t_L g2510 ( 
.A(n_1280),
.Y(n_2510)
);

BUFx3_ASAP7_75t_L g2511 ( 
.A(n_349),
.Y(n_2511)
);

CKINVDCx20_ASAP7_75t_R g2512 ( 
.A(n_255),
.Y(n_2512)
);

CKINVDCx5p33_ASAP7_75t_R g2513 ( 
.A(n_936),
.Y(n_2513)
);

CKINVDCx5p33_ASAP7_75t_R g2514 ( 
.A(n_89),
.Y(n_2514)
);

CKINVDCx5p33_ASAP7_75t_R g2515 ( 
.A(n_1360),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_1400),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_351),
.Y(n_2517)
);

CKINVDCx20_ASAP7_75t_R g2518 ( 
.A(n_1489),
.Y(n_2518)
);

CKINVDCx5p33_ASAP7_75t_R g2519 ( 
.A(n_513),
.Y(n_2519)
);

INVx2_ASAP7_75t_L g2520 ( 
.A(n_68),
.Y(n_2520)
);

CKINVDCx5p33_ASAP7_75t_R g2521 ( 
.A(n_358),
.Y(n_2521)
);

BUFx3_ASAP7_75t_L g2522 ( 
.A(n_1035),
.Y(n_2522)
);

CKINVDCx5p33_ASAP7_75t_R g2523 ( 
.A(n_629),
.Y(n_2523)
);

CKINVDCx20_ASAP7_75t_R g2524 ( 
.A(n_1363),
.Y(n_2524)
);

CKINVDCx5p33_ASAP7_75t_R g2525 ( 
.A(n_1042),
.Y(n_2525)
);

CKINVDCx5p33_ASAP7_75t_R g2526 ( 
.A(n_532),
.Y(n_2526)
);

INVx1_ASAP7_75t_SL g2527 ( 
.A(n_510),
.Y(n_2527)
);

CKINVDCx5p33_ASAP7_75t_R g2528 ( 
.A(n_1630),
.Y(n_2528)
);

CKINVDCx5p33_ASAP7_75t_R g2529 ( 
.A(n_1602),
.Y(n_2529)
);

CKINVDCx5p33_ASAP7_75t_R g2530 ( 
.A(n_110),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_1213),
.Y(n_2531)
);

CKINVDCx5p33_ASAP7_75t_R g2532 ( 
.A(n_20),
.Y(n_2532)
);

BUFx5_ASAP7_75t_L g2533 ( 
.A(n_1442),
.Y(n_2533)
);

INVxp67_ASAP7_75t_L g2534 ( 
.A(n_884),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_253),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_1688),
.Y(n_2536)
);

INVx1_ASAP7_75t_SL g2537 ( 
.A(n_1723),
.Y(n_2537)
);

CKINVDCx5p33_ASAP7_75t_R g2538 ( 
.A(n_449),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_702),
.Y(n_2539)
);

INVx2_ASAP7_75t_L g2540 ( 
.A(n_1127),
.Y(n_2540)
);

CKINVDCx5p33_ASAP7_75t_R g2541 ( 
.A(n_201),
.Y(n_2541)
);

CKINVDCx5p33_ASAP7_75t_R g2542 ( 
.A(n_228),
.Y(n_2542)
);

CKINVDCx5p33_ASAP7_75t_R g2543 ( 
.A(n_1356),
.Y(n_2543)
);

CKINVDCx20_ASAP7_75t_R g2544 ( 
.A(n_83),
.Y(n_2544)
);

CKINVDCx5p33_ASAP7_75t_R g2545 ( 
.A(n_396),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_624),
.Y(n_2546)
);

INVxp67_ASAP7_75t_L g2547 ( 
.A(n_333),
.Y(n_2547)
);

INVx1_ASAP7_75t_SL g2548 ( 
.A(n_627),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_609),
.Y(n_2549)
);

CKINVDCx5p33_ASAP7_75t_R g2550 ( 
.A(n_825),
.Y(n_2550)
);

CKINVDCx16_ASAP7_75t_R g2551 ( 
.A(n_1328),
.Y(n_2551)
);

CKINVDCx5p33_ASAP7_75t_R g2552 ( 
.A(n_1317),
.Y(n_2552)
);

CKINVDCx5p33_ASAP7_75t_R g2553 ( 
.A(n_633),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_1597),
.Y(n_2554)
);

BUFx6f_ASAP7_75t_L g2555 ( 
.A(n_1672),
.Y(n_2555)
);

CKINVDCx5p33_ASAP7_75t_R g2556 ( 
.A(n_1578),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_1100),
.Y(n_2557)
);

CKINVDCx5p33_ASAP7_75t_R g2558 ( 
.A(n_1040),
.Y(n_2558)
);

INVx2_ASAP7_75t_L g2559 ( 
.A(n_724),
.Y(n_2559)
);

CKINVDCx5p33_ASAP7_75t_R g2560 ( 
.A(n_450),
.Y(n_2560)
);

CKINVDCx5p33_ASAP7_75t_R g2561 ( 
.A(n_1616),
.Y(n_2561)
);

INVx1_ASAP7_75t_SL g2562 ( 
.A(n_1613),
.Y(n_2562)
);

CKINVDCx5p33_ASAP7_75t_R g2563 ( 
.A(n_28),
.Y(n_2563)
);

CKINVDCx5p33_ASAP7_75t_R g2564 ( 
.A(n_1657),
.Y(n_2564)
);

CKINVDCx5p33_ASAP7_75t_R g2565 ( 
.A(n_389),
.Y(n_2565)
);

CKINVDCx5p33_ASAP7_75t_R g2566 ( 
.A(n_1161),
.Y(n_2566)
);

CKINVDCx5p33_ASAP7_75t_R g2567 ( 
.A(n_606),
.Y(n_2567)
);

INVx2_ASAP7_75t_SL g2568 ( 
.A(n_979),
.Y(n_2568)
);

CKINVDCx5p33_ASAP7_75t_R g2569 ( 
.A(n_1084),
.Y(n_2569)
);

CKINVDCx20_ASAP7_75t_R g2570 ( 
.A(n_1342),
.Y(n_2570)
);

CKINVDCx5p33_ASAP7_75t_R g2571 ( 
.A(n_99),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_1702),
.Y(n_2572)
);

CKINVDCx20_ASAP7_75t_R g2573 ( 
.A(n_372),
.Y(n_2573)
);

INVx2_ASAP7_75t_L g2574 ( 
.A(n_1421),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_874),
.Y(n_2575)
);

CKINVDCx20_ASAP7_75t_R g2576 ( 
.A(n_475),
.Y(n_2576)
);

CKINVDCx5p33_ASAP7_75t_R g2577 ( 
.A(n_1470),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_921),
.Y(n_2578)
);

CKINVDCx5p33_ASAP7_75t_R g2579 ( 
.A(n_1705),
.Y(n_2579)
);

CKINVDCx5p33_ASAP7_75t_R g2580 ( 
.A(n_276),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_457),
.Y(n_2581)
);

CKINVDCx5p33_ASAP7_75t_R g2582 ( 
.A(n_726),
.Y(n_2582)
);

CKINVDCx5p33_ASAP7_75t_R g2583 ( 
.A(n_1027),
.Y(n_2583)
);

BUFx5_ASAP7_75t_L g2584 ( 
.A(n_311),
.Y(n_2584)
);

CKINVDCx5p33_ASAP7_75t_R g2585 ( 
.A(n_847),
.Y(n_2585)
);

BUFx6f_ASAP7_75t_L g2586 ( 
.A(n_179),
.Y(n_2586)
);

CKINVDCx5p33_ASAP7_75t_R g2587 ( 
.A(n_1349),
.Y(n_2587)
);

CKINVDCx16_ASAP7_75t_R g2588 ( 
.A(n_1303),
.Y(n_2588)
);

CKINVDCx5p33_ASAP7_75t_R g2589 ( 
.A(n_1093),
.Y(n_2589)
);

CKINVDCx5p33_ASAP7_75t_R g2590 ( 
.A(n_882),
.Y(n_2590)
);

CKINVDCx5p33_ASAP7_75t_R g2591 ( 
.A(n_944),
.Y(n_2591)
);

CKINVDCx5p33_ASAP7_75t_R g2592 ( 
.A(n_633),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_242),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_1021),
.Y(n_2594)
);

CKINVDCx5p33_ASAP7_75t_R g2595 ( 
.A(n_1293),
.Y(n_2595)
);

CKINVDCx5p33_ASAP7_75t_R g2596 ( 
.A(n_544),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_820),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_1035),
.Y(n_2598)
);

CKINVDCx5p33_ASAP7_75t_R g2599 ( 
.A(n_668),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_280),
.Y(n_2600)
);

CKINVDCx5p33_ASAP7_75t_R g2601 ( 
.A(n_63),
.Y(n_2601)
);

CKINVDCx5p33_ASAP7_75t_R g2602 ( 
.A(n_95),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_1661),
.Y(n_2603)
);

CKINVDCx20_ASAP7_75t_R g2604 ( 
.A(n_719),
.Y(n_2604)
);

CKINVDCx5p33_ASAP7_75t_R g2605 ( 
.A(n_1721),
.Y(n_2605)
);

INVx1_ASAP7_75t_SL g2606 ( 
.A(n_1499),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_1305),
.Y(n_2607)
);

CKINVDCx5p33_ASAP7_75t_R g2608 ( 
.A(n_1012),
.Y(n_2608)
);

CKINVDCx5p33_ASAP7_75t_R g2609 ( 
.A(n_566),
.Y(n_2609)
);

BUFx3_ASAP7_75t_L g2610 ( 
.A(n_564),
.Y(n_2610)
);

CKINVDCx5p33_ASAP7_75t_R g2611 ( 
.A(n_411),
.Y(n_2611)
);

CKINVDCx5p33_ASAP7_75t_R g2612 ( 
.A(n_1718),
.Y(n_2612)
);

BUFx3_ASAP7_75t_L g2613 ( 
.A(n_318),
.Y(n_2613)
);

CKINVDCx5p33_ASAP7_75t_R g2614 ( 
.A(n_1300),
.Y(n_2614)
);

CKINVDCx20_ASAP7_75t_R g2615 ( 
.A(n_1496),
.Y(n_2615)
);

CKINVDCx20_ASAP7_75t_R g2616 ( 
.A(n_1055),
.Y(n_2616)
);

CKINVDCx5p33_ASAP7_75t_R g2617 ( 
.A(n_123),
.Y(n_2617)
);

CKINVDCx16_ASAP7_75t_R g2618 ( 
.A(n_252),
.Y(n_2618)
);

CKINVDCx5p33_ASAP7_75t_R g2619 ( 
.A(n_924),
.Y(n_2619)
);

CKINVDCx5p33_ASAP7_75t_R g2620 ( 
.A(n_1424),
.Y(n_2620)
);

CKINVDCx5p33_ASAP7_75t_R g2621 ( 
.A(n_1690),
.Y(n_2621)
);

CKINVDCx5p33_ASAP7_75t_R g2622 ( 
.A(n_416),
.Y(n_2622)
);

CKINVDCx5p33_ASAP7_75t_R g2623 ( 
.A(n_891),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_1171),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_1494),
.Y(n_2625)
);

HB1xp67_ASAP7_75t_L g2626 ( 
.A(n_1386),
.Y(n_2626)
);

CKINVDCx16_ASAP7_75t_R g2627 ( 
.A(n_1487),
.Y(n_2627)
);

INVx2_ASAP7_75t_L g2628 ( 
.A(n_422),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_1692),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_1587),
.Y(n_2630)
);

CKINVDCx5p33_ASAP7_75t_R g2631 ( 
.A(n_1004),
.Y(n_2631)
);

CKINVDCx20_ASAP7_75t_R g2632 ( 
.A(n_1022),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_1033),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_136),
.Y(n_2634)
);

CKINVDCx5p33_ASAP7_75t_R g2635 ( 
.A(n_1148),
.Y(n_2635)
);

BUFx10_ASAP7_75t_L g2636 ( 
.A(n_478),
.Y(n_2636)
);

CKINVDCx5p33_ASAP7_75t_R g2637 ( 
.A(n_1458),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_987),
.Y(n_2638)
);

INVx1_ASAP7_75t_SL g2639 ( 
.A(n_642),
.Y(n_2639)
);

CKINVDCx5p33_ASAP7_75t_R g2640 ( 
.A(n_426),
.Y(n_2640)
);

CKINVDCx5p33_ASAP7_75t_R g2641 ( 
.A(n_587),
.Y(n_2641)
);

CKINVDCx5p33_ASAP7_75t_R g2642 ( 
.A(n_25),
.Y(n_2642)
);

CKINVDCx5p33_ASAP7_75t_R g2643 ( 
.A(n_1590),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_1058),
.Y(n_2644)
);

INVx1_ASAP7_75t_SL g2645 ( 
.A(n_1525),
.Y(n_2645)
);

INVx3_ASAP7_75t_L g2646 ( 
.A(n_846),
.Y(n_2646)
);

CKINVDCx5p33_ASAP7_75t_R g2647 ( 
.A(n_1724),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_184),
.Y(n_2648)
);

CKINVDCx5p33_ASAP7_75t_R g2649 ( 
.A(n_1714),
.Y(n_2649)
);

CKINVDCx5p33_ASAP7_75t_R g2650 ( 
.A(n_1609),
.Y(n_2650)
);

CKINVDCx5p33_ASAP7_75t_R g2651 ( 
.A(n_895),
.Y(n_2651)
);

INVx2_ASAP7_75t_SL g2652 ( 
.A(n_282),
.Y(n_2652)
);

HB1xp67_ASAP7_75t_L g2653 ( 
.A(n_790),
.Y(n_2653)
);

CKINVDCx5p33_ASAP7_75t_R g2654 ( 
.A(n_1698),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_1010),
.Y(n_2655)
);

INVx2_ASAP7_75t_SL g2656 ( 
.A(n_1512),
.Y(n_2656)
);

CKINVDCx5p33_ASAP7_75t_R g2657 ( 
.A(n_1147),
.Y(n_2657)
);

CKINVDCx5p33_ASAP7_75t_R g2658 ( 
.A(n_1524),
.Y(n_2658)
);

CKINVDCx5p33_ASAP7_75t_R g2659 ( 
.A(n_637),
.Y(n_2659)
);

CKINVDCx5p33_ASAP7_75t_R g2660 ( 
.A(n_137),
.Y(n_2660)
);

CKINVDCx5p33_ASAP7_75t_R g2661 ( 
.A(n_103),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_757),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_931),
.Y(n_2663)
);

CKINVDCx5p33_ASAP7_75t_R g2664 ( 
.A(n_1423),
.Y(n_2664)
);

INVx2_ASAP7_75t_L g2665 ( 
.A(n_1456),
.Y(n_2665)
);

CKINVDCx5p33_ASAP7_75t_R g2666 ( 
.A(n_587),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_284),
.Y(n_2667)
);

CKINVDCx5p33_ASAP7_75t_R g2668 ( 
.A(n_1580),
.Y(n_2668)
);

CKINVDCx5p33_ASAP7_75t_R g2669 ( 
.A(n_688),
.Y(n_2669)
);

CKINVDCx5p33_ASAP7_75t_R g2670 ( 
.A(n_26),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_487),
.Y(n_2671)
);

CKINVDCx5p33_ASAP7_75t_R g2672 ( 
.A(n_383),
.Y(n_2672)
);

CKINVDCx5p33_ASAP7_75t_R g2673 ( 
.A(n_88),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_1732),
.Y(n_2674)
);

BUFx3_ASAP7_75t_L g2675 ( 
.A(n_281),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_379),
.Y(n_2676)
);

CKINVDCx5p33_ASAP7_75t_R g2677 ( 
.A(n_222),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_1640),
.Y(n_2678)
);

CKINVDCx5p33_ASAP7_75t_R g2679 ( 
.A(n_805),
.Y(n_2679)
);

CKINVDCx20_ASAP7_75t_R g2680 ( 
.A(n_1468),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_226),
.Y(n_2681)
);

CKINVDCx5p33_ASAP7_75t_R g2682 ( 
.A(n_1492),
.Y(n_2682)
);

CKINVDCx5p33_ASAP7_75t_R g2683 ( 
.A(n_79),
.Y(n_2683)
);

INVx2_ASAP7_75t_L g2684 ( 
.A(n_29),
.Y(n_2684)
);

INVx2_ASAP7_75t_SL g2685 ( 
.A(n_1052),
.Y(n_2685)
);

CKINVDCx5p33_ASAP7_75t_R g2686 ( 
.A(n_1014),
.Y(n_2686)
);

BUFx6f_ASAP7_75t_L g2687 ( 
.A(n_434),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_605),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_1173),
.Y(n_2689)
);

INVx2_ASAP7_75t_L g2690 ( 
.A(n_419),
.Y(n_2690)
);

CKINVDCx5p33_ASAP7_75t_R g2691 ( 
.A(n_1610),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_1712),
.Y(n_2692)
);

BUFx2_ASAP7_75t_L g2693 ( 
.A(n_858),
.Y(n_2693)
);

BUFx3_ASAP7_75t_L g2694 ( 
.A(n_779),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_1514),
.Y(n_2695)
);

CKINVDCx5p33_ASAP7_75t_R g2696 ( 
.A(n_993),
.Y(n_2696)
);

CKINVDCx5p33_ASAP7_75t_R g2697 ( 
.A(n_1504),
.Y(n_2697)
);

CKINVDCx5p33_ASAP7_75t_R g2698 ( 
.A(n_1709),
.Y(n_2698)
);

CKINVDCx5p33_ASAP7_75t_R g2699 ( 
.A(n_978),
.Y(n_2699)
);

CKINVDCx20_ASAP7_75t_R g2700 ( 
.A(n_778),
.Y(n_2700)
);

CKINVDCx5p33_ASAP7_75t_R g2701 ( 
.A(n_1667),
.Y(n_2701)
);

CKINVDCx20_ASAP7_75t_R g2702 ( 
.A(n_941),
.Y(n_2702)
);

CKINVDCx5p33_ASAP7_75t_R g2703 ( 
.A(n_78),
.Y(n_2703)
);

CKINVDCx5p33_ASAP7_75t_R g2704 ( 
.A(n_1449),
.Y(n_2704)
);

CKINVDCx20_ASAP7_75t_R g2705 ( 
.A(n_1668),
.Y(n_2705)
);

INVx2_ASAP7_75t_SL g2706 ( 
.A(n_128),
.Y(n_2706)
);

CKINVDCx5p33_ASAP7_75t_R g2707 ( 
.A(n_1225),
.Y(n_2707)
);

CKINVDCx20_ASAP7_75t_R g2708 ( 
.A(n_1023),
.Y(n_2708)
);

BUFx6f_ASAP7_75t_L g2709 ( 
.A(n_1153),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_869),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_98),
.Y(n_2711)
);

CKINVDCx5p33_ASAP7_75t_R g2712 ( 
.A(n_623),
.Y(n_2712)
);

CKINVDCx20_ASAP7_75t_R g2713 ( 
.A(n_1323),
.Y(n_2713)
);

CKINVDCx5p33_ASAP7_75t_R g2714 ( 
.A(n_1676),
.Y(n_2714)
);

INVx1_ASAP7_75t_SL g2715 ( 
.A(n_155),
.Y(n_2715)
);

CKINVDCx5p33_ASAP7_75t_R g2716 ( 
.A(n_1552),
.Y(n_2716)
);

CKINVDCx5p33_ASAP7_75t_R g2717 ( 
.A(n_115),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_839),
.Y(n_2718)
);

CKINVDCx5p33_ASAP7_75t_R g2719 ( 
.A(n_1675),
.Y(n_2719)
);

CKINVDCx20_ASAP7_75t_R g2720 ( 
.A(n_1098),
.Y(n_2720)
);

CKINVDCx5p33_ASAP7_75t_R g2721 ( 
.A(n_132),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_1392),
.Y(n_2722)
);

CKINVDCx5p33_ASAP7_75t_R g2723 ( 
.A(n_519),
.Y(n_2723)
);

CKINVDCx20_ASAP7_75t_R g2724 ( 
.A(n_1045),
.Y(n_2724)
);

CKINVDCx5p33_ASAP7_75t_R g2725 ( 
.A(n_572),
.Y(n_2725)
);

CKINVDCx5p33_ASAP7_75t_R g2726 ( 
.A(n_608),
.Y(n_2726)
);

INVx2_ASAP7_75t_SL g2727 ( 
.A(n_1555),
.Y(n_2727)
);

INVx2_ASAP7_75t_L g2728 ( 
.A(n_1485),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_998),
.Y(n_2729)
);

BUFx6f_ASAP7_75t_L g2730 ( 
.A(n_1000),
.Y(n_2730)
);

CKINVDCx5p33_ASAP7_75t_R g2731 ( 
.A(n_1641),
.Y(n_2731)
);

CKINVDCx14_ASAP7_75t_R g2732 ( 
.A(n_569),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_865),
.Y(n_2733)
);

INVx1_ASAP7_75t_SL g2734 ( 
.A(n_1582),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_1652),
.Y(n_2735)
);

CKINVDCx16_ASAP7_75t_R g2736 ( 
.A(n_1699),
.Y(n_2736)
);

BUFx2_ASAP7_75t_L g2737 ( 
.A(n_702),
.Y(n_2737)
);

BUFx8_ASAP7_75t_SL g2738 ( 
.A(n_87),
.Y(n_2738)
);

BUFx3_ASAP7_75t_L g2739 ( 
.A(n_878),
.Y(n_2739)
);

CKINVDCx5p33_ASAP7_75t_R g2740 ( 
.A(n_600),
.Y(n_2740)
);

CKINVDCx5p33_ASAP7_75t_R g2741 ( 
.A(n_753),
.Y(n_2741)
);

CKINVDCx5p33_ASAP7_75t_R g2742 ( 
.A(n_252),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_1528),
.Y(n_2743)
);

CKINVDCx5p33_ASAP7_75t_R g2744 ( 
.A(n_1660),
.Y(n_2744)
);

BUFx3_ASAP7_75t_L g2745 ( 
.A(n_1684),
.Y(n_2745)
);

CKINVDCx5p33_ASAP7_75t_R g2746 ( 
.A(n_222),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_1495),
.Y(n_2747)
);

CKINVDCx5p33_ASAP7_75t_R g2748 ( 
.A(n_441),
.Y(n_2748)
);

CKINVDCx5p33_ASAP7_75t_R g2749 ( 
.A(n_1383),
.Y(n_2749)
);

CKINVDCx5p33_ASAP7_75t_R g2750 ( 
.A(n_918),
.Y(n_2750)
);

CKINVDCx5p33_ASAP7_75t_R g2751 ( 
.A(n_1261),
.Y(n_2751)
);

CKINVDCx20_ASAP7_75t_R g2752 ( 
.A(n_48),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_173),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_1088),
.Y(n_2754)
);

CKINVDCx5p33_ASAP7_75t_R g2755 ( 
.A(n_1588),
.Y(n_2755)
);

BUFx3_ASAP7_75t_L g2756 ( 
.A(n_1624),
.Y(n_2756)
);

CKINVDCx5p33_ASAP7_75t_R g2757 ( 
.A(n_196),
.Y(n_2757)
);

BUFx3_ASAP7_75t_L g2758 ( 
.A(n_1346),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_1643),
.Y(n_2759)
);

CKINVDCx20_ASAP7_75t_R g2760 ( 
.A(n_1571),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_1254),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_203),
.Y(n_2762)
);

CKINVDCx5p33_ASAP7_75t_R g2763 ( 
.A(n_299),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_549),
.Y(n_2764)
);

CKINVDCx5p33_ASAP7_75t_R g2765 ( 
.A(n_290),
.Y(n_2765)
);

INVx2_ASAP7_75t_SL g2766 ( 
.A(n_1070),
.Y(n_2766)
);

CKINVDCx5p33_ASAP7_75t_R g2767 ( 
.A(n_1619),
.Y(n_2767)
);

BUFx3_ASAP7_75t_L g2768 ( 
.A(n_80),
.Y(n_2768)
);

CKINVDCx5p33_ASAP7_75t_R g2769 ( 
.A(n_782),
.Y(n_2769)
);

CKINVDCx5p33_ASAP7_75t_R g2770 ( 
.A(n_883),
.Y(n_2770)
);

INVx2_ASAP7_75t_L g2771 ( 
.A(n_994),
.Y(n_2771)
);

CKINVDCx5p33_ASAP7_75t_R g2772 ( 
.A(n_1628),
.Y(n_2772)
);

CKINVDCx5p33_ASAP7_75t_R g2773 ( 
.A(n_815),
.Y(n_2773)
);

CKINVDCx5p33_ASAP7_75t_R g2774 ( 
.A(n_1024),
.Y(n_2774)
);

CKINVDCx5p33_ASAP7_75t_R g2775 ( 
.A(n_1634),
.Y(n_2775)
);

CKINVDCx20_ASAP7_75t_R g2776 ( 
.A(n_1333),
.Y(n_2776)
);

CKINVDCx16_ASAP7_75t_R g2777 ( 
.A(n_1013),
.Y(n_2777)
);

CKINVDCx5p33_ASAP7_75t_R g2778 ( 
.A(n_949),
.Y(n_2778)
);

CKINVDCx5p33_ASAP7_75t_R g2779 ( 
.A(n_202),
.Y(n_2779)
);

CKINVDCx5p33_ASAP7_75t_R g2780 ( 
.A(n_1716),
.Y(n_2780)
);

BUFx3_ASAP7_75t_L g2781 ( 
.A(n_427),
.Y(n_2781)
);

CKINVDCx5p33_ASAP7_75t_R g2782 ( 
.A(n_127),
.Y(n_2782)
);

CKINVDCx5p33_ASAP7_75t_R g2783 ( 
.A(n_1480),
.Y(n_2783)
);

INVx3_ASAP7_75t_L g2784 ( 
.A(n_1092),
.Y(n_2784)
);

CKINVDCx5p33_ASAP7_75t_R g2785 ( 
.A(n_1101),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_543),
.Y(n_2786)
);

BUFx6f_ASAP7_75t_L g2787 ( 
.A(n_1564),
.Y(n_2787)
);

CKINVDCx5p33_ASAP7_75t_R g2788 ( 
.A(n_717),
.Y(n_2788)
);

CKINVDCx5p33_ASAP7_75t_R g2789 ( 
.A(n_1680),
.Y(n_2789)
);

BUFx2_ASAP7_75t_L g2790 ( 
.A(n_70),
.Y(n_2790)
);

CKINVDCx5p33_ASAP7_75t_R g2791 ( 
.A(n_862),
.Y(n_2791)
);

CKINVDCx5p33_ASAP7_75t_R g2792 ( 
.A(n_1002),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_914),
.Y(n_2793)
);

BUFx10_ASAP7_75t_L g2794 ( 
.A(n_1042),
.Y(n_2794)
);

CKINVDCx20_ASAP7_75t_R g2795 ( 
.A(n_349),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_450),
.Y(n_2796)
);

CKINVDCx5p33_ASAP7_75t_R g2797 ( 
.A(n_284),
.Y(n_2797)
);

CKINVDCx5p33_ASAP7_75t_R g2798 ( 
.A(n_1096),
.Y(n_2798)
);

CKINVDCx5p33_ASAP7_75t_R g2799 ( 
.A(n_682),
.Y(n_2799)
);

INVx2_ASAP7_75t_L g2800 ( 
.A(n_438),
.Y(n_2800)
);

CKINVDCx20_ASAP7_75t_R g2801 ( 
.A(n_1531),
.Y(n_2801)
);

CKINVDCx5p33_ASAP7_75t_R g2802 ( 
.A(n_1041),
.Y(n_2802)
);

BUFx6f_ASAP7_75t_L g2803 ( 
.A(n_901),
.Y(n_2803)
);

CKINVDCx5p33_ASAP7_75t_R g2804 ( 
.A(n_11),
.Y(n_2804)
);

CKINVDCx5p33_ASAP7_75t_R g2805 ( 
.A(n_1029),
.Y(n_2805)
);

INVx1_ASAP7_75t_SL g2806 ( 
.A(n_195),
.Y(n_2806)
);

CKINVDCx5p33_ASAP7_75t_R g2807 ( 
.A(n_1431),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_1009),
.Y(n_2808)
);

CKINVDCx5p33_ASAP7_75t_R g2809 ( 
.A(n_370),
.Y(n_2809)
);

CKINVDCx5p33_ASAP7_75t_R g2810 ( 
.A(n_142),
.Y(n_2810)
);

CKINVDCx5p33_ASAP7_75t_R g2811 ( 
.A(n_1687),
.Y(n_2811)
);

CKINVDCx5p33_ASAP7_75t_R g2812 ( 
.A(n_756),
.Y(n_2812)
);

CKINVDCx20_ASAP7_75t_R g2813 ( 
.A(n_312),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_265),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_896),
.Y(n_2815)
);

BUFx5_ASAP7_75t_L g2816 ( 
.A(n_875),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_1568),
.Y(n_2817)
);

CKINVDCx5p33_ASAP7_75t_R g2818 ( 
.A(n_2194),
.Y(n_2818)
);

HB1xp67_ASAP7_75t_L g2819 ( 
.A(n_1880),
.Y(n_2819)
);

INVxp67_ASAP7_75t_SL g2820 ( 
.A(n_1778),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2259),
.Y(n_2821)
);

INVxp33_ASAP7_75t_L g2822 ( 
.A(n_1817),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2259),
.Y(n_2823)
);

INVxp67_ASAP7_75t_SL g2824 ( 
.A(n_2199),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2259),
.Y(n_2825)
);

INVxp67_ASAP7_75t_L g2826 ( 
.A(n_1802),
.Y(n_2826)
);

CKINVDCx20_ASAP7_75t_R g2827 ( 
.A(n_1793),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2259),
.Y(n_2828)
);

CKINVDCx20_ASAP7_75t_R g2829 ( 
.A(n_1796),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2259),
.Y(n_2830)
);

INVxp67_ASAP7_75t_SL g2831 ( 
.A(n_2205),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2584),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2584),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2584),
.Y(n_2834)
);

INVxp67_ASAP7_75t_L g2835 ( 
.A(n_1836),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2584),
.Y(n_2836)
);

INVxp67_ASAP7_75t_SL g2837 ( 
.A(n_2626),
.Y(n_2837)
);

INVxp67_ASAP7_75t_SL g2838 ( 
.A(n_1741),
.Y(n_2838)
);

CKINVDCx16_ASAP7_75t_R g2839 ( 
.A(n_1885),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2584),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2816),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2816),
.Y(n_2842)
);

INVxp67_ASAP7_75t_SL g2843 ( 
.A(n_1927),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2816),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2816),
.Y(n_2845)
);

CKINVDCx5p33_ASAP7_75t_R g2846 ( 
.A(n_2283),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2816),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_1739),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_1739),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2646),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2646),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2041),
.Y(n_2852)
);

INVxp33_ASAP7_75t_SL g2853 ( 
.A(n_2295),
.Y(n_2853)
);

CKINVDCx16_ASAP7_75t_R g2854 ( 
.A(n_1944),
.Y(n_2854)
);

CKINVDCx5p33_ASAP7_75t_R g2855 ( 
.A(n_2501),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2041),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2041),
.Y(n_2857)
);

INVxp67_ASAP7_75t_L g2858 ( 
.A(n_2306),
.Y(n_2858)
);

INVx3_ASAP7_75t_L g2859 ( 
.A(n_2115),
.Y(n_2859)
);

INVxp33_ASAP7_75t_L g2860 ( 
.A(n_2653),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2115),
.Y(n_2861)
);

CKINVDCx5p33_ASAP7_75t_R g2862 ( 
.A(n_2738),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2115),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2245),
.Y(n_2864)
);

BUFx3_ASAP7_75t_L g2865 ( 
.A(n_1822),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2245),
.Y(n_2866)
);

CKINVDCx16_ASAP7_75t_R g2867 ( 
.A(n_2014),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2245),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2392),
.Y(n_2869)
);

INVxp67_ASAP7_75t_L g2870 ( 
.A(n_2693),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2392),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2392),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2586),
.Y(n_2873)
);

BUFx2_ASAP7_75t_L g2874 ( 
.A(n_2737),
.Y(n_2874)
);

INVxp67_ASAP7_75t_SL g2875 ( 
.A(n_2784),
.Y(n_2875)
);

HB1xp67_ASAP7_75t_L g2876 ( 
.A(n_2132),
.Y(n_2876)
);

INVxp67_ASAP7_75t_SL g2877 ( 
.A(n_2784),
.Y(n_2877)
);

BUFx3_ASAP7_75t_L g2878 ( 
.A(n_1822),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2586),
.Y(n_2879)
);

INVxp67_ASAP7_75t_SL g2880 ( 
.A(n_1763),
.Y(n_2880)
);

INVxp33_ASAP7_75t_L g2881 ( 
.A(n_2790),
.Y(n_2881)
);

INVxp67_ASAP7_75t_SL g2882 ( 
.A(n_1894),
.Y(n_2882)
);

INVxp67_ASAP7_75t_L g2883 ( 
.A(n_1764),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2586),
.Y(n_2884)
);

INVxp67_ASAP7_75t_SL g2885 ( 
.A(n_1953),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2687),
.Y(n_2886)
);

INVx2_ASAP7_75t_L g2887 ( 
.A(n_2803),
.Y(n_2887)
);

INVxp67_ASAP7_75t_SL g2888 ( 
.A(n_1968),
.Y(n_2888)
);

INVxp33_ASAP7_75t_SL g2889 ( 
.A(n_1747),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2687),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2687),
.Y(n_2891)
);

CKINVDCx5p33_ASAP7_75t_R g2892 ( 
.A(n_1738),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2730),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2730),
.Y(n_2894)
);

BUFx8_ASAP7_75t_SL g2895 ( 
.A(n_1749),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2730),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2803),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2803),
.Y(n_2898)
);

BUFx10_ASAP7_75t_L g2899 ( 
.A(n_1753),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_1744),
.Y(n_2900)
);

CKINVDCx14_ASAP7_75t_R g2901 ( 
.A(n_2425),
.Y(n_2901)
);

NOR2xp67_ASAP7_75t_L g2902 ( 
.A(n_1879),
.B(n_0),
.Y(n_2902)
);

INVx2_ASAP7_75t_L g2903 ( 
.A(n_1998),
.Y(n_2903)
);

CKINVDCx5p33_ASAP7_75t_R g2904 ( 
.A(n_1740),
.Y(n_2904)
);

INVxp67_ASAP7_75t_SL g2905 ( 
.A(n_1989),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_1998),
.Y(n_2906)
);

INVx2_ASAP7_75t_L g2907 ( 
.A(n_1998),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_1835),
.Y(n_2908)
);

INVxp67_ASAP7_75t_SL g2909 ( 
.A(n_2037),
.Y(n_2909)
);

CKINVDCx14_ASAP7_75t_R g2910 ( 
.A(n_2732),
.Y(n_2910)
);

NOR2xp67_ASAP7_75t_L g2911 ( 
.A(n_2196),
.B(n_0),
.Y(n_2911)
);

INVx2_ASAP7_75t_L g2912 ( 
.A(n_1998),
.Y(n_2912)
);

CKINVDCx5p33_ASAP7_75t_R g2913 ( 
.A(n_1742),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_1873),
.Y(n_2914)
);

BUFx6f_ASAP7_75t_L g2915 ( 
.A(n_1891),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_1984),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2038),
.Y(n_2917)
);

INVxp67_ASAP7_75t_SL g2918 ( 
.A(n_2377),
.Y(n_2918)
);

BUFx8_ASAP7_75t_SL g2919 ( 
.A(n_1786),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2133),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2208),
.Y(n_2921)
);

CKINVDCx16_ASAP7_75t_R g2922 ( 
.A(n_2149),
.Y(n_2922)
);

INVx2_ASAP7_75t_L g2923 ( 
.A(n_1998),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2269),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2315),
.Y(n_2925)
);

CKINVDCx5p33_ASAP7_75t_R g2926 ( 
.A(n_1746),
.Y(n_2926)
);

INVxp67_ASAP7_75t_SL g2927 ( 
.A(n_2510),
.Y(n_2927)
);

INVxp67_ASAP7_75t_SL g2928 ( 
.A(n_2745),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2373),
.Y(n_2929)
);

INVxp67_ASAP7_75t_SL g2930 ( 
.A(n_2756),
.Y(n_2930)
);

INVxp33_ASAP7_75t_SL g2931 ( 
.A(n_1755),
.Y(n_2931)
);

CKINVDCx20_ASAP7_75t_R g2932 ( 
.A(n_1863),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2380),
.Y(n_2933)
);

INVxp67_ASAP7_75t_L g2934 ( 
.A(n_1764),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2401),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2458),
.Y(n_2936)
);

BUFx2_ASAP7_75t_SL g2937 ( 
.A(n_1965),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2499),
.Y(n_2938)
);

CKINVDCx5p33_ASAP7_75t_R g2939 ( 
.A(n_1750),
.Y(n_2939)
);

BUFx3_ASAP7_75t_L g2940 ( 
.A(n_2758),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2511),
.Y(n_2941)
);

INVxp67_ASAP7_75t_L g2942 ( 
.A(n_1783),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2522),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2610),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2613),
.Y(n_2945)
);

CKINVDCx5p33_ASAP7_75t_R g2946 ( 
.A(n_1751),
.Y(n_2946)
);

INVx1_ASAP7_75t_L g2947 ( 
.A(n_2675),
.Y(n_2947)
);

INVxp33_ASAP7_75t_L g2948 ( 
.A(n_1743),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2694),
.Y(n_2949)
);

INVxp33_ASAP7_75t_SL g2950 ( 
.A(n_1760),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2739),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2768),
.Y(n_2952)
);

BUFx5_ASAP7_75t_L g2953 ( 
.A(n_1748),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2781),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2814),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2815),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_1745),
.Y(n_2957)
);

INVxp67_ASAP7_75t_L g2958 ( 
.A(n_1783),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_1766),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_1774),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_1782),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2808),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_1785),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_1791),
.Y(n_2964)
);

INVxp67_ASAP7_75t_SL g2965 ( 
.A(n_1871),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_1815),
.Y(n_2966)
);

INVxp67_ASAP7_75t_SL g2967 ( 
.A(n_2120),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_1833),
.Y(n_2968)
);

BUFx3_ASAP7_75t_L g2969 ( 
.A(n_1754),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_1838),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_1842),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_1849),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_1852),
.Y(n_2973)
);

BUFx6f_ASAP7_75t_L g2974 ( 
.A(n_1891),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_1853),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_1892),
.Y(n_2976)
);

BUFx6f_ASAP7_75t_L g2977 ( 
.A(n_1891),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_1900),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_1901),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_1923),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_1925),
.Y(n_2981)
);

INVxp67_ASAP7_75t_SL g2982 ( 
.A(n_1759),
.Y(n_2982)
);

INVxp33_ASAP7_75t_L g2983 ( 
.A(n_1934),
.Y(n_2983)
);

CKINVDCx20_ASAP7_75t_R g2984 ( 
.A(n_1966),
.Y(n_2984)
);

CKINVDCx5p33_ASAP7_75t_R g2985 ( 
.A(n_1756),
.Y(n_2985)
);

HB1xp67_ASAP7_75t_L g2986 ( 
.A(n_2190),
.Y(n_2986)
);

CKINVDCx5p33_ASAP7_75t_R g2987 ( 
.A(n_1757),
.Y(n_2987)
);

CKINVDCx16_ASAP7_75t_R g2988 ( 
.A(n_2242),
.Y(n_2988)
);

CKINVDCx14_ASAP7_75t_R g2989 ( 
.A(n_1902),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_1958),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_1970),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_1971),
.Y(n_2992)
);

INVxp67_ASAP7_75t_SL g2993 ( 
.A(n_1787),
.Y(n_2993)
);

INVx2_ASAP7_75t_L g2994 ( 
.A(n_2284),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_1974),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_1980),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_1987),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_1992),
.Y(n_2998)
);

INVxp67_ASAP7_75t_SL g2999 ( 
.A(n_1789),
.Y(n_2999)
);

CKINVDCx5p33_ASAP7_75t_R g3000 ( 
.A(n_1758),
.Y(n_3000)
);

CKINVDCx20_ASAP7_75t_R g3001 ( 
.A(n_1977),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_1993),
.Y(n_3002)
);

INVxp33_ASAP7_75t_SL g3003 ( 
.A(n_1761),
.Y(n_3003)
);

INVxp67_ASAP7_75t_SL g3004 ( 
.A(n_1795),
.Y(n_3004)
);

INVxp67_ASAP7_75t_SL g3005 ( 
.A(n_1799),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_1999),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2010),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2022),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2023),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2044),
.Y(n_3010)
);

CKINVDCx5p33_ASAP7_75t_R g3011 ( 
.A(n_1768),
.Y(n_3011)
);

INVx2_ASAP7_75t_SL g3012 ( 
.A(n_2069),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2047),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2063),
.Y(n_3014)
);

CKINVDCx5p33_ASAP7_75t_R g3015 ( 
.A(n_1770),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2064),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2072),
.Y(n_3017)
);

INVx1_ASAP7_75t_SL g3018 ( 
.A(n_1855),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2074),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2082),
.Y(n_3020)
);

INVxp67_ASAP7_75t_SL g3021 ( 
.A(n_1803),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2085),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2095),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2099),
.Y(n_3024)
);

INVxp33_ASAP7_75t_L g3025 ( 
.A(n_2108),
.Y(n_3025)
);

INVxp33_ASAP7_75t_L g3026 ( 
.A(n_2109),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2111),
.Y(n_3027)
);

INVx2_ASAP7_75t_L g3028 ( 
.A(n_2284),
.Y(n_3028)
);

CKINVDCx20_ASAP7_75t_R g3029 ( 
.A(n_1983),
.Y(n_3029)
);

INVxp33_ASAP7_75t_SL g3030 ( 
.A(n_1762),
.Y(n_3030)
);

INVxp33_ASAP7_75t_SL g3031 ( 
.A(n_1765),
.Y(n_3031)
);

CKINVDCx5p33_ASAP7_75t_R g3032 ( 
.A(n_1773),
.Y(n_3032)
);

INVxp67_ASAP7_75t_SL g3033 ( 
.A(n_1807),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2124),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2134),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2147),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_2157),
.Y(n_3037)
);

CKINVDCx5p33_ASAP7_75t_R g3038 ( 
.A(n_1776),
.Y(n_3038)
);

CKINVDCx5p33_ASAP7_75t_R g3039 ( 
.A(n_1777),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2167),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2173),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2224),
.Y(n_3042)
);

INVxp33_ASAP7_75t_SL g3043 ( 
.A(n_1769),
.Y(n_3043)
);

INVx2_ASAP7_75t_L g3044 ( 
.A(n_2284),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2227),
.Y(n_3045)
);

CKINVDCx20_ASAP7_75t_R g3046 ( 
.A(n_2040),
.Y(n_3046)
);

CKINVDCx20_ASAP7_75t_R g3047 ( 
.A(n_2801),
.Y(n_3047)
);

INVxp67_ASAP7_75t_SL g3048 ( 
.A(n_1818),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_2230),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2233),
.Y(n_3050)
);

CKINVDCx5p33_ASAP7_75t_R g3051 ( 
.A(n_1784),
.Y(n_3051)
);

CKINVDCx5p33_ASAP7_75t_R g3052 ( 
.A(n_1788),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2243),
.Y(n_3053)
);

CKINVDCx5p33_ASAP7_75t_R g3054 ( 
.A(n_1790),
.Y(n_3054)
);

INVxp67_ASAP7_75t_L g3055 ( 
.A(n_2069),
.Y(n_3055)
);

CKINVDCx5p33_ASAP7_75t_R g3056 ( 
.A(n_1798),
.Y(n_3056)
);

INVxp67_ASAP7_75t_SL g3057 ( 
.A(n_1825),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_2262),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2263),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_2264),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2271),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_2272),
.Y(n_3062)
);

CKINVDCx16_ASAP7_75t_R g3063 ( 
.A(n_2381),
.Y(n_3063)
);

BUFx2_ASAP7_75t_L g3064 ( 
.A(n_2435),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2277),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2291),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2304),
.Y(n_3067)
);

INVx2_ASAP7_75t_L g3068 ( 
.A(n_2284),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2310),
.Y(n_3069)
);

CKINVDCx16_ASAP7_75t_R g3070 ( 
.A(n_2446),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2318),
.Y(n_3071)
);

BUFx6f_ASAP7_75t_L g3072 ( 
.A(n_1981),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2321),
.Y(n_3073)
);

CKINVDCx16_ASAP7_75t_R g3074 ( 
.A(n_2618),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_2326),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2333),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2337),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2343),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2887),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2852),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2856),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2892),
.B(n_1991),
.Y(n_3082)
);

INVx2_ASAP7_75t_L g3083 ( 
.A(n_2915),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_L g3084 ( 
.A(n_2904),
.B(n_2002),
.Y(n_3084)
);

AOI22xp5_ASAP7_75t_L g3085 ( 
.A1(n_2853),
.A2(n_2223),
.B1(n_2355),
.B2(n_2169),
.Y(n_3085)
);

INVx5_ASAP7_75t_L g3086 ( 
.A(n_2899),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2857),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2861),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_2863),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2864),
.Y(n_3090)
);

AND2x2_ASAP7_75t_L g3091 ( 
.A(n_2901),
.B(n_2777),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2866),
.Y(n_3092)
);

CKINVDCx5p33_ASAP7_75t_R g3093 ( 
.A(n_2913),
.Y(n_3093)
);

OAI22xp5_ASAP7_75t_L g3094 ( 
.A1(n_2838),
.A2(n_2056),
.B1(n_2191),
.B2(n_1809),
.Y(n_3094)
);

AND2x4_ASAP7_75t_L g3095 ( 
.A(n_2969),
.B(n_1920),
.Y(n_3095)
);

AND2x2_ASAP7_75t_L g3096 ( 
.A(n_2910),
.B(n_2254),
.Y(n_3096)
);

BUFx2_ASAP7_75t_L g3097 ( 
.A(n_2865),
.Y(n_3097)
);

INVx2_ASAP7_75t_L g3098 ( 
.A(n_2915),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2868),
.Y(n_3099)
);

INVx3_ASAP7_75t_L g3100 ( 
.A(n_2859),
.Y(n_3100)
);

AND2x2_ASAP7_75t_L g3101 ( 
.A(n_2989),
.B(n_2393),
.Y(n_3101)
);

AND2x6_ASAP7_75t_L g3102 ( 
.A(n_2878),
.B(n_1752),
.Y(n_3102)
);

BUFx6f_ASAP7_75t_L g3103 ( 
.A(n_2915),
.Y(n_3103)
);

BUFx2_ASAP7_75t_L g3104 ( 
.A(n_2819),
.Y(n_3104)
);

INVx3_ASAP7_75t_L g3105 ( 
.A(n_2859),
.Y(n_3105)
);

AND2x2_ASAP7_75t_L g3106 ( 
.A(n_2880),
.B(n_2551),
.Y(n_3106)
);

BUFx6f_ASAP7_75t_L g3107 ( 
.A(n_2974),
.Y(n_3107)
);

AND2x6_ASAP7_75t_L g3108 ( 
.A(n_2900),
.B(n_1812),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_2869),
.Y(n_3109)
);

OAI22x1_ASAP7_75t_L g3110 ( 
.A1(n_2874),
.A2(n_1906),
.B1(n_2036),
.B2(n_1935),
.Y(n_3110)
);

AND2x4_ASAP7_75t_L g3111 ( 
.A(n_2843),
.B(n_2882),
.Y(n_3111)
);

AND2x4_ASAP7_75t_L g3112 ( 
.A(n_2885),
.B(n_2076),
.Y(n_3112)
);

BUFx2_ASAP7_75t_L g3113 ( 
.A(n_2876),
.Y(n_3113)
);

INVx2_ASAP7_75t_L g3114 ( 
.A(n_2974),
.Y(n_3114)
);

BUFx6f_ASAP7_75t_L g3115 ( 
.A(n_2974),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_2871),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_2872),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_L g3118 ( 
.A(n_2926),
.B(n_2055),
.Y(n_3118)
);

INVx3_ASAP7_75t_L g3119 ( 
.A(n_2940),
.Y(n_3119)
);

INVx2_ASAP7_75t_L g3120 ( 
.A(n_2977),
.Y(n_3120)
);

OA21x2_ASAP7_75t_L g3121 ( 
.A1(n_2821),
.A2(n_2825),
.B(n_2823),
.Y(n_3121)
);

BUFx6f_ASAP7_75t_L g3122 ( 
.A(n_2977),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_2873),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_2879),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_L g3125 ( 
.A(n_2939),
.B(n_2141),
.Y(n_3125)
);

HB1xp67_ASAP7_75t_L g3126 ( 
.A(n_2986),
.Y(n_3126)
);

AND2x4_ASAP7_75t_L g3127 ( 
.A(n_2888),
.B(n_2091),
.Y(n_3127)
);

INVx3_ASAP7_75t_L g3128 ( 
.A(n_2977),
.Y(n_3128)
);

BUFx6f_ASAP7_75t_L g3129 ( 
.A(n_3072),
.Y(n_3129)
);

INVx2_ASAP7_75t_L g3130 ( 
.A(n_3072),
.Y(n_3130)
);

BUFx12f_ASAP7_75t_L g3131 ( 
.A(n_2818),
.Y(n_3131)
);

BUFx6f_ASAP7_75t_L g3132 ( 
.A(n_3072),
.Y(n_3132)
);

AND2x2_ASAP7_75t_L g3133 ( 
.A(n_2905),
.B(n_2588),
.Y(n_3133)
);

INVxp67_ASAP7_75t_L g3134 ( 
.A(n_3064),
.Y(n_3134)
);

INVx4_ASAP7_75t_L g3135 ( 
.A(n_2946),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_2884),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2886),
.Y(n_3137)
);

BUFx6f_ASAP7_75t_L g3138 ( 
.A(n_2890),
.Y(n_3138)
);

INVx2_ASAP7_75t_SL g3139 ( 
.A(n_2899),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2891),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_2893),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_2894),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_2896),
.Y(n_3143)
);

HB1xp67_ASAP7_75t_L g3144 ( 
.A(n_2839),
.Y(n_3144)
);

CKINVDCx5p33_ASAP7_75t_R g3145 ( 
.A(n_2985),
.Y(n_3145)
);

OA21x2_ASAP7_75t_L g3146 ( 
.A1(n_2828),
.A2(n_1830),
.B(n_1827),
.Y(n_3146)
);

BUFx12f_ASAP7_75t_L g3147 ( 
.A(n_2846),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_2897),
.Y(n_3148)
);

CKINVDCx5p33_ASAP7_75t_R g3149 ( 
.A(n_2987),
.Y(n_3149)
);

BUFx6f_ASAP7_75t_L g3150 ( 
.A(n_2898),
.Y(n_3150)
);

OAI21x1_ASAP7_75t_L g3151 ( 
.A1(n_2903),
.A2(n_1872),
.B(n_1834),
.Y(n_3151)
);

CKINVDCx5p33_ASAP7_75t_R g3152 ( 
.A(n_3000),
.Y(n_3152)
);

BUFx3_ASAP7_75t_L g3153 ( 
.A(n_2908),
.Y(n_3153)
);

INVxp67_ASAP7_75t_L g3154 ( 
.A(n_3012),
.Y(n_3154)
);

INVx2_ASAP7_75t_L g3155 ( 
.A(n_2830),
.Y(n_3155)
);

INVx3_ASAP7_75t_L g3156 ( 
.A(n_2914),
.Y(n_3156)
);

BUFx12f_ASAP7_75t_L g3157 ( 
.A(n_2855),
.Y(n_3157)
);

AND2x4_ASAP7_75t_L g3158 ( 
.A(n_2909),
.B(n_2252),
.Y(n_3158)
);

INVx1_ASAP7_75t_L g3159 ( 
.A(n_2832),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_2833),
.Y(n_3160)
);

BUFx6f_ASAP7_75t_L g3161 ( 
.A(n_2955),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_L g3162 ( 
.A(n_3011),
.B(n_2308),
.Y(n_3162)
);

BUFx12f_ASAP7_75t_L g3163 ( 
.A(n_2862),
.Y(n_3163)
);

INVx2_ASAP7_75t_L g3164 ( 
.A(n_2834),
.Y(n_3164)
);

OA21x2_ASAP7_75t_L g3165 ( 
.A1(n_2836),
.A2(n_1843),
.B(n_1832),
.Y(n_3165)
);

AOI22xp5_ASAP7_75t_L g3166 ( 
.A1(n_2854),
.A2(n_2736),
.B1(n_2627),
.B2(n_2193),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_2840),
.Y(n_3167)
);

AND2x4_ASAP7_75t_L g3168 ( 
.A(n_2918),
.B(n_2443),
.Y(n_3168)
);

OA21x2_ASAP7_75t_L g3169 ( 
.A1(n_2841),
.A2(n_1851),
.B(n_1848),
.Y(n_3169)
);

CKINVDCx5p33_ASAP7_75t_R g3170 ( 
.A(n_3015),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_L g3171 ( 
.A(n_3032),
.B(n_2485),
.Y(n_3171)
);

BUFx6f_ASAP7_75t_L g3172 ( 
.A(n_2956),
.Y(n_3172)
);

BUFx6f_ASAP7_75t_L g3173 ( 
.A(n_2957),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_2842),
.Y(n_3174)
);

AND2x6_ASAP7_75t_L g3175 ( 
.A(n_2916),
.B(n_2917),
.Y(n_3175)
);

OAI22x1_ASAP7_75t_SL g3176 ( 
.A1(n_3018),
.A2(n_1859),
.B1(n_1882),
.B2(n_1794),
.Y(n_3176)
);

AND2x6_ASAP7_75t_L g3177 ( 
.A(n_2920),
.B(n_2049),
.Y(n_3177)
);

INVx2_ASAP7_75t_L g3178 ( 
.A(n_2844),
.Y(n_3178)
);

OAI21x1_ASAP7_75t_L g3179 ( 
.A1(n_2906),
.A2(n_1893),
.B(n_1890),
.Y(n_3179)
);

AND2x6_ASAP7_75t_L g3180 ( 
.A(n_2921),
.B(n_2924),
.Y(n_3180)
);

BUFx3_ASAP7_75t_L g3181 ( 
.A(n_2925),
.Y(n_3181)
);

INVx3_ASAP7_75t_L g3182 ( 
.A(n_2929),
.Y(n_3182)
);

CKINVDCx5p33_ASAP7_75t_R g3183 ( 
.A(n_3038),
.Y(n_3183)
);

BUFx6f_ASAP7_75t_L g3184 ( 
.A(n_2959),
.Y(n_3184)
);

BUFx6f_ASAP7_75t_L g3185 ( 
.A(n_2960),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_L g3186 ( 
.A(n_3039),
.B(n_2504),
.Y(n_3186)
);

BUFx12f_ASAP7_75t_L g3187 ( 
.A(n_3051),
.Y(n_3187)
);

AOI22xp5_ASAP7_75t_L g3188 ( 
.A1(n_2867),
.A2(n_2215),
.B1(n_2367),
.B2(n_2353),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_2845),
.Y(n_3189)
);

OAI22xp5_ASAP7_75t_L g3190 ( 
.A1(n_2881),
.A2(n_2534),
.B1(n_2547),
.B2(n_2398),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_2847),
.Y(n_3191)
);

NAND2xp33_ASAP7_75t_L g3192 ( 
.A(n_3052),
.B(n_1771),
.Y(n_3192)
);

NOR2xp33_ASAP7_75t_L g3193 ( 
.A(n_2889),
.B(n_2931),
.Y(n_3193)
);

NAND2xp5_ASAP7_75t_L g3194 ( 
.A(n_3054),
.B(n_2656),
.Y(n_3194)
);

BUFx6f_ASAP7_75t_L g3195 ( 
.A(n_2961),
.Y(n_3195)
);

INVx2_ASAP7_75t_L g3196 ( 
.A(n_2953),
.Y(n_3196)
);

INVx1_ASAP7_75t_L g3197 ( 
.A(n_2848),
.Y(n_3197)
);

BUFx3_ASAP7_75t_L g3198 ( 
.A(n_2933),
.Y(n_3198)
);

OAI21x1_ASAP7_75t_L g3199 ( 
.A1(n_2907),
.A2(n_1904),
.B(n_1895),
.Y(n_3199)
);

OA21x2_ASAP7_75t_L g3200 ( 
.A1(n_2875),
.A2(n_1905),
.B(n_1883),
.Y(n_3200)
);

BUFx6f_ASAP7_75t_L g3201 ( 
.A(n_2962),
.Y(n_3201)
);

INVx2_ASAP7_75t_L g3202 ( 
.A(n_2953),
.Y(n_3202)
);

OAI22x1_ASAP7_75t_R g3203 ( 
.A1(n_2827),
.A2(n_1959),
.B1(n_1978),
.B2(n_1954),
.Y(n_3203)
);

BUFx6f_ASAP7_75t_L g3204 ( 
.A(n_2963),
.Y(n_3204)
);

INVx2_ASAP7_75t_L g3205 ( 
.A(n_2953),
.Y(n_3205)
);

AND2x4_ASAP7_75t_L g3206 ( 
.A(n_2927),
.B(n_2496),
.Y(n_3206)
);

BUFx3_ASAP7_75t_L g3207 ( 
.A(n_2935),
.Y(n_3207)
);

AND2x4_ASAP7_75t_L g3208 ( 
.A(n_2928),
.B(n_2537),
.Y(n_3208)
);

OAI22x1_ASAP7_75t_SL g3209 ( 
.A1(n_2829),
.A2(n_2025),
.B1(n_2061),
.B2(n_2015),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_2849),
.Y(n_3210)
);

NOR2xp33_ASAP7_75t_L g3211 ( 
.A(n_2950),
.B(n_2562),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_2850),
.Y(n_3212)
);

BUFx6f_ASAP7_75t_L g3213 ( 
.A(n_2964),
.Y(n_3213)
);

INVx6_ASAP7_75t_L g3214 ( 
.A(n_2922),
.Y(n_3214)
);

INVx2_ASAP7_75t_L g3215 ( 
.A(n_2953),
.Y(n_3215)
);

INVx3_ASAP7_75t_L g3216 ( 
.A(n_2936),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_2851),
.Y(n_3217)
);

INVx1_ASAP7_75t_L g3218 ( 
.A(n_2966),
.Y(n_3218)
);

AND2x4_ASAP7_75t_L g3219 ( 
.A(n_2930),
.B(n_2606),
.Y(n_3219)
);

AND2x2_ASAP7_75t_L g3220 ( 
.A(n_2965),
.B(n_2645),
.Y(n_3220)
);

INVx2_ASAP7_75t_L g3221 ( 
.A(n_2953),
.Y(n_3221)
);

INVx2_ASAP7_75t_L g3222 ( 
.A(n_2968),
.Y(n_3222)
);

BUFx6f_ASAP7_75t_L g3223 ( 
.A(n_2970),
.Y(n_3223)
);

NOR2xp33_ASAP7_75t_L g3224 ( 
.A(n_3003),
.B(n_2734),
.Y(n_3224)
);

HB1xp67_ASAP7_75t_L g3225 ( 
.A(n_2988),
.Y(n_3225)
);

BUFx12f_ASAP7_75t_L g3226 ( 
.A(n_3056),
.Y(n_3226)
);

INVx2_ASAP7_75t_L g3227 ( 
.A(n_2971),
.Y(n_3227)
);

BUFx12f_ASAP7_75t_L g3228 ( 
.A(n_3063),
.Y(n_3228)
);

CKINVDCx6p67_ASAP7_75t_R g3229 ( 
.A(n_3070),
.Y(n_3229)
);

OAI21x1_ASAP7_75t_L g3230 ( 
.A1(n_2912),
.A2(n_1940),
.B(n_1929),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_2972),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_2973),
.Y(n_3232)
);

AND2x4_ASAP7_75t_L g3233 ( 
.A(n_2820),
.B(n_2727),
.Y(n_3233)
);

OA21x2_ASAP7_75t_L g3234 ( 
.A1(n_2877),
.A2(n_2993),
.B(n_2982),
.Y(n_3234)
);

BUFx6f_ASAP7_75t_L g3235 ( 
.A(n_2975),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_2976),
.Y(n_3236)
);

OAI21x1_ASAP7_75t_L g3237 ( 
.A1(n_2923),
.A2(n_3028),
.B(n_2994),
.Y(n_3237)
);

INVxp67_ASAP7_75t_L g3238 ( 
.A(n_2938),
.Y(n_3238)
);

BUFx2_ASAP7_75t_L g3239 ( 
.A(n_3074),
.Y(n_3239)
);

NAND2xp5_ASAP7_75t_L g3240 ( 
.A(n_2967),
.B(n_2766),
.Y(n_3240)
);

NOR2xp33_ASAP7_75t_L g3241 ( 
.A(n_3030),
.B(n_1924),
.Y(n_3241)
);

BUFx6f_ASAP7_75t_L g3242 ( 
.A(n_2978),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_2979),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_2980),
.Y(n_3244)
);

OAI22xp5_ASAP7_75t_L g3245 ( 
.A1(n_2826),
.A2(n_1772),
.B1(n_1780),
.B2(n_1775),
.Y(n_3245)
);

INVx3_ASAP7_75t_L g3246 ( 
.A(n_2941),
.Y(n_3246)
);

BUFx6f_ASAP7_75t_L g3247 ( 
.A(n_2981),
.Y(n_3247)
);

INVx2_ASAP7_75t_L g3248 ( 
.A(n_2990),
.Y(n_3248)
);

OAI22xp5_ASAP7_75t_L g3249 ( 
.A1(n_2835),
.A2(n_1792),
.B1(n_1797),
.B2(n_1781),
.Y(n_3249)
);

INVx2_ASAP7_75t_L g3250 ( 
.A(n_2991),
.Y(n_3250)
);

INVx4_ASAP7_75t_L g3251 ( 
.A(n_3044),
.Y(n_3251)
);

OA21x2_ASAP7_75t_L g3252 ( 
.A1(n_2999),
.A2(n_1943),
.B(n_1938),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_L g3253 ( 
.A(n_3004),
.B(n_1986),
.Y(n_3253)
);

BUFx6f_ASAP7_75t_L g3254 ( 
.A(n_2992),
.Y(n_3254)
);

INVx2_ASAP7_75t_L g3255 ( 
.A(n_2995),
.Y(n_3255)
);

AND2x2_ASAP7_75t_L g3256 ( 
.A(n_2824),
.B(n_2050),
.Y(n_3256)
);

NAND2xp5_ASAP7_75t_L g3257 ( 
.A(n_3005),
.B(n_3021),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_2996),
.Y(n_3258)
);

BUFx6f_ASAP7_75t_L g3259 ( 
.A(n_2997),
.Y(n_3259)
);

NAND2xp5_ASAP7_75t_L g3260 ( 
.A(n_3033),
.B(n_2024),
.Y(n_3260)
);

BUFx2_ASAP7_75t_L g3261 ( 
.A(n_2883),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_2998),
.Y(n_3262)
);

INVx3_ASAP7_75t_L g3263 ( 
.A(n_2943),
.Y(n_3263)
);

AOI22xp5_ASAP7_75t_L g3264 ( 
.A1(n_2831),
.A2(n_2412),
.B1(n_2495),
.B2(n_2390),
.Y(n_3264)
);

INVx3_ASAP7_75t_L g3265 ( 
.A(n_2944),
.Y(n_3265)
);

INVx3_ASAP7_75t_L g3266 ( 
.A(n_2945),
.Y(n_3266)
);

BUFx2_ASAP7_75t_L g3267 ( 
.A(n_2934),
.Y(n_3267)
);

BUFx6f_ASAP7_75t_L g3268 ( 
.A(n_3002),
.Y(n_3268)
);

INVx3_ASAP7_75t_L g3269 ( 
.A(n_2947),
.Y(n_3269)
);

INVx2_ASAP7_75t_L g3270 ( 
.A(n_3006),
.Y(n_3270)
);

HB1xp67_ASAP7_75t_L g3271 ( 
.A(n_2942),
.Y(n_3271)
);

BUFx8_ASAP7_75t_L g3272 ( 
.A(n_2949),
.Y(n_3272)
);

INVx2_ASAP7_75t_SL g3273 ( 
.A(n_2951),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_3007),
.Y(n_3274)
);

INVx3_ASAP7_75t_L g3275 ( 
.A(n_2952),
.Y(n_3275)
);

AOI22x1_ASAP7_75t_SL g3276 ( 
.A1(n_2932),
.A2(n_2139),
.B1(n_2143),
.B2(n_2089),
.Y(n_3276)
);

BUFx3_ASAP7_75t_L g3277 ( 
.A(n_2954),
.Y(n_3277)
);

CKINVDCx11_ASAP7_75t_R g3278 ( 
.A(n_2984),
.Y(n_3278)
);

BUFx8_ASAP7_75t_SL g3279 ( 
.A(n_2895),
.Y(n_3279)
);

BUFx6f_ASAP7_75t_L g3280 ( 
.A(n_3008),
.Y(n_3280)
);

CKINVDCx16_ASAP7_75t_R g3281 ( 
.A(n_3001),
.Y(n_3281)
);

AOI22xp5_ASAP7_75t_L g3282 ( 
.A1(n_2837),
.A2(n_2507),
.B1(n_2524),
.B2(n_2518),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_3009),
.Y(n_3283)
);

INVx2_ASAP7_75t_L g3284 ( 
.A(n_3010),
.Y(n_3284)
);

INVx2_ASAP7_75t_L g3285 ( 
.A(n_3013),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_3014),
.Y(n_3286)
);

OAI21x1_ASAP7_75t_L g3287 ( 
.A1(n_3068),
.A2(n_2138),
.B(n_2027),
.Y(n_3287)
);

INVx3_ASAP7_75t_L g3288 ( 
.A(n_3016),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_3017),
.Y(n_3289)
);

INVx2_ASAP7_75t_L g3290 ( 
.A(n_3019),
.Y(n_3290)
);

OAI21x1_ASAP7_75t_L g3291 ( 
.A1(n_3048),
.A2(n_2164),
.B(n_2153),
.Y(n_3291)
);

AND2x2_ASAP7_75t_L g3292 ( 
.A(n_3220),
.B(n_2858),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_3218),
.Y(n_3293)
);

INVx1_ASAP7_75t_L g3294 ( 
.A(n_3231),
.Y(n_3294)
);

AND2x6_ASAP7_75t_L g3295 ( 
.A(n_3091),
.B(n_1981),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_3232),
.Y(n_3296)
);

INVxp67_ASAP7_75t_L g3297 ( 
.A(n_3271),
.Y(n_3297)
);

INVx2_ASAP7_75t_L g3298 ( 
.A(n_3083),
.Y(n_3298)
);

INVx1_ASAP7_75t_L g3299 ( 
.A(n_3236),
.Y(n_3299)
);

INVx2_ASAP7_75t_L g3300 ( 
.A(n_3098),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_3243),
.Y(n_3301)
);

BUFx6f_ASAP7_75t_L g3302 ( 
.A(n_3103),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_L g3303 ( 
.A(n_3234),
.B(n_3057),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_L g3304 ( 
.A(n_3106),
.B(n_3031),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_3244),
.Y(n_3305)
);

BUFx6f_ASAP7_75t_L g3306 ( 
.A(n_3107),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_3258),
.Y(n_3307)
);

INVx2_ASAP7_75t_L g3308 ( 
.A(n_3114),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_3262),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_3274),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_3283),
.Y(n_3311)
);

INVx2_ASAP7_75t_L g3312 ( 
.A(n_3120),
.Y(n_3312)
);

INVx2_ASAP7_75t_L g3313 ( 
.A(n_3130),
.Y(n_3313)
);

BUFx6f_ASAP7_75t_L g3314 ( 
.A(n_3115),
.Y(n_3314)
);

NOR2xp33_ASAP7_75t_L g3315 ( 
.A(n_3211),
.B(n_3043),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_3286),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_3289),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3161),
.Y(n_3318)
);

INVx2_ASAP7_75t_L g3319 ( 
.A(n_3128),
.Y(n_3319)
);

AND2x4_ASAP7_75t_L g3320 ( 
.A(n_3119),
.B(n_2870),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_3172),
.Y(n_3321)
);

INVx1_ASAP7_75t_L g3322 ( 
.A(n_3173),
.Y(n_3322)
);

INVx2_ASAP7_75t_SL g3323 ( 
.A(n_3214),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_3184),
.Y(n_3324)
);

OA21x2_ASAP7_75t_L g3325 ( 
.A1(n_3237),
.A2(n_2258),
.B(n_2251),
.Y(n_3325)
);

HB1xp67_ASAP7_75t_L g3326 ( 
.A(n_3104),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_3185),
.Y(n_3327)
);

INVx2_ASAP7_75t_L g3328 ( 
.A(n_3122),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_SL g3329 ( 
.A(n_3224),
.B(n_2958),
.Y(n_3329)
);

AND2x4_ASAP7_75t_L g3330 ( 
.A(n_3097),
.B(n_3020),
.Y(n_3330)
);

OA21x2_ASAP7_75t_L g3331 ( 
.A1(n_3151),
.A2(n_3199),
.B(n_3179),
.Y(n_3331)
);

NAND2xp33_ASAP7_75t_SL g3332 ( 
.A(n_3094),
.B(n_2822),
.Y(n_3332)
);

INVx2_ASAP7_75t_L g3333 ( 
.A(n_3129),
.Y(n_3333)
);

HB1xp67_ASAP7_75t_L g3334 ( 
.A(n_3113),
.Y(n_3334)
);

AND2x2_ASAP7_75t_L g3335 ( 
.A(n_3133),
.B(n_2860),
.Y(n_3335)
);

INVx1_ASAP7_75t_L g3336 ( 
.A(n_3195),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_3201),
.Y(n_3337)
);

INVx2_ASAP7_75t_L g3338 ( 
.A(n_3132),
.Y(n_3338)
);

INVx1_ASAP7_75t_L g3339 ( 
.A(n_3204),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_3213),
.Y(n_3340)
);

INVx2_ASAP7_75t_L g3341 ( 
.A(n_3080),
.Y(n_3341)
);

OA21x2_ASAP7_75t_L g3342 ( 
.A1(n_3230),
.A2(n_2281),
.B(n_2275),
.Y(n_3342)
);

INVx2_ASAP7_75t_L g3343 ( 
.A(n_3081),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_3223),
.Y(n_3344)
);

INVx2_ASAP7_75t_L g3345 ( 
.A(n_3087),
.Y(n_3345)
);

AND2x2_ASAP7_75t_L g3346 ( 
.A(n_3112),
.B(n_2937),
.Y(n_3346)
);

NAND2xp5_ASAP7_75t_L g3347 ( 
.A(n_3127),
.B(n_1800),
.Y(n_3347)
);

INVx1_ASAP7_75t_L g3348 ( 
.A(n_3235),
.Y(n_3348)
);

INVx1_ASAP7_75t_L g3349 ( 
.A(n_3242),
.Y(n_3349)
);

INVx2_ASAP7_75t_L g3350 ( 
.A(n_3088),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_L g3351 ( 
.A(n_3158),
.B(n_1804),
.Y(n_3351)
);

INVx3_ASAP7_75t_L g3352 ( 
.A(n_3247),
.Y(n_3352)
);

INVx2_ASAP7_75t_L g3353 ( 
.A(n_3089),
.Y(n_3353)
);

INVxp67_ASAP7_75t_L g3354 ( 
.A(n_3261),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_L g3355 ( 
.A(n_3168),
.B(n_1805),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_3254),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_3259),
.Y(n_3357)
);

INVx1_ASAP7_75t_L g3358 ( 
.A(n_3268),
.Y(n_3358)
);

INVx2_ASAP7_75t_L g3359 ( 
.A(n_3090),
.Y(n_3359)
);

BUFx6f_ASAP7_75t_L g3360 ( 
.A(n_3138),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_3280),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3159),
.Y(n_3362)
);

AND2x4_ASAP7_75t_L g3363 ( 
.A(n_3111),
.B(n_3022),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_3160),
.Y(n_3364)
);

INVx2_ASAP7_75t_L g3365 ( 
.A(n_3092),
.Y(n_3365)
);

INVx1_ASAP7_75t_L g3366 ( 
.A(n_3167),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_3174),
.Y(n_3367)
);

NOR2x1_ASAP7_75t_L g3368 ( 
.A(n_3082),
.B(n_2570),
.Y(n_3368)
);

INVx2_ASAP7_75t_L g3369 ( 
.A(n_3099),
.Y(n_3369)
);

INVx2_ASAP7_75t_L g3370 ( 
.A(n_3109),
.Y(n_3370)
);

INVx2_ASAP7_75t_L g3371 ( 
.A(n_3116),
.Y(n_3371)
);

OAI21x1_ASAP7_75t_L g3372 ( 
.A1(n_3287),
.A2(n_2508),
.B(n_2462),
.Y(n_3372)
);

INVx1_ASAP7_75t_L g3373 ( 
.A(n_3189),
.Y(n_3373)
);

AO21x2_ASAP7_75t_L g3374 ( 
.A1(n_3084),
.A2(n_1946),
.B(n_1945),
.Y(n_3374)
);

AND2x2_ASAP7_75t_L g3375 ( 
.A(n_3206),
.B(n_2948),
.Y(n_3375)
);

AND2x4_ASAP7_75t_L g3376 ( 
.A(n_3095),
.B(n_3023),
.Y(n_3376)
);

BUFx6f_ASAP7_75t_L g3377 ( 
.A(n_3150),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_3191),
.Y(n_3378)
);

AND2x2_ASAP7_75t_L g3379 ( 
.A(n_3208),
.B(n_2983),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_3155),
.Y(n_3380)
);

NAND2xp5_ASAP7_75t_L g3381 ( 
.A(n_3219),
.B(n_3251),
.Y(n_3381)
);

INVx2_ASAP7_75t_L g3382 ( 
.A(n_3117),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_L g3383 ( 
.A(n_3241),
.B(n_1808),
.Y(n_3383)
);

CKINVDCx5p33_ASAP7_75t_R g3384 ( 
.A(n_3279),
.Y(n_3384)
);

BUFx6f_ASAP7_75t_L g3385 ( 
.A(n_3153),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_3164),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_3178),
.Y(n_3387)
);

NOR2xp33_ASAP7_75t_L g3388 ( 
.A(n_3118),
.B(n_3055),
.Y(n_3388)
);

INVx3_ASAP7_75t_L g3389 ( 
.A(n_3100),
.Y(n_3389)
);

INVxp33_ASAP7_75t_SL g3390 ( 
.A(n_3188),
.Y(n_3390)
);

BUFx6f_ASAP7_75t_L g3391 ( 
.A(n_3181),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_SL g3392 ( 
.A(n_3086),
.B(n_2615),
.Y(n_3392)
);

INVx2_ASAP7_75t_L g3393 ( 
.A(n_3123),
.Y(n_3393)
);

INVx2_ASAP7_75t_L g3394 ( 
.A(n_3124),
.Y(n_3394)
);

INVx2_ASAP7_75t_L g3395 ( 
.A(n_3136),
.Y(n_3395)
);

INVx1_ASAP7_75t_L g3396 ( 
.A(n_3198),
.Y(n_3396)
);

INVx2_ASAP7_75t_L g3397 ( 
.A(n_3137),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_L g3398 ( 
.A(n_3125),
.B(n_3162),
.Y(n_3398)
);

INVx1_ASAP7_75t_L g3399 ( 
.A(n_3207),
.Y(n_3399)
);

INVx2_ASAP7_75t_L g3400 ( 
.A(n_3140),
.Y(n_3400)
);

HB1xp67_ASAP7_75t_L g3401 ( 
.A(n_3126),
.Y(n_3401)
);

INVx1_ASAP7_75t_L g3402 ( 
.A(n_3277),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_3197),
.Y(n_3403)
);

INVx2_ASAP7_75t_L g3404 ( 
.A(n_3141),
.Y(n_3404)
);

INVx3_ASAP7_75t_L g3405 ( 
.A(n_3105),
.Y(n_3405)
);

INVx2_ASAP7_75t_L g3406 ( 
.A(n_3142),
.Y(n_3406)
);

INVx2_ASAP7_75t_L g3407 ( 
.A(n_3143),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_SL g3408 ( 
.A(n_3193),
.B(n_2680),
.Y(n_3408)
);

INVx1_ASAP7_75t_L g3409 ( 
.A(n_3210),
.Y(n_3409)
);

HB1xp67_ASAP7_75t_L g3410 ( 
.A(n_3144),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_3212),
.Y(n_3411)
);

NAND2xp5_ASAP7_75t_L g3412 ( 
.A(n_3171),
.B(n_1811),
.Y(n_3412)
);

INVx6_ASAP7_75t_L g3413 ( 
.A(n_3272),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_L g3414 ( 
.A(n_3186),
.B(n_1813),
.Y(n_3414)
);

AND2x2_ASAP7_75t_L g3415 ( 
.A(n_3096),
.B(n_3025),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_3217),
.Y(n_3416)
);

OA21x2_ASAP7_75t_L g3417 ( 
.A1(n_3291),
.A2(n_2574),
.B(n_2540),
.Y(n_3417)
);

INVx2_ASAP7_75t_L g3418 ( 
.A(n_3148),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_SL g3419 ( 
.A(n_3101),
.B(n_2705),
.Y(n_3419)
);

INVx2_ASAP7_75t_L g3420 ( 
.A(n_3222),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_3227),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_3248),
.Y(n_3422)
);

AND2x4_ASAP7_75t_L g3423 ( 
.A(n_3239),
.B(n_3024),
.Y(n_3423)
);

AND2x2_ASAP7_75t_L g3424 ( 
.A(n_3256),
.B(n_3026),
.Y(n_3424)
);

INVx1_ASAP7_75t_L g3425 ( 
.A(n_3250),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_3255),
.Y(n_3426)
);

BUFx6f_ASAP7_75t_L g3427 ( 
.A(n_3121),
.Y(n_3427)
);

INVx2_ASAP7_75t_L g3428 ( 
.A(n_3270),
.Y(n_3428)
);

INVx3_ASAP7_75t_L g3429 ( 
.A(n_3288),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_3284),
.Y(n_3430)
);

INVx2_ASAP7_75t_L g3431 ( 
.A(n_3285),
.Y(n_3431)
);

NAND2xp5_ASAP7_75t_L g3432 ( 
.A(n_3194),
.B(n_1816),
.Y(n_3432)
);

INVx2_ASAP7_75t_L g3433 ( 
.A(n_3290),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_3273),
.Y(n_3434)
);

CKINVDCx5p33_ASAP7_75t_R g3435 ( 
.A(n_3093),
.Y(n_3435)
);

INVx1_ASAP7_75t_L g3436 ( 
.A(n_3156),
.Y(n_3436)
);

INVx1_ASAP7_75t_L g3437 ( 
.A(n_3182),
.Y(n_3437)
);

BUFx2_ASAP7_75t_L g3438 ( 
.A(n_3225),
.Y(n_3438)
);

AND2x2_ASAP7_75t_L g3439 ( 
.A(n_3233),
.B(n_3154),
.Y(n_3439)
);

INVx2_ASAP7_75t_L g3440 ( 
.A(n_3079),
.Y(n_3440)
);

NAND2xp5_ASAP7_75t_SL g3441 ( 
.A(n_3145),
.B(n_2713),
.Y(n_3441)
);

INVx3_ASAP7_75t_L g3442 ( 
.A(n_3216),
.Y(n_3442)
);

INVx2_ASAP7_75t_L g3443 ( 
.A(n_3246),
.Y(n_3443)
);

AND2x6_ASAP7_75t_L g3444 ( 
.A(n_3166),
.B(n_1981),
.Y(n_3444)
);

INVx2_ASAP7_75t_L g3445 ( 
.A(n_3263),
.Y(n_3445)
);

INVx2_ASAP7_75t_L g3446 ( 
.A(n_3265),
.Y(n_3446)
);

BUFx4f_ASAP7_75t_L g3447 ( 
.A(n_3229),
.Y(n_3447)
);

INVx2_ASAP7_75t_L g3448 ( 
.A(n_3266),
.Y(n_3448)
);

INVx1_ASAP7_75t_L g3449 ( 
.A(n_3269),
.Y(n_3449)
);

INVx1_ASAP7_75t_L g3450 ( 
.A(n_3275),
.Y(n_3450)
);

INVx1_ASAP7_75t_L g3451 ( 
.A(n_3196),
.Y(n_3451)
);

OAI21x1_ASAP7_75t_L g3452 ( 
.A1(n_3200),
.A2(n_2665),
.B(n_2629),
.Y(n_3452)
);

AOI22xp5_ASAP7_75t_L g3453 ( 
.A1(n_3085),
.A2(n_2720),
.B1(n_2776),
.B2(n_2760),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_3202),
.Y(n_3454)
);

INVx2_ASAP7_75t_L g3455 ( 
.A(n_3205),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_3215),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_3221),
.Y(n_3457)
);

INVx3_ASAP7_75t_L g3458 ( 
.A(n_3146),
.Y(n_3458)
);

INVx2_ASAP7_75t_L g3459 ( 
.A(n_3165),
.Y(n_3459)
);

INVx2_ASAP7_75t_L g3460 ( 
.A(n_3169),
.Y(n_3460)
);

INVx2_ASAP7_75t_L g3461 ( 
.A(n_3252),
.Y(n_3461)
);

AND2x2_ASAP7_75t_L g3462 ( 
.A(n_3267),
.B(n_3027),
.Y(n_3462)
);

INVx1_ASAP7_75t_L g3463 ( 
.A(n_3238),
.Y(n_3463)
);

INVx2_ASAP7_75t_L g3464 ( 
.A(n_3257),
.Y(n_3464)
);

INVx2_ASAP7_75t_L g3465 ( 
.A(n_3253),
.Y(n_3465)
);

INVx2_ASAP7_75t_L g3466 ( 
.A(n_3260),
.Y(n_3466)
);

BUFx6f_ASAP7_75t_L g3467 ( 
.A(n_3175),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_3240),
.Y(n_3468)
);

CKINVDCx16_ASAP7_75t_R g3469 ( 
.A(n_3203),
.Y(n_3469)
);

INVx2_ASAP7_75t_L g3470 ( 
.A(n_3175),
.Y(n_3470)
);

INVx3_ASAP7_75t_L g3471 ( 
.A(n_3180),
.Y(n_3471)
);

NAND2xp5_ASAP7_75t_L g3472 ( 
.A(n_3180),
.B(n_3135),
.Y(n_3472)
);

NAND2xp5_ASAP7_75t_L g3473 ( 
.A(n_3192),
.B(n_1819),
.Y(n_3473)
);

INVx1_ASAP7_75t_L g3474 ( 
.A(n_3108),
.Y(n_3474)
);

INVx2_ASAP7_75t_L g3475 ( 
.A(n_3108),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_L g3476 ( 
.A(n_3149),
.B(n_1824),
.Y(n_3476)
);

INVx1_ASAP7_75t_L g3477 ( 
.A(n_3177),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_3177),
.Y(n_3478)
);

OAI21x1_ASAP7_75t_L g3479 ( 
.A1(n_3245),
.A2(n_2728),
.B(n_1951),
.Y(n_3479)
);

HB1xp67_ASAP7_75t_L g3480 ( 
.A(n_3134),
.Y(n_3480)
);

BUFx2_ASAP7_75t_L g3481 ( 
.A(n_3102),
.Y(n_3481)
);

CKINVDCx20_ASAP7_75t_R g3482 ( 
.A(n_3281),
.Y(n_3482)
);

INVx2_ASAP7_75t_L g3483 ( 
.A(n_3110),
.Y(n_3483)
);

BUFx6f_ASAP7_75t_L g3484 ( 
.A(n_3102),
.Y(n_3484)
);

HB1xp67_ASAP7_75t_L g3485 ( 
.A(n_3249),
.Y(n_3485)
);

INVx2_ASAP7_75t_L g3486 ( 
.A(n_3152),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3190),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_3170),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_L g3489 ( 
.A(n_3183),
.B(n_1829),
.Y(n_3489)
);

INVxp67_ASAP7_75t_L g3490 ( 
.A(n_3264),
.Y(n_3490)
);

INVx2_ASAP7_75t_L g3491 ( 
.A(n_3139),
.Y(n_3491)
);

INVx3_ASAP7_75t_L g3492 ( 
.A(n_3228),
.Y(n_3492)
);

INVx2_ASAP7_75t_L g3493 ( 
.A(n_3187),
.Y(n_3493)
);

INVx2_ASAP7_75t_L g3494 ( 
.A(n_3226),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3282),
.Y(n_3495)
);

INVx1_ASAP7_75t_L g3496 ( 
.A(n_3176),
.Y(n_3496)
);

OAI21x1_ASAP7_75t_L g3497 ( 
.A1(n_3131),
.A2(n_1952),
.B(n_1947),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_3147),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_L g3499 ( 
.A(n_3157),
.B(n_1840),
.Y(n_3499)
);

INVx1_ASAP7_75t_L g3500 ( 
.A(n_3163),
.Y(n_3500)
);

INVx2_ASAP7_75t_L g3501 ( 
.A(n_3276),
.Y(n_3501)
);

INVx3_ASAP7_75t_L g3502 ( 
.A(n_3278),
.Y(n_3502)
);

INVx2_ASAP7_75t_L g3503 ( 
.A(n_3209),
.Y(n_3503)
);

BUFx6f_ASAP7_75t_L g3504 ( 
.A(n_3103),
.Y(n_3504)
);

AND2x2_ASAP7_75t_L g3505 ( 
.A(n_3220),
.B(n_3034),
.Y(n_3505)
);

INVx3_ASAP7_75t_L g3506 ( 
.A(n_3103),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_3218),
.Y(n_3507)
);

INVx2_ASAP7_75t_L g3508 ( 
.A(n_3083),
.Y(n_3508)
);

INVx2_ASAP7_75t_L g3509 ( 
.A(n_3083),
.Y(n_3509)
);

BUFx8_ASAP7_75t_L g3510 ( 
.A(n_3239),
.Y(n_3510)
);

INVx1_ASAP7_75t_L g3511 ( 
.A(n_3218),
.Y(n_3511)
);

INVx2_ASAP7_75t_L g3512 ( 
.A(n_3083),
.Y(n_3512)
);

INVx2_ASAP7_75t_L g3513 ( 
.A(n_3083),
.Y(n_3513)
);

BUFx6f_ASAP7_75t_L g3514 ( 
.A(n_3103),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_L g3515 ( 
.A(n_3234),
.B(n_1841),
.Y(n_3515)
);

BUFx6f_ASAP7_75t_L g3516 ( 
.A(n_3103),
.Y(n_3516)
);

INVx2_ASAP7_75t_L g3517 ( 
.A(n_3083),
.Y(n_3517)
);

INVx1_ASAP7_75t_L g3518 ( 
.A(n_3218),
.Y(n_3518)
);

INVx2_ASAP7_75t_L g3519 ( 
.A(n_3420),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_SL g3520 ( 
.A(n_3346),
.B(n_3029),
.Y(n_3520)
);

AND2x2_ASAP7_75t_L g3521 ( 
.A(n_3375),
.B(n_3046),
.Y(n_3521)
);

BUFx3_ASAP7_75t_L g3522 ( 
.A(n_3385),
.Y(n_3522)
);

INVx4_ASAP7_75t_L g3523 ( 
.A(n_3360),
.Y(n_3523)
);

INVx3_ASAP7_75t_L g3524 ( 
.A(n_3302),
.Y(n_3524)
);

OAI22xp33_ASAP7_75t_L g3525 ( 
.A1(n_3495),
.A2(n_3047),
.B1(n_2902),
.B2(n_2911),
.Y(n_3525)
);

INVx4_ASAP7_75t_SL g3526 ( 
.A(n_3413),
.Y(n_3526)
);

NAND2xp5_ASAP7_75t_L g3527 ( 
.A(n_3398),
.B(n_1961),
.Y(n_3527)
);

CKINVDCx5p33_ASAP7_75t_R g3528 ( 
.A(n_3435),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_3293),
.Y(n_3529)
);

INVx2_ASAP7_75t_L g3530 ( 
.A(n_3428),
.Y(n_3530)
);

BUFx6f_ASAP7_75t_L g3531 ( 
.A(n_3302),
.Y(n_3531)
);

AND2x2_ASAP7_75t_L g3532 ( 
.A(n_3379),
.B(n_3035),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_3294),
.Y(n_3533)
);

BUFx3_ASAP7_75t_L g3534 ( 
.A(n_3385),
.Y(n_3534)
);

NAND2xp5_ASAP7_75t_L g3535 ( 
.A(n_3464),
.B(n_1963),
.Y(n_3535)
);

OR2x6_ASAP7_75t_L g3536 ( 
.A(n_3323),
.B(n_2182),
.Y(n_3536)
);

AND2x2_ASAP7_75t_L g3537 ( 
.A(n_3424),
.B(n_3036),
.Y(n_3537)
);

INVxp67_ASAP7_75t_SL g3538 ( 
.A(n_3427),
.Y(n_3538)
);

BUFx3_ASAP7_75t_L g3539 ( 
.A(n_3391),
.Y(n_3539)
);

CKINVDCx5p33_ASAP7_75t_R g3540 ( 
.A(n_3384),
.Y(n_3540)
);

NOR2xp33_ASAP7_75t_L g3541 ( 
.A(n_3315),
.B(n_2919),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_L g3542 ( 
.A(n_3468),
.B(n_1979),
.Y(n_3542)
);

INVx5_ASAP7_75t_L g3543 ( 
.A(n_3484),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3296),
.Y(n_3544)
);

AND2x2_ASAP7_75t_L g3545 ( 
.A(n_3335),
.B(n_3037),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_3299),
.Y(n_3546)
);

INVx5_ASAP7_75t_L g3547 ( 
.A(n_3484),
.Y(n_3547)
);

INVx2_ASAP7_75t_SL g3548 ( 
.A(n_3320),
.Y(n_3548)
);

BUFx4f_ASAP7_75t_L g3549 ( 
.A(n_3492),
.Y(n_3549)
);

INVx4_ASAP7_75t_L g3550 ( 
.A(n_3360),
.Y(n_3550)
);

AND2x2_ASAP7_75t_L g3551 ( 
.A(n_3292),
.B(n_3040),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_SL g3552 ( 
.A(n_3304),
.B(n_1844),
.Y(n_3552)
);

AND2x6_ASAP7_75t_L g3553 ( 
.A(n_3415),
.B(n_2344),
.Y(n_3553)
);

INVx1_ASAP7_75t_L g3554 ( 
.A(n_3301),
.Y(n_3554)
);

BUFx4f_ASAP7_75t_L g3555 ( 
.A(n_3502),
.Y(n_3555)
);

NAND2xp5_ASAP7_75t_L g3556 ( 
.A(n_3465),
.B(n_3466),
.Y(n_3556)
);

INVx2_ASAP7_75t_L g3557 ( 
.A(n_3431),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_L g3558 ( 
.A(n_3505),
.B(n_2000),
.Y(n_3558)
);

NAND2xp5_ASAP7_75t_L g3559 ( 
.A(n_3362),
.B(n_2006),
.Y(n_3559)
);

INVx2_ASAP7_75t_L g3560 ( 
.A(n_3433),
.Y(n_3560)
);

INVx4_ASAP7_75t_L g3561 ( 
.A(n_3377),
.Y(n_3561)
);

INVx1_ASAP7_75t_L g3562 ( 
.A(n_3305),
.Y(n_3562)
);

AND2x2_ASAP7_75t_L g3563 ( 
.A(n_3462),
.B(n_3041),
.Y(n_3563)
);

AOI22xp33_ASAP7_75t_L g3564 ( 
.A1(n_3461),
.A2(n_2008),
.B1(n_2012),
.B2(n_2007),
.Y(n_3564)
);

AOI22xp33_ASAP7_75t_L g3565 ( 
.A1(n_3487),
.A2(n_2035),
.B1(n_2042),
.B2(n_2016),
.Y(n_3565)
);

NOR2xp33_ASAP7_75t_L g3566 ( 
.A(n_3388),
.B(n_2053),
.Y(n_3566)
);

BUFx6f_ASAP7_75t_L g3567 ( 
.A(n_3306),
.Y(n_3567)
);

NOR2xp33_ASAP7_75t_L g3568 ( 
.A(n_3383),
.B(n_2075),
.Y(n_3568)
);

CKINVDCx6p67_ASAP7_75t_R g3569 ( 
.A(n_3469),
.Y(n_3569)
);

INVxp67_ASAP7_75t_SL g3570 ( 
.A(n_3427),
.Y(n_3570)
);

INVx4_ASAP7_75t_L g3571 ( 
.A(n_3377),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3307),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_3309),
.Y(n_3573)
);

BUFx2_ASAP7_75t_L g3574 ( 
.A(n_3326),
.Y(n_3574)
);

AND2x4_ASAP7_75t_L g3575 ( 
.A(n_3352),
.B(n_3042),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_3310),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3311),
.Y(n_3577)
);

NAND2xp33_ASAP7_75t_L g3578 ( 
.A(n_3368),
.B(n_1846),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_SL g3579 ( 
.A(n_3381),
.B(n_1854),
.Y(n_3579)
);

NOR2xp33_ASAP7_75t_L g3580 ( 
.A(n_3329),
.B(n_2158),
.Y(n_3580)
);

INVx2_ASAP7_75t_L g3581 ( 
.A(n_3455),
.Y(n_3581)
);

OR2x2_ASAP7_75t_L g3582 ( 
.A(n_3334),
.B(n_2183),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_3316),
.Y(n_3583)
);

AOI22xp33_ASAP7_75t_L g3584 ( 
.A1(n_3303),
.A2(n_2060),
.B1(n_2077),
.B2(n_2046),
.Y(n_3584)
);

BUFx6f_ASAP7_75t_L g3585 ( 
.A(n_3306),
.Y(n_3585)
);

NAND2xp33_ASAP7_75t_L g3586 ( 
.A(n_3470),
.B(n_1857),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_3364),
.B(n_2081),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_3317),
.Y(n_3588)
);

OR2x2_ASAP7_75t_L g3589 ( 
.A(n_3401),
.B(n_2239),
.Y(n_3589)
);

BUFx2_ASAP7_75t_L g3590 ( 
.A(n_3438),
.Y(n_3590)
);

INVx1_ASAP7_75t_L g3591 ( 
.A(n_3507),
.Y(n_3591)
);

INVx2_ASAP7_75t_L g3592 ( 
.A(n_3440),
.Y(n_3592)
);

AND2x4_ASAP7_75t_L g3593 ( 
.A(n_3389),
.B(n_3045),
.Y(n_3593)
);

CKINVDCx20_ASAP7_75t_R g3594 ( 
.A(n_3482),
.Y(n_3594)
);

AND2x4_ASAP7_75t_L g3595 ( 
.A(n_3405),
.B(n_3049),
.Y(n_3595)
);

BUFx2_ASAP7_75t_L g3596 ( 
.A(n_3410),
.Y(n_3596)
);

INVx6_ASAP7_75t_L g3597 ( 
.A(n_3510),
.Y(n_3597)
);

INVx4_ASAP7_75t_L g3598 ( 
.A(n_3391),
.Y(n_3598)
);

INVx5_ASAP7_75t_L g3599 ( 
.A(n_3314),
.Y(n_3599)
);

NOR2x1p5_ASAP7_75t_L g3600 ( 
.A(n_3475),
.B(n_3474),
.Y(n_3600)
);

INVx3_ASAP7_75t_L g3601 ( 
.A(n_3314),
.Y(n_3601)
);

BUFx3_ASAP7_75t_L g3602 ( 
.A(n_3504),
.Y(n_3602)
);

INVx1_ASAP7_75t_SL g3603 ( 
.A(n_3439),
.Y(n_3603)
);

INVx2_ASAP7_75t_L g3604 ( 
.A(n_3380),
.Y(n_3604)
);

INVx4_ASAP7_75t_SL g3605 ( 
.A(n_3444),
.Y(n_3605)
);

INVx6_ASAP7_75t_L g3606 ( 
.A(n_3504),
.Y(n_3606)
);

INVxp67_ASAP7_75t_SL g3607 ( 
.A(n_3429),
.Y(n_3607)
);

NOR2xp33_ASAP7_75t_L g3608 ( 
.A(n_3297),
.B(n_2303),
.Y(n_3608)
);

OAI22xp5_ASAP7_75t_L g3609 ( 
.A1(n_3485),
.A2(n_2097),
.B1(n_2123),
.B2(n_2094),
.Y(n_3609)
);

CKINVDCx20_ASAP7_75t_R g3610 ( 
.A(n_3447),
.Y(n_3610)
);

INVx2_ASAP7_75t_L g3611 ( 
.A(n_3386),
.Y(n_3611)
);

NAND2xp5_ASAP7_75t_L g3612 ( 
.A(n_3366),
.B(n_2127),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_L g3613 ( 
.A(n_3367),
.B(n_2129),
.Y(n_3613)
);

INVx3_ASAP7_75t_L g3614 ( 
.A(n_3514),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_L g3615 ( 
.A(n_3373),
.B(n_2145),
.Y(n_3615)
);

OR2x6_ASAP7_75t_L g3616 ( 
.A(n_3493),
.B(n_1779),
.Y(n_3616)
);

NAND2xp5_ASAP7_75t_SL g3617 ( 
.A(n_3376),
.B(n_1858),
.Y(n_3617)
);

BUFx10_ASAP7_75t_L g3618 ( 
.A(n_3498),
.Y(n_3618)
);

INVx2_ASAP7_75t_L g3619 ( 
.A(n_3387),
.Y(n_3619)
);

BUFx4f_ASAP7_75t_L g3620 ( 
.A(n_3500),
.Y(n_3620)
);

INVx1_ASAP7_75t_L g3621 ( 
.A(n_3511),
.Y(n_3621)
);

NAND2xp5_ASAP7_75t_L g3622 ( 
.A(n_3378),
.B(n_2146),
.Y(n_3622)
);

NOR2xp33_ASAP7_75t_L g3623 ( 
.A(n_3476),
.B(n_2374),
.Y(n_3623)
);

INVx6_ASAP7_75t_L g3624 ( 
.A(n_3514),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_L g3625 ( 
.A(n_3412),
.B(n_2152),
.Y(n_3625)
);

NAND2xp5_ASAP7_75t_L g3626 ( 
.A(n_3414),
.B(n_2155),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_SL g3627 ( 
.A(n_3467),
.B(n_1860),
.Y(n_3627)
);

OR2x2_ASAP7_75t_L g3628 ( 
.A(n_3490),
.B(n_2394),
.Y(n_3628)
);

INVx2_ASAP7_75t_L g3629 ( 
.A(n_3341),
.Y(n_3629)
);

INVx2_ASAP7_75t_L g3630 ( 
.A(n_3343),
.Y(n_3630)
);

INVx2_ASAP7_75t_L g3631 ( 
.A(n_3345),
.Y(n_3631)
);

BUFx10_ASAP7_75t_L g3632 ( 
.A(n_3423),
.Y(n_3632)
);

INVx4_ASAP7_75t_L g3633 ( 
.A(n_3467),
.Y(n_3633)
);

INVx1_ASAP7_75t_L g3634 ( 
.A(n_3518),
.Y(n_3634)
);

INVx2_ASAP7_75t_L g3635 ( 
.A(n_3350),
.Y(n_3635)
);

INVx1_ASAP7_75t_L g3636 ( 
.A(n_3403),
.Y(n_3636)
);

OR2x2_ASAP7_75t_L g3637 ( 
.A(n_3354),
.B(n_2416),
.Y(n_3637)
);

INVx2_ASAP7_75t_L g3638 ( 
.A(n_3353),
.Y(n_3638)
);

INVx3_ASAP7_75t_L g3639 ( 
.A(n_3516),
.Y(n_3639)
);

AND2x2_ASAP7_75t_L g3640 ( 
.A(n_3330),
.B(n_3050),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3409),
.Y(n_3641)
);

INVx2_ASAP7_75t_SL g3642 ( 
.A(n_3363),
.Y(n_3642)
);

INVx2_ASAP7_75t_L g3643 ( 
.A(n_3359),
.Y(n_3643)
);

INVx4_ASAP7_75t_SL g3644 ( 
.A(n_3444),
.Y(n_3644)
);

AND2x2_ASAP7_75t_L g3645 ( 
.A(n_3481),
.B(n_3053),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_3411),
.Y(n_3646)
);

NAND2xp5_ASAP7_75t_L g3647 ( 
.A(n_3432),
.B(n_2170),
.Y(n_3647)
);

NOR2xp33_ASAP7_75t_L g3648 ( 
.A(n_3489),
.B(n_3480),
.Y(n_3648)
);

AND2x6_ASAP7_75t_L g3649 ( 
.A(n_3477),
.B(n_2357),
.Y(n_3649)
);

OR2x6_ASAP7_75t_L g3650 ( 
.A(n_3494),
.B(n_3497),
.Y(n_3650)
);

INVx1_ASAP7_75t_L g3651 ( 
.A(n_3416),
.Y(n_3651)
);

NOR2xp33_ASAP7_75t_L g3652 ( 
.A(n_3478),
.B(n_2463),
.Y(n_3652)
);

BUFx2_ASAP7_75t_L g3653 ( 
.A(n_3444),
.Y(n_3653)
);

INVx1_ASAP7_75t_L g3654 ( 
.A(n_3421),
.Y(n_3654)
);

NAND2xp5_ASAP7_75t_L g3655 ( 
.A(n_3451),
.B(n_2178),
.Y(n_3655)
);

AND2x2_ASAP7_75t_SL g3656 ( 
.A(n_3453),
.B(n_2413),
.Y(n_3656)
);

INVx1_ASAP7_75t_L g3657 ( 
.A(n_3422),
.Y(n_3657)
);

BUFx10_ASAP7_75t_L g3658 ( 
.A(n_3488),
.Y(n_3658)
);

NAND2xp5_ASAP7_75t_L g3659 ( 
.A(n_3454),
.B(n_2181),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_L g3660 ( 
.A(n_3456),
.B(n_2189),
.Y(n_3660)
);

AND2x6_ASAP7_75t_L g3661 ( 
.A(n_3501),
.B(n_2360),
.Y(n_3661)
);

AND2x2_ASAP7_75t_L g3662 ( 
.A(n_3463),
.B(n_3058),
.Y(n_3662)
);

NAND2xp5_ASAP7_75t_SL g3663 ( 
.A(n_3347),
.B(n_1865),
.Y(n_3663)
);

INVx3_ASAP7_75t_L g3664 ( 
.A(n_3516),
.Y(n_3664)
);

INVx1_ASAP7_75t_L g3665 ( 
.A(n_3425),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_SL g3666 ( 
.A(n_3351),
.B(n_1866),
.Y(n_3666)
);

OR2x2_ASAP7_75t_L g3667 ( 
.A(n_3483),
.B(n_2468),
.Y(n_3667)
);

INVx1_ASAP7_75t_L g3668 ( 
.A(n_3426),
.Y(n_3668)
);

BUFx2_ASAP7_75t_L g3669 ( 
.A(n_3332),
.Y(n_3669)
);

BUFx6f_ASAP7_75t_L g3670 ( 
.A(n_3506),
.Y(n_3670)
);

INVx2_ASAP7_75t_L g3671 ( 
.A(n_3365),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_L g3672 ( 
.A(n_3457),
.B(n_2195),
.Y(n_3672)
);

NOR2xp33_ASAP7_75t_L g3673 ( 
.A(n_3408),
.B(n_2527),
.Y(n_3673)
);

INVx2_ASAP7_75t_L g3674 ( 
.A(n_3369),
.Y(n_3674)
);

INVx2_ASAP7_75t_L g3675 ( 
.A(n_3370),
.Y(n_3675)
);

NOR2xp33_ASAP7_75t_L g3676 ( 
.A(n_3355),
.B(n_2548),
.Y(n_3676)
);

INVx1_ASAP7_75t_L g3677 ( 
.A(n_3430),
.Y(n_3677)
);

INVx2_ASAP7_75t_L g3678 ( 
.A(n_3371),
.Y(n_3678)
);

AND2x2_ASAP7_75t_L g3679 ( 
.A(n_3442),
.B(n_3059),
.Y(n_3679)
);

INVx2_ASAP7_75t_L g3680 ( 
.A(n_3382),
.Y(n_3680)
);

INVx1_ASAP7_75t_L g3681 ( 
.A(n_3393),
.Y(n_3681)
);

AND2x2_ASAP7_75t_L g3682 ( 
.A(n_3491),
.B(n_3396),
.Y(n_3682)
);

INVx2_ASAP7_75t_L g3683 ( 
.A(n_3394),
.Y(n_3683)
);

BUFx3_ASAP7_75t_L g3684 ( 
.A(n_3318),
.Y(n_3684)
);

INVx4_ASAP7_75t_SL g3685 ( 
.A(n_3295),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_SL g3686 ( 
.A(n_3472),
.B(n_1867),
.Y(n_3686)
);

INVx1_ASAP7_75t_L g3687 ( 
.A(n_3395),
.Y(n_3687)
);

INVx4_ASAP7_75t_L g3688 ( 
.A(n_3471),
.Y(n_3688)
);

BUFx4f_ASAP7_75t_L g3689 ( 
.A(n_3295),
.Y(n_3689)
);

INVx1_ASAP7_75t_L g3690 ( 
.A(n_3397),
.Y(n_3690)
);

INVx5_ASAP7_75t_L g3691 ( 
.A(n_3295),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_3400),
.Y(n_3692)
);

INVx4_ASAP7_75t_L g3693 ( 
.A(n_3443),
.Y(n_3693)
);

BUFx10_ASAP7_75t_L g3694 ( 
.A(n_3496),
.Y(n_3694)
);

AND2x4_ASAP7_75t_L g3695 ( 
.A(n_3321),
.B(n_3060),
.Y(n_3695)
);

INVx1_ASAP7_75t_L g3696 ( 
.A(n_3404),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_3406),
.Y(n_3697)
);

NAND2xp5_ASAP7_75t_L g3698 ( 
.A(n_3458),
.B(n_2201),
.Y(n_3698)
);

AO22x2_ASAP7_75t_L g3699 ( 
.A1(n_3503),
.A2(n_2715),
.B1(n_2806),
.B2(n_2639),
.Y(n_3699)
);

INVx2_ASAP7_75t_L g3700 ( 
.A(n_3407),
.Y(n_3700)
);

INVx1_ASAP7_75t_L g3701 ( 
.A(n_3418),
.Y(n_3701)
);

AOI22xp5_ASAP7_75t_L g3702 ( 
.A1(n_3374),
.A2(n_1886),
.B1(n_1897),
.B2(n_1878),
.Y(n_3702)
);

BUFx6f_ASAP7_75t_L g3703 ( 
.A(n_3328),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_3298),
.Y(n_3704)
);

NOR2xp33_ASAP7_75t_L g3705 ( 
.A(n_3486),
.B(n_1801),
.Y(n_3705)
);

INVx4_ASAP7_75t_L g3706 ( 
.A(n_3445),
.Y(n_3706)
);

NAND2xp5_ASAP7_75t_L g3707 ( 
.A(n_3515),
.B(n_2207),
.Y(n_3707)
);

INVx1_ASAP7_75t_L g3708 ( 
.A(n_3300),
.Y(n_3708)
);

AOI22xp33_ASAP7_75t_L g3709 ( 
.A1(n_3459),
.A2(n_3460),
.B1(n_3479),
.B2(n_3390),
.Y(n_3709)
);

NOR2xp33_ASAP7_75t_R g3710 ( 
.A(n_3499),
.B(n_1898),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_SL g3711 ( 
.A(n_3399),
.B(n_1908),
.Y(n_3711)
);

INVx4_ASAP7_75t_L g3712 ( 
.A(n_3446),
.Y(n_3712)
);

BUFx6f_ASAP7_75t_L g3713 ( 
.A(n_3333),
.Y(n_3713)
);

NAND2xp5_ASAP7_75t_SL g3714 ( 
.A(n_3402),
.B(n_3434),
.Y(n_3714)
);

INVx2_ASAP7_75t_L g3715 ( 
.A(n_3308),
.Y(n_3715)
);

INVx2_ASAP7_75t_L g3716 ( 
.A(n_3312),
.Y(n_3716)
);

INVx2_ASAP7_75t_L g3717 ( 
.A(n_3313),
.Y(n_3717)
);

NOR2xp33_ASAP7_75t_L g3718 ( 
.A(n_3419),
.B(n_1806),
.Y(n_3718)
);

NAND2xp5_ASAP7_75t_SL g3719 ( 
.A(n_3448),
.B(n_1909),
.Y(n_3719)
);

NAND2xp5_ASAP7_75t_L g3720 ( 
.A(n_3473),
.B(n_2214),
.Y(n_3720)
);

BUFx6f_ASAP7_75t_L g3721 ( 
.A(n_3338),
.Y(n_3721)
);

NOR2xp33_ASAP7_75t_L g3722 ( 
.A(n_3441),
.B(n_1810),
.Y(n_3722)
);

INVx2_ASAP7_75t_L g3723 ( 
.A(n_3508),
.Y(n_3723)
);

BUFx3_ASAP7_75t_L g3724 ( 
.A(n_3322),
.Y(n_3724)
);

AOI22xp33_ASAP7_75t_SL g3725 ( 
.A1(n_3436),
.A2(n_2211),
.B1(n_2226),
.B2(n_2160),
.Y(n_3725)
);

BUFx3_ASAP7_75t_L g3726 ( 
.A(n_3324),
.Y(n_3726)
);

NOR2xp33_ASAP7_75t_L g3727 ( 
.A(n_3392),
.B(n_1814),
.Y(n_3727)
);

AO22x2_ASAP7_75t_L g3728 ( 
.A1(n_3437),
.A2(n_2029),
.B1(n_2162),
.B2(n_1973),
.Y(n_3728)
);

BUFx3_ASAP7_75t_L g3729 ( 
.A(n_3327),
.Y(n_3729)
);

INVx4_ASAP7_75t_L g3730 ( 
.A(n_3336),
.Y(n_3730)
);

INVx3_ASAP7_75t_L g3731 ( 
.A(n_3509),
.Y(n_3731)
);

NAND3xp33_ASAP7_75t_L g3732 ( 
.A(n_3449),
.B(n_1821),
.C(n_1820),
.Y(n_3732)
);

INVx4_ASAP7_75t_L g3733 ( 
.A(n_3337),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_3512),
.Y(n_3734)
);

INVx3_ASAP7_75t_L g3735 ( 
.A(n_3513),
.Y(n_3735)
);

INVx2_ASAP7_75t_L g3736 ( 
.A(n_3517),
.Y(n_3736)
);

AOI22xp33_ASAP7_75t_L g3737 ( 
.A1(n_3325),
.A2(n_2225),
.B1(n_2238),
.B2(n_2216),
.Y(n_3737)
);

INVx2_ASAP7_75t_L g3738 ( 
.A(n_3319),
.Y(n_3738)
);

NAND2xp5_ASAP7_75t_SL g3739 ( 
.A(n_3450),
.B(n_1913),
.Y(n_3739)
);

INVx2_ASAP7_75t_L g3740 ( 
.A(n_3331),
.Y(n_3740)
);

BUFx6f_ASAP7_75t_SL g3741 ( 
.A(n_3339),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3340),
.Y(n_3742)
);

BUFx4f_ASAP7_75t_L g3743 ( 
.A(n_3344),
.Y(n_3743)
);

CKINVDCx5p33_ASAP7_75t_R g3744 ( 
.A(n_3348),
.Y(n_3744)
);

INVx4_ASAP7_75t_L g3745 ( 
.A(n_3349),
.Y(n_3745)
);

INVx2_ASAP7_75t_L g3746 ( 
.A(n_3342),
.Y(n_3746)
);

INVx6_ASAP7_75t_L g3747 ( 
.A(n_3356),
.Y(n_3747)
);

INVx2_ASAP7_75t_L g3748 ( 
.A(n_3417),
.Y(n_3748)
);

BUFx3_ASAP7_75t_L g3749 ( 
.A(n_3357),
.Y(n_3749)
);

OAI22xp5_ASAP7_75t_L g3750 ( 
.A1(n_3358),
.A2(n_2261),
.B1(n_2267),
.B2(n_2247),
.Y(n_3750)
);

AOI22xp33_ASAP7_75t_L g3751 ( 
.A1(n_3452),
.A2(n_2286),
.B1(n_2293),
.B2(n_2289),
.Y(n_3751)
);

AOI22xp33_ASAP7_75t_L g3752 ( 
.A1(n_3372),
.A2(n_2298),
.B1(n_2338),
.B2(n_2325),
.Y(n_3752)
);

AND2x4_ASAP7_75t_L g3753 ( 
.A(n_3361),
.B(n_3061),
.Y(n_3753)
);

INVx2_ASAP7_75t_L g3754 ( 
.A(n_3420),
.Y(n_3754)
);

OAI22xp33_ASAP7_75t_L g3755 ( 
.A1(n_3495),
.A2(n_2455),
.B1(n_2349),
.B2(n_2371),
.Y(n_3755)
);

NAND2xp5_ASAP7_75t_L g3756 ( 
.A(n_3398),
.B(n_2340),
.Y(n_3756)
);

BUFx2_ASAP7_75t_L g3757 ( 
.A(n_3326),
.Y(n_3757)
);

BUFx3_ASAP7_75t_L g3758 ( 
.A(n_3385),
.Y(n_3758)
);

INVx4_ASAP7_75t_L g3759 ( 
.A(n_3360),
.Y(n_3759)
);

INVx5_ASAP7_75t_L g3760 ( 
.A(n_3484),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3293),
.Y(n_3761)
);

INVx4_ASAP7_75t_SL g3762 ( 
.A(n_3413),
.Y(n_3762)
);

NAND2xp5_ASAP7_75t_L g3763 ( 
.A(n_3398),
.B(n_2383),
.Y(n_3763)
);

AND2x2_ASAP7_75t_L g3764 ( 
.A(n_3375),
.B(n_3062),
.Y(n_3764)
);

INVx3_ASAP7_75t_L g3765 ( 
.A(n_3302),
.Y(n_3765)
);

INVxp67_ASAP7_75t_L g3766 ( 
.A(n_3375),
.Y(n_3766)
);

INVx2_ASAP7_75t_L g3767 ( 
.A(n_3420),
.Y(n_3767)
);

NOR2xp33_ASAP7_75t_L g3768 ( 
.A(n_3315),
.B(n_1823),
.Y(n_3768)
);

NOR2xp33_ASAP7_75t_L g3769 ( 
.A(n_3315),
.B(n_1826),
.Y(n_3769)
);

NAND2xp5_ASAP7_75t_SL g3770 ( 
.A(n_3346),
.B(n_1914),
.Y(n_3770)
);

BUFx6f_ASAP7_75t_L g3771 ( 
.A(n_3302),
.Y(n_3771)
);

AND2x2_ASAP7_75t_SL g3772 ( 
.A(n_3469),
.B(n_1767),
.Y(n_3772)
);

INVx2_ASAP7_75t_L g3773 ( 
.A(n_3420),
.Y(n_3773)
);

NOR2xp33_ASAP7_75t_L g3774 ( 
.A(n_3315),
.B(n_1828),
.Y(n_3774)
);

OAI22xp5_ASAP7_75t_L g3775 ( 
.A1(n_3398),
.A2(n_2395),
.B1(n_2430),
.B2(n_2386),
.Y(n_3775)
);

INVx1_ASAP7_75t_L g3776 ( 
.A(n_3293),
.Y(n_3776)
);

NOR2xp33_ASAP7_75t_L g3777 ( 
.A(n_3315),
.B(n_1831),
.Y(n_3777)
);

NOR2xp33_ASAP7_75t_L g3778 ( 
.A(n_3315),
.B(n_1837),
.Y(n_3778)
);

BUFx2_ASAP7_75t_L g3779 ( 
.A(n_3326),
.Y(n_3779)
);

AND2x2_ASAP7_75t_L g3780 ( 
.A(n_3375),
.B(n_3065),
.Y(n_3780)
);

NAND2xp5_ASAP7_75t_L g3781 ( 
.A(n_3398),
.B(n_2434),
.Y(n_3781)
);

NOR2xp33_ASAP7_75t_L g3782 ( 
.A(n_3315),
.B(n_1839),
.Y(n_3782)
);

NAND2xp5_ASAP7_75t_SL g3783 ( 
.A(n_3346),
.B(n_1915),
.Y(n_3783)
);

OR2x2_ASAP7_75t_L g3784 ( 
.A(n_3375),
.B(n_3066),
.Y(n_3784)
);

OAI21xp33_ASAP7_75t_SL g3785 ( 
.A1(n_3303),
.A2(n_2438),
.B(n_2347),
.Y(n_3785)
);

INVx4_ASAP7_75t_L g3786 ( 
.A(n_3360),
.Y(n_3786)
);

INVx2_ASAP7_75t_SL g3787 ( 
.A(n_3375),
.Y(n_3787)
);

OR2x6_ASAP7_75t_L g3788 ( 
.A(n_3323),
.B(n_2447),
.Y(n_3788)
);

BUFx3_ASAP7_75t_L g3789 ( 
.A(n_3385),
.Y(n_3789)
);

AOI22xp5_ASAP7_75t_L g3790 ( 
.A1(n_3315),
.A2(n_1919),
.B1(n_1921),
.B2(n_1918),
.Y(n_3790)
);

NAND2xp5_ASAP7_75t_L g3791 ( 
.A(n_3398),
.B(n_2439),
.Y(n_3791)
);

AND2x2_ASAP7_75t_L g3792 ( 
.A(n_3375),
.B(n_3067),
.Y(n_3792)
);

AND2x2_ASAP7_75t_L g3793 ( 
.A(n_3375),
.B(n_3069),
.Y(n_3793)
);

NOR2xp33_ASAP7_75t_SL g3794 ( 
.A(n_3447),
.B(n_2244),
.Y(n_3794)
);

NOR2xp33_ASAP7_75t_L g3795 ( 
.A(n_3315),
.B(n_1845),
.Y(n_3795)
);

INVxp67_ASAP7_75t_SL g3796 ( 
.A(n_3427),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_L g3797 ( 
.A(n_3398),
.B(n_2442),
.Y(n_3797)
);

BUFx2_ASAP7_75t_L g3798 ( 
.A(n_3326),
.Y(n_3798)
);

NAND2xp5_ASAP7_75t_L g3799 ( 
.A(n_3398),
.B(n_2452),
.Y(n_3799)
);

NAND2xp5_ASAP7_75t_L g3800 ( 
.A(n_3398),
.B(n_2459),
.Y(n_3800)
);

INVxp67_ASAP7_75t_SL g3801 ( 
.A(n_3427),
.Y(n_3801)
);

INVx3_ASAP7_75t_L g3802 ( 
.A(n_3302),
.Y(n_3802)
);

NAND2xp5_ASAP7_75t_L g3803 ( 
.A(n_3398),
.B(n_2467),
.Y(n_3803)
);

INVx1_ASAP7_75t_L g3804 ( 
.A(n_3293),
.Y(n_3804)
);

INVx4_ASAP7_75t_L g3805 ( 
.A(n_3360),
.Y(n_3805)
);

NAND2xp5_ASAP7_75t_SL g3806 ( 
.A(n_3346),
.B(n_1930),
.Y(n_3806)
);

INVx1_ASAP7_75t_L g3807 ( 
.A(n_3293),
.Y(n_3807)
);

BUFx2_ASAP7_75t_L g3808 ( 
.A(n_3326),
.Y(n_3808)
);

INVx5_ASAP7_75t_L g3809 ( 
.A(n_3484),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_L g3810 ( 
.A(n_3398),
.B(n_2470),
.Y(n_3810)
);

INVx4_ASAP7_75t_L g3811 ( 
.A(n_3360),
.Y(n_3811)
);

INVx2_ASAP7_75t_SL g3812 ( 
.A(n_3375),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3293),
.Y(n_3813)
);

NAND2xp5_ASAP7_75t_SL g3814 ( 
.A(n_3346),
.B(n_1931),
.Y(n_3814)
);

INVx1_ASAP7_75t_L g3815 ( 
.A(n_3293),
.Y(n_3815)
);

NOR2xp33_ASAP7_75t_L g3816 ( 
.A(n_3315),
.B(n_1847),
.Y(n_3816)
);

NAND2xp5_ASAP7_75t_L g3817 ( 
.A(n_3398),
.B(n_2484),
.Y(n_3817)
);

HB1xp67_ASAP7_75t_L g3818 ( 
.A(n_3375),
.Y(n_3818)
);

O2A1O1Ixp5_ASAP7_75t_L g3819 ( 
.A1(n_3707),
.A2(n_2531),
.B(n_2536),
.C(n_2516),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_3568),
.B(n_2554),
.Y(n_3820)
);

INVx2_ASAP7_75t_SL g3821 ( 
.A(n_3590),
.Y(n_3821)
);

NAND2xp5_ASAP7_75t_SL g3822 ( 
.A(n_3623),
.B(n_1936),
.Y(n_3822)
);

INVx2_ASAP7_75t_L g3823 ( 
.A(n_3519),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_SL g3824 ( 
.A(n_3648),
.B(n_1937),
.Y(n_3824)
);

NAND2xp5_ASAP7_75t_SL g3825 ( 
.A(n_3556),
.B(n_3768),
.Y(n_3825)
);

NOR2xp33_ASAP7_75t_L g3826 ( 
.A(n_3566),
.B(n_2280),
.Y(n_3826)
);

A2O1A1Ixp33_ASAP7_75t_L g3827 ( 
.A1(n_3769),
.A2(n_2572),
.B(n_2603),
.C(n_2557),
.Y(n_3827)
);

INVx1_ASAP7_75t_L g3828 ( 
.A(n_3529),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_SL g3829 ( 
.A(n_3774),
.B(n_1948),
.Y(n_3829)
);

NAND2xp5_ASAP7_75t_L g3830 ( 
.A(n_3777),
.B(n_2607),
.Y(n_3830)
);

HB1xp67_ASAP7_75t_L g3831 ( 
.A(n_3574),
.Y(n_3831)
);

AND2x2_ASAP7_75t_L g3832 ( 
.A(n_3563),
.B(n_2232),
.Y(n_3832)
);

NAND2xp5_ASAP7_75t_SL g3833 ( 
.A(n_3778),
.B(n_1949),
.Y(n_3833)
);

NAND2xp5_ASAP7_75t_L g3834 ( 
.A(n_3782),
.B(n_2624),
.Y(n_3834)
);

AND2x6_ASAP7_75t_L g3835 ( 
.A(n_3537),
.B(n_2625),
.Y(n_3835)
);

INVx3_ASAP7_75t_L g3836 ( 
.A(n_3531),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_L g3837 ( 
.A(n_3795),
.B(n_2630),
.Y(n_3837)
);

INVx1_ASAP7_75t_L g3838 ( 
.A(n_3533),
.Y(n_3838)
);

NAND2x1p5_ASAP7_75t_L g3839 ( 
.A(n_3633),
.B(n_3071),
.Y(n_3839)
);

INVxp33_ASAP7_75t_SL g3840 ( 
.A(n_3528),
.Y(n_3840)
);

NAND2xp5_ASAP7_75t_SL g3841 ( 
.A(n_3816),
.B(n_1955),
.Y(n_3841)
);

NAND2xp5_ASAP7_75t_SL g3842 ( 
.A(n_3603),
.B(n_3787),
.Y(n_3842)
);

AND2x2_ASAP7_75t_L g3843 ( 
.A(n_3551),
.B(n_2232),
.Y(n_3843)
);

INVx1_ASAP7_75t_L g3844 ( 
.A(n_3544),
.Y(n_3844)
);

NAND2xp5_ASAP7_75t_L g3845 ( 
.A(n_3538),
.B(n_2674),
.Y(n_3845)
);

NAND2xp5_ASAP7_75t_L g3846 ( 
.A(n_3570),
.B(n_2678),
.Y(n_3846)
);

INVx2_ASAP7_75t_L g3847 ( 
.A(n_3530),
.Y(n_3847)
);

INVx2_ASAP7_75t_L g3848 ( 
.A(n_3557),
.Y(n_3848)
);

NOR2x1p5_ASAP7_75t_L g3849 ( 
.A(n_3569),
.B(n_1850),
.Y(n_3849)
);

NOR2xp33_ASAP7_75t_L g3850 ( 
.A(n_3628),
.B(n_2327),
.Y(n_3850)
);

AOI22xp5_ASAP7_75t_L g3851 ( 
.A1(n_3669),
.A2(n_2692),
.B1(n_2695),
.B2(n_2689),
.Y(n_3851)
);

INVxp67_ASAP7_75t_L g3852 ( 
.A(n_3608),
.Y(n_3852)
);

NOR2xp33_ASAP7_75t_L g3853 ( 
.A(n_3766),
.B(n_2492),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_3546),
.Y(n_3854)
);

HB1xp67_ASAP7_75t_L g3855 ( 
.A(n_3757),
.Y(n_3855)
);

CKINVDCx5p33_ASAP7_75t_R g3856 ( 
.A(n_3540),
.Y(n_3856)
);

NOR3xp33_ASAP7_75t_L g3857 ( 
.A(n_3673),
.B(n_3075),
.C(n_3073),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_L g3858 ( 
.A(n_3796),
.B(n_2722),
.Y(n_3858)
);

INVx2_ASAP7_75t_L g3859 ( 
.A(n_3560),
.Y(n_3859)
);

NAND2xp5_ASAP7_75t_L g3860 ( 
.A(n_3801),
.B(n_2735),
.Y(n_3860)
);

NOR2xp33_ASAP7_75t_L g3861 ( 
.A(n_3812),
.B(n_2512),
.Y(n_3861)
);

INVx1_ASAP7_75t_SL g3862 ( 
.A(n_3779),
.Y(n_3862)
);

NAND2xp5_ASAP7_75t_L g3863 ( 
.A(n_3527),
.B(n_2743),
.Y(n_3863)
);

NAND2xp5_ASAP7_75t_L g3864 ( 
.A(n_3756),
.B(n_3763),
.Y(n_3864)
);

INVx1_ASAP7_75t_L g3865 ( 
.A(n_3554),
.Y(n_3865)
);

AOI22xp33_ASAP7_75t_L g3866 ( 
.A1(n_3775),
.A2(n_2754),
.B1(n_2759),
.B2(n_2747),
.Y(n_3866)
);

AOI21xp5_ASAP7_75t_L g3867 ( 
.A1(n_3698),
.A2(n_2817),
.B(n_2761),
.Y(n_3867)
);

INVx1_ASAP7_75t_L g3868 ( 
.A(n_3562),
.Y(n_3868)
);

NOR2xp67_ASAP7_75t_L g3869 ( 
.A(n_3691),
.B(n_3076),
.Y(n_3869)
);

NOR2xp33_ASAP7_75t_SL g3870 ( 
.A(n_3656),
.B(n_2544),
.Y(n_3870)
);

OR2x2_ASAP7_75t_L g3871 ( 
.A(n_3582),
.B(n_3077),
.Y(n_3871)
);

NOR2xp33_ASAP7_75t_L g3872 ( 
.A(n_3676),
.B(n_2573),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_SL g3873 ( 
.A(n_3705),
.B(n_1957),
.Y(n_3873)
);

NAND2xp5_ASAP7_75t_SL g3874 ( 
.A(n_3781),
.B(n_1964),
.Y(n_3874)
);

NAND2xp5_ASAP7_75t_L g3875 ( 
.A(n_3791),
.B(n_1969),
.Y(n_3875)
);

NAND2xp5_ASAP7_75t_L g3876 ( 
.A(n_3797),
.B(n_1976),
.Y(n_3876)
);

BUFx12f_ASAP7_75t_L g3877 ( 
.A(n_3632),
.Y(n_3877)
);

NAND2xp5_ASAP7_75t_L g3878 ( 
.A(n_3799),
.B(n_1990),
.Y(n_3878)
);

NAND2xp5_ASAP7_75t_L g3879 ( 
.A(n_3800),
.B(n_1994),
.Y(n_3879)
);

NOR2xp33_ASAP7_75t_SL g3880 ( 
.A(n_3610),
.B(n_2576),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_3572),
.Y(n_3881)
);

AO22x1_ASAP7_75t_L g3882 ( 
.A1(n_3580),
.A2(n_1861),
.B1(n_1862),
.B2(n_1856),
.Y(n_3882)
);

NOR3xp33_ASAP7_75t_L g3883 ( 
.A(n_3520),
.B(n_3078),
.C(n_2471),
.Y(n_3883)
);

NAND2xp5_ASAP7_75t_L g3884 ( 
.A(n_3803),
.B(n_1996),
.Y(n_3884)
);

INVx2_ASAP7_75t_L g3885 ( 
.A(n_3754),
.Y(n_3885)
);

INVxp67_ASAP7_75t_SL g3886 ( 
.A(n_3818),
.Y(n_3886)
);

NAND2xp5_ASAP7_75t_SL g3887 ( 
.A(n_3810),
.B(n_2009),
.Y(n_3887)
);

NOR2xp33_ASAP7_75t_L g3888 ( 
.A(n_3637),
.B(n_2604),
.Y(n_3888)
);

NAND2xp5_ASAP7_75t_L g3889 ( 
.A(n_3817),
.B(n_2011),
.Y(n_3889)
);

NOR3xp33_ASAP7_75t_L g3890 ( 
.A(n_3722),
.B(n_2497),
.C(n_2465),
.Y(n_3890)
);

AND2x2_ASAP7_75t_L g3891 ( 
.A(n_3545),
.B(n_2372),
.Y(n_3891)
);

INVx1_ASAP7_75t_L g3892 ( 
.A(n_3573),
.Y(n_3892)
);

NAND2x1p5_ASAP7_75t_L g3893 ( 
.A(n_3598),
.B(n_2273),
.Y(n_3893)
);

NAND2xp33_ASAP7_75t_L g3894 ( 
.A(n_3710),
.B(n_2284),
.Y(n_3894)
);

INVx2_ASAP7_75t_L g3895 ( 
.A(n_3767),
.Y(n_3895)
);

NOR2xp33_ASAP7_75t_L g3896 ( 
.A(n_3541),
.B(n_2616),
.Y(n_3896)
);

NOR2xp33_ASAP7_75t_L g3897 ( 
.A(n_3798),
.B(n_2632),
.Y(n_3897)
);

NAND2xp5_ASAP7_75t_L g3898 ( 
.A(n_3542),
.B(n_2017),
.Y(n_3898)
);

NOR2xp33_ASAP7_75t_L g3899 ( 
.A(n_3808),
.B(n_2700),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_L g3900 ( 
.A(n_3532),
.B(n_2020),
.Y(n_3900)
);

HB1xp67_ASAP7_75t_L g3901 ( 
.A(n_3596),
.Y(n_3901)
);

NAND2xp5_ASAP7_75t_L g3902 ( 
.A(n_3764),
.B(n_2021),
.Y(n_3902)
);

AOI22xp33_ASAP7_75t_L g3903 ( 
.A1(n_3565),
.A2(n_2533),
.B1(n_2391),
.B2(n_2494),
.Y(n_3903)
);

INVx2_ASAP7_75t_L g3904 ( 
.A(n_3773),
.Y(n_3904)
);

INVx1_ASAP7_75t_L g3905 ( 
.A(n_3576),
.Y(n_3905)
);

BUFx6f_ASAP7_75t_L g3906 ( 
.A(n_3531),
.Y(n_3906)
);

NOR3xp33_ASAP7_75t_L g3907 ( 
.A(n_3525),
.B(n_2568),
.C(n_2509),
.Y(n_3907)
);

AOI22xp5_ASAP7_75t_L g3908 ( 
.A1(n_3718),
.A2(n_2030),
.B1(n_2032),
.B2(n_2028),
.Y(n_3908)
);

NAND2xp5_ASAP7_75t_L g3909 ( 
.A(n_3780),
.B(n_2034),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3577),
.Y(n_3910)
);

AND2x2_ASAP7_75t_SL g3911 ( 
.A(n_3794),
.B(n_1903),
.Y(n_3911)
);

NAND2xp5_ASAP7_75t_L g3912 ( 
.A(n_3792),
.B(n_2051),
.Y(n_3912)
);

INVx2_ASAP7_75t_L g3913 ( 
.A(n_3581),
.Y(n_3913)
);

INVx1_ASAP7_75t_L g3914 ( 
.A(n_3583),
.Y(n_3914)
);

INVx2_ASAP7_75t_L g3915 ( 
.A(n_3588),
.Y(n_3915)
);

AOI22xp33_ASAP7_75t_L g3916 ( 
.A1(n_3584),
.A2(n_2533),
.B1(n_2391),
.B2(n_2494),
.Y(n_3916)
);

NOR2xp33_ASAP7_75t_L g3917 ( 
.A(n_3589),
.B(n_2702),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3591),
.Y(n_3918)
);

INVx2_ASAP7_75t_L g3919 ( 
.A(n_3621),
.Y(n_3919)
);

NAND2xp5_ASAP7_75t_SL g3920 ( 
.A(n_3793),
.B(n_2054),
.Y(n_3920)
);

INVx2_ASAP7_75t_L g3921 ( 
.A(n_3634),
.Y(n_3921)
);

INVx2_ASAP7_75t_L g3922 ( 
.A(n_3636),
.Y(n_3922)
);

CKINVDCx5p33_ASAP7_75t_R g3923 ( 
.A(n_3594),
.Y(n_3923)
);

NAND2x1p5_ASAP7_75t_L g3924 ( 
.A(n_3522),
.B(n_2273),
.Y(n_3924)
);

INVx2_ASAP7_75t_L g3925 ( 
.A(n_3641),
.Y(n_3925)
);

NAND2xp5_ASAP7_75t_L g3926 ( 
.A(n_3535),
.B(n_2062),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3646),
.Y(n_3927)
);

INVx2_ASAP7_75t_L g3928 ( 
.A(n_3651),
.Y(n_3928)
);

OAI22xp5_ASAP7_75t_L g3929 ( 
.A1(n_3709),
.A2(n_2724),
.B1(n_2752),
.B2(n_2708),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_SL g3930 ( 
.A(n_3658),
.B(n_2065),
.Y(n_3930)
);

O2A1O1Ixp5_ASAP7_75t_L g3931 ( 
.A1(n_3720),
.A2(n_1916),
.B(n_1917),
.C(n_1911),
.Y(n_3931)
);

NOR2xp33_ASAP7_75t_L g3932 ( 
.A(n_3652),
.B(n_2795),
.Y(n_3932)
);

NOR2xp33_ASAP7_75t_L g3933 ( 
.A(n_3521),
.B(n_2813),
.Y(n_3933)
);

INVx1_ASAP7_75t_L g3934 ( 
.A(n_3761),
.Y(n_3934)
);

INVx1_ASAP7_75t_L g3935 ( 
.A(n_3776),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_3804),
.Y(n_3936)
);

INVx2_ASAP7_75t_L g3937 ( 
.A(n_3807),
.Y(n_3937)
);

INVxp67_ASAP7_75t_L g3938 ( 
.A(n_3645),
.Y(n_3938)
);

NAND2xp5_ASAP7_75t_L g3939 ( 
.A(n_3625),
.B(n_2068),
.Y(n_3939)
);

NAND2xp5_ASAP7_75t_L g3940 ( 
.A(n_3626),
.B(n_2071),
.Y(n_3940)
);

NAND2xp5_ASAP7_75t_L g3941 ( 
.A(n_3647),
.B(n_2080),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_SL g3942 ( 
.A(n_3691),
.B(n_2083),
.Y(n_3942)
);

INVx2_ASAP7_75t_L g3943 ( 
.A(n_3813),
.Y(n_3943)
);

NAND2xp5_ASAP7_75t_SL g3944 ( 
.A(n_3815),
.B(n_2098),
.Y(n_3944)
);

NAND2xp5_ASAP7_75t_SL g3945 ( 
.A(n_3543),
.B(n_2101),
.Y(n_3945)
);

NAND2xp5_ASAP7_75t_L g3946 ( 
.A(n_3558),
.B(n_2102),
.Y(n_3946)
);

INVx1_ASAP7_75t_L g3947 ( 
.A(n_3654),
.Y(n_3947)
);

NAND2xp5_ASAP7_75t_L g3948 ( 
.A(n_3564),
.B(n_2104),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_L g3949 ( 
.A(n_3679),
.B(n_2105),
.Y(n_3949)
);

O2A1O1Ixp5_ASAP7_75t_L g3950 ( 
.A1(n_3686),
.A2(n_2058),
.B(n_2103),
.C(n_2045),
.Y(n_3950)
);

OR2x6_ASAP7_75t_L g3951 ( 
.A(n_3597),
.B(n_2652),
.Y(n_3951)
);

AOI22xp5_ASAP7_75t_L g3952 ( 
.A1(n_3785),
.A2(n_2107),
.B1(n_2110),
.B2(n_2106),
.Y(n_3952)
);

NAND2xp5_ASAP7_75t_SL g3953 ( 
.A(n_3543),
.B(n_2116),
.Y(n_3953)
);

NOR2xp33_ASAP7_75t_L g3954 ( 
.A(n_3784),
.B(n_1864),
.Y(n_3954)
);

NAND2xp5_ASAP7_75t_SL g3955 ( 
.A(n_3547),
.B(n_2118),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_L g3956 ( 
.A(n_3662),
.B(n_2121),
.Y(n_3956)
);

NAND2xp5_ASAP7_75t_SL g3957 ( 
.A(n_3547),
.B(n_2130),
.Y(n_3957)
);

INVxp67_ASAP7_75t_SL g3958 ( 
.A(n_3567),
.Y(n_3958)
);

AND2x4_ASAP7_75t_L g3959 ( 
.A(n_3534),
.B(n_2384),
.Y(n_3959)
);

INVx2_ASAP7_75t_L g3960 ( 
.A(n_3715),
.Y(n_3960)
);

O2A1O1Ixp5_ASAP7_75t_L g3961 ( 
.A1(n_3748),
.A2(n_2136),
.B(n_2218),
.C(n_2142),
.Y(n_3961)
);

INVx2_ASAP7_75t_L g3962 ( 
.A(n_3716),
.Y(n_3962)
);

AND2x4_ASAP7_75t_L g3963 ( 
.A(n_3539),
.B(n_2419),
.Y(n_3963)
);

NAND2xp5_ASAP7_75t_SL g3964 ( 
.A(n_3760),
.B(n_2135),
.Y(n_3964)
);

CKINVDCx5p33_ASAP7_75t_R g3965 ( 
.A(n_3555),
.Y(n_3965)
);

INVx1_ASAP7_75t_L g3966 ( 
.A(n_3657),
.Y(n_3966)
);

OAI221xp5_ASAP7_75t_L g3967 ( 
.A1(n_3609),
.A2(n_2706),
.B1(n_2685),
.B2(n_2423),
.C(n_2428),
.Y(n_3967)
);

O2A1O1Ixp33_ASAP7_75t_L g3968 ( 
.A1(n_3755),
.A2(n_2422),
.B(n_2448),
.C(n_2420),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_L g3969 ( 
.A(n_3607),
.B(n_2140),
.Y(n_3969)
);

BUFx12f_ASAP7_75t_L g3970 ( 
.A(n_3618),
.Y(n_3970)
);

INVx2_ASAP7_75t_L g3971 ( 
.A(n_3717),
.Y(n_3971)
);

INVxp67_ASAP7_75t_L g3972 ( 
.A(n_3640),
.Y(n_3972)
);

NAND2xp5_ASAP7_75t_L g3973 ( 
.A(n_3629),
.B(n_2148),
.Y(n_3973)
);

INVxp33_ASAP7_75t_L g3974 ( 
.A(n_3667),
.Y(n_3974)
);

NOR2xp33_ASAP7_75t_L g3975 ( 
.A(n_3790),
.B(n_1868),
.Y(n_3975)
);

NAND2xp5_ASAP7_75t_SL g3976 ( 
.A(n_3760),
.B(n_2151),
.Y(n_3976)
);

NAND2xp33_ASAP7_75t_L g3977 ( 
.A(n_3649),
.B(n_2533),
.Y(n_3977)
);

INVx1_ASAP7_75t_L g3978 ( 
.A(n_3665),
.Y(n_3978)
);

AOI22xp5_ASAP7_75t_L g3979 ( 
.A1(n_3578),
.A2(n_2163),
.B1(n_2165),
.B2(n_2161),
.Y(n_3979)
);

NAND2xp5_ASAP7_75t_L g3980 ( 
.A(n_3630),
.B(n_2166),
.Y(n_3980)
);

NAND3xp33_ASAP7_75t_L g3981 ( 
.A(n_3725),
.B(n_1870),
.C(n_1869),
.Y(n_3981)
);

INVxp67_ASAP7_75t_L g3982 ( 
.A(n_3642),
.Y(n_3982)
);

INVxp33_ASAP7_75t_L g3983 ( 
.A(n_3567),
.Y(n_3983)
);

NAND2xp5_ASAP7_75t_L g3984 ( 
.A(n_3631),
.B(n_2168),
.Y(n_3984)
);

INVx2_ASAP7_75t_L g3985 ( 
.A(n_3723),
.Y(n_3985)
);

NOR2xp33_ASAP7_75t_L g3986 ( 
.A(n_3727),
.B(n_3552),
.Y(n_3986)
);

INVx2_ASAP7_75t_L g3987 ( 
.A(n_3736),
.Y(n_3987)
);

INVx2_ASAP7_75t_SL g3988 ( 
.A(n_3606),
.Y(n_3988)
);

INVx2_ASAP7_75t_L g3989 ( 
.A(n_3604),
.Y(n_3989)
);

NAND2xp5_ASAP7_75t_SL g3990 ( 
.A(n_3809),
.B(n_2172),
.Y(n_3990)
);

AND2x2_ASAP7_75t_L g3991 ( 
.A(n_3758),
.B(n_2372),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_3668),
.Y(n_3992)
);

NAND2xp5_ASAP7_75t_L g3993 ( 
.A(n_3635),
.B(n_2179),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_L g3994 ( 
.A(n_3638),
.B(n_2180),
.Y(n_3994)
);

AND2x4_ASAP7_75t_SL g3995 ( 
.A(n_3523),
.B(n_2636),
.Y(n_3995)
);

NAND2xp5_ASAP7_75t_SL g3996 ( 
.A(n_3809),
.B(n_3653),
.Y(n_3996)
);

NAND2xp5_ASAP7_75t_L g3997 ( 
.A(n_3643),
.B(n_2185),
.Y(n_3997)
);

INVx1_ASAP7_75t_L g3998 ( 
.A(n_3677),
.Y(n_3998)
);

AND2x2_ASAP7_75t_L g3999 ( 
.A(n_3789),
.B(n_2636),
.Y(n_3999)
);

INVx1_ASAP7_75t_L g4000 ( 
.A(n_3681),
.Y(n_4000)
);

NAND2xp5_ASAP7_75t_L g4001 ( 
.A(n_3671),
.B(n_2197),
.Y(n_4001)
);

NAND2x1p5_ASAP7_75t_L g4002 ( 
.A(n_3550),
.B(n_3561),
.Y(n_4002)
);

INVx2_ASAP7_75t_SL g4003 ( 
.A(n_3624),
.Y(n_4003)
);

INVx4_ASAP7_75t_L g4004 ( 
.A(n_3599),
.Y(n_4004)
);

NAND3xp33_ASAP7_75t_L g4005 ( 
.A(n_3732),
.B(n_1875),
.C(n_1874),
.Y(n_4005)
);

NOR2xp33_ASAP7_75t_L g4006 ( 
.A(n_3770),
.B(n_1876),
.Y(n_4006)
);

AND2x2_ASAP7_75t_L g4007 ( 
.A(n_3548),
.B(n_2794),
.Y(n_4007)
);

AND2x4_ASAP7_75t_L g4008 ( 
.A(n_3526),
.B(n_2451),
.Y(n_4008)
);

NAND2xp5_ASAP7_75t_L g4009 ( 
.A(n_3674),
.B(n_2203),
.Y(n_4009)
);

NOR2xp33_ASAP7_75t_L g4010 ( 
.A(n_3783),
.B(n_1877),
.Y(n_4010)
);

O2A1O1Ixp33_ASAP7_75t_L g4011 ( 
.A1(n_3559),
.A2(n_3612),
.B(n_3613),
.C(n_3587),
.Y(n_4011)
);

INVx2_ASAP7_75t_L g4012 ( 
.A(n_3611),
.Y(n_4012)
);

NOR2xp33_ASAP7_75t_SL g4013 ( 
.A(n_3549),
.B(n_2794),
.Y(n_4013)
);

INVx2_ASAP7_75t_SL g4014 ( 
.A(n_3599),
.Y(n_4014)
);

AND2x2_ASAP7_75t_L g4015 ( 
.A(n_3682),
.B(n_1881),
.Y(n_4015)
);

INVx1_ASAP7_75t_L g4016 ( 
.A(n_3687),
.Y(n_4016)
);

NOR2xp67_ASAP7_75t_L g4017 ( 
.A(n_3571),
.B(n_2206),
.Y(n_4017)
);

NAND2xp5_ASAP7_75t_L g4018 ( 
.A(n_3675),
.B(n_3678),
.Y(n_4018)
);

NAND2xp5_ASAP7_75t_L g4019 ( 
.A(n_3680),
.B(n_2209),
.Y(n_4019)
);

INVxp67_ASAP7_75t_L g4020 ( 
.A(n_3806),
.Y(n_4020)
);

AOI22xp5_ASAP7_75t_L g4021 ( 
.A1(n_3690),
.A2(n_2213),
.B1(n_2220),
.B2(n_2210),
.Y(n_4021)
);

OAI22xp5_ASAP7_75t_L g4022 ( 
.A1(n_3737),
.A2(n_2228),
.B1(n_2231),
.B2(n_2221),
.Y(n_4022)
);

NAND2xp5_ASAP7_75t_SL g4023 ( 
.A(n_3689),
.B(n_2234),
.Y(n_4023)
);

INVx1_ASAP7_75t_L g4024 ( 
.A(n_3692),
.Y(n_4024)
);

NAND2xp5_ASAP7_75t_SL g4025 ( 
.A(n_3688),
.B(n_3605),
.Y(n_4025)
);

INVx1_ASAP7_75t_L g4026 ( 
.A(n_3696),
.Y(n_4026)
);

INVx1_ASAP7_75t_L g4027 ( 
.A(n_3697),
.Y(n_4027)
);

INVx2_ASAP7_75t_L g4028 ( 
.A(n_3619),
.Y(n_4028)
);

AND2x4_ASAP7_75t_L g4029 ( 
.A(n_3762),
.B(n_2461),
.Y(n_4029)
);

NOR2xp33_ASAP7_75t_L g4030 ( 
.A(n_3814),
.B(n_1884),
.Y(n_4030)
);

AOI22xp5_ASAP7_75t_L g4031 ( 
.A1(n_3701),
.A2(n_2240),
.B1(n_2246),
.B2(n_2237),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_L g4032 ( 
.A(n_3683),
.B(n_2257),
.Y(n_4032)
);

INVx2_ASAP7_75t_L g4033 ( 
.A(n_3700),
.Y(n_4033)
);

NAND2xp5_ASAP7_75t_L g4034 ( 
.A(n_3592),
.B(n_2260),
.Y(n_4034)
);

NAND2xp5_ASAP7_75t_SL g4035 ( 
.A(n_3644),
.B(n_2266),
.Y(n_4035)
);

NAND2xp33_ASAP7_75t_L g4036 ( 
.A(n_3649),
.B(n_2533),
.Y(n_4036)
);

INVxp67_ASAP7_75t_L g4037 ( 
.A(n_3585),
.Y(n_4037)
);

NAND2xp5_ASAP7_75t_L g4038 ( 
.A(n_3615),
.B(n_2268),
.Y(n_4038)
);

INVx1_ASAP7_75t_L g4039 ( 
.A(n_3704),
.Y(n_4039)
);

INVx2_ASAP7_75t_L g4040 ( 
.A(n_3708),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_L g4041 ( 
.A(n_3622),
.B(n_3734),
.Y(n_4041)
);

INVx1_ASAP7_75t_L g4042 ( 
.A(n_3738),
.Y(n_4042)
);

AND2x2_ASAP7_75t_L g4043 ( 
.A(n_3593),
.B(n_1887),
.Y(n_4043)
);

INVx1_ASAP7_75t_L g4044 ( 
.A(n_3731),
.Y(n_4044)
);

NOR2xp33_ASAP7_75t_L g4045 ( 
.A(n_3663),
.B(n_1888),
.Y(n_4045)
);

INVx1_ASAP7_75t_L g4046 ( 
.A(n_3735),
.Y(n_4046)
);

INVx2_ASAP7_75t_L g4047 ( 
.A(n_3595),
.Y(n_4047)
);

AND2x2_ASAP7_75t_L g4048 ( 
.A(n_3536),
.B(n_1889),
.Y(n_4048)
);

INVx2_ASAP7_75t_L g4049 ( 
.A(n_3695),
.Y(n_4049)
);

AOI22xp33_ASAP7_75t_L g4050 ( 
.A1(n_3553),
.A2(n_2533),
.B1(n_2391),
.B2(n_2494),
.Y(n_4050)
);

NAND2xp5_ASAP7_75t_L g4051 ( 
.A(n_3740),
.B(n_2276),
.Y(n_4051)
);

NAND2xp5_ASAP7_75t_L g4052 ( 
.A(n_3655),
.B(n_2288),
.Y(n_4052)
);

NAND2xp5_ASAP7_75t_L g4053 ( 
.A(n_3659),
.B(n_2296),
.Y(n_4053)
);

INVxp67_ASAP7_75t_L g4054 ( 
.A(n_3585),
.Y(n_4054)
);

BUFx5_ASAP7_75t_L g4055 ( 
.A(n_3742),
.Y(n_4055)
);

A2O1A1Ixp33_ASAP7_75t_L g4056 ( 
.A1(n_3702),
.A2(n_2474),
.B(n_2475),
.C(n_2466),
.Y(n_4056)
);

INVx1_ASAP7_75t_L g4057 ( 
.A(n_3753),
.Y(n_4057)
);

INVx1_ASAP7_75t_L g4058 ( 
.A(n_3660),
.Y(n_4058)
);

BUFx3_ASAP7_75t_L g4059 ( 
.A(n_3771),
.Y(n_4059)
);

INVx2_ASAP7_75t_SL g4060 ( 
.A(n_3771),
.Y(n_4060)
);

INVx2_ASAP7_75t_L g4061 ( 
.A(n_3746),
.Y(n_4061)
);

NAND2xp5_ASAP7_75t_L g4062 ( 
.A(n_3672),
.B(n_3579),
.Y(n_4062)
);

NOR2xp67_ASAP7_75t_L g4063 ( 
.A(n_3759),
.B(n_2301),
.Y(n_4063)
);

INVx2_ASAP7_75t_SL g4064 ( 
.A(n_3575),
.Y(n_4064)
);

NAND2xp5_ASAP7_75t_L g4065 ( 
.A(n_3553),
.B(n_2312),
.Y(n_4065)
);

NAND2xp5_ASAP7_75t_SL g4066 ( 
.A(n_3693),
.B(n_2313),
.Y(n_4066)
);

A2O1A1Ixp33_ASAP7_75t_L g4067 ( 
.A1(n_3586),
.A2(n_2486),
.B(n_2493),
.C(n_2477),
.Y(n_4067)
);

INVx2_ASAP7_75t_L g4068 ( 
.A(n_3706),
.Y(n_4068)
);

INVx1_ASAP7_75t_L g4069 ( 
.A(n_3600),
.Y(n_4069)
);

INVx2_ASAP7_75t_L g4070 ( 
.A(n_3712),
.Y(n_4070)
);

NAND2xp5_ASAP7_75t_L g4071 ( 
.A(n_3666),
.B(n_2316),
.Y(n_4071)
);

NAND2xp5_ASAP7_75t_L g4072 ( 
.A(n_3714),
.B(n_3739),
.Y(n_4072)
);

NOR2xp33_ASAP7_75t_L g4073 ( 
.A(n_3744),
.B(n_1896),
.Y(n_4073)
);

INVx4_ASAP7_75t_L g4074 ( 
.A(n_3786),
.Y(n_4074)
);

A2O1A1Ixp33_ASAP7_75t_L g4075 ( 
.A1(n_3751),
.A2(n_2517),
.B(n_2535),
.C(n_2500),
.Y(n_4075)
);

INVx2_ASAP7_75t_L g4076 ( 
.A(n_3703),
.Y(n_4076)
);

AOI22xp5_ASAP7_75t_L g4077 ( 
.A1(n_3711),
.A2(n_2319),
.B1(n_2323),
.B2(n_2322),
.Y(n_4077)
);

NAND3xp33_ASAP7_75t_L g4078 ( 
.A(n_3617),
.B(n_1907),
.C(n_1899),
.Y(n_4078)
);

NAND2xp5_ASAP7_75t_SL g4079 ( 
.A(n_3743),
.B(n_2324),
.Y(n_4079)
);

INVx2_ASAP7_75t_L g4080 ( 
.A(n_3703),
.Y(n_4080)
);

NAND2xp5_ASAP7_75t_L g4081 ( 
.A(n_3627),
.B(n_2328),
.Y(n_4081)
);

INVx1_ASAP7_75t_L g4082 ( 
.A(n_3684),
.Y(n_4082)
);

NOR2xp33_ASAP7_75t_L g4083 ( 
.A(n_3730),
.B(n_1910),
.Y(n_4083)
);

OAI21xp5_ASAP7_75t_L g4084 ( 
.A1(n_3752),
.A2(n_2331),
.B(n_2330),
.Y(n_4084)
);

AOI22xp5_ASAP7_75t_L g4085 ( 
.A1(n_3719),
.A2(n_2334),
.B1(n_2346),
.B2(n_2339),
.Y(n_4085)
);

NAND2xp5_ASAP7_75t_L g4086 ( 
.A(n_3685),
.B(n_2348),
.Y(n_4086)
);

NAND2xp5_ASAP7_75t_SL g4087 ( 
.A(n_3772),
.B(n_2350),
.Y(n_4087)
);

INVx1_ASAP7_75t_L g4088 ( 
.A(n_3724),
.Y(n_4088)
);

NOR2xp33_ASAP7_75t_L g4089 ( 
.A(n_3733),
.B(n_1912),
.Y(n_4089)
);

INVx1_ASAP7_75t_L g4090 ( 
.A(n_3726),
.Y(n_4090)
);

INVxp67_ASAP7_75t_L g4091 ( 
.A(n_3602),
.Y(n_4091)
);

INVxp67_ASAP7_75t_SL g4092 ( 
.A(n_3524),
.Y(n_4092)
);

NAND2xp5_ASAP7_75t_L g4093 ( 
.A(n_3745),
.B(n_2352),
.Y(n_4093)
);

INVx1_ASAP7_75t_L g4094 ( 
.A(n_3729),
.Y(n_4094)
);

INVx5_ASAP7_75t_L g4095 ( 
.A(n_3650),
.Y(n_4095)
);

INVx2_ASAP7_75t_L g4096 ( 
.A(n_3713),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_SL g4097 ( 
.A(n_3620),
.B(n_2354),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_L g4098 ( 
.A(n_3713),
.B(n_2356),
.Y(n_4098)
);

NAND2xp5_ASAP7_75t_L g4099 ( 
.A(n_3721),
.B(n_2361),
.Y(n_4099)
);

INVx1_ASAP7_75t_L g4100 ( 
.A(n_3749),
.Y(n_4100)
);

INVx2_ASAP7_75t_L g4101 ( 
.A(n_3721),
.Y(n_4101)
);

NAND2xp5_ASAP7_75t_L g4102 ( 
.A(n_3728),
.B(n_2363),
.Y(n_4102)
);

AOI22xp5_ASAP7_75t_L g4103 ( 
.A1(n_3750),
.A2(n_2364),
.B1(n_2378),
.B2(n_2376),
.Y(n_4103)
);

BUFx6f_ASAP7_75t_L g4104 ( 
.A(n_3670),
.Y(n_4104)
);

NOR2xp33_ASAP7_75t_L g4105 ( 
.A(n_3805),
.B(n_1922),
.Y(n_4105)
);

BUFx3_ASAP7_75t_L g4106 ( 
.A(n_3601),
.Y(n_4106)
);

NAND2xp5_ASAP7_75t_L g4107 ( 
.A(n_3811),
.B(n_2382),
.Y(n_4107)
);

AOI22xp5_ASAP7_75t_L g4108 ( 
.A1(n_3747),
.A2(n_2385),
.B1(n_2389),
.B2(n_2387),
.Y(n_4108)
);

NAND2xp5_ASAP7_75t_SL g4109 ( 
.A(n_3670),
.B(n_2397),
.Y(n_4109)
);

NAND2xp5_ASAP7_75t_SL g4110 ( 
.A(n_3614),
.B(n_2405),
.Y(n_4110)
);

NAND2xp5_ASAP7_75t_SL g4111 ( 
.A(n_3639),
.B(n_2406),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_SL g4112 ( 
.A(n_3664),
.B(n_2407),
.Y(n_4112)
);

NOR2xp33_ASAP7_75t_L g4113 ( 
.A(n_3765),
.B(n_3802),
.Y(n_4113)
);

NAND2x1_ASAP7_75t_L g4114 ( 
.A(n_3788),
.B(n_2273),
.Y(n_4114)
);

INVx2_ASAP7_75t_SL g4115 ( 
.A(n_3616),
.Y(n_4115)
);

INVx2_ASAP7_75t_L g4116 ( 
.A(n_3741),
.Y(n_4116)
);

NAND2xp5_ASAP7_75t_SL g4117 ( 
.A(n_3694),
.B(n_2421),
.Y(n_4117)
);

INVx1_ASAP7_75t_L g4118 ( 
.A(n_3699),
.Y(n_4118)
);

CKINVDCx5p33_ASAP7_75t_R g4119 ( 
.A(n_3661),
.Y(n_4119)
);

INVx1_ASAP7_75t_L g4120 ( 
.A(n_3661),
.Y(n_4120)
);

BUFx2_ASAP7_75t_L g4121 ( 
.A(n_3590),
.Y(n_4121)
);

INVx2_ASAP7_75t_L g4122 ( 
.A(n_3519),
.Y(n_4122)
);

INVx1_ASAP7_75t_L g4123 ( 
.A(n_3529),
.Y(n_4123)
);

NAND2xp5_ASAP7_75t_SL g4124 ( 
.A(n_3623),
.B(n_2424),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_3529),
.Y(n_4125)
);

INVx2_ASAP7_75t_L g4126 ( 
.A(n_3519),
.Y(n_4126)
);

INVx1_ASAP7_75t_L g4127 ( 
.A(n_3529),
.Y(n_4127)
);

INVx1_ASAP7_75t_L g4128 ( 
.A(n_3529),
.Y(n_4128)
);

NAND2xp5_ASAP7_75t_L g4129 ( 
.A(n_3568),
.B(n_2429),
.Y(n_4129)
);

NAND2xp33_ASAP7_75t_L g4130 ( 
.A(n_3710),
.B(n_2432),
.Y(n_4130)
);

NAND2xp5_ASAP7_75t_SL g4131 ( 
.A(n_3623),
.B(n_2436),
.Y(n_4131)
);

NOR2xp67_ASAP7_75t_L g4132 ( 
.A(n_3540),
.B(n_2441),
.Y(n_4132)
);

NAND2xp5_ASAP7_75t_SL g4133 ( 
.A(n_3623),
.B(n_2449),
.Y(n_4133)
);

INVx1_ASAP7_75t_L g4134 ( 
.A(n_3529),
.Y(n_4134)
);

NAND2xp5_ASAP7_75t_L g4135 ( 
.A(n_3568),
.B(n_2450),
.Y(n_4135)
);

NAND2xp5_ASAP7_75t_SL g4136 ( 
.A(n_3623),
.B(n_2454),
.Y(n_4136)
);

INVx1_ASAP7_75t_L g4137 ( 
.A(n_3529),
.Y(n_4137)
);

NAND2xp5_ASAP7_75t_SL g4138 ( 
.A(n_3623),
.B(n_2456),
.Y(n_4138)
);

AND2x4_ASAP7_75t_L g4139 ( 
.A(n_3522),
.B(n_2539),
.Y(n_4139)
);

AOI22xp33_ASAP7_75t_L g4140 ( 
.A1(n_3566),
.A2(n_2709),
.B1(n_2787),
.B2(n_2555),
.Y(n_4140)
);

AOI22xp5_ASAP7_75t_L g4141 ( 
.A1(n_3768),
.A2(n_2472),
.B1(n_2479),
.B2(n_2457),
.Y(n_4141)
);

NAND2xp5_ASAP7_75t_L g4142 ( 
.A(n_3568),
.B(n_2488),
.Y(n_4142)
);

OR2x2_ASAP7_75t_L g4143 ( 
.A(n_3628),
.B(n_1926),
.Y(n_4143)
);

INVx2_ASAP7_75t_L g4144 ( 
.A(n_3519),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_3529),
.Y(n_4145)
);

CKINVDCx5p33_ASAP7_75t_R g4146 ( 
.A(n_3528),
.Y(n_4146)
);

INVx2_ASAP7_75t_L g4147 ( 
.A(n_3519),
.Y(n_4147)
);

NAND2xp5_ASAP7_75t_L g4148 ( 
.A(n_3568),
.B(n_2489),
.Y(n_4148)
);

NAND2xp5_ASAP7_75t_SL g4149 ( 
.A(n_3623),
.B(n_2503),
.Y(n_4149)
);

INVx2_ASAP7_75t_L g4150 ( 
.A(n_3519),
.Y(n_4150)
);

AOI21xp5_ASAP7_75t_L g4151 ( 
.A1(n_3538),
.A2(n_2709),
.B(n_2555),
.Y(n_4151)
);

INVx1_ASAP7_75t_L g4152 ( 
.A(n_3529),
.Y(n_4152)
);

NAND2xp5_ASAP7_75t_L g4153 ( 
.A(n_3568),
.B(n_2506),
.Y(n_4153)
);

NAND2xp5_ASAP7_75t_SL g4154 ( 
.A(n_3623),
.B(n_2515),
.Y(n_4154)
);

NAND2xp5_ASAP7_75t_L g4155 ( 
.A(n_3568),
.B(n_2528),
.Y(n_4155)
);

NAND2xp33_ASAP7_75t_L g4156 ( 
.A(n_3710),
.B(n_2529),
.Y(n_4156)
);

NAND2xp5_ASAP7_75t_L g4157 ( 
.A(n_3568),
.B(n_2543),
.Y(n_4157)
);

NAND2xp5_ASAP7_75t_L g4158 ( 
.A(n_3568),
.B(n_2552),
.Y(n_4158)
);

INVxp67_ASAP7_75t_L g4159 ( 
.A(n_3608),
.Y(n_4159)
);

INVx2_ASAP7_75t_L g4160 ( 
.A(n_3519),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_SL g4161 ( 
.A(n_3623),
.B(n_2556),
.Y(n_4161)
);

NAND2xp5_ASAP7_75t_L g4162 ( 
.A(n_3568),
.B(n_2561),
.Y(n_4162)
);

NAND2xp5_ASAP7_75t_SL g4163 ( 
.A(n_3623),
.B(n_2564),
.Y(n_4163)
);

NOR2xp33_ASAP7_75t_L g4164 ( 
.A(n_3566),
.B(n_1928),
.Y(n_4164)
);

NAND3xp33_ASAP7_75t_L g4165 ( 
.A(n_3566),
.B(n_1933),
.C(n_1932),
.Y(n_4165)
);

AND2x2_ASAP7_75t_L g4166 ( 
.A(n_3566),
.B(n_1939),
.Y(n_4166)
);

NAND2xp5_ASAP7_75t_SL g4167 ( 
.A(n_3623),
.B(n_2566),
.Y(n_4167)
);

NAND2xp5_ASAP7_75t_L g4168 ( 
.A(n_3568),
.B(n_2569),
.Y(n_4168)
);

NAND2xp5_ASAP7_75t_SL g4169 ( 
.A(n_3623),
.B(n_2577),
.Y(n_4169)
);

INVx1_ASAP7_75t_L g4170 ( 
.A(n_3529),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_3529),
.Y(n_4171)
);

NAND2x1p5_ASAP7_75t_L g4172 ( 
.A(n_3633),
.B(n_2555),
.Y(n_4172)
);

NAND2xp5_ASAP7_75t_SL g4173 ( 
.A(n_3623),
.B(n_2579),
.Y(n_4173)
);

NAND2xp5_ASAP7_75t_L g4174 ( 
.A(n_3568),
.B(n_2587),
.Y(n_4174)
);

INVx1_ASAP7_75t_L g4175 ( 
.A(n_3529),
.Y(n_4175)
);

NAND2xp5_ASAP7_75t_L g4176 ( 
.A(n_3568),
.B(n_2589),
.Y(n_4176)
);

INVx1_ASAP7_75t_L g4177 ( 
.A(n_3529),
.Y(n_4177)
);

OR2x2_ASAP7_75t_L g4178 ( 
.A(n_3862),
.B(n_1941),
.Y(n_4178)
);

INVx1_ASAP7_75t_L g4179 ( 
.A(n_3828),
.Y(n_4179)
);

NAND2xp5_ASAP7_75t_L g4180 ( 
.A(n_3864),
.B(n_4164),
.Y(n_4180)
);

NAND2xp5_ASAP7_75t_L g4181 ( 
.A(n_3825),
.B(n_2595),
.Y(n_4181)
);

NAND2xp5_ASAP7_75t_L g4182 ( 
.A(n_3852),
.B(n_4159),
.Y(n_4182)
);

INVx2_ASAP7_75t_SL g4183 ( 
.A(n_4121),
.Y(n_4183)
);

INVx2_ASAP7_75t_L g4184 ( 
.A(n_4061),
.Y(n_4184)
);

INVx1_ASAP7_75t_L g4185 ( 
.A(n_3838),
.Y(n_4185)
);

NAND2xp5_ASAP7_75t_L g4186 ( 
.A(n_3986),
.B(n_2605),
.Y(n_4186)
);

NAND2xp5_ASAP7_75t_L g4187 ( 
.A(n_3826),
.B(n_2612),
.Y(n_4187)
);

BUFx6f_ASAP7_75t_L g4188 ( 
.A(n_3906),
.Y(n_4188)
);

INVx1_ASAP7_75t_L g4189 ( 
.A(n_3844),
.Y(n_4189)
);

BUFx6f_ASAP7_75t_L g4190 ( 
.A(n_3906),
.Y(n_4190)
);

INVx2_ASAP7_75t_L g4191 ( 
.A(n_3915),
.Y(n_4191)
);

INVx2_ASAP7_75t_L g4192 ( 
.A(n_3919),
.Y(n_4192)
);

INVx4_ASAP7_75t_L g4193 ( 
.A(n_4104),
.Y(n_4193)
);

NAND2xp5_ASAP7_75t_L g4194 ( 
.A(n_4166),
.B(n_2614),
.Y(n_4194)
);

INVx2_ASAP7_75t_L g4195 ( 
.A(n_3921),
.Y(n_4195)
);

AOI22xp33_ASAP7_75t_L g4196 ( 
.A1(n_3872),
.A2(n_3932),
.B1(n_3830),
.B2(n_3837),
.Y(n_4196)
);

AOI22xp33_ASAP7_75t_L g4197 ( 
.A1(n_3834),
.A2(n_2787),
.B1(n_2709),
.B2(n_2621),
.Y(n_4197)
);

NAND2xp5_ASAP7_75t_L g4198 ( 
.A(n_4058),
.B(n_2620),
.Y(n_4198)
);

NOR2xp33_ASAP7_75t_L g4199 ( 
.A(n_3850),
.B(n_1942),
.Y(n_4199)
);

NAND2xp5_ASAP7_75t_L g4200 ( 
.A(n_3820),
.B(n_2635),
.Y(n_4200)
);

AOI22xp5_ASAP7_75t_L g4201 ( 
.A1(n_3896),
.A2(n_2643),
.B1(n_2647),
.B2(n_2637),
.Y(n_4201)
);

NOR2xp33_ASAP7_75t_L g4202 ( 
.A(n_3888),
.B(n_1950),
.Y(n_4202)
);

NAND3xp33_ASAP7_75t_SL g4203 ( 
.A(n_3870),
.B(n_1960),
.C(n_1956),
.Y(n_4203)
);

NAND2xp5_ASAP7_75t_L g4204 ( 
.A(n_4129),
.B(n_4135),
.Y(n_4204)
);

AOI22xp33_ASAP7_75t_L g4205 ( 
.A1(n_3975),
.A2(n_2787),
.B1(n_2650),
.B2(n_2654),
.Y(n_4205)
);

INVx1_ASAP7_75t_L g4206 ( 
.A(n_3854),
.Y(n_4206)
);

INVx5_ASAP7_75t_L g4207 ( 
.A(n_3970),
.Y(n_4207)
);

BUFx6f_ASAP7_75t_SL g4208 ( 
.A(n_3821),
.Y(n_4208)
);

CKINVDCx20_ASAP7_75t_R g4209 ( 
.A(n_3923),
.Y(n_4209)
);

NAND2xp5_ASAP7_75t_L g4210 ( 
.A(n_4142),
.B(n_2649),
.Y(n_4210)
);

AOI22xp33_ASAP7_75t_L g4211 ( 
.A1(n_3890),
.A2(n_2658),
.B1(n_2664),
.B2(n_2657),
.Y(n_4211)
);

INVx3_ASAP7_75t_L g4212 ( 
.A(n_4004),
.Y(n_4212)
);

NOR2xp33_ASAP7_75t_R g4213 ( 
.A(n_4146),
.B(n_2668),
.Y(n_4213)
);

INVx2_ASAP7_75t_SL g4214 ( 
.A(n_3831),
.Y(n_4214)
);

OR2x2_ASAP7_75t_L g4215 ( 
.A(n_3871),
.B(n_1962),
.Y(n_4215)
);

BUFx3_ASAP7_75t_L g4216 ( 
.A(n_4059),
.Y(n_4216)
);

NAND2xp5_ASAP7_75t_L g4217 ( 
.A(n_4148),
.B(n_2682),
.Y(n_4217)
);

CKINVDCx5p33_ASAP7_75t_R g4218 ( 
.A(n_3856),
.Y(n_4218)
);

INVx5_ASAP7_75t_L g4219 ( 
.A(n_3877),
.Y(n_4219)
);

BUFx3_ASAP7_75t_L g4220 ( 
.A(n_4104),
.Y(n_4220)
);

INVx1_ASAP7_75t_L g4221 ( 
.A(n_3865),
.Y(n_4221)
);

AOI22xp5_ASAP7_75t_L g4222 ( 
.A1(n_4153),
.A2(n_2697),
.B1(n_2698),
.B2(n_2691),
.Y(n_4222)
);

BUFx12f_ASAP7_75t_L g4223 ( 
.A(n_3965),
.Y(n_4223)
);

INVx1_ASAP7_75t_SL g4224 ( 
.A(n_3901),
.Y(n_4224)
);

BUFx4f_ASAP7_75t_L g4225 ( 
.A(n_4002),
.Y(n_4225)
);

INVx1_ASAP7_75t_L g4226 ( 
.A(n_3868),
.Y(n_4226)
);

CKINVDCx5p33_ASAP7_75t_R g4227 ( 
.A(n_3840),
.Y(n_4227)
);

NOR2xp33_ASAP7_75t_L g4228 ( 
.A(n_3917),
.B(n_1967),
.Y(n_4228)
);

INVx1_ASAP7_75t_L g4229 ( 
.A(n_3881),
.Y(n_4229)
);

BUFx6f_ASAP7_75t_L g4230 ( 
.A(n_4060),
.Y(n_4230)
);

NAND2xp5_ASAP7_75t_L g4231 ( 
.A(n_4155),
.B(n_2701),
.Y(n_4231)
);

BUFx4f_ASAP7_75t_L g4232 ( 
.A(n_3835),
.Y(n_4232)
);

INVx1_ASAP7_75t_L g4233 ( 
.A(n_3892),
.Y(n_4233)
);

NAND2xp5_ASAP7_75t_SL g4234 ( 
.A(n_3911),
.B(n_2704),
.Y(n_4234)
);

NAND2xp5_ASAP7_75t_L g4235 ( 
.A(n_4157),
.B(n_2707),
.Y(n_4235)
);

NAND2xp5_ASAP7_75t_L g4236 ( 
.A(n_4158),
.B(n_2714),
.Y(n_4236)
);

INVx5_ASAP7_75t_L g4237 ( 
.A(n_3951),
.Y(n_4237)
);

NAND2xp5_ASAP7_75t_L g4238 ( 
.A(n_4162),
.B(n_2716),
.Y(n_4238)
);

NOR2xp33_ASAP7_75t_L g4239 ( 
.A(n_3933),
.B(n_1972),
.Y(n_4239)
);

INVx1_ASAP7_75t_SL g4240 ( 
.A(n_3855),
.Y(n_4240)
);

INVx1_ASAP7_75t_L g4241 ( 
.A(n_3905),
.Y(n_4241)
);

NAND3xp33_ASAP7_75t_SL g4242 ( 
.A(n_4168),
.B(n_1982),
.C(n_1975),
.Y(n_4242)
);

INVx1_ASAP7_75t_L g4243 ( 
.A(n_3910),
.Y(n_4243)
);

INVx1_ASAP7_75t_L g4244 ( 
.A(n_3914),
.Y(n_4244)
);

INVx3_ASAP7_75t_L g4245 ( 
.A(n_4074),
.Y(n_4245)
);

NOR2xp33_ASAP7_75t_L g4246 ( 
.A(n_3929),
.B(n_1985),
.Y(n_4246)
);

NAND2xp5_ASAP7_75t_L g4247 ( 
.A(n_4174),
.B(n_2719),
.Y(n_4247)
);

NAND2xp5_ASAP7_75t_L g4248 ( 
.A(n_4176),
.B(n_2731),
.Y(n_4248)
);

BUFx2_ASAP7_75t_L g4249 ( 
.A(n_4037),
.Y(n_4249)
);

INVx4_ASAP7_75t_L g4250 ( 
.A(n_3836),
.Y(n_4250)
);

INVx2_ASAP7_75t_L g4251 ( 
.A(n_3922),
.Y(n_4251)
);

AND2x4_ASAP7_75t_SL g4252 ( 
.A(n_4116),
.B(n_4076),
.Y(n_4252)
);

INVxp67_ASAP7_75t_L g4253 ( 
.A(n_3861),
.Y(n_4253)
);

INVx2_ASAP7_75t_SL g4254 ( 
.A(n_4106),
.Y(n_4254)
);

NAND2xp5_ASAP7_75t_SL g4255 ( 
.A(n_3938),
.B(n_2744),
.Y(n_4255)
);

INVx3_ASAP7_75t_L g4256 ( 
.A(n_3988),
.Y(n_4256)
);

NAND2xp5_ASAP7_75t_L g4257 ( 
.A(n_3918),
.B(n_2749),
.Y(n_4257)
);

BUFx6f_ASAP7_75t_L g4258 ( 
.A(n_4014),
.Y(n_4258)
);

NOR2xp33_ASAP7_75t_L g4259 ( 
.A(n_3897),
.B(n_1988),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_3927),
.Y(n_4260)
);

INVx2_ASAP7_75t_SL g4261 ( 
.A(n_4003),
.Y(n_4261)
);

NAND2xp5_ASAP7_75t_L g4262 ( 
.A(n_3934),
.B(n_2751),
.Y(n_4262)
);

INVx2_ASAP7_75t_L g4263 ( 
.A(n_3925),
.Y(n_4263)
);

INVx1_ASAP7_75t_L g4264 ( 
.A(n_3935),
.Y(n_4264)
);

INVx5_ASAP7_75t_L g4265 ( 
.A(n_3951),
.Y(n_4265)
);

OR2x2_ASAP7_75t_L g4266 ( 
.A(n_4143),
.B(n_3972),
.Y(n_4266)
);

NOR2xp33_ASAP7_75t_SL g4267 ( 
.A(n_3880),
.B(n_2755),
.Y(n_4267)
);

INVx3_ASAP7_75t_SL g4268 ( 
.A(n_4119),
.Y(n_4268)
);

INVx4_ASAP7_75t_L g4269 ( 
.A(n_4095),
.Y(n_4269)
);

NAND2xp5_ASAP7_75t_L g4270 ( 
.A(n_3936),
.B(n_2767),
.Y(n_4270)
);

NAND2xp5_ASAP7_75t_L g4271 ( 
.A(n_4123),
.B(n_2772),
.Y(n_4271)
);

NAND2xp5_ASAP7_75t_SL g4272 ( 
.A(n_4055),
.B(n_2775),
.Y(n_4272)
);

NAND2xp5_ASAP7_75t_L g4273 ( 
.A(n_4125),
.B(n_2780),
.Y(n_4273)
);

INVxp67_ASAP7_75t_L g4274 ( 
.A(n_3991),
.Y(n_4274)
);

NAND2xp5_ASAP7_75t_L g4275 ( 
.A(n_4127),
.B(n_4128),
.Y(n_4275)
);

NAND2xp5_ASAP7_75t_L g4276 ( 
.A(n_4134),
.B(n_2783),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_4137),
.Y(n_4277)
);

INVx2_ASAP7_75t_L g4278 ( 
.A(n_3928),
.Y(n_4278)
);

OR2x2_ASAP7_75t_L g4279 ( 
.A(n_3886),
.B(n_1995),
.Y(n_4279)
);

NAND2xp5_ASAP7_75t_L g4280 ( 
.A(n_4145),
.B(n_2785),
.Y(n_4280)
);

NAND2xp5_ASAP7_75t_L g4281 ( 
.A(n_4152),
.B(n_2789),
.Y(n_4281)
);

OR2x2_ASAP7_75t_L g4282 ( 
.A(n_3899),
.B(n_1997),
.Y(n_4282)
);

INVxp67_ASAP7_75t_L g4283 ( 
.A(n_3999),
.Y(n_4283)
);

NAND2xp5_ASAP7_75t_L g4284 ( 
.A(n_4170),
.B(n_4171),
.Y(n_4284)
);

INVx1_ASAP7_75t_L g4285 ( 
.A(n_4175),
.Y(n_4285)
);

NAND2xp5_ASAP7_75t_L g4286 ( 
.A(n_4177),
.B(n_2798),
.Y(n_4286)
);

NAND3xp33_ASAP7_75t_SL g4287 ( 
.A(n_4013),
.B(n_2003),
.C(n_2001),
.Y(n_4287)
);

INVx2_ASAP7_75t_L g4288 ( 
.A(n_3937),
.Y(n_4288)
);

AOI21xp5_ASAP7_75t_L g4289 ( 
.A1(n_4011),
.A2(n_2811),
.B(n_2807),
.Y(n_4289)
);

NAND2xp5_ASAP7_75t_SL g4290 ( 
.A(n_4055),
.B(n_3943),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_3947),
.Y(n_4291)
);

INVx2_ASAP7_75t_SL g4292 ( 
.A(n_3959),
.Y(n_4292)
);

NAND2xp5_ASAP7_75t_SL g4293 ( 
.A(n_4055),
.B(n_2004),
.Y(n_4293)
);

INVx1_ASAP7_75t_L g4294 ( 
.A(n_3966),
.Y(n_4294)
);

NAND2xp5_ASAP7_75t_SL g4295 ( 
.A(n_4055),
.B(n_2005),
.Y(n_4295)
);

NAND2xp5_ASAP7_75t_L g4296 ( 
.A(n_3954),
.B(n_2013),
.Y(n_4296)
);

INVx2_ASAP7_75t_L g4297 ( 
.A(n_3823),
.Y(n_4297)
);

INVx1_ASAP7_75t_L g4298 ( 
.A(n_3978),
.Y(n_4298)
);

NAND2xp5_ASAP7_75t_L g4299 ( 
.A(n_4041),
.B(n_2018),
.Y(n_4299)
);

NOR2xp33_ASAP7_75t_L g4300 ( 
.A(n_3974),
.B(n_2019),
.Y(n_4300)
);

NAND2xp5_ASAP7_75t_L g4301 ( 
.A(n_3900),
.B(n_3902),
.Y(n_4301)
);

NAND2x1p5_ASAP7_75t_L g4302 ( 
.A(n_4095),
.B(n_2546),
.Y(n_4302)
);

CKINVDCx6p67_ASAP7_75t_R g4303 ( 
.A(n_4095),
.Y(n_4303)
);

AND2x4_ASAP7_75t_L g4304 ( 
.A(n_4047),
.B(n_2549),
.Y(n_4304)
);

INVx1_ASAP7_75t_L g4305 ( 
.A(n_3992),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_3998),
.Y(n_4306)
);

OAI21x1_ASAP7_75t_L g4307 ( 
.A1(n_3961),
.A2(n_2578),
.B(n_2575),
.Y(n_4307)
);

INVx3_ASAP7_75t_L g4308 ( 
.A(n_4080),
.Y(n_4308)
);

AOI22xp5_ASAP7_75t_L g4309 ( 
.A1(n_4020),
.A2(n_4124),
.B1(n_4131),
.B2(n_3822),
.Y(n_4309)
);

NAND2xp5_ASAP7_75t_SL g4310 ( 
.A(n_3909),
.B(n_2026),
.Y(n_4310)
);

NAND2xp5_ASAP7_75t_L g4311 ( 
.A(n_3912),
.B(n_2031),
.Y(n_4311)
);

NAND2xp5_ASAP7_75t_SL g4312 ( 
.A(n_3949),
.B(n_2033),
.Y(n_4312)
);

INVx1_ASAP7_75t_L g4313 ( 
.A(n_4039),
.Y(n_4313)
);

BUFx4f_ASAP7_75t_L g4314 ( 
.A(n_3835),
.Y(n_4314)
);

INVx1_ASAP7_75t_L g4315 ( 
.A(n_4000),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_4016),
.Y(n_4316)
);

INVx2_ASAP7_75t_L g4317 ( 
.A(n_3847),
.Y(n_4317)
);

NAND2xp5_ASAP7_75t_L g4318 ( 
.A(n_3875),
.B(n_2039),
.Y(n_4318)
);

NOR3xp33_ASAP7_75t_SL g4319 ( 
.A(n_3981),
.B(n_2048),
.C(n_2043),
.Y(n_4319)
);

INVx1_ASAP7_75t_L g4320 ( 
.A(n_4024),
.Y(n_4320)
);

NAND2xp5_ASAP7_75t_SL g4321 ( 
.A(n_3956),
.B(n_2052),
.Y(n_4321)
);

NAND2xp5_ASAP7_75t_L g4322 ( 
.A(n_3876),
.B(n_2057),
.Y(n_4322)
);

AND2x2_ASAP7_75t_L g4323 ( 
.A(n_3891),
.B(n_2059),
.Y(n_4323)
);

NOR2xp33_ASAP7_75t_L g4324 ( 
.A(n_3853),
.B(n_2066),
.Y(n_4324)
);

INVx2_ASAP7_75t_L g4325 ( 
.A(n_3848),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_4026),
.Y(n_4326)
);

AOI21xp5_ASAP7_75t_L g4327 ( 
.A1(n_4062),
.A2(n_2593),
.B(n_2581),
.Y(n_4327)
);

INVx1_ASAP7_75t_L g4328 ( 
.A(n_4027),
.Y(n_4328)
);

NAND2xp5_ASAP7_75t_SL g4329 ( 
.A(n_4083),
.B(n_2067),
.Y(n_4329)
);

BUFx6f_ASAP7_75t_L g4330 ( 
.A(n_3963),
.Y(n_4330)
);

CKINVDCx5p33_ASAP7_75t_R g4331 ( 
.A(n_3849),
.Y(n_4331)
);

INVxp33_ASAP7_75t_SL g4332 ( 
.A(n_4073),
.Y(n_4332)
);

INVx3_ASAP7_75t_L g4333 ( 
.A(n_4096),
.Y(n_4333)
);

INVx8_ASAP7_75t_L g4334 ( 
.A(n_3835),
.Y(n_4334)
);

NAND2xp5_ASAP7_75t_SL g4335 ( 
.A(n_4089),
.B(n_2070),
.Y(n_4335)
);

INVx1_ASAP7_75t_L g4336 ( 
.A(n_4018),
.Y(n_4336)
);

INVx4_ASAP7_75t_L g4337 ( 
.A(n_4139),
.Y(n_4337)
);

AND2x2_ASAP7_75t_L g4338 ( 
.A(n_3832),
.B(n_2073),
.Y(n_4338)
);

CKINVDCx16_ASAP7_75t_R g4339 ( 
.A(n_3843),
.Y(n_4339)
);

NOR2xp33_ASAP7_75t_L g4340 ( 
.A(n_3824),
.B(n_2078),
.Y(n_4340)
);

NAND2xp5_ASAP7_75t_SL g4341 ( 
.A(n_4072),
.B(n_2079),
.Y(n_4341)
);

BUFx6f_ASAP7_75t_L g4342 ( 
.A(n_4008),
.Y(n_4342)
);

INVx1_ASAP7_75t_L g4343 ( 
.A(n_4040),
.Y(n_4343)
);

INVx3_ASAP7_75t_L g4344 ( 
.A(n_4101),
.Y(n_4344)
);

NOR2x2_ASAP7_75t_L g4345 ( 
.A(n_4049),
.B(n_2222),
.Y(n_4345)
);

NAND2xp5_ASAP7_75t_SL g4346 ( 
.A(n_4068),
.B(n_2084),
.Y(n_4346)
);

BUFx8_ASAP7_75t_L g4347 ( 
.A(n_4115),
.Y(n_4347)
);

INVx2_ASAP7_75t_L g4348 ( 
.A(n_3859),
.Y(n_4348)
);

NAND2xp5_ASAP7_75t_L g4349 ( 
.A(n_3878),
.B(n_2086),
.Y(n_4349)
);

INVx1_ASAP7_75t_L g4350 ( 
.A(n_3885),
.Y(n_4350)
);

INVx3_ASAP7_75t_L g4351 ( 
.A(n_4070),
.Y(n_4351)
);

INVx2_ASAP7_75t_L g4352 ( 
.A(n_3895),
.Y(n_4352)
);

INVxp67_ASAP7_75t_SL g4353 ( 
.A(n_3842),
.Y(n_4353)
);

INVx2_ASAP7_75t_L g4354 ( 
.A(n_3904),
.Y(n_4354)
);

NAND2xp5_ASAP7_75t_SL g4355 ( 
.A(n_4165),
.B(n_2087),
.Y(n_4355)
);

AND2x4_ASAP7_75t_L g4356 ( 
.A(n_4064),
.B(n_2594),
.Y(n_4356)
);

INVx1_ASAP7_75t_L g4357 ( 
.A(n_3913),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_3960),
.Y(n_4358)
);

NAND2xp5_ASAP7_75t_L g4359 ( 
.A(n_3879),
.B(n_2088),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_3962),
.Y(n_4360)
);

INVx1_ASAP7_75t_L g4361 ( 
.A(n_3971),
.Y(n_4361)
);

INVx1_ASAP7_75t_L g4362 ( 
.A(n_3985),
.Y(n_4362)
);

NAND2xp5_ASAP7_75t_L g4363 ( 
.A(n_3884),
.B(n_2090),
.Y(n_4363)
);

INVxp67_ASAP7_75t_L g4364 ( 
.A(n_4007),
.Y(n_4364)
);

INVx1_ASAP7_75t_L g4365 ( 
.A(n_3987),
.Y(n_4365)
);

NAND2xp5_ASAP7_75t_SL g4366 ( 
.A(n_4006),
.B(n_2092),
.Y(n_4366)
);

INVx1_ASAP7_75t_L g4367 ( 
.A(n_4122),
.Y(n_4367)
);

INVx2_ASAP7_75t_L g4368 ( 
.A(n_4126),
.Y(n_4368)
);

BUFx3_ASAP7_75t_L g4369 ( 
.A(n_4082),
.Y(n_4369)
);

BUFx6f_ASAP7_75t_L g4370 ( 
.A(n_4029),
.Y(n_4370)
);

INVx1_ASAP7_75t_L g4371 ( 
.A(n_4144),
.Y(n_4371)
);

INVx3_ASAP7_75t_L g4372 ( 
.A(n_4088),
.Y(n_4372)
);

NAND2xp5_ASAP7_75t_L g4373 ( 
.A(n_3889),
.B(n_2093),
.Y(n_4373)
);

NAND2xp5_ASAP7_75t_SL g4374 ( 
.A(n_4010),
.B(n_2096),
.Y(n_4374)
);

BUFx3_ASAP7_75t_L g4375 ( 
.A(n_4090),
.Y(n_4375)
);

AOI21xp5_ASAP7_75t_L g4376 ( 
.A1(n_3845),
.A2(n_2598),
.B(n_2597),
.Y(n_4376)
);

INVx1_ASAP7_75t_L g4377 ( 
.A(n_4147),
.Y(n_4377)
);

INVx2_ASAP7_75t_L g4378 ( 
.A(n_4150),
.Y(n_4378)
);

NAND2xp5_ASAP7_75t_L g4379 ( 
.A(n_3939),
.B(n_2100),
.Y(n_4379)
);

CKINVDCx5p33_ASAP7_75t_R g4380 ( 
.A(n_3982),
.Y(n_4380)
);

NAND2xp5_ASAP7_75t_SL g4381 ( 
.A(n_4030),
.B(n_2112),
.Y(n_4381)
);

BUFx3_ASAP7_75t_L g4382 ( 
.A(n_4094),
.Y(n_4382)
);

INVx1_ASAP7_75t_L g4383 ( 
.A(n_4160),
.Y(n_4383)
);

AND2x4_ASAP7_75t_L g4384 ( 
.A(n_4057),
.B(n_2600),
.Y(n_4384)
);

INVx3_ASAP7_75t_L g4385 ( 
.A(n_4100),
.Y(n_4385)
);

NAND2xp5_ASAP7_75t_SL g4386 ( 
.A(n_4045),
.B(n_2113),
.Y(n_4386)
);

NAND2xp5_ASAP7_75t_L g4387 ( 
.A(n_3940),
.B(n_2114),
.Y(n_4387)
);

INVx2_ASAP7_75t_SL g4388 ( 
.A(n_4120),
.Y(n_4388)
);

INVx1_ASAP7_75t_L g4389 ( 
.A(n_4033),
.Y(n_4389)
);

AOI22xp5_ASAP7_75t_L g4390 ( 
.A1(n_4133),
.A2(n_2119),
.B1(n_2122),
.B2(n_2117),
.Y(n_4390)
);

NAND2xp5_ASAP7_75t_SL g4391 ( 
.A(n_3946),
.B(n_2125),
.Y(n_4391)
);

CKINVDCx5p33_ASAP7_75t_R g4392 ( 
.A(n_4091),
.Y(n_4392)
);

NAND2xp5_ASAP7_75t_L g4393 ( 
.A(n_3941),
.B(n_2126),
.Y(n_4393)
);

INVx3_ASAP7_75t_L g4394 ( 
.A(n_4069),
.Y(n_4394)
);

AND2x4_ASAP7_75t_L g4395 ( 
.A(n_3958),
.B(n_2633),
.Y(n_4395)
);

NAND2xp5_ASAP7_75t_L g4396 ( 
.A(n_4015),
.B(n_3898),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_3989),
.Y(n_4397)
);

BUFx5_ASAP7_75t_L g4398 ( 
.A(n_4042),
.Y(n_4398)
);

AOI21xp5_ASAP7_75t_L g4399 ( 
.A1(n_3846),
.A2(n_2638),
.B(n_2634),
.Y(n_4399)
);

INVx2_ASAP7_75t_L g4400 ( 
.A(n_4012),
.Y(n_4400)
);

AND2x2_ASAP7_75t_L g4401 ( 
.A(n_4043),
.B(n_2128),
.Y(n_4401)
);

NAND2xp5_ASAP7_75t_L g4402 ( 
.A(n_4136),
.B(n_2131),
.Y(n_4402)
);

INVx2_ASAP7_75t_L g4403 ( 
.A(n_4028),
.Y(n_4403)
);

INVx3_ASAP7_75t_L g4404 ( 
.A(n_3839),
.Y(n_4404)
);

CKINVDCx5p33_ASAP7_75t_R g4405 ( 
.A(n_4086),
.Y(n_4405)
);

INVx1_ASAP7_75t_L g4406 ( 
.A(n_4044),
.Y(n_4406)
);

AND2x2_ASAP7_75t_L g4407 ( 
.A(n_3857),
.B(n_2137),
.Y(n_4407)
);

NAND2xp5_ASAP7_75t_L g4408 ( 
.A(n_4138),
.B(n_2144),
.Y(n_4408)
);

INVx1_ASAP7_75t_L g4409 ( 
.A(n_4046),
.Y(n_4409)
);

HB1xp67_ASAP7_75t_L g4410 ( 
.A(n_4054),
.Y(n_4410)
);

BUFx6f_ASAP7_75t_L g4411 ( 
.A(n_3996),
.Y(n_4411)
);

AOI22xp5_ASAP7_75t_L g4412 ( 
.A1(n_4149),
.A2(n_4161),
.B1(n_4163),
.B2(n_4154),
.Y(n_4412)
);

OR2x2_ASAP7_75t_SL g4413 ( 
.A(n_4078),
.B(n_2644),
.Y(n_4413)
);

INVxp67_ASAP7_75t_L g4414 ( 
.A(n_4118),
.Y(n_4414)
);

NAND2xp5_ASAP7_75t_L g4415 ( 
.A(n_4167),
.B(n_2150),
.Y(n_4415)
);

NAND2xp5_ASAP7_75t_L g4416 ( 
.A(n_4169),
.B(n_2154),
.Y(n_4416)
);

INVx2_ASAP7_75t_SL g4417 ( 
.A(n_3995),
.Y(n_4417)
);

NOR2xp33_ASAP7_75t_L g4418 ( 
.A(n_4173),
.B(n_2156),
.Y(n_4418)
);

NAND2xp5_ASAP7_75t_L g4419 ( 
.A(n_3863),
.B(n_2159),
.Y(n_4419)
);

INVx1_ASAP7_75t_L g4420 ( 
.A(n_3858),
.Y(n_4420)
);

INVx1_ASAP7_75t_SL g4421 ( 
.A(n_3983),
.Y(n_4421)
);

CKINVDCx20_ASAP7_75t_R g4422 ( 
.A(n_3930),
.Y(n_4422)
);

INVx4_ASAP7_75t_L g4423 ( 
.A(n_3924),
.Y(n_4423)
);

NAND2xp5_ASAP7_75t_SL g4424 ( 
.A(n_4093),
.B(n_2171),
.Y(n_4424)
);

INVx1_ASAP7_75t_L g4425 ( 
.A(n_3860),
.Y(n_4425)
);

NAND2xp5_ASAP7_75t_SL g4426 ( 
.A(n_4071),
.B(n_2174),
.Y(n_4426)
);

BUFx3_ASAP7_75t_L g4427 ( 
.A(n_4113),
.Y(n_4427)
);

INVx1_ASAP7_75t_L g4428 ( 
.A(n_3931),
.Y(n_4428)
);

NAND2xp5_ASAP7_75t_SL g4429 ( 
.A(n_4038),
.B(n_2175),
.Y(n_4429)
);

NAND2xp5_ASAP7_75t_L g4430 ( 
.A(n_3829),
.B(n_2176),
.Y(n_4430)
);

INVx2_ASAP7_75t_SL g4431 ( 
.A(n_4048),
.Y(n_4431)
);

NAND2xp5_ASAP7_75t_SL g4432 ( 
.A(n_3907),
.B(n_2177),
.Y(n_4432)
);

INVx1_ASAP7_75t_L g4433 ( 
.A(n_3973),
.Y(n_4433)
);

INVx3_ASAP7_75t_L g4434 ( 
.A(n_4114),
.Y(n_4434)
);

INVx2_ASAP7_75t_SL g4435 ( 
.A(n_4098),
.Y(n_4435)
);

BUFx6f_ASAP7_75t_L g4436 ( 
.A(n_4025),
.Y(n_4436)
);

INVx2_ASAP7_75t_L g4437 ( 
.A(n_4051),
.Y(n_4437)
);

AND2x4_ASAP7_75t_L g4438 ( 
.A(n_4092),
.B(n_2648),
.Y(n_4438)
);

AOI22xp33_ASAP7_75t_L g4439 ( 
.A1(n_3833),
.A2(n_2250),
.B1(n_2256),
.B2(n_2248),
.Y(n_4439)
);

NAND3xp33_ASAP7_75t_L g4440 ( 
.A(n_4141),
.B(n_2186),
.C(n_2184),
.Y(n_4440)
);

INVx1_ASAP7_75t_L g4441 ( 
.A(n_3980),
.Y(n_4441)
);

NAND2xp5_ASAP7_75t_SL g4442 ( 
.A(n_4065),
.B(n_2187),
.Y(n_4442)
);

HB1xp67_ASAP7_75t_L g4443 ( 
.A(n_3869),
.Y(n_4443)
);

INVx2_ASAP7_75t_L g4444 ( 
.A(n_3950),
.Y(n_4444)
);

NAND2xp5_ASAP7_75t_L g4445 ( 
.A(n_3841),
.B(n_2188),
.Y(n_4445)
);

AOI22xp33_ASAP7_75t_L g4446 ( 
.A1(n_3873),
.A2(n_2329),
.B1(n_2351),
.B2(n_2294),
.Y(n_4446)
);

INVx1_ASAP7_75t_L g4447 ( 
.A(n_3984),
.Y(n_4447)
);

INVx1_ASAP7_75t_L g4448 ( 
.A(n_3993),
.Y(n_4448)
);

NAND2xp5_ASAP7_75t_L g4449 ( 
.A(n_3926),
.B(n_2192),
.Y(n_4449)
);

INVx4_ASAP7_75t_L g4450 ( 
.A(n_4172),
.Y(n_4450)
);

AND2x4_ASAP7_75t_L g4451 ( 
.A(n_4132),
.B(n_2655),
.Y(n_4451)
);

BUFx6f_ASAP7_75t_L g4452 ( 
.A(n_4099),
.Y(n_4452)
);

AOI22xp5_ASAP7_75t_L g4453 ( 
.A1(n_3920),
.A2(n_4156),
.B1(n_4130),
.B2(n_3883),
.Y(n_4453)
);

NAND2xp5_ASAP7_75t_L g4454 ( 
.A(n_4052),
.B(n_2198),
.Y(n_4454)
);

INVx2_ASAP7_75t_L g4455 ( 
.A(n_3994),
.Y(n_4455)
);

A2O1A1Ixp33_ASAP7_75t_L g4456 ( 
.A1(n_4056),
.A2(n_2667),
.B(n_2671),
.C(n_2663),
.Y(n_4456)
);

INVx1_ASAP7_75t_L g4457 ( 
.A(n_3997),
.Y(n_4457)
);

INVx4_ASAP7_75t_L g4458 ( 
.A(n_3893),
.Y(n_4458)
);

NAND3xp33_ASAP7_75t_SL g4459 ( 
.A(n_3851),
.B(n_2202),
.C(n_2200),
.Y(n_4459)
);

INVx3_ASAP7_75t_L g4460 ( 
.A(n_4107),
.Y(n_4460)
);

NOR2xp33_ASAP7_75t_L g4461 ( 
.A(n_4105),
.B(n_2204),
.Y(n_4461)
);

AOI22xp5_ASAP7_75t_L g4462 ( 
.A1(n_3874),
.A2(n_2217),
.B1(n_2219),
.B2(n_2212),
.Y(n_4462)
);

NAND2xp5_ASAP7_75t_L g4463 ( 
.A(n_4053),
.B(n_2229),
.Y(n_4463)
);

AOI22xp33_ASAP7_75t_L g4464 ( 
.A1(n_3948),
.A2(n_2399),
.B1(n_2426),
.B2(n_2368),
.Y(n_4464)
);

NOR2xp33_ASAP7_75t_L g4465 ( 
.A(n_4087),
.B(n_2235),
.Y(n_4465)
);

AOI22xp5_ASAP7_75t_L g4466 ( 
.A1(n_3887),
.A2(n_3944),
.B1(n_3908),
.B2(n_4023),
.Y(n_4466)
);

OR2x6_ASAP7_75t_L g4467 ( 
.A(n_3968),
.B(n_2676),
.Y(n_4467)
);

INVx1_ASAP7_75t_L g4468 ( 
.A(n_4001),
.Y(n_4468)
);

BUFx3_ASAP7_75t_L g4469 ( 
.A(n_4102),
.Y(n_4469)
);

CKINVDCx5p33_ASAP7_75t_R g4470 ( 
.A(n_4108),
.Y(n_4470)
);

INVx4_ASAP7_75t_L g4471 ( 
.A(n_4035),
.Y(n_4471)
);

INVx1_ASAP7_75t_L g4472 ( 
.A(n_4179),
.Y(n_4472)
);

INVx2_ASAP7_75t_L g4473 ( 
.A(n_4185),
.Y(n_4473)
);

CKINVDCx14_ASAP7_75t_R g4474 ( 
.A(n_4209),
.Y(n_4474)
);

BUFx2_ASAP7_75t_L g4475 ( 
.A(n_4183),
.Y(n_4475)
);

NOR2xp33_ASAP7_75t_L g4476 ( 
.A(n_4332),
.B(n_4097),
.Y(n_4476)
);

HB1xp67_ASAP7_75t_L g4477 ( 
.A(n_4224),
.Y(n_4477)
);

NAND2xp5_ASAP7_75t_L g4478 ( 
.A(n_4180),
.B(n_3882),
.Y(n_4478)
);

INVx2_ASAP7_75t_SL g4479 ( 
.A(n_4216),
.Y(n_4479)
);

BUFx3_ASAP7_75t_L g4480 ( 
.A(n_4220),
.Y(n_4480)
);

NOR2xp33_ASAP7_75t_L g4481 ( 
.A(n_4253),
.B(n_4079),
.Y(n_4481)
);

BUFx4f_ASAP7_75t_L g4482 ( 
.A(n_4188),
.Y(n_4482)
);

OR2x6_ASAP7_75t_L g4483 ( 
.A(n_4334),
.B(n_4109),
.Y(n_4483)
);

INVx3_ASAP7_75t_L g4484 ( 
.A(n_4193),
.Y(n_4484)
);

INVx2_ASAP7_75t_L g4485 ( 
.A(n_4189),
.Y(n_4485)
);

INVx4_ASAP7_75t_L g4486 ( 
.A(n_4188),
.Y(n_4486)
);

NAND2xp5_ASAP7_75t_L g4487 ( 
.A(n_4196),
.B(n_3969),
.Y(n_4487)
);

NOR2xp33_ASAP7_75t_L g4488 ( 
.A(n_4182),
.B(n_4117),
.Y(n_4488)
);

CKINVDCx20_ASAP7_75t_R g4489 ( 
.A(n_4218),
.Y(n_4489)
);

AND2x2_ASAP7_75t_L g4490 ( 
.A(n_4323),
.B(n_4338),
.Y(n_4490)
);

NAND2xp5_ASAP7_75t_SL g4491 ( 
.A(n_4339),
.B(n_4017),
.Y(n_4491)
);

OR2x6_ASAP7_75t_L g4492 ( 
.A(n_4334),
.B(n_3942),
.Y(n_4492)
);

NAND2xp5_ASAP7_75t_L g4493 ( 
.A(n_4301),
.B(n_4081),
.Y(n_4493)
);

BUFx6f_ASAP7_75t_L g4494 ( 
.A(n_4190),
.Y(n_4494)
);

OAI21xp5_ASAP7_75t_L g4495 ( 
.A1(n_4204),
.A2(n_3819),
.B(n_4084),
.Y(n_4495)
);

INVx2_ASAP7_75t_L g4496 ( 
.A(n_4206),
.Y(n_4496)
);

INVx2_ASAP7_75t_L g4497 ( 
.A(n_4221),
.Y(n_4497)
);

BUFx6f_ASAP7_75t_L g4498 ( 
.A(n_4190),
.Y(n_4498)
);

BUFx2_ASAP7_75t_L g4499 ( 
.A(n_4380),
.Y(n_4499)
);

INVxp67_ASAP7_75t_SL g4500 ( 
.A(n_4214),
.Y(n_4500)
);

NAND2xp5_ASAP7_75t_L g4501 ( 
.A(n_4420),
.B(n_4009),
.Y(n_4501)
);

INVx1_ASAP7_75t_L g4502 ( 
.A(n_4226),
.Y(n_4502)
);

INVx1_ASAP7_75t_L g4503 ( 
.A(n_4229),
.Y(n_4503)
);

BUFx6f_ASAP7_75t_L g4504 ( 
.A(n_4230),
.Y(n_4504)
);

NOR2xp33_ASAP7_75t_L g4505 ( 
.A(n_4199),
.B(n_3945),
.Y(n_4505)
);

HB1xp67_ASAP7_75t_L g4506 ( 
.A(n_4240),
.Y(n_4506)
);

AND2x4_ASAP7_75t_L g4507 ( 
.A(n_4337),
.B(n_4110),
.Y(n_4507)
);

AND2x2_ASAP7_75t_L g4508 ( 
.A(n_4401),
.B(n_3952),
.Y(n_4508)
);

NAND2xp5_ASAP7_75t_L g4509 ( 
.A(n_4425),
.B(n_4336),
.Y(n_4509)
);

BUFx2_ASAP7_75t_L g4510 ( 
.A(n_4392),
.Y(n_4510)
);

BUFx2_ASAP7_75t_L g4511 ( 
.A(n_4249),
.Y(n_4511)
);

OAI22xp5_ASAP7_75t_L g4512 ( 
.A1(n_4396),
.A2(n_4140),
.B1(n_4019),
.B2(n_4034),
.Y(n_4512)
);

NOR2xp33_ASAP7_75t_L g4513 ( 
.A(n_4202),
.B(n_3953),
.Y(n_4513)
);

INVx2_ASAP7_75t_L g4514 ( 
.A(n_4233),
.Y(n_4514)
);

NAND2xp5_ASAP7_75t_L g4515 ( 
.A(n_4461),
.B(n_4032),
.Y(n_4515)
);

INVxp67_ASAP7_75t_SL g4516 ( 
.A(n_4410),
.Y(n_4516)
);

CKINVDCx5p33_ASAP7_75t_R g4517 ( 
.A(n_4227),
.Y(n_4517)
);

AOI22xp5_ASAP7_75t_L g4518 ( 
.A1(n_4228),
.A2(n_4005),
.B1(n_4063),
.B2(n_4077),
.Y(n_4518)
);

NAND2xp5_ASAP7_75t_L g4519 ( 
.A(n_4433),
.B(n_4021),
.Y(n_4519)
);

BUFx4f_ASAP7_75t_L g4520 ( 
.A(n_4223),
.Y(n_4520)
);

NAND2xp5_ASAP7_75t_L g4521 ( 
.A(n_4441),
.B(n_4031),
.Y(n_4521)
);

BUFx2_ASAP7_75t_L g4522 ( 
.A(n_4421),
.Y(n_4522)
);

NAND2xp5_ASAP7_75t_SL g4523 ( 
.A(n_4267),
.B(n_4103),
.Y(n_4523)
);

HB1xp67_ASAP7_75t_L g4524 ( 
.A(n_4208),
.Y(n_4524)
);

BUFx2_ASAP7_75t_L g4525 ( 
.A(n_4427),
.Y(n_4525)
);

AND2x4_ASAP7_75t_L g4526 ( 
.A(n_4254),
.B(n_4111),
.Y(n_4526)
);

INVx2_ASAP7_75t_L g4527 ( 
.A(n_4241),
.Y(n_4527)
);

NAND2xp5_ASAP7_75t_L g4528 ( 
.A(n_4447),
.B(n_4066),
.Y(n_4528)
);

INVx1_ASAP7_75t_L g4529 ( 
.A(n_4243),
.Y(n_4529)
);

INVx1_ASAP7_75t_L g4530 ( 
.A(n_4244),
.Y(n_4530)
);

AND2x2_ASAP7_75t_L g4531 ( 
.A(n_4246),
.B(n_3955),
.Y(n_4531)
);

HB1xp67_ASAP7_75t_L g4532 ( 
.A(n_4230),
.Y(n_4532)
);

BUFx6f_ASAP7_75t_L g4533 ( 
.A(n_4258),
.Y(n_4533)
);

NAND2xp5_ASAP7_75t_L g4534 ( 
.A(n_4448),
.B(n_4112),
.Y(n_4534)
);

BUFx3_ASAP7_75t_L g4535 ( 
.A(n_4347),
.Y(n_4535)
);

AOI21xp33_ASAP7_75t_L g4536 ( 
.A1(n_4239),
.A2(n_4022),
.B(n_3894),
.Y(n_4536)
);

INVx1_ASAP7_75t_L g4537 ( 
.A(n_4260),
.Y(n_4537)
);

AOI21xp5_ASAP7_75t_L g4538 ( 
.A1(n_4272),
.A2(n_4036),
.B(n_3977),
.Y(n_4538)
);

NAND2xp5_ASAP7_75t_SL g4539 ( 
.A(n_4470),
.B(n_4085),
.Y(n_4539)
);

NAND2xp5_ASAP7_75t_L g4540 ( 
.A(n_4457),
.B(n_3957),
.Y(n_4540)
);

INVx1_ASAP7_75t_L g4541 ( 
.A(n_4264),
.Y(n_4541)
);

NAND2xp5_ASAP7_75t_SL g4542 ( 
.A(n_4266),
.B(n_4452),
.Y(n_4542)
);

AND2x4_ASAP7_75t_L g4543 ( 
.A(n_4292),
.B(n_3964),
.Y(n_4543)
);

INVx1_ASAP7_75t_L g4544 ( 
.A(n_4277),
.Y(n_4544)
);

INVx2_ASAP7_75t_SL g4545 ( 
.A(n_4258),
.Y(n_4545)
);

INVx2_ASAP7_75t_L g4546 ( 
.A(n_4285),
.Y(n_4546)
);

CKINVDCx5p33_ASAP7_75t_R g4547 ( 
.A(n_4405),
.Y(n_4547)
);

INVx4_ASAP7_75t_L g4548 ( 
.A(n_4225),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_4291),
.Y(n_4549)
);

INVx1_ASAP7_75t_L g4550 ( 
.A(n_4294),
.Y(n_4550)
);

INVx1_ASAP7_75t_SL g4551 ( 
.A(n_4345),
.Y(n_4551)
);

BUFx3_ASAP7_75t_L g4552 ( 
.A(n_4252),
.Y(n_4552)
);

INVx2_ASAP7_75t_L g4553 ( 
.A(n_4298),
.Y(n_4553)
);

NAND2xp5_ASAP7_75t_L g4554 ( 
.A(n_4468),
.B(n_3976),
.Y(n_4554)
);

NAND2xp5_ASAP7_75t_L g4555 ( 
.A(n_4455),
.B(n_3990),
.Y(n_4555)
);

INVx2_ASAP7_75t_L g4556 ( 
.A(n_4305),
.Y(n_4556)
);

INVx3_ASAP7_75t_L g4557 ( 
.A(n_4245),
.Y(n_4557)
);

INVx2_ASAP7_75t_SL g4558 ( 
.A(n_4342),
.Y(n_4558)
);

NAND2xp5_ASAP7_75t_L g4559 ( 
.A(n_4299),
.B(n_4067),
.Y(n_4559)
);

AOI22xp33_ASAP7_75t_L g4560 ( 
.A1(n_4259),
.A2(n_3967),
.B1(n_4050),
.B2(n_3866),
.Y(n_4560)
);

INVx3_ASAP7_75t_L g4561 ( 
.A(n_4250),
.Y(n_4561)
);

INVx1_ASAP7_75t_L g4562 ( 
.A(n_4306),
.Y(n_4562)
);

NAND2xp5_ASAP7_75t_SL g4563 ( 
.A(n_4452),
.B(n_3979),
.Y(n_4563)
);

AND2x2_ASAP7_75t_L g4564 ( 
.A(n_4407),
.B(n_3827),
.Y(n_4564)
);

NOR2x1p5_ASAP7_75t_L g4565 ( 
.A(n_4203),
.B(n_2236),
.Y(n_4565)
);

NAND2xp5_ASAP7_75t_L g4566 ( 
.A(n_4324),
.B(n_3867),
.Y(n_4566)
);

INVx2_ASAP7_75t_L g4567 ( 
.A(n_4313),
.Y(n_4567)
);

NOR2xp67_ASAP7_75t_L g4568 ( 
.A(n_4471),
.B(n_4364),
.Y(n_4568)
);

BUFx3_ASAP7_75t_L g4569 ( 
.A(n_4342),
.Y(n_4569)
);

NAND2xp5_ASAP7_75t_SL g4570 ( 
.A(n_4309),
.B(n_3903),
.Y(n_4570)
);

NAND2xp5_ASAP7_75t_L g4571 ( 
.A(n_4296),
.B(n_4075),
.Y(n_4571)
);

INVx2_ASAP7_75t_L g4572 ( 
.A(n_4315),
.Y(n_4572)
);

CKINVDCx5p33_ASAP7_75t_R g4573 ( 
.A(n_4213),
.Y(n_4573)
);

NAND2xp5_ASAP7_75t_L g4574 ( 
.A(n_4186),
.B(n_4437),
.Y(n_4574)
);

CKINVDCx5p33_ASAP7_75t_R g4575 ( 
.A(n_4331),
.Y(n_4575)
);

AOI22xp5_ASAP7_75t_L g4576 ( 
.A1(n_4422),
.A2(n_3916),
.B1(n_2249),
.B2(n_2253),
.Y(n_4576)
);

NAND2xp5_ASAP7_75t_L g4577 ( 
.A(n_4187),
.B(n_4435),
.Y(n_4577)
);

NAND2xp5_ASAP7_75t_L g4578 ( 
.A(n_4194),
.B(n_4151),
.Y(n_4578)
);

NAND2xp5_ASAP7_75t_L g4579 ( 
.A(n_4198),
.B(n_2688),
.Y(n_4579)
);

AOI22xp5_ASAP7_75t_L g4580 ( 
.A1(n_4340),
.A2(n_2255),
.B1(n_2265),
.B2(n_2241),
.Y(n_4580)
);

HB1xp67_ASAP7_75t_L g4581 ( 
.A(n_4369),
.Y(n_4581)
);

INVx4_ASAP7_75t_L g4582 ( 
.A(n_4370),
.Y(n_4582)
);

OR2x2_ASAP7_75t_SL g4583 ( 
.A(n_4287),
.B(n_2431),
.Y(n_4583)
);

AOI22xp33_ASAP7_75t_L g4584 ( 
.A1(n_4459),
.A2(n_2711),
.B1(n_2718),
.B2(n_2710),
.Y(n_4584)
);

NOR2xp33_ASAP7_75t_L g4585 ( 
.A(n_4282),
.B(n_2270),
.Y(n_4585)
);

INVx3_ASAP7_75t_L g4586 ( 
.A(n_4436),
.Y(n_4586)
);

INVx1_ASAP7_75t_L g4587 ( 
.A(n_4275),
.Y(n_4587)
);

OR2x6_ASAP7_75t_L g4588 ( 
.A(n_4370),
.B(n_2729),
.Y(n_4588)
);

INVx2_ASAP7_75t_L g4589 ( 
.A(n_4316),
.Y(n_4589)
);

INVx4_ASAP7_75t_L g4590 ( 
.A(n_4303),
.Y(n_4590)
);

AND2x2_ASAP7_75t_L g4591 ( 
.A(n_4215),
.B(n_2274),
.Y(n_4591)
);

AND2x2_ASAP7_75t_L g4592 ( 
.A(n_4395),
.B(n_2278),
.Y(n_4592)
);

NAND2xp5_ASAP7_75t_L g4593 ( 
.A(n_4311),
.B(n_2733),
.Y(n_4593)
);

INVx2_ASAP7_75t_L g4594 ( 
.A(n_4320),
.Y(n_4594)
);

BUFx4f_ASAP7_75t_L g4595 ( 
.A(n_4268),
.Y(n_4595)
);

NAND2xp5_ASAP7_75t_L g4596 ( 
.A(n_4284),
.B(n_2753),
.Y(n_4596)
);

AND2x4_ASAP7_75t_L g4597 ( 
.A(n_4375),
.B(n_2762),
.Y(n_4597)
);

OAI22xp5_ASAP7_75t_L g4598 ( 
.A1(n_4412),
.A2(n_2282),
.B1(n_2285),
.B2(n_2279),
.Y(n_4598)
);

INVx1_ASAP7_75t_L g4599 ( 
.A(n_4326),
.Y(n_4599)
);

AND2x2_ASAP7_75t_L g4600 ( 
.A(n_4353),
.B(n_2287),
.Y(n_4600)
);

INVx1_ASAP7_75t_L g4601 ( 
.A(n_4328),
.Y(n_4601)
);

INVx2_ASAP7_75t_L g4602 ( 
.A(n_4184),
.Y(n_4602)
);

NAND2xp5_ASAP7_75t_L g4603 ( 
.A(n_4318),
.B(n_2764),
.Y(n_4603)
);

NAND2xp5_ASAP7_75t_L g4604 ( 
.A(n_4322),
.B(n_4349),
.Y(n_4604)
);

NAND2xp5_ASAP7_75t_L g4605 ( 
.A(n_4359),
.B(n_4363),
.Y(n_4605)
);

NOR2xp33_ASAP7_75t_L g4606 ( 
.A(n_4373),
.B(n_4379),
.Y(n_4606)
);

O2A1O1Ixp33_ASAP7_75t_L g4607 ( 
.A1(n_4386),
.A2(n_2793),
.B(n_2796),
.C(n_2786),
.Y(n_4607)
);

CKINVDCx16_ASAP7_75t_R g4608 ( 
.A(n_4330),
.Y(n_4608)
);

INVx1_ASAP7_75t_L g4609 ( 
.A(n_4191),
.Y(n_4609)
);

BUFx6f_ASAP7_75t_L g4610 ( 
.A(n_4330),
.Y(n_4610)
);

INVx2_ASAP7_75t_L g4611 ( 
.A(n_4192),
.Y(n_4611)
);

INVx1_ASAP7_75t_L g4612 ( 
.A(n_4195),
.Y(n_4612)
);

INVx3_ASAP7_75t_L g4613 ( 
.A(n_4436),
.Y(n_4613)
);

INVx2_ASAP7_75t_L g4614 ( 
.A(n_4251),
.Y(n_4614)
);

HB1xp67_ASAP7_75t_L g4615 ( 
.A(n_4382),
.Y(n_4615)
);

NAND2xp5_ASAP7_75t_L g4616 ( 
.A(n_4387),
.B(n_2290),
.Y(n_4616)
);

NAND2xp5_ASAP7_75t_L g4617 ( 
.A(n_4393),
.B(n_4460),
.Y(n_4617)
);

INVx3_ASAP7_75t_L g4618 ( 
.A(n_4269),
.Y(n_4618)
);

INVx4_ASAP7_75t_SL g4619 ( 
.A(n_4411),
.Y(n_4619)
);

INVx1_ASAP7_75t_L g4620 ( 
.A(n_4263),
.Y(n_4620)
);

BUFx6f_ASAP7_75t_L g4621 ( 
.A(n_4411),
.Y(n_4621)
);

INVx2_ASAP7_75t_SL g4622 ( 
.A(n_4237),
.Y(n_4622)
);

HB1xp67_ASAP7_75t_L g4623 ( 
.A(n_4261),
.Y(n_4623)
);

BUFx3_ASAP7_75t_L g4624 ( 
.A(n_4219),
.Y(n_4624)
);

AND2x4_ASAP7_75t_L g4625 ( 
.A(n_4256),
.B(n_4417),
.Y(n_4625)
);

INVx5_ASAP7_75t_L g4626 ( 
.A(n_4207),
.Y(n_4626)
);

BUFx6f_ASAP7_75t_L g4627 ( 
.A(n_4219),
.Y(n_4627)
);

INVx1_ASAP7_75t_L g4628 ( 
.A(n_4278),
.Y(n_4628)
);

INVx4_ASAP7_75t_L g4629 ( 
.A(n_4237),
.Y(n_4629)
);

NAND2xp5_ASAP7_75t_L g4630 ( 
.A(n_4419),
.B(n_2292),
.Y(n_4630)
);

AO22x1_ASAP7_75t_L g4631 ( 
.A1(n_4265),
.A2(n_4465),
.B1(n_4418),
.B2(n_4404),
.Y(n_4631)
);

AND2x2_ASAP7_75t_L g4632 ( 
.A(n_4274),
.B(n_2297),
.Y(n_4632)
);

CKINVDCx5p33_ASAP7_75t_R g4633 ( 
.A(n_4207),
.Y(n_4633)
);

NAND2xp5_ASAP7_75t_SL g4634 ( 
.A(n_4283),
.B(n_2300),
.Y(n_4634)
);

NAND2xp5_ASAP7_75t_L g4635 ( 
.A(n_4454),
.B(n_2302),
.Y(n_4635)
);

BUFx6f_ASAP7_75t_L g4636 ( 
.A(n_4265),
.Y(n_4636)
);

NOR2xp33_ASAP7_75t_L g4637 ( 
.A(n_4463),
.B(n_2305),
.Y(n_4637)
);

CKINVDCx5p33_ASAP7_75t_R g4638 ( 
.A(n_4431),
.Y(n_4638)
);

OR2x2_ASAP7_75t_L g4639 ( 
.A(n_4279),
.B(n_2307),
.Y(n_4639)
);

AND2x6_ASAP7_75t_L g4640 ( 
.A(n_4453),
.B(n_2482),
.Y(n_4640)
);

NAND2xp5_ASAP7_75t_L g4641 ( 
.A(n_4449),
.B(n_2309),
.Y(n_4641)
);

NAND2xp5_ASAP7_75t_SL g4642 ( 
.A(n_4232),
.B(n_2311),
.Y(n_4642)
);

INVxp67_ASAP7_75t_SL g4643 ( 
.A(n_4372),
.Y(n_4643)
);

BUFx6f_ASAP7_75t_L g4644 ( 
.A(n_4212),
.Y(n_4644)
);

AOI22xp33_ASAP7_75t_L g4645 ( 
.A1(n_4366),
.A2(n_2520),
.B1(n_2559),
.B2(n_2490),
.Y(n_4645)
);

NAND2xp5_ASAP7_75t_L g4646 ( 
.A(n_4200),
.B(n_2314),
.Y(n_4646)
);

BUFx6f_ASAP7_75t_L g4647 ( 
.A(n_4384),
.Y(n_4647)
);

NAND2xp5_ASAP7_75t_L g4648 ( 
.A(n_4288),
.B(n_2317),
.Y(n_4648)
);

CKINVDCx5p33_ASAP7_75t_R g4649 ( 
.A(n_4469),
.Y(n_4649)
);

NAND2xp5_ASAP7_75t_SL g4650 ( 
.A(n_4314),
.B(n_2320),
.Y(n_4650)
);

INVx2_ASAP7_75t_L g4651 ( 
.A(n_4400),
.Y(n_4651)
);

BUFx6f_ASAP7_75t_L g4652 ( 
.A(n_4356),
.Y(n_4652)
);

INVx2_ASAP7_75t_SL g4653 ( 
.A(n_4394),
.Y(n_4653)
);

INVx3_ASAP7_75t_L g4654 ( 
.A(n_4385),
.Y(n_4654)
);

BUFx3_ASAP7_75t_L g4655 ( 
.A(n_4304),
.Y(n_4655)
);

INVx1_ASAP7_75t_L g4656 ( 
.A(n_4343),
.Y(n_4656)
);

NAND2xp5_ASAP7_75t_L g4657 ( 
.A(n_4210),
.B(n_4217),
.Y(n_4657)
);

INVx3_ASAP7_75t_L g4658 ( 
.A(n_4308),
.Y(n_4658)
);

NAND2xp5_ASAP7_75t_L g4659 ( 
.A(n_4231),
.B(n_4235),
.Y(n_4659)
);

HB1xp67_ASAP7_75t_L g4660 ( 
.A(n_4414),
.Y(n_4660)
);

INVx2_ASAP7_75t_L g4661 ( 
.A(n_4403),
.Y(n_4661)
);

OR2x2_ASAP7_75t_L g4662 ( 
.A(n_4178),
.B(n_2332),
.Y(n_4662)
);

BUFx3_ASAP7_75t_L g4663 ( 
.A(n_4388),
.Y(n_4663)
);

BUFx6f_ASAP7_75t_L g4664 ( 
.A(n_4438),
.Y(n_4664)
);

NAND2xp5_ASAP7_75t_L g4665 ( 
.A(n_4236),
.B(n_2335),
.Y(n_4665)
);

NAND2x1p5_ASAP7_75t_L g4666 ( 
.A(n_4333),
.B(n_2628),
.Y(n_4666)
);

AOI22xp5_ASAP7_75t_L g4667 ( 
.A1(n_4300),
.A2(n_2336),
.B1(n_2342),
.B2(n_2341),
.Y(n_4667)
);

INVx6_ASAP7_75t_L g4668 ( 
.A(n_4423),
.Y(n_4668)
);

INVx2_ASAP7_75t_L g4669 ( 
.A(n_4297),
.Y(n_4669)
);

INVx1_ASAP7_75t_L g4670 ( 
.A(n_4397),
.Y(n_4670)
);

NAND2xp5_ASAP7_75t_L g4671 ( 
.A(n_4238),
.B(n_2345),
.Y(n_4671)
);

BUFx2_ASAP7_75t_L g4672 ( 
.A(n_4344),
.Y(n_4672)
);

INVx1_ASAP7_75t_L g4673 ( 
.A(n_4350),
.Y(n_4673)
);

NAND2xp5_ASAP7_75t_L g4674 ( 
.A(n_4247),
.B(n_2358),
.Y(n_4674)
);

AND2x2_ASAP7_75t_L g4675 ( 
.A(n_4467),
.B(n_2359),
.Y(n_4675)
);

INVx1_ASAP7_75t_L g4676 ( 
.A(n_4357),
.Y(n_4676)
);

A2O1A1Ixp33_ASAP7_75t_L g4677 ( 
.A1(n_4466),
.A2(n_2681),
.B(n_2684),
.C(n_2662),
.Y(n_4677)
);

INVx2_ASAP7_75t_L g4678 ( 
.A(n_4317),
.Y(n_4678)
);

NAND2xp5_ASAP7_75t_L g4679 ( 
.A(n_4248),
.B(n_2362),
.Y(n_4679)
);

AOI22xp33_ASAP7_75t_L g4680 ( 
.A1(n_4374),
.A2(n_2771),
.B1(n_2800),
.B2(n_2690),
.Y(n_4680)
);

AOI21xp5_ASAP7_75t_L g4681 ( 
.A1(n_4293),
.A2(n_1061),
.B(n_1060),
.Y(n_4681)
);

NAND2xp5_ASAP7_75t_L g4682 ( 
.A(n_4329),
.B(n_2365),
.Y(n_4682)
);

AND2x2_ASAP7_75t_L g4683 ( 
.A(n_4467),
.B(n_2366),
.Y(n_4683)
);

INVx1_ASAP7_75t_L g4684 ( 
.A(n_4358),
.Y(n_4684)
);

INVx1_ASAP7_75t_L g4685 ( 
.A(n_4360),
.Y(n_4685)
);

INVx1_ASAP7_75t_L g4686 ( 
.A(n_4361),
.Y(n_4686)
);

A2O1A1Ixp33_ASAP7_75t_L g4687 ( 
.A1(n_4381),
.A2(n_4440),
.B(n_4242),
.C(n_4335),
.Y(n_4687)
);

INVx8_ASAP7_75t_L g4688 ( 
.A(n_4451),
.Y(n_4688)
);

NAND2x1_ASAP7_75t_L g4689 ( 
.A(n_4362),
.B(n_2299),
.Y(n_4689)
);

OR2x6_ASAP7_75t_L g4690 ( 
.A(n_4302),
.B(n_1062),
.Y(n_4690)
);

INVxp67_ASAP7_75t_L g4691 ( 
.A(n_4406),
.Y(n_4691)
);

AND2x4_ASAP7_75t_L g4692 ( 
.A(n_4409),
.B(n_1063),
.Y(n_4692)
);

INVx2_ASAP7_75t_L g4693 ( 
.A(n_4325),
.Y(n_4693)
);

INVx3_ASAP7_75t_L g4694 ( 
.A(n_4351),
.Y(n_4694)
);

BUFx2_ASAP7_75t_L g4695 ( 
.A(n_4413),
.Y(n_4695)
);

OR2x2_ASAP7_75t_L g4696 ( 
.A(n_4257),
.B(n_2369),
.Y(n_4696)
);

AND2x4_ASAP7_75t_L g4697 ( 
.A(n_4443),
.B(n_1064),
.Y(n_4697)
);

BUFx6f_ASAP7_75t_L g4698 ( 
.A(n_4348),
.Y(n_4698)
);

AND2x2_ASAP7_75t_L g4699 ( 
.A(n_4352),
.B(n_4354),
.Y(n_4699)
);

AND2x2_ASAP7_75t_SL g4700 ( 
.A(n_4205),
.B(n_1),
.Y(n_4700)
);

INVx1_ASAP7_75t_L g4701 ( 
.A(n_4365),
.Y(n_4701)
);

BUFx6f_ASAP7_75t_L g4702 ( 
.A(n_4368),
.Y(n_4702)
);

CKINVDCx5p33_ASAP7_75t_R g4703 ( 
.A(n_4319),
.Y(n_4703)
);

AND2x2_ASAP7_75t_L g4704 ( 
.A(n_4378),
.B(n_2370),
.Y(n_4704)
);

HB1xp67_ASAP7_75t_L g4705 ( 
.A(n_4367),
.Y(n_4705)
);

AND2x2_ASAP7_75t_L g4706 ( 
.A(n_4371),
.B(n_2375),
.Y(n_4706)
);

NAND2xp5_ASAP7_75t_SL g4707 ( 
.A(n_4430),
.B(n_4445),
.Y(n_4707)
);

AND2x4_ASAP7_75t_L g4708 ( 
.A(n_4377),
.B(n_1066),
.Y(n_4708)
);

AND2x2_ASAP7_75t_L g4709 ( 
.A(n_4383),
.B(n_2379),
.Y(n_4709)
);

AOI22xp5_ASAP7_75t_L g4710 ( 
.A1(n_4234),
.A2(n_2396),
.B1(n_2400),
.B2(n_2388),
.Y(n_4710)
);

INVx2_ASAP7_75t_L g4711 ( 
.A(n_4389),
.Y(n_4711)
);

NAND2xp5_ASAP7_75t_L g4712 ( 
.A(n_4327),
.B(n_4262),
.Y(n_4712)
);

AND2x2_ASAP7_75t_L g4713 ( 
.A(n_4390),
.B(n_2402),
.Y(n_4713)
);

NOR2xp33_ASAP7_75t_L g4714 ( 
.A(n_4310),
.B(n_2403),
.Y(n_4714)
);

NAND2xp5_ASAP7_75t_L g4715 ( 
.A(n_4270),
.B(n_2404),
.Y(n_4715)
);

CKINVDCx5p33_ASAP7_75t_R g4716 ( 
.A(n_4442),
.Y(n_4716)
);

NAND2xp5_ASAP7_75t_L g4717 ( 
.A(n_4271),
.B(n_2408),
.Y(n_4717)
);

HB1xp67_ASAP7_75t_L g4718 ( 
.A(n_4273),
.Y(n_4718)
);

INVx1_ASAP7_75t_L g4719 ( 
.A(n_4398),
.Y(n_4719)
);

BUFx6f_ASAP7_75t_L g4720 ( 
.A(n_4450),
.Y(n_4720)
);

BUFx6f_ASAP7_75t_L g4721 ( 
.A(n_4458),
.Y(n_4721)
);

OR2x6_ASAP7_75t_L g4722 ( 
.A(n_4434),
.B(n_1067),
.Y(n_4722)
);

AND2x2_ASAP7_75t_L g4723 ( 
.A(n_4276),
.B(n_2409),
.Y(n_4723)
);

NAND2xp5_ASAP7_75t_SL g4724 ( 
.A(n_4181),
.B(n_2410),
.Y(n_4724)
);

INVx2_ASAP7_75t_L g4725 ( 
.A(n_4398),
.Y(n_4725)
);

NAND2xp33_ASAP7_75t_L g4726 ( 
.A(n_4398),
.B(n_2411),
.Y(n_4726)
);

NAND2xp5_ASAP7_75t_L g4727 ( 
.A(n_4280),
.B(n_2414),
.Y(n_4727)
);

INVx2_ASAP7_75t_L g4728 ( 
.A(n_4444),
.Y(n_4728)
);

AND2x2_ASAP7_75t_L g4729 ( 
.A(n_4281),
.B(n_2415),
.Y(n_4729)
);

HB1xp67_ASAP7_75t_L g4730 ( 
.A(n_4286),
.Y(n_4730)
);

INVx2_ASAP7_75t_L g4731 ( 
.A(n_4428),
.Y(n_4731)
);

INVx2_ASAP7_75t_L g4732 ( 
.A(n_4307),
.Y(n_4732)
);

CKINVDCx20_ASAP7_75t_R g4733 ( 
.A(n_4321),
.Y(n_4733)
);

NAND2xp5_ASAP7_75t_L g4734 ( 
.A(n_4312),
.B(n_2417),
.Y(n_4734)
);

INVxp67_ASAP7_75t_L g4735 ( 
.A(n_4432),
.Y(n_4735)
);

INVx1_ASAP7_75t_L g4736 ( 
.A(n_4376),
.Y(n_4736)
);

INVx3_ASAP7_75t_L g4737 ( 
.A(n_4402),
.Y(n_4737)
);

BUFx4f_ASAP7_75t_L g4738 ( 
.A(n_4346),
.Y(n_4738)
);

INVx1_ASAP7_75t_L g4739 ( 
.A(n_4399),
.Y(n_4739)
);

INVx3_ASAP7_75t_L g4740 ( 
.A(n_4408),
.Y(n_4740)
);

INVx2_ASAP7_75t_L g4741 ( 
.A(n_4290),
.Y(n_4741)
);

AND2x4_ASAP7_75t_L g4742 ( 
.A(n_4255),
.B(n_1069),
.Y(n_4742)
);

INVx2_ASAP7_75t_L g4743 ( 
.A(n_4295),
.Y(n_4743)
);

INVx3_ASAP7_75t_L g4744 ( 
.A(n_4415),
.Y(n_4744)
);

INVx2_ASAP7_75t_L g4745 ( 
.A(n_4341),
.Y(n_4745)
);

NAND2x1_ASAP7_75t_L g4746 ( 
.A(n_4197),
.B(n_1072),
.Y(n_4746)
);

BUFx6f_ASAP7_75t_L g4747 ( 
.A(n_4355),
.Y(n_4747)
);

BUFx3_ASAP7_75t_L g4748 ( 
.A(n_4416),
.Y(n_4748)
);

INVx2_ASAP7_75t_L g4749 ( 
.A(n_4391),
.Y(n_4749)
);

NAND2xp5_ASAP7_75t_L g4750 ( 
.A(n_4429),
.B(n_2418),
.Y(n_4750)
);

AND2x4_ASAP7_75t_L g4751 ( 
.A(n_4426),
.B(n_1073),
.Y(n_4751)
);

HB1xp67_ASAP7_75t_L g4752 ( 
.A(n_4456),
.Y(n_4752)
);

NAND3xp33_ASAP7_75t_L g4753 ( 
.A(n_4201),
.B(n_2433),
.C(n_2427),
.Y(n_4753)
);

INVx2_ASAP7_75t_L g4754 ( 
.A(n_4424),
.Y(n_4754)
);

NAND2xp5_ASAP7_75t_L g4755 ( 
.A(n_4222),
.B(n_2437),
.Y(n_4755)
);

INVx3_ASAP7_75t_L g4756 ( 
.A(n_4464),
.Y(n_4756)
);

INVx3_ASAP7_75t_L g4757 ( 
.A(n_4211),
.Y(n_4757)
);

BUFx6f_ASAP7_75t_L g4758 ( 
.A(n_4439),
.Y(n_4758)
);

INVx1_ASAP7_75t_L g4759 ( 
.A(n_4446),
.Y(n_4759)
);

OR2x2_ASAP7_75t_L g4760 ( 
.A(n_4462),
.B(n_2440),
.Y(n_4760)
);

INVx1_ASAP7_75t_L g4761 ( 
.A(n_4289),
.Y(n_4761)
);

NAND2xp5_ASAP7_75t_L g4762 ( 
.A(n_4180),
.B(n_2444),
.Y(n_4762)
);

INVx1_ASAP7_75t_L g4763 ( 
.A(n_4179),
.Y(n_4763)
);

BUFx6f_ASAP7_75t_L g4764 ( 
.A(n_4188),
.Y(n_4764)
);

INVx1_ASAP7_75t_L g4765 ( 
.A(n_4179),
.Y(n_4765)
);

NAND2xp5_ASAP7_75t_L g4766 ( 
.A(n_4180),
.B(n_2445),
.Y(n_4766)
);

CKINVDCx20_ASAP7_75t_R g4767 ( 
.A(n_4209),
.Y(n_4767)
);

INVx1_ASAP7_75t_L g4768 ( 
.A(n_4179),
.Y(n_4768)
);

INVx1_ASAP7_75t_SL g4769 ( 
.A(n_4224),
.Y(n_4769)
);

BUFx6f_ASAP7_75t_L g4770 ( 
.A(n_4188),
.Y(n_4770)
);

INVx2_ASAP7_75t_L g4771 ( 
.A(n_4179),
.Y(n_4771)
);

AOI221x1_ASAP7_75t_L g4772 ( 
.A1(n_4495),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.C(n_4),
.Y(n_4772)
);

INVx2_ASAP7_75t_L g4773 ( 
.A(n_4473),
.Y(n_4773)
);

INVx2_ASAP7_75t_L g4774 ( 
.A(n_4485),
.Y(n_4774)
);

AOI21x1_ASAP7_75t_L g4775 ( 
.A1(n_4761),
.A2(n_1076),
.B(n_1075),
.Y(n_4775)
);

NAND2xp5_ASAP7_75t_L g4776 ( 
.A(n_4606),
.B(n_2453),
.Y(n_4776)
);

NAND2xp5_ASAP7_75t_L g4777 ( 
.A(n_4587),
.B(n_2460),
.Y(n_4777)
);

NOR2x1_ASAP7_75t_L g4778 ( 
.A(n_4489),
.B(n_2464),
.Y(n_4778)
);

INVx5_ASAP7_75t_L g4779 ( 
.A(n_4636),
.Y(n_4779)
);

OAI21x1_ASAP7_75t_L g4780 ( 
.A1(n_4732),
.A2(n_1079),
.B(n_1077),
.Y(n_4780)
);

NOR4xp25_ASAP7_75t_L g4781 ( 
.A(n_4570),
.B(n_5),
.C(n_3),
.D(n_4),
.Y(n_4781)
);

A2O1A1Ixp33_ASAP7_75t_L g4782 ( 
.A1(n_4505),
.A2(n_2473),
.B(n_2476),
.C(n_2469),
.Y(n_4782)
);

OAI21x1_ASAP7_75t_L g4783 ( 
.A1(n_4731),
.A2(n_1085),
.B(n_1082),
.Y(n_4783)
);

OAI21x1_ASAP7_75t_L g4784 ( 
.A1(n_4538),
.A2(n_1087),
.B(n_1086),
.Y(n_4784)
);

OAI22xp5_ASAP7_75t_L g4785 ( 
.A1(n_4478),
.A2(n_2480),
.B1(n_2481),
.B2(n_2478),
.Y(n_4785)
);

NAND2xp5_ASAP7_75t_L g4786 ( 
.A(n_4493),
.B(n_2483),
.Y(n_4786)
);

OAI21x1_ASAP7_75t_L g4787 ( 
.A1(n_4728),
.A2(n_1094),
.B(n_1091),
.Y(n_4787)
);

AOI21xp5_ASAP7_75t_L g4788 ( 
.A1(n_4566),
.A2(n_1099),
.B(n_1095),
.Y(n_4788)
);

OAI21x1_ASAP7_75t_L g4789 ( 
.A1(n_4725),
.A2(n_1104),
.B(n_1103),
.Y(n_4789)
);

CKINVDCx8_ASAP7_75t_R g4790 ( 
.A(n_4608),
.Y(n_4790)
);

AOI21xp5_ASAP7_75t_L g4791 ( 
.A1(n_4712),
.A2(n_4536),
.B(n_4657),
.Y(n_4791)
);

AOI21xp5_ASAP7_75t_SL g4792 ( 
.A1(n_4687),
.A2(n_2491),
.B(n_2487),
.Y(n_4792)
);

AO31x2_ASAP7_75t_L g4793 ( 
.A1(n_4512),
.A2(n_1108),
.A3(n_1110),
.B(n_1105),
.Y(n_4793)
);

A2O1A1Ixp33_ASAP7_75t_L g4794 ( 
.A1(n_4513),
.A2(n_2502),
.B(n_2505),
.C(n_2498),
.Y(n_4794)
);

OAI21x1_ASAP7_75t_L g4795 ( 
.A1(n_4719),
.A2(n_1113),
.B(n_1111),
.Y(n_4795)
);

BUFx6f_ASAP7_75t_L g4796 ( 
.A(n_4482),
.Y(n_4796)
);

NAND2xp5_ASAP7_75t_L g4797 ( 
.A(n_4509),
.B(n_2513),
.Y(n_4797)
);

INVx1_ASAP7_75t_L g4798 ( 
.A(n_4496),
.Y(n_4798)
);

OAI21x1_ASAP7_75t_L g4799 ( 
.A1(n_4578),
.A2(n_1117),
.B(n_1115),
.Y(n_4799)
);

INVx1_ASAP7_75t_L g4800 ( 
.A(n_4497),
.Y(n_4800)
);

NAND2xp5_ASAP7_75t_L g4801 ( 
.A(n_4574),
.B(n_4604),
.Y(n_4801)
);

NAND2xp5_ASAP7_75t_L g4802 ( 
.A(n_4605),
.B(n_2514),
.Y(n_4802)
);

OAI21x1_ASAP7_75t_SL g4803 ( 
.A1(n_4487),
.A2(n_5),
.B(n_6),
.Y(n_4803)
);

NAND2xp5_ASAP7_75t_L g4804 ( 
.A(n_4515),
.B(n_4718),
.Y(n_4804)
);

NAND2xp5_ASAP7_75t_L g4805 ( 
.A(n_4730),
.B(n_2519),
.Y(n_4805)
);

OR2x6_ASAP7_75t_L g4806 ( 
.A(n_4688),
.B(n_1118),
.Y(n_4806)
);

INVx2_ASAP7_75t_SL g4807 ( 
.A(n_4533),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_4514),
.Y(n_4808)
);

AOI21xp33_ASAP7_75t_L g4809 ( 
.A1(n_4585),
.A2(n_2523),
.B(n_2521),
.Y(n_4809)
);

NAND2xp5_ASAP7_75t_SL g4810 ( 
.A(n_4488),
.B(n_2525),
.Y(n_4810)
);

OAI21xp5_ASAP7_75t_L g4811 ( 
.A1(n_4637),
.A2(n_2530),
.B(n_2526),
.Y(n_4811)
);

AOI21xp5_ASAP7_75t_L g4812 ( 
.A1(n_4659),
.A2(n_1120),
.B(n_1119),
.Y(n_4812)
);

OAI21x1_ASAP7_75t_L g4813 ( 
.A1(n_4681),
.A2(n_1122),
.B(n_1121),
.Y(n_4813)
);

OAI21x1_ASAP7_75t_L g4814 ( 
.A1(n_4741),
.A2(n_1125),
.B(n_1124),
.Y(n_4814)
);

AND2x2_ASAP7_75t_L g4815 ( 
.A(n_4490),
.B(n_2532),
.Y(n_4815)
);

INVx2_ASAP7_75t_L g4816 ( 
.A(n_4527),
.Y(n_4816)
);

AND2x4_ASAP7_75t_L g4817 ( 
.A(n_4619),
.B(n_1126),
.Y(n_4817)
);

INVx2_ASAP7_75t_L g4818 ( 
.A(n_4546),
.Y(n_4818)
);

OAI21x1_ASAP7_75t_L g4819 ( 
.A1(n_4736),
.A2(n_1130),
.B(n_1129),
.Y(n_4819)
);

AND2x2_ASAP7_75t_L g4820 ( 
.A(n_4704),
.B(n_4600),
.Y(n_4820)
);

NAND2xp5_ASAP7_75t_L g4821 ( 
.A(n_4762),
.B(n_2538),
.Y(n_4821)
);

OAI22x1_ASAP7_75t_L g4822 ( 
.A1(n_4695),
.A2(n_2542),
.B1(n_2545),
.B2(n_2541),
.Y(n_4822)
);

OAI22xp5_ASAP7_75t_L g4823 ( 
.A1(n_4539),
.A2(n_2553),
.B1(n_2558),
.B2(n_2550),
.Y(n_4823)
);

OAI22xp5_ASAP7_75t_L g4824 ( 
.A1(n_4560),
.A2(n_2563),
.B1(n_2565),
.B2(n_2560),
.Y(n_4824)
);

HB1xp67_ASAP7_75t_L g4825 ( 
.A(n_4477),
.Y(n_4825)
);

AOI221x1_ASAP7_75t_L g4826 ( 
.A1(n_4677),
.A2(n_4598),
.B1(n_4739),
.B2(n_4559),
.C(n_4757),
.Y(n_4826)
);

AOI21xp5_ASAP7_75t_L g4827 ( 
.A1(n_4571),
.A2(n_1136),
.B(n_1132),
.Y(n_4827)
);

AOI21xp5_ASAP7_75t_L g4828 ( 
.A1(n_4707),
.A2(n_1138),
.B(n_1137),
.Y(n_4828)
);

INVx1_ASAP7_75t_L g4829 ( 
.A(n_4553),
.Y(n_4829)
);

INVx3_ASAP7_75t_L g4830 ( 
.A(n_4548),
.Y(n_4830)
);

AOI22xp5_ASAP7_75t_L g4831 ( 
.A1(n_4531),
.A2(n_2571),
.B1(n_2580),
.B2(n_2567),
.Y(n_4831)
);

AOI21xp5_ASAP7_75t_L g4832 ( 
.A1(n_4523),
.A2(n_1140),
.B(n_1139),
.Y(n_4832)
);

CKINVDCx5p33_ASAP7_75t_R g4833 ( 
.A(n_4767),
.Y(n_4833)
);

AOI21xp5_ASAP7_75t_L g4834 ( 
.A1(n_4726),
.A2(n_1142),
.B(n_1141),
.Y(n_4834)
);

OAI21x1_ASAP7_75t_L g4835 ( 
.A1(n_4746),
.A2(n_1144),
.B(n_1143),
.Y(n_4835)
);

A2O1A1Ixp33_ASAP7_75t_L g4836 ( 
.A1(n_4564),
.A2(n_2583),
.B(n_2585),
.C(n_2582),
.Y(n_4836)
);

AND2x4_ASAP7_75t_L g4837 ( 
.A(n_4480),
.B(n_1149),
.Y(n_4837)
);

AOI22xp5_ASAP7_75t_L g4838 ( 
.A1(n_4703),
.A2(n_2591),
.B1(n_2592),
.B2(n_2590),
.Y(n_4838)
);

AOI21xp5_ASAP7_75t_SL g4839 ( 
.A1(n_4722),
.A2(n_2599),
.B(n_2596),
.Y(n_4839)
);

OAI21xp5_ASAP7_75t_L g4840 ( 
.A1(n_4766),
.A2(n_2602),
.B(n_2601),
.Y(n_4840)
);

NAND2xp5_ASAP7_75t_L g4841 ( 
.A(n_4577),
.B(n_4501),
.Y(n_4841)
);

OA21x2_ASAP7_75t_L g4842 ( 
.A1(n_4596),
.A2(n_2609),
.B(n_2608),
.Y(n_4842)
);

OAI21x1_ASAP7_75t_L g4843 ( 
.A1(n_4743),
.A2(n_1151),
.B(n_1150),
.Y(n_4843)
);

BUFx2_ASAP7_75t_L g4844 ( 
.A(n_4525),
.Y(n_4844)
);

INVxp67_ASAP7_75t_L g4845 ( 
.A(n_4506),
.Y(n_4845)
);

OAI21x1_ASAP7_75t_L g4846 ( 
.A1(n_4689),
.A2(n_1156),
.B(n_1155),
.Y(n_4846)
);

OAI21x1_ASAP7_75t_L g4847 ( 
.A1(n_4670),
.A2(n_1158),
.B(n_1157),
.Y(n_4847)
);

AO31x2_ASAP7_75t_L g4848 ( 
.A1(n_4472),
.A2(n_1160),
.A3(n_1162),
.B(n_1159),
.Y(n_4848)
);

CKINVDCx6p67_ASAP7_75t_R g4849 ( 
.A(n_4626),
.Y(n_4849)
);

NAND2xp5_ASAP7_75t_L g4850 ( 
.A(n_4617),
.B(n_2611),
.Y(n_4850)
);

BUFx6f_ASAP7_75t_L g4851 ( 
.A(n_4533),
.Y(n_4851)
);

NOR2x1_ASAP7_75t_SL g4852 ( 
.A(n_4722),
.B(n_1163),
.Y(n_4852)
);

OAI21xp5_ASAP7_75t_L g4853 ( 
.A1(n_4665),
.A2(n_2619),
.B(n_2617),
.Y(n_4853)
);

OAI21xp5_ASAP7_75t_L g4854 ( 
.A1(n_4671),
.A2(n_2623),
.B(n_2622),
.Y(n_4854)
);

AO31x2_ASAP7_75t_L g4855 ( 
.A1(n_4502),
.A2(n_4503),
.A3(n_4530),
.B(n_4529),
.Y(n_4855)
);

BUFx6f_ASAP7_75t_L g4856 ( 
.A(n_4504),
.Y(n_4856)
);

OA21x2_ASAP7_75t_L g4857 ( 
.A1(n_4528),
.A2(n_4554),
.B(n_4540),
.Y(n_4857)
);

NAND3xp33_ASAP7_75t_L g4858 ( 
.A(n_4584),
.B(n_2640),
.C(n_2631),
.Y(n_4858)
);

NAND2xp5_ASAP7_75t_SL g4859 ( 
.A(n_4748),
.B(n_2641),
.Y(n_4859)
);

AND2x4_ASAP7_75t_L g4860 ( 
.A(n_4479),
.B(n_1165),
.Y(n_4860)
);

NAND2xp5_ASAP7_75t_L g4861 ( 
.A(n_4737),
.B(n_2642),
.Y(n_4861)
);

NAND2xp5_ASAP7_75t_L g4862 ( 
.A(n_4740),
.B(n_2651),
.Y(n_4862)
);

OAI22x1_ASAP7_75t_L g4863 ( 
.A1(n_4745),
.A2(n_2660),
.B1(n_2661),
.B2(n_2659),
.Y(n_4863)
);

AO21x2_ASAP7_75t_L g4864 ( 
.A1(n_4518),
.A2(n_1169),
.B(n_1166),
.Y(n_4864)
);

NOR2xp33_ASAP7_75t_L g4865 ( 
.A(n_4769),
.B(n_2666),
.Y(n_4865)
);

OA21x2_ASAP7_75t_L g4866 ( 
.A1(n_4534),
.A2(n_2670),
.B(n_2669),
.Y(n_4866)
);

NAND2xp5_ASAP7_75t_L g4867 ( 
.A(n_4744),
.B(n_2672),
.Y(n_4867)
);

OAI21x1_ASAP7_75t_L g4868 ( 
.A1(n_4673),
.A2(n_1172),
.B(n_1170),
.Y(n_4868)
);

INVx1_ASAP7_75t_L g4869 ( 
.A(n_4556),
.Y(n_4869)
);

NAND2xp5_ASAP7_75t_L g4870 ( 
.A(n_4476),
.B(n_2673),
.Y(n_4870)
);

AOI21xp5_ASAP7_75t_L g4871 ( 
.A1(n_4519),
.A2(n_1178),
.B(n_1175),
.Y(n_4871)
);

AOI21xp5_ASAP7_75t_L g4872 ( 
.A1(n_4521),
.A2(n_1181),
.B(n_1179),
.Y(n_4872)
);

NOR2xp67_ASAP7_75t_SL g4873 ( 
.A(n_4626),
.B(n_2677),
.Y(n_4873)
);

BUFx3_ASAP7_75t_L g4874 ( 
.A(n_4504),
.Y(n_4874)
);

OAI21xp33_ASAP7_75t_L g4875 ( 
.A1(n_4580),
.A2(n_2683),
.B(n_2679),
.Y(n_4875)
);

NOR2xp33_ASAP7_75t_L g4876 ( 
.A(n_4522),
.B(n_2686),
.Y(n_4876)
);

A2O1A1Ixp33_ASAP7_75t_L g4877 ( 
.A1(n_4714),
.A2(n_2699),
.B(n_2703),
.C(n_2696),
.Y(n_4877)
);

INVx2_ASAP7_75t_L g4878 ( 
.A(n_4567),
.Y(n_4878)
);

A2O1A1Ixp33_ASAP7_75t_L g4879 ( 
.A1(n_4481),
.A2(n_2717),
.B(n_2721),
.C(n_2712),
.Y(n_4879)
);

INVx1_ASAP7_75t_L g4880 ( 
.A(n_4572),
.Y(n_4880)
);

INVx1_ASAP7_75t_L g4881 ( 
.A(n_4589),
.Y(n_4881)
);

INVx3_ASAP7_75t_L g4882 ( 
.A(n_4668),
.Y(n_4882)
);

OAI21x1_ASAP7_75t_L g4883 ( 
.A1(n_4676),
.A2(n_1185),
.B(n_1183),
.Y(n_4883)
);

CKINVDCx5p33_ASAP7_75t_R g4884 ( 
.A(n_4517),
.Y(n_4884)
);

AND2x2_ASAP7_75t_L g4885 ( 
.A(n_4591),
.B(n_2723),
.Y(n_4885)
);

OAI21x1_ASAP7_75t_L g4886 ( 
.A1(n_4684),
.A2(n_1191),
.B(n_1188),
.Y(n_4886)
);

INVx6_ASAP7_75t_SL g4887 ( 
.A(n_4588),
.Y(n_4887)
);

OAI21x1_ASAP7_75t_L g4888 ( 
.A1(n_4685),
.A2(n_1196),
.B(n_1194),
.Y(n_4888)
);

OAI21xp5_ASAP7_75t_L g4889 ( 
.A1(n_4674),
.A2(n_2726),
.B(n_2725),
.Y(n_4889)
);

INVx3_ASAP7_75t_L g4890 ( 
.A(n_4552),
.Y(n_4890)
);

AO31x2_ASAP7_75t_L g4891 ( 
.A1(n_4537),
.A2(n_1198),
.A3(n_1199),
.B(n_1197),
.Y(n_4891)
);

INVxp67_ASAP7_75t_L g4892 ( 
.A(n_4511),
.Y(n_4892)
);

AO31x2_ASAP7_75t_L g4893 ( 
.A1(n_4541),
.A2(n_1207),
.A3(n_1208),
.B(n_1201),
.Y(n_4893)
);

NAND2xp5_ASAP7_75t_L g4894 ( 
.A(n_4723),
.B(n_2740),
.Y(n_4894)
);

AND2x4_ASAP7_75t_L g4895 ( 
.A(n_4569),
.B(n_1210),
.Y(n_4895)
);

AOI21xp5_ASAP7_75t_L g4896 ( 
.A1(n_4631),
.A2(n_1212),
.B(n_1211),
.Y(n_4896)
);

OR2x2_ASAP7_75t_L g4897 ( 
.A(n_4542),
.B(n_2741),
.Y(n_4897)
);

AND2x2_ASAP7_75t_L g4898 ( 
.A(n_4706),
.B(n_2742),
.Y(n_4898)
);

OAI21x1_ASAP7_75t_L g4899 ( 
.A1(n_4686),
.A2(n_1215),
.B(n_1214),
.Y(n_4899)
);

INVx5_ASAP7_75t_L g4900 ( 
.A(n_4636),
.Y(n_4900)
);

AOI21xp5_ASAP7_75t_L g4901 ( 
.A1(n_4563),
.A2(n_1217),
.B(n_1216),
.Y(n_4901)
);

OAI21x1_ASAP7_75t_L g4902 ( 
.A1(n_4701),
.A2(n_1221),
.B(n_1218),
.Y(n_4902)
);

AND2x2_ASAP7_75t_L g4903 ( 
.A(n_4709),
.B(n_2746),
.Y(n_4903)
);

OAI21x1_ASAP7_75t_L g4904 ( 
.A1(n_4711),
.A2(n_1226),
.B(n_1224),
.Y(n_4904)
);

AO21x1_ASAP7_75t_L g4905 ( 
.A1(n_4755),
.A2(n_6),
.B(n_7),
.Y(n_4905)
);

NOR2xp33_ASAP7_75t_L g4906 ( 
.A(n_4551),
.B(n_4547),
.Y(n_4906)
);

INVx1_ASAP7_75t_L g4907 ( 
.A(n_4594),
.Y(n_4907)
);

NOR2xp67_ASAP7_75t_SL g4908 ( 
.A(n_4627),
.B(n_4624),
.Y(n_4908)
);

NAND2xp5_ASAP7_75t_L g4909 ( 
.A(n_4729),
.B(n_2748),
.Y(n_4909)
);

OAI21x1_ASAP7_75t_L g4910 ( 
.A1(n_4656),
.A2(n_1228),
.B(n_1227),
.Y(n_4910)
);

AND2x4_ASAP7_75t_L g4911 ( 
.A(n_4622),
.B(n_4545),
.Y(n_4911)
);

NAND2xp5_ASAP7_75t_L g4912 ( 
.A(n_4700),
.B(n_2750),
.Y(n_4912)
);

AOI21xp5_ASAP7_75t_L g4913 ( 
.A1(n_4724),
.A2(n_1234),
.B(n_1233),
.Y(n_4913)
);

OAI21x1_ASAP7_75t_L g4914 ( 
.A1(n_4544),
.A2(n_1240),
.B(n_1235),
.Y(n_4914)
);

A2O1A1Ixp33_ASAP7_75t_L g4915 ( 
.A1(n_4753),
.A2(n_4713),
.B(n_4749),
.C(n_4508),
.Y(n_4915)
);

OAI21xp33_ASAP7_75t_L g4916 ( 
.A1(n_4667),
.A2(n_2763),
.B(n_2757),
.Y(n_4916)
);

AOI21xp5_ASAP7_75t_L g4917 ( 
.A1(n_4679),
.A2(n_1246),
.B(n_1242),
.Y(n_4917)
);

NAND2xp5_ASAP7_75t_L g4918 ( 
.A(n_4593),
.B(n_2765),
.Y(n_4918)
);

OAI21x1_ASAP7_75t_L g4919 ( 
.A1(n_4549),
.A2(n_4562),
.B(n_4550),
.Y(n_4919)
);

AND2x4_ASAP7_75t_L g4920 ( 
.A(n_4558),
.B(n_1248),
.Y(n_4920)
);

AOI21xp5_ASAP7_75t_L g4921 ( 
.A1(n_4579),
.A2(n_1252),
.B(n_1250),
.Y(n_4921)
);

AO31x2_ASAP7_75t_L g4922 ( 
.A1(n_4599),
.A2(n_1256),
.A3(n_1257),
.B(n_1253),
.Y(n_4922)
);

OA22x2_ASAP7_75t_L g4923 ( 
.A1(n_4588),
.A2(n_2770),
.B1(n_2773),
.B2(n_2769),
.Y(n_4923)
);

AO21x2_ASAP7_75t_L g4924 ( 
.A1(n_4603),
.A2(n_1259),
.B(n_1258),
.Y(n_4924)
);

OAI21x1_ASAP7_75t_L g4925 ( 
.A1(n_4601),
.A2(n_1264),
.B(n_1263),
.Y(n_4925)
);

AOI21xp5_ASAP7_75t_L g4926 ( 
.A1(n_4646),
.A2(n_1266),
.B(n_1265),
.Y(n_4926)
);

AOI21xp5_ASAP7_75t_L g4927 ( 
.A1(n_4555),
.A2(n_1269),
.B(n_1268),
.Y(n_4927)
);

OAI21x1_ASAP7_75t_L g4928 ( 
.A1(n_4763),
.A2(n_1272),
.B(n_1271),
.Y(n_4928)
);

INVx1_ASAP7_75t_L g4929 ( 
.A(n_4771),
.Y(n_4929)
);

NAND2xp5_ASAP7_75t_SL g4930 ( 
.A(n_4649),
.B(n_2774),
.Y(n_4930)
);

INVx1_ASAP7_75t_L g4931 ( 
.A(n_4765),
.Y(n_4931)
);

NOR2x1_ASAP7_75t_SL g4932 ( 
.A(n_4483),
.B(n_1273),
.Y(n_4932)
);

AO21x1_ASAP7_75t_L g4933 ( 
.A1(n_4607),
.A2(n_7),
.B(n_8),
.Y(n_4933)
);

OAI22xp5_ASAP7_75t_L g4934 ( 
.A1(n_4568),
.A2(n_2779),
.B1(n_2782),
.B2(n_2778),
.Y(n_4934)
);

AOI21xp5_ASAP7_75t_L g4935 ( 
.A1(n_4754),
.A2(n_1275),
.B(n_1274),
.Y(n_4935)
);

NAND2xp5_ASAP7_75t_L g4936 ( 
.A(n_4699),
.B(n_2788),
.Y(n_4936)
);

AO31x2_ASAP7_75t_L g4937 ( 
.A1(n_4768),
.A2(n_4759),
.A3(n_4612),
.B(n_4620),
.Y(n_4937)
);

AND2x4_ASAP7_75t_L g4938 ( 
.A(n_4582),
.B(n_1276),
.Y(n_4938)
);

NAND2xp5_ASAP7_75t_L g4939 ( 
.A(n_4616),
.B(n_2791),
.Y(n_4939)
);

INVx6_ASAP7_75t_L g4940 ( 
.A(n_4627),
.Y(n_4940)
);

NAND2xp5_ASAP7_75t_L g4941 ( 
.A(n_4635),
.B(n_2792),
.Y(n_4941)
);

OAI21x1_ASAP7_75t_L g4942 ( 
.A1(n_4609),
.A2(n_1278),
.B(n_1277),
.Y(n_4942)
);

AO31x2_ASAP7_75t_L g4943 ( 
.A1(n_4628),
.A2(n_1284),
.A3(n_1285),
.B(n_1282),
.Y(n_4943)
);

AOI21xp5_ASAP7_75t_L g4944 ( 
.A1(n_4715),
.A2(n_1288),
.B(n_1286),
.Y(n_4944)
);

INVx2_ASAP7_75t_L g4945 ( 
.A(n_4611),
.Y(n_4945)
);

NAND2xp5_ASAP7_75t_SL g4946 ( 
.A(n_4738),
.B(n_2797),
.Y(n_4946)
);

OAI22xp5_ASAP7_75t_L g4947 ( 
.A1(n_4733),
.A2(n_2802),
.B1(n_2804),
.B2(n_2799),
.Y(n_4947)
);

AOI21x1_ASAP7_75t_L g4948 ( 
.A1(n_4752),
.A2(n_1290),
.B(n_1289),
.Y(n_4948)
);

NOR2xp33_ASAP7_75t_L g4949 ( 
.A(n_4499),
.B(n_2805),
.Y(n_4949)
);

NAND2x1_ASAP7_75t_L g4950 ( 
.A(n_4640),
.B(n_1291),
.Y(n_4950)
);

INVx1_ASAP7_75t_L g4951 ( 
.A(n_4705),
.Y(n_4951)
);

AOI21xp5_ASAP7_75t_L g4952 ( 
.A1(n_4717),
.A2(n_1295),
.B(n_1294),
.Y(n_4952)
);

AOI21xp5_ASAP7_75t_L g4953 ( 
.A1(n_4727),
.A2(n_1298),
.B(n_1297),
.Y(n_4953)
);

HB1xp67_ASAP7_75t_L g4954 ( 
.A(n_4475),
.Y(n_4954)
);

AOI22xp33_ASAP7_75t_SL g4955 ( 
.A1(n_4640),
.A2(n_2810),
.B1(n_2812),
.B2(n_2809),
.Y(n_4955)
);

OAI21x1_ASAP7_75t_L g4956 ( 
.A1(n_4602),
.A2(n_1301),
.B(n_1299),
.Y(n_4956)
);

NAND2xp5_ASAP7_75t_L g4957 ( 
.A(n_4641),
.B(n_8),
.Y(n_4957)
);

AOI221xp5_ASAP7_75t_SL g4958 ( 
.A1(n_4583),
.A2(n_12),
.B1(n_9),
.B2(n_11),
.C(n_13),
.Y(n_4958)
);

OAI21x1_ASAP7_75t_L g4959 ( 
.A1(n_4651),
.A2(n_1304),
.B(n_1302),
.Y(n_4959)
);

AO22x2_ASAP7_75t_L g4960 ( 
.A1(n_4760),
.A2(n_15),
.B1(n_9),
.B2(n_14),
.Y(n_4960)
);

OAI21xp5_ASAP7_75t_L g4961 ( 
.A1(n_4630),
.A2(n_16),
.B(n_17),
.Y(n_4961)
);

NAND2xp5_ASAP7_75t_L g4962 ( 
.A(n_4638),
.B(n_4581),
.Y(n_4962)
);

CKINVDCx12_ASAP7_75t_R g4963 ( 
.A(n_4690),
.Y(n_4963)
);

BUFx6f_ASAP7_75t_L g4964 ( 
.A(n_4494),
.Y(n_4964)
);

OAI21xp5_ASAP7_75t_L g4965 ( 
.A1(n_4696),
.A2(n_18),
.B(n_19),
.Y(n_4965)
);

OAI22xp5_ASAP7_75t_L g4966 ( 
.A1(n_4516),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_4966)
);

NAND2xp5_ASAP7_75t_L g4967 ( 
.A(n_4615),
.B(n_21),
.Y(n_4967)
);

NAND3x1_ASAP7_75t_L g4968 ( 
.A(n_4675),
.B(n_21),
.C(n_22),
.Y(n_4968)
);

AOI21xp5_ASAP7_75t_L g4969 ( 
.A1(n_4643),
.A2(n_4756),
.B(n_4734),
.Y(n_4969)
);

OAI21xp5_ASAP7_75t_L g4970 ( 
.A1(n_4682),
.A2(n_22),
.B(n_23),
.Y(n_4970)
);

NAND2xp5_ASAP7_75t_L g4971 ( 
.A(n_4500),
.B(n_23),
.Y(n_4971)
);

NOR2xp33_ASAP7_75t_L g4972 ( 
.A(n_4510),
.B(n_1306),
.Y(n_4972)
);

AND2x4_ASAP7_75t_L g4973 ( 
.A(n_4586),
.B(n_1308),
.Y(n_4973)
);

NAND2xp5_ASAP7_75t_L g4974 ( 
.A(n_4614),
.B(n_24),
.Y(n_4974)
);

INVx1_ASAP7_75t_SL g4975 ( 
.A(n_4623),
.Y(n_4975)
);

OAI21xp5_ASAP7_75t_L g4976 ( 
.A1(n_4750),
.A2(n_4640),
.B(n_4735),
.Y(n_4976)
);

NOR2xp33_ASAP7_75t_L g4977 ( 
.A(n_4573),
.B(n_1309),
.Y(n_4977)
);

OAI21xp5_ASAP7_75t_L g4978 ( 
.A1(n_4710),
.A2(n_25),
.B(n_26),
.Y(n_4978)
);

AOI21xp5_ASAP7_75t_L g4979 ( 
.A1(n_4751),
.A2(n_4742),
.B(n_4758),
.Y(n_4979)
);

AOI21xp5_ASAP7_75t_L g4980 ( 
.A1(n_4758),
.A2(n_1312),
.B(n_1311),
.Y(n_4980)
);

INVx1_ASAP7_75t_L g4981 ( 
.A(n_4661),
.Y(n_4981)
);

INVx4_ASAP7_75t_L g4982 ( 
.A(n_4494),
.Y(n_4982)
);

OAI22xp5_ASAP7_75t_L g4983 ( 
.A1(n_4660),
.A2(n_4691),
.B1(n_4716),
.B2(n_4653),
.Y(n_4983)
);

AO31x2_ASAP7_75t_L g4984 ( 
.A1(n_4669),
.A2(n_1315),
.A3(n_1318),
.B(n_1314),
.Y(n_4984)
);

INVx3_ASAP7_75t_L g4985 ( 
.A(n_4644),
.Y(n_4985)
);

OAI21x1_ASAP7_75t_L g4986 ( 
.A1(n_4678),
.A2(n_1321),
.B(n_1319),
.Y(n_4986)
);

NAND2xp5_ASAP7_75t_L g4987 ( 
.A(n_4592),
.B(n_27),
.Y(n_4987)
);

AO21x1_ASAP7_75t_L g4988 ( 
.A1(n_4708),
.A2(n_27),
.B(n_28),
.Y(n_4988)
);

OAI21xp5_ASAP7_75t_L g4989 ( 
.A1(n_4648),
.A2(n_29),
.B(n_30),
.Y(n_4989)
);

AND2x2_ASAP7_75t_L g4990 ( 
.A(n_4632),
.B(n_30),
.Y(n_4990)
);

AND3x4_ASAP7_75t_L g4991 ( 
.A(n_4535),
.B(n_31),
.C(n_32),
.Y(n_4991)
);

AO31x2_ASAP7_75t_L g4992 ( 
.A1(n_4693),
.A2(n_1324),
.A3(n_1325),
.B(n_1322),
.Y(n_4992)
);

NOR2x1_ASAP7_75t_SL g4993 ( 
.A(n_4483),
.B(n_1326),
.Y(n_4993)
);

INVx2_ASAP7_75t_SL g4994 ( 
.A(n_4498),
.Y(n_4994)
);

NAND2xp5_ASAP7_75t_L g4995 ( 
.A(n_4683),
.B(n_31),
.Y(n_4995)
);

INVx2_ASAP7_75t_SL g4996 ( 
.A(n_4498),
.Y(n_4996)
);

HB1xp67_ASAP7_75t_L g4997 ( 
.A(n_4532),
.Y(n_4997)
);

NOR2xp33_ASAP7_75t_L g4998 ( 
.A(n_4747),
.B(n_1329),
.Y(n_4998)
);

OAI21x1_ASAP7_75t_L g4999 ( 
.A1(n_4666),
.A2(n_1331),
.B(n_1330),
.Y(n_4999)
);

OAI21x1_ASAP7_75t_L g5000 ( 
.A1(n_4618),
.A2(n_1335),
.B(n_1332),
.Y(n_5000)
);

AO31x2_ASAP7_75t_L g5001 ( 
.A1(n_4672),
.A2(n_1340),
.A3(n_1341),
.B(n_1338),
.Y(n_5001)
);

NAND2xp5_ASAP7_75t_L g5002 ( 
.A(n_4652),
.B(n_32),
.Y(n_5002)
);

OAI21x1_ASAP7_75t_L g5003 ( 
.A1(n_4654),
.A2(n_1345),
.B(n_1343),
.Y(n_5003)
);

A2O1A1Ixp33_ASAP7_75t_L g5004 ( 
.A1(n_4576),
.A2(n_36),
.B(n_33),
.C(n_35),
.Y(n_5004)
);

AO31x2_ASAP7_75t_L g5005 ( 
.A1(n_4629),
.A2(n_1348),
.A3(n_1350),
.B(n_1347),
.Y(n_5005)
);

NAND2x1p5_ASAP7_75t_L g5006 ( 
.A(n_4779),
.B(n_4595),
.Y(n_5006)
);

AND2x4_ASAP7_75t_L g5007 ( 
.A(n_4844),
.B(n_4524),
.Y(n_5007)
);

BUFx2_ASAP7_75t_L g5008 ( 
.A(n_4825),
.Y(n_5008)
);

NOR2xp67_ASAP7_75t_SL g5009 ( 
.A(n_4792),
.B(n_4633),
.Y(n_5009)
);

NAND3xp33_ASAP7_75t_L g5010 ( 
.A(n_4961),
.B(n_4680),
.C(n_4645),
.Y(n_5010)
);

OAI22xp5_ASAP7_75t_L g5011 ( 
.A1(n_4915),
.A2(n_4655),
.B1(n_4663),
.B2(n_4747),
.Y(n_5011)
);

NAND2xp5_ASAP7_75t_L g5012 ( 
.A(n_4801),
.B(n_4697),
.Y(n_5012)
);

INVx2_ASAP7_75t_L g5013 ( 
.A(n_4773),
.Y(n_5013)
);

INVx2_ASAP7_75t_L g5014 ( 
.A(n_4774),
.Y(n_5014)
);

HB1xp67_ASAP7_75t_L g5015 ( 
.A(n_4951),
.Y(n_5015)
);

AND2x2_ASAP7_75t_L g5016 ( 
.A(n_4820),
.B(n_4565),
.Y(n_5016)
);

INVx5_ASAP7_75t_L g5017 ( 
.A(n_4796),
.Y(n_5017)
);

OR2x6_ASAP7_75t_L g5018 ( 
.A(n_4806),
.B(n_4688),
.Y(n_5018)
);

BUFx10_ASAP7_75t_L g5019 ( 
.A(n_4884),
.Y(n_5019)
);

HB1xp67_ASAP7_75t_L g5020 ( 
.A(n_4855),
.Y(n_5020)
);

HB1xp67_ASAP7_75t_L g5021 ( 
.A(n_4855),
.Y(n_5021)
);

INVxp67_ASAP7_75t_SL g5022 ( 
.A(n_4857),
.Y(n_5022)
);

BUFx6f_ASAP7_75t_L g5023 ( 
.A(n_4796),
.Y(n_5023)
);

NAND2x1_ASAP7_75t_L g5024 ( 
.A(n_4969),
.B(n_4690),
.Y(n_5024)
);

OAI21xp33_ASAP7_75t_L g5025 ( 
.A1(n_4965),
.A2(n_4662),
.B(n_4639),
.Y(n_5025)
);

BUFx2_ASAP7_75t_L g5026 ( 
.A(n_4954),
.Y(n_5026)
);

INVx1_ASAP7_75t_L g5027 ( 
.A(n_4937),
.Y(n_5027)
);

AO32x2_ASAP7_75t_L g5028 ( 
.A1(n_4966),
.A2(n_4590),
.A3(n_4486),
.B1(n_4491),
.B2(n_4597),
.Y(n_5028)
);

INVx2_ASAP7_75t_SL g5029 ( 
.A(n_4779),
.Y(n_5029)
);

A2O1A1Ixp33_ASAP7_75t_L g5030 ( 
.A1(n_4978),
.A2(n_4692),
.B(n_4543),
.C(n_4507),
.Y(n_5030)
);

INVx2_ASAP7_75t_SL g5031 ( 
.A(n_4900),
.Y(n_5031)
);

BUFx2_ASAP7_75t_L g5032 ( 
.A(n_4892),
.Y(n_5032)
);

INVx3_ASAP7_75t_L g5033 ( 
.A(n_4882),
.Y(n_5033)
);

INVx3_ASAP7_75t_L g5034 ( 
.A(n_4790),
.Y(n_5034)
);

AND2x4_ASAP7_75t_L g5035 ( 
.A(n_4900),
.B(n_4621),
.Y(n_5035)
);

NOR2xp33_ASAP7_75t_L g5036 ( 
.A(n_4962),
.B(n_4474),
.Y(n_5036)
);

NOR2xp67_ASAP7_75t_L g5037 ( 
.A(n_4830),
.B(n_4557),
.Y(n_5037)
);

NAND2x1p5_ASAP7_75t_L g5038 ( 
.A(n_4908),
.B(n_4520),
.Y(n_5038)
);

AND2x2_ASAP7_75t_L g5039 ( 
.A(n_4804),
.B(n_4698),
.Y(n_5039)
);

NAND2xp5_ASAP7_75t_L g5040 ( 
.A(n_4841),
.B(n_4698),
.Y(n_5040)
);

INVx3_ASAP7_75t_L g5041 ( 
.A(n_4982),
.Y(n_5041)
);

NAND2xp5_ASAP7_75t_L g5042 ( 
.A(n_4845),
.B(n_4702),
.Y(n_5042)
);

NOR2xp67_ASAP7_75t_SL g5043 ( 
.A(n_4839),
.B(n_4610),
.Y(n_5043)
);

BUFx10_ASAP7_75t_L g5044 ( 
.A(n_4833),
.Y(n_5044)
);

AND2x2_ASAP7_75t_L g5045 ( 
.A(n_4990),
.B(n_4702),
.Y(n_5045)
);

INVx1_ASAP7_75t_L g5046 ( 
.A(n_4937),
.Y(n_5046)
);

AND2x2_ASAP7_75t_L g5047 ( 
.A(n_4816),
.B(n_4818),
.Y(n_5047)
);

INVx1_ASAP7_75t_L g5048 ( 
.A(n_4931),
.Y(n_5048)
);

NOR2xp33_ASAP7_75t_SL g5049 ( 
.A(n_4906),
.B(n_4575),
.Y(n_5049)
);

INVx2_ASAP7_75t_L g5050 ( 
.A(n_4878),
.Y(n_5050)
);

CKINVDCx5p33_ASAP7_75t_R g5051 ( 
.A(n_4849),
.Y(n_5051)
);

A2O1A1Ixp33_ASAP7_75t_SL g5052 ( 
.A1(n_4970),
.A2(n_4613),
.B(n_4484),
.C(n_4561),
.Y(n_5052)
);

AND2x2_ASAP7_75t_L g5053 ( 
.A(n_4945),
.B(n_4658),
.Y(n_5053)
);

INVx1_ASAP7_75t_SL g5054 ( 
.A(n_4975),
.Y(n_5054)
);

NAND2xp5_ASAP7_75t_L g5055 ( 
.A(n_4791),
.B(n_4979),
.Y(n_5055)
);

BUFx6f_ASAP7_75t_L g5056 ( 
.A(n_4851),
.Y(n_5056)
);

INVx2_ASAP7_75t_L g5057 ( 
.A(n_4919),
.Y(n_5057)
);

HB1xp67_ASAP7_75t_L g5058 ( 
.A(n_4997),
.Y(n_5058)
);

NAND2xp5_ASAP7_75t_SL g5059 ( 
.A(n_4976),
.B(n_4664),
.Y(n_5059)
);

INVxp67_ASAP7_75t_L g5060 ( 
.A(n_4815),
.Y(n_5060)
);

INVx2_ASAP7_75t_SL g5061 ( 
.A(n_4940),
.Y(n_5061)
);

INVx2_ASAP7_75t_L g5062 ( 
.A(n_4798),
.Y(n_5062)
);

NOR2xp33_ASAP7_75t_L g5063 ( 
.A(n_4870),
.B(n_4652),
.Y(n_5063)
);

OR2x6_ASAP7_75t_L g5064 ( 
.A(n_4806),
.B(n_4492),
.Y(n_5064)
);

INVx1_ASAP7_75t_L g5065 ( 
.A(n_4800),
.Y(n_5065)
);

NAND2xp5_ASAP7_75t_SL g5066 ( 
.A(n_4776),
.B(n_4664),
.Y(n_5066)
);

AND2x2_ASAP7_75t_L g5067 ( 
.A(n_4960),
.B(n_4634),
.Y(n_5067)
);

INVx2_ASAP7_75t_L g5068 ( 
.A(n_4808),
.Y(n_5068)
);

AOI22xp5_ASAP7_75t_L g5069 ( 
.A1(n_4963),
.A2(n_4912),
.B1(n_4810),
.B2(n_4811),
.Y(n_5069)
);

OAI22xp5_ASAP7_75t_L g5070 ( 
.A1(n_4831),
.A2(n_4492),
.B1(n_4650),
.B2(n_4642),
.Y(n_5070)
);

BUFx12f_ASAP7_75t_L g5071 ( 
.A(n_4851),
.Y(n_5071)
);

NAND2xp5_ASAP7_75t_L g5072 ( 
.A(n_4981),
.B(n_4694),
.Y(n_5072)
);

BUFx2_ASAP7_75t_L g5073 ( 
.A(n_4887),
.Y(n_5073)
);

INVx2_ASAP7_75t_L g5074 ( 
.A(n_4829),
.Y(n_5074)
);

INVx3_ASAP7_75t_L g5075 ( 
.A(n_4874),
.Y(n_5075)
);

AND2x2_ASAP7_75t_L g5076 ( 
.A(n_4869),
.B(n_4526),
.Y(n_5076)
);

INVx2_ASAP7_75t_L g5077 ( 
.A(n_4880),
.Y(n_5077)
);

AND2x4_ASAP7_75t_L g5078 ( 
.A(n_4890),
.B(n_4985),
.Y(n_5078)
);

NAND2xp5_ASAP7_75t_L g5079 ( 
.A(n_4881),
.B(n_4647),
.Y(n_5079)
);

AOI21xp5_ASAP7_75t_L g5080 ( 
.A1(n_4834),
.A2(n_4721),
.B(n_4720),
.Y(n_5080)
);

AOI21xp33_ASAP7_75t_L g5081 ( 
.A1(n_4842),
.A2(n_4647),
.B(n_4625),
.Y(n_5081)
);

INVx1_ASAP7_75t_L g5082 ( 
.A(n_4907),
.Y(n_5082)
);

INVx1_ASAP7_75t_L g5083 ( 
.A(n_4929),
.Y(n_5083)
);

NAND2xp5_ASAP7_75t_SL g5084 ( 
.A(n_4983),
.B(n_4621),
.Y(n_5084)
);

AOI22xp5_ASAP7_75t_L g5085 ( 
.A1(n_4989),
.A2(n_4610),
.B1(n_4644),
.B2(n_4720),
.Y(n_5085)
);

NAND2xp5_ASAP7_75t_L g5086 ( 
.A(n_4786),
.B(n_4764),
.Y(n_5086)
);

OR2x2_ASAP7_75t_L g5087 ( 
.A(n_4936),
.B(n_4897),
.Y(n_5087)
);

INVx1_ASAP7_75t_L g5088 ( 
.A(n_4974),
.Y(n_5088)
);

CKINVDCx20_ASAP7_75t_R g5089 ( 
.A(n_4977),
.Y(n_5089)
);

AOI21xp5_ASAP7_75t_L g5090 ( 
.A1(n_4826),
.A2(n_4721),
.B(n_4764),
.Y(n_5090)
);

AND2x4_ASAP7_75t_L g5091 ( 
.A(n_4807),
.B(n_4770),
.Y(n_5091)
);

AOI21xp5_ASAP7_75t_L g5092 ( 
.A1(n_4788),
.A2(n_4770),
.B(n_1354),
.Y(n_5092)
);

INVx1_ASAP7_75t_L g5093 ( 
.A(n_4793),
.Y(n_5093)
);

BUFx6f_ASAP7_75t_L g5094 ( 
.A(n_4856),
.Y(n_5094)
);

INVx2_ASAP7_75t_L g5095 ( 
.A(n_4787),
.Y(n_5095)
);

AND2x4_ASAP7_75t_L g5096 ( 
.A(n_4911),
.B(n_1351),
.Y(n_5096)
);

NAND2xp5_ASAP7_75t_L g5097 ( 
.A(n_4802),
.B(n_33),
.Y(n_5097)
);

INVx1_ASAP7_75t_SL g5098 ( 
.A(n_4856),
.Y(n_5098)
);

INVx2_ASAP7_75t_L g5099 ( 
.A(n_4984),
.Y(n_5099)
);

NAND2xp5_ASAP7_75t_L g5100 ( 
.A(n_4797),
.B(n_35),
.Y(n_5100)
);

HB1xp67_ASAP7_75t_L g5101 ( 
.A(n_4864),
.Y(n_5101)
);

AOI22xp33_ASAP7_75t_SL g5102 ( 
.A1(n_4852),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_5102)
);

INVx2_ASAP7_75t_L g5103 ( 
.A(n_4984),
.Y(n_5103)
);

NAND2xp5_ASAP7_75t_SL g5104 ( 
.A(n_4957),
.B(n_1359),
.Y(n_5104)
);

INVx1_ASAP7_75t_L g5105 ( 
.A(n_4793),
.Y(n_5105)
);

HB1xp67_ASAP7_75t_L g5106 ( 
.A(n_4971),
.Y(n_5106)
);

NAND2xp5_ASAP7_75t_L g5107 ( 
.A(n_4958),
.B(n_37),
.Y(n_5107)
);

A2O1A1Ixp33_ASAP7_75t_L g5108 ( 
.A1(n_4836),
.A2(n_40),
.B(n_38),
.C(n_39),
.Y(n_5108)
);

AND2x2_ASAP7_75t_L g5109 ( 
.A(n_4866),
.B(n_4998),
.Y(n_5109)
);

OAI21xp33_ASAP7_75t_L g5110 ( 
.A1(n_4809),
.A2(n_39),
.B(n_41),
.Y(n_5110)
);

HB1xp67_ASAP7_75t_L g5111 ( 
.A(n_4967),
.Y(n_5111)
);

AOI21xp5_ASAP7_75t_L g5112 ( 
.A1(n_4772),
.A2(n_1365),
.B(n_1362),
.Y(n_5112)
);

BUFx6f_ASAP7_75t_L g5113 ( 
.A(n_4964),
.Y(n_5113)
);

OAI21x1_ASAP7_75t_SL g5114 ( 
.A1(n_4988),
.A2(n_41),
.B(n_43),
.Y(n_5114)
);

INVx2_ASAP7_75t_L g5115 ( 
.A(n_4992),
.Y(n_5115)
);

BUFx8_ASAP7_75t_L g5116 ( 
.A(n_4964),
.Y(n_5116)
);

BUFx12f_ASAP7_75t_L g5117 ( 
.A(n_4837),
.Y(n_5117)
);

A2O1A1Ixp33_ASAP7_75t_L g5118 ( 
.A1(n_5004),
.A2(n_47),
.B(n_45),
.C(n_46),
.Y(n_5118)
);

NOR2xp33_ASAP7_75t_L g5119 ( 
.A(n_4949),
.B(n_1366),
.Y(n_5119)
);

INVx3_ASAP7_75t_L g5120 ( 
.A(n_4994),
.Y(n_5120)
);

NAND2xp5_ASAP7_75t_L g5121 ( 
.A(n_4850),
.B(n_45),
.Y(n_5121)
);

NAND2xp5_ASAP7_75t_SL g5122 ( 
.A(n_4896),
.B(n_1373),
.Y(n_5122)
);

NAND2xp5_ASAP7_75t_L g5123 ( 
.A(n_4777),
.B(n_46),
.Y(n_5123)
);

OAI22xp5_ASAP7_75t_L g5124 ( 
.A1(n_4955),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_5124)
);

OAI21x1_ASAP7_75t_L g5125 ( 
.A1(n_4784),
.A2(n_1376),
.B(n_1374),
.Y(n_5125)
);

AOI22xp5_ASAP7_75t_L g5126 ( 
.A1(n_4946),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_5126)
);

NOR2x1_ASAP7_75t_SL g5127 ( 
.A(n_4924),
.B(n_1377),
.Y(n_5127)
);

AOI22xp33_ASAP7_75t_L g5128 ( 
.A1(n_4905),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_5128)
);

INVx2_ASAP7_75t_L g5129 ( 
.A(n_4992),
.Y(n_5129)
);

INVx1_ASAP7_75t_L g5130 ( 
.A(n_5001),
.Y(n_5130)
);

AOI222xp33_ASAP7_75t_L g5131 ( 
.A1(n_4875),
.A2(n_54),
.B1(n_57),
.B2(n_52),
.C1(n_53),
.C2(n_55),
.Y(n_5131)
);

CKINVDCx11_ASAP7_75t_R g5132 ( 
.A(n_4817),
.Y(n_5132)
);

CKINVDCx20_ASAP7_75t_R g5133 ( 
.A(n_4930),
.Y(n_5133)
);

INVx3_ASAP7_75t_L g5134 ( 
.A(n_4996),
.Y(n_5134)
);

AOI21xp5_ASAP7_75t_L g5135 ( 
.A1(n_4812),
.A2(n_1380),
.B(n_1378),
.Y(n_5135)
);

AOI21xp5_ASAP7_75t_L g5136 ( 
.A1(n_4871),
.A2(n_1384),
.B(n_1382),
.Y(n_5136)
);

NOR2xp67_ASAP7_75t_SL g5137 ( 
.A(n_4980),
.B(n_4872),
.Y(n_5137)
);

INVx1_ASAP7_75t_L g5138 ( 
.A(n_5001),
.Y(n_5138)
);

CKINVDCx5p33_ASAP7_75t_R g5139 ( 
.A(n_4822),
.Y(n_5139)
);

AND2x2_ASAP7_75t_L g5140 ( 
.A(n_4995),
.B(n_1385),
.Y(n_5140)
);

NAND2xp5_ASAP7_75t_L g5141 ( 
.A(n_4821),
.B(n_53),
.Y(n_5141)
);

INVx1_ASAP7_75t_L g5142 ( 
.A(n_4943),
.Y(n_5142)
);

AND2x2_ASAP7_75t_L g5143 ( 
.A(n_4972),
.B(n_1387),
.Y(n_5143)
);

BUFx6f_ASAP7_75t_L g5144 ( 
.A(n_4895),
.Y(n_5144)
);

INVx5_ASAP7_75t_L g5145 ( 
.A(n_4973),
.Y(n_5145)
);

INVx1_ASAP7_75t_L g5146 ( 
.A(n_4943),
.Y(n_5146)
);

AOI22xp33_ASAP7_75t_L g5147 ( 
.A1(n_4933),
.A2(n_57),
.B1(n_54),
.B2(n_55),
.Y(n_5147)
);

BUFx2_ASAP7_75t_L g5148 ( 
.A(n_4860),
.Y(n_5148)
);

NAND2xp5_ASAP7_75t_L g5149 ( 
.A(n_4781),
.B(n_58),
.Y(n_5149)
);

OAI22xp5_ASAP7_75t_SL g5150 ( 
.A1(n_4991),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_5150)
);

AND2x4_ASAP7_75t_L g5151 ( 
.A(n_4938),
.B(n_1389),
.Y(n_5151)
);

AND2x2_ASAP7_75t_L g5152 ( 
.A(n_4898),
.B(n_1390),
.Y(n_5152)
);

INVx2_ASAP7_75t_L g5153 ( 
.A(n_4783),
.Y(n_5153)
);

NOR2xp33_ASAP7_75t_L g5154 ( 
.A(n_4859),
.B(n_1396),
.Y(n_5154)
);

AOI21xp5_ASAP7_75t_L g5155 ( 
.A1(n_4944),
.A2(n_1401),
.B(n_1399),
.Y(n_5155)
);

NAND2x1p5_ASAP7_75t_L g5156 ( 
.A(n_4950),
.B(n_1402),
.Y(n_5156)
);

INVx2_ASAP7_75t_SL g5157 ( 
.A(n_4920),
.Y(n_5157)
);

INVx3_ASAP7_75t_SL g5158 ( 
.A(n_4923),
.Y(n_5158)
);

INVx4_ASAP7_75t_L g5159 ( 
.A(n_4903),
.Y(n_5159)
);

INVx2_ASAP7_75t_L g5160 ( 
.A(n_4956),
.Y(n_5160)
);

INVx5_ASAP7_75t_L g5161 ( 
.A(n_4885),
.Y(n_5161)
);

INVx3_ASAP7_75t_L g5162 ( 
.A(n_4846),
.Y(n_5162)
);

INVx1_ASAP7_75t_L g5163 ( 
.A(n_4848),
.Y(n_5163)
);

INVx1_ASAP7_75t_SL g5164 ( 
.A(n_4805),
.Y(n_5164)
);

AOI22xp5_ASAP7_75t_L g5165 ( 
.A1(n_4968),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_5165)
);

OA21x2_ASAP7_75t_L g5166 ( 
.A1(n_4799),
.A2(n_63),
.B(n_64),
.Y(n_5166)
);

NAND3xp33_ASAP7_75t_L g5167 ( 
.A(n_4877),
.B(n_64),
.C(n_66),
.Y(n_5167)
);

OR2x2_ASAP7_75t_L g5168 ( 
.A(n_4987),
.B(n_67),
.Y(n_5168)
);

NAND2xp5_ASAP7_75t_L g5169 ( 
.A(n_4918),
.B(n_68),
.Y(n_5169)
);

INVx2_ASAP7_75t_SL g5170 ( 
.A(n_5056),
.Y(n_5170)
);

INVx2_ASAP7_75t_L g5171 ( 
.A(n_5062),
.Y(n_5171)
);

AND2x2_ASAP7_75t_L g5172 ( 
.A(n_5039),
.B(n_5002),
.Y(n_5172)
);

INVx1_ASAP7_75t_L g5173 ( 
.A(n_5048),
.Y(n_5173)
);

BUFx12f_ASAP7_75t_L g5174 ( 
.A(n_5044),
.Y(n_5174)
);

AND2x4_ASAP7_75t_L g5175 ( 
.A(n_5026),
.B(n_4932),
.Y(n_5175)
);

NOR2x2_ASAP7_75t_L g5176 ( 
.A(n_5064),
.B(n_4778),
.Y(n_5176)
);

O2A1O1Ixp5_ASAP7_75t_L g5177 ( 
.A1(n_5112),
.A2(n_4901),
.B(n_4832),
.C(n_4927),
.Y(n_5177)
);

A2O1A1Ixp33_ASAP7_75t_L g5178 ( 
.A1(n_5025),
.A2(n_4913),
.B(n_4953),
.C(n_4952),
.Y(n_5178)
);

AOI21xp5_ASAP7_75t_SL g5179 ( 
.A1(n_5118),
.A2(n_4993),
.B(n_4926),
.Y(n_5179)
);

NAND2xp5_ASAP7_75t_L g5180 ( 
.A(n_5008),
.B(n_4876),
.Y(n_5180)
);

AND2x4_ASAP7_75t_L g5181 ( 
.A(n_5058),
.B(n_5005),
.Y(n_5181)
);

NOR2xp67_ASAP7_75t_L g5182 ( 
.A(n_5161),
.B(n_4861),
.Y(n_5182)
);

INVx1_ASAP7_75t_L g5183 ( 
.A(n_5015),
.Y(n_5183)
);

OR2x2_ASAP7_75t_L g5184 ( 
.A(n_5106),
.B(n_4862),
.Y(n_5184)
);

AOI21x1_ASAP7_75t_SL g5185 ( 
.A1(n_5149),
.A2(n_4867),
.B(n_4939),
.Y(n_5185)
);

BUFx6f_ASAP7_75t_L g5186 ( 
.A(n_5023),
.Y(n_5186)
);

NOR2xp33_ASAP7_75t_L g5187 ( 
.A(n_5012),
.B(n_5159),
.Y(n_5187)
);

AND2x2_ASAP7_75t_L g5188 ( 
.A(n_5045),
.B(n_5005),
.Y(n_5188)
);

HB1xp67_ASAP7_75t_L g5189 ( 
.A(n_5020),
.Y(n_5189)
);

AND2x2_ASAP7_75t_L g5190 ( 
.A(n_5076),
.B(n_4863),
.Y(n_5190)
);

O2A1O1Ixp5_ASAP7_75t_L g5191 ( 
.A1(n_5024),
.A2(n_4827),
.B(n_4917),
.C(n_4828),
.Y(n_5191)
);

AND2x2_ASAP7_75t_L g5192 ( 
.A(n_5016),
.B(n_4848),
.Y(n_5192)
);

INVx1_ASAP7_75t_L g5193 ( 
.A(n_5021),
.Y(n_5193)
);

HB1xp67_ASAP7_75t_L g5194 ( 
.A(n_5055),
.Y(n_5194)
);

AND2x2_ASAP7_75t_L g5195 ( 
.A(n_5067),
.B(n_4891),
.Y(n_5195)
);

AND2x4_ASAP7_75t_L g5196 ( 
.A(n_5007),
.B(n_4891),
.Y(n_5196)
);

NAND3xp33_ASAP7_75t_L g5197 ( 
.A(n_5131),
.B(n_4794),
.C(n_4782),
.Y(n_5197)
);

INVx2_ASAP7_75t_L g5198 ( 
.A(n_5068),
.Y(n_5198)
);

OA21x2_ASAP7_75t_L g5199 ( 
.A1(n_5130),
.A2(n_4819),
.B(n_4914),
.Y(n_5199)
);

AND2x2_ASAP7_75t_L g5200 ( 
.A(n_5111),
.B(n_4893),
.Y(n_5200)
);

O2A1O1Ixp33_ASAP7_75t_L g5201 ( 
.A1(n_5108),
.A2(n_4879),
.B(n_4824),
.C(n_4823),
.Y(n_5201)
);

INVx2_ASAP7_75t_L g5202 ( 
.A(n_5074),
.Y(n_5202)
);

OR2x6_ASAP7_75t_L g5203 ( 
.A(n_5064),
.B(n_5000),
.Y(n_5203)
);

CKINVDCx5p33_ASAP7_75t_R g5204 ( 
.A(n_5019),
.Y(n_5204)
);

A2O1A1Ixp33_ASAP7_75t_L g5205 ( 
.A1(n_5110),
.A2(n_4921),
.B(n_4935),
.C(n_4916),
.Y(n_5205)
);

NAND2xp5_ASAP7_75t_L g5206 ( 
.A(n_5088),
.B(n_4941),
.Y(n_5206)
);

INVx2_ASAP7_75t_L g5207 ( 
.A(n_5077),
.Y(n_5207)
);

NAND2x1p5_ASAP7_75t_L g5208 ( 
.A(n_5145),
.B(n_5161),
.Y(n_5208)
);

NOR2xp67_ASAP7_75t_L g5209 ( 
.A(n_5087),
.B(n_4865),
.Y(n_5209)
);

INVx1_ASAP7_75t_L g5210 ( 
.A(n_5065),
.Y(n_5210)
);

HB1xp67_ASAP7_75t_L g5211 ( 
.A(n_5082),
.Y(n_5211)
);

NAND2xp5_ASAP7_75t_L g5212 ( 
.A(n_5047),
.B(n_4894),
.Y(n_5212)
);

OR2x2_ASAP7_75t_L g5213 ( 
.A(n_5083),
.B(n_4893),
.Y(n_5213)
);

AND2x2_ASAP7_75t_L g5214 ( 
.A(n_5109),
.B(n_5053),
.Y(n_5214)
);

AND2x2_ASAP7_75t_L g5215 ( 
.A(n_5032),
.B(n_4922),
.Y(n_5215)
);

AND2x2_ASAP7_75t_L g5216 ( 
.A(n_5060),
.B(n_5040),
.Y(n_5216)
);

AND2x2_ASAP7_75t_L g5217 ( 
.A(n_5059),
.B(n_4922),
.Y(n_5217)
);

NOR2xp33_ASAP7_75t_SL g5218 ( 
.A(n_5051),
.B(n_4873),
.Y(n_5218)
);

OA21x2_ASAP7_75t_L g5219 ( 
.A1(n_5138),
.A2(n_4928),
.B(n_4925),
.Y(n_5219)
);

A2O1A1Ixp33_ASAP7_75t_L g5220 ( 
.A1(n_5119),
.A2(n_5167),
.B(n_5030),
.C(n_5069),
.Y(n_5220)
);

NAND2xp5_ASAP7_75t_L g5221 ( 
.A(n_5054),
.B(n_4909),
.Y(n_5221)
);

A2O1A1Ixp33_ASAP7_75t_L g5222 ( 
.A1(n_5165),
.A2(n_4840),
.B(n_4854),
.C(n_4853),
.Y(n_5222)
);

AND2x2_ASAP7_75t_SL g5223 ( 
.A(n_5147),
.B(n_4803),
.Y(n_5223)
);

AND2x2_ASAP7_75t_L g5224 ( 
.A(n_5148),
.B(n_4847),
.Y(n_5224)
);

AOI21xp5_ASAP7_75t_L g5225 ( 
.A1(n_5022),
.A2(n_4813),
.B(n_4835),
.Y(n_5225)
);

NOR2xp67_ASAP7_75t_L g5226 ( 
.A(n_5041),
.B(n_5080),
.Y(n_5226)
);

O2A1O1Ixp33_ASAP7_75t_L g5227 ( 
.A1(n_5052),
.A2(n_4889),
.B(n_4785),
.C(n_4947),
.Y(n_5227)
);

INVx2_ASAP7_75t_L g5228 ( 
.A(n_5013),
.Y(n_5228)
);

AND2x2_ASAP7_75t_L g5229 ( 
.A(n_5014),
.B(n_4868),
.Y(n_5229)
);

INVx1_ASAP7_75t_L g5230 ( 
.A(n_5027),
.Y(n_5230)
);

NAND2xp5_ASAP7_75t_L g5231 ( 
.A(n_5050),
.B(n_4838),
.Y(n_5231)
);

A2O1A1Ixp33_ASAP7_75t_L g5232 ( 
.A1(n_5136),
.A2(n_4858),
.B(n_4888),
.C(n_4886),
.Y(n_5232)
);

OR2x6_ASAP7_75t_L g5233 ( 
.A(n_5018),
.B(n_5003),
.Y(n_5233)
);

AOI21xp5_ASAP7_75t_L g5234 ( 
.A1(n_5122),
.A2(n_4899),
.B(n_4883),
.Y(n_5234)
);

OR2x6_ASAP7_75t_SL g5235 ( 
.A(n_5139),
.B(n_4934),
.Y(n_5235)
);

AND2x2_ASAP7_75t_L g5236 ( 
.A(n_5164),
.B(n_4902),
.Y(n_5236)
);

OR2x2_ASAP7_75t_L g5237 ( 
.A(n_5046),
.B(n_4843),
.Y(n_5237)
);

OAI22xp5_ASAP7_75t_SL g5238 ( 
.A1(n_5150),
.A2(n_4948),
.B1(n_4910),
.B2(n_4775),
.Y(n_5238)
);

INVx1_ASAP7_75t_L g5239 ( 
.A(n_5057),
.Y(n_5239)
);

AOI21xp5_ASAP7_75t_SL g5240 ( 
.A1(n_5018),
.A2(n_5011),
.B(n_5092),
.Y(n_5240)
);

OA21x2_ASAP7_75t_L g5241 ( 
.A1(n_5090),
.A2(n_4942),
.B(n_4795),
.Y(n_5241)
);

NAND2xp5_ASAP7_75t_L g5242 ( 
.A(n_5066),
.B(n_4904),
.Y(n_5242)
);

NAND2xp5_ASAP7_75t_L g5243 ( 
.A(n_5086),
.B(n_4814),
.Y(n_5243)
);

INVx1_ASAP7_75t_L g5244 ( 
.A(n_5163),
.Y(n_5244)
);

INVx1_ASAP7_75t_L g5245 ( 
.A(n_5142),
.Y(n_5245)
);

AND2x2_ASAP7_75t_L g5246 ( 
.A(n_5084),
.B(n_4789),
.Y(n_5246)
);

AND2x2_ASAP7_75t_L g5247 ( 
.A(n_5042),
.B(n_4959),
.Y(n_5247)
);

NAND2xp5_ASAP7_75t_L g5248 ( 
.A(n_5072),
.B(n_69),
.Y(n_5248)
);

INVx1_ASAP7_75t_L g5249 ( 
.A(n_5146),
.Y(n_5249)
);

OR2x6_ASAP7_75t_SL g5250 ( 
.A(n_5168),
.B(n_4999),
.Y(n_5250)
);

AND2x2_ASAP7_75t_L g5251 ( 
.A(n_5079),
.B(n_4986),
.Y(n_5251)
);

NAND2xp5_ASAP7_75t_L g5252 ( 
.A(n_5107),
.B(n_71),
.Y(n_5252)
);

OA21x2_ASAP7_75t_L g5253 ( 
.A1(n_5093),
.A2(n_4780),
.B(n_71),
.Y(n_5253)
);

AND2x2_ASAP7_75t_L g5254 ( 
.A(n_5140),
.B(n_72),
.Y(n_5254)
);

INVx2_ASAP7_75t_L g5255 ( 
.A(n_5099),
.Y(n_5255)
);

NAND2xp5_ASAP7_75t_L g5256 ( 
.A(n_5097),
.B(n_5121),
.Y(n_5256)
);

OR2x2_ASAP7_75t_L g5257 ( 
.A(n_5105),
.B(n_72),
.Y(n_5257)
);

A2O1A1Ixp33_ASAP7_75t_L g5258 ( 
.A1(n_5010),
.A2(n_75),
.B(n_73),
.C(n_74),
.Y(n_5258)
);

BUFx2_ASAP7_75t_L g5259 ( 
.A(n_5071),
.Y(n_5259)
);

INVxp67_ASAP7_75t_SL g5260 ( 
.A(n_5101),
.Y(n_5260)
);

AND2x2_ASAP7_75t_L g5261 ( 
.A(n_5028),
.B(n_73),
.Y(n_5261)
);

INVx2_ASAP7_75t_L g5262 ( 
.A(n_5103),
.Y(n_5262)
);

A2O1A1Ixp33_ASAP7_75t_L g5263 ( 
.A1(n_5135),
.A2(n_78),
.B(n_75),
.C(n_77),
.Y(n_5263)
);

INVx1_ASAP7_75t_L g5264 ( 
.A(n_5115),
.Y(n_5264)
);

INVx1_ASAP7_75t_L g5265 ( 
.A(n_5129),
.Y(n_5265)
);

O2A1O1Ixp33_ASAP7_75t_L g5266 ( 
.A1(n_5124),
.A2(n_81),
.B(n_77),
.C(n_80),
.Y(n_5266)
);

INVx1_ASAP7_75t_L g5267 ( 
.A(n_5153),
.Y(n_5267)
);

O2A1O1Ixp5_ASAP7_75t_L g5268 ( 
.A1(n_5137),
.A2(n_83),
.B(n_81),
.C(n_82),
.Y(n_5268)
);

INVx3_ASAP7_75t_L g5269 ( 
.A(n_5056),
.Y(n_5269)
);

OAI22xp5_ASAP7_75t_L g5270 ( 
.A1(n_5158),
.A2(n_89),
.B1(n_84),
.B2(n_85),
.Y(n_5270)
);

OR2x2_ASAP7_75t_L g5271 ( 
.A(n_5100),
.B(n_84),
.Y(n_5271)
);

AND2x2_ASAP7_75t_L g5272 ( 
.A(n_5028),
.B(n_5063),
.Y(n_5272)
);

INVx1_ASAP7_75t_L g5273 ( 
.A(n_5095),
.Y(n_5273)
);

INVx1_ASAP7_75t_L g5274 ( 
.A(n_5160),
.Y(n_5274)
);

NAND2xp5_ASAP7_75t_L g5275 ( 
.A(n_5141),
.B(n_90),
.Y(n_5275)
);

NAND2xp5_ASAP7_75t_L g5276 ( 
.A(n_5123),
.B(n_91),
.Y(n_5276)
);

OAI22xp5_ASAP7_75t_L g5277 ( 
.A1(n_5085),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.Y(n_5277)
);

INVx1_ASAP7_75t_L g5278 ( 
.A(n_5166),
.Y(n_5278)
);

INVxp67_ASAP7_75t_L g5279 ( 
.A(n_5120),
.Y(n_5279)
);

AND2x2_ASAP7_75t_L g5280 ( 
.A(n_5036),
.B(n_94),
.Y(n_5280)
);

OR2x2_ASAP7_75t_L g5281 ( 
.A(n_5169),
.B(n_95),
.Y(n_5281)
);

O2A1O1Ixp33_ASAP7_75t_L g5282 ( 
.A1(n_5114),
.A2(n_98),
.B(n_96),
.C(n_97),
.Y(n_5282)
);

BUFx10_ASAP7_75t_L g5283 ( 
.A(n_5035),
.Y(n_5283)
);

A2O1A1Ixp33_ASAP7_75t_SL g5284 ( 
.A1(n_5009),
.A2(n_101),
.B(n_96),
.C(n_100),
.Y(n_5284)
);

NOR2xp33_ASAP7_75t_R g5285 ( 
.A(n_5089),
.B(n_1404),
.Y(n_5285)
);

NAND2xp5_ASAP7_75t_L g5286 ( 
.A(n_5128),
.B(n_100),
.Y(n_5286)
);

NOR2xp33_ASAP7_75t_L g5287 ( 
.A(n_5049),
.B(n_102),
.Y(n_5287)
);

HB1xp67_ASAP7_75t_L g5288 ( 
.A(n_5162),
.Y(n_5288)
);

OR2x2_ASAP7_75t_L g5289 ( 
.A(n_5034),
.B(n_103),
.Y(n_5289)
);

NAND2xp5_ASAP7_75t_L g5290 ( 
.A(n_5157),
.B(n_104),
.Y(n_5290)
);

INVx3_ASAP7_75t_SL g5291 ( 
.A(n_5017),
.Y(n_5291)
);

INVx2_ASAP7_75t_L g5292 ( 
.A(n_5134),
.Y(n_5292)
);

INVx1_ASAP7_75t_L g5293 ( 
.A(n_5127),
.Y(n_5293)
);

OR2x2_ASAP7_75t_L g5294 ( 
.A(n_5075),
.B(n_104),
.Y(n_5294)
);

INVx1_ASAP7_75t_L g5295 ( 
.A(n_5125),
.Y(n_5295)
);

NAND2xp5_ASAP7_75t_L g5296 ( 
.A(n_5145),
.B(n_106),
.Y(n_5296)
);

INVx3_ASAP7_75t_L g5297 ( 
.A(n_5094),
.Y(n_5297)
);

AOI21xp5_ASAP7_75t_L g5298 ( 
.A1(n_5155),
.A2(n_1408),
.B(n_1407),
.Y(n_5298)
);

AND2x4_ASAP7_75t_L g5299 ( 
.A(n_5078),
.B(n_1409),
.Y(n_5299)
);

BUFx6f_ASAP7_75t_L g5300 ( 
.A(n_5023),
.Y(n_5300)
);

INVx1_ASAP7_75t_L g5301 ( 
.A(n_5029),
.Y(n_5301)
);

AND2x2_ASAP7_75t_L g5302 ( 
.A(n_5152),
.B(n_5098),
.Y(n_5302)
);

OA21x2_ASAP7_75t_L g5303 ( 
.A1(n_5104),
.A2(n_106),
.B(n_107),
.Y(n_5303)
);

OA22x2_ASAP7_75t_L g5304 ( 
.A1(n_5126),
.A2(n_111),
.B1(n_108),
.B2(n_109),
.Y(n_5304)
);

INVx1_ASAP7_75t_L g5305 ( 
.A(n_5031),
.Y(n_5305)
);

AOI21xp5_ASAP7_75t_SL g5306 ( 
.A1(n_5070),
.A2(n_1414),
.B(n_1410),
.Y(n_5306)
);

NAND4xp25_ASAP7_75t_L g5307 ( 
.A(n_5081),
.B(n_113),
.C(n_108),
.D(n_112),
.Y(n_5307)
);

OAI22xp5_ASAP7_75t_SL g5308 ( 
.A1(n_5102),
.A2(n_114),
.B1(n_112),
.B2(n_113),
.Y(n_5308)
);

CKINVDCx16_ASAP7_75t_R g5309 ( 
.A(n_5117),
.Y(n_5309)
);

NAND2xp5_ASAP7_75t_L g5310 ( 
.A(n_5143),
.B(n_114),
.Y(n_5310)
);

A2O1A1Ixp33_ASAP7_75t_L g5311 ( 
.A1(n_5154),
.A2(n_5043),
.B(n_5151),
.C(n_5037),
.Y(n_5311)
);

OAI22xp5_ASAP7_75t_L g5312 ( 
.A1(n_5038),
.A2(n_5133),
.B1(n_5006),
.B2(n_5017),
.Y(n_5312)
);

NOR2x2_ASAP7_75t_L g5313 ( 
.A(n_5132),
.B(n_115),
.Y(n_5313)
);

AOI21xp5_ASAP7_75t_L g5314 ( 
.A1(n_5156),
.A2(n_1418),
.B(n_1416),
.Y(n_5314)
);

NAND2xp5_ASAP7_75t_L g5315 ( 
.A(n_5144),
.B(n_116),
.Y(n_5315)
);

NAND2x1p5_ASAP7_75t_L g5316 ( 
.A(n_5144),
.B(n_1427),
.Y(n_5316)
);

INVx2_ASAP7_75t_L g5317 ( 
.A(n_5094),
.Y(n_5317)
);

BUFx4f_ASAP7_75t_SL g5318 ( 
.A(n_5174),
.Y(n_5318)
);

AND2x2_ASAP7_75t_L g5319 ( 
.A(n_5214),
.B(n_5073),
.Y(n_5319)
);

HB1xp67_ASAP7_75t_L g5320 ( 
.A(n_5194),
.Y(n_5320)
);

INVx2_ASAP7_75t_L g5321 ( 
.A(n_5173),
.Y(n_5321)
);

INVx1_ASAP7_75t_L g5322 ( 
.A(n_5211),
.Y(n_5322)
);

INVx2_ASAP7_75t_L g5323 ( 
.A(n_5171),
.Y(n_5323)
);

INVx2_ASAP7_75t_L g5324 ( 
.A(n_5198),
.Y(n_5324)
);

AND2x4_ASAP7_75t_L g5325 ( 
.A(n_5183),
.B(n_5091),
.Y(n_5325)
);

CKINVDCx5p33_ASAP7_75t_R g5326 ( 
.A(n_5204),
.Y(n_5326)
);

INVxp67_ASAP7_75t_L g5327 ( 
.A(n_5209),
.Y(n_5327)
);

INVx3_ASAP7_75t_L g5328 ( 
.A(n_5208),
.Y(n_5328)
);

INVx1_ASAP7_75t_L g5329 ( 
.A(n_5210),
.Y(n_5329)
);

NAND2xp5_ASAP7_75t_L g5330 ( 
.A(n_5200),
.B(n_5033),
.Y(n_5330)
);

INVx1_ASAP7_75t_L g5331 ( 
.A(n_5230),
.Y(n_5331)
);

NAND2xp5_ASAP7_75t_L g5332 ( 
.A(n_5202),
.B(n_5113),
.Y(n_5332)
);

HB1xp67_ASAP7_75t_L g5333 ( 
.A(n_5189),
.Y(n_5333)
);

CKINVDCx6p67_ASAP7_75t_R g5334 ( 
.A(n_5291),
.Y(n_5334)
);

AND2x2_ASAP7_75t_L g5335 ( 
.A(n_5272),
.B(n_5061),
.Y(n_5335)
);

INVx3_ASAP7_75t_L g5336 ( 
.A(n_5283),
.Y(n_5336)
);

NAND2x1p5_ASAP7_75t_L g5337 ( 
.A(n_5182),
.B(n_5236),
.Y(n_5337)
);

INVx1_ASAP7_75t_L g5338 ( 
.A(n_5244),
.Y(n_5338)
);

INVx1_ASAP7_75t_L g5339 ( 
.A(n_5245),
.Y(n_5339)
);

INVx1_ASAP7_75t_L g5340 ( 
.A(n_5249),
.Y(n_5340)
);

BUFx3_ASAP7_75t_L g5341 ( 
.A(n_5186),
.Y(n_5341)
);

BUFx6f_ASAP7_75t_L g5342 ( 
.A(n_5186),
.Y(n_5342)
);

INVx1_ASAP7_75t_L g5343 ( 
.A(n_5193),
.Y(n_5343)
);

AND2x2_ASAP7_75t_L g5344 ( 
.A(n_5216),
.B(n_5113),
.Y(n_5344)
);

INVx1_ASAP7_75t_L g5345 ( 
.A(n_5207),
.Y(n_5345)
);

HB1xp67_ASAP7_75t_L g5346 ( 
.A(n_5181),
.Y(n_5346)
);

INVx2_ASAP7_75t_L g5347 ( 
.A(n_5228),
.Y(n_5347)
);

INVx1_ASAP7_75t_L g5348 ( 
.A(n_5213),
.Y(n_5348)
);

AO21x2_ASAP7_75t_L g5349 ( 
.A1(n_5278),
.A2(n_5096),
.B(n_5116),
.Y(n_5349)
);

INVx1_ASAP7_75t_L g5350 ( 
.A(n_5239),
.Y(n_5350)
);

OAI21x1_ASAP7_75t_L g5351 ( 
.A1(n_5225),
.A2(n_1430),
.B(n_1428),
.Y(n_5351)
);

OAI21x1_ASAP7_75t_L g5352 ( 
.A1(n_5234),
.A2(n_1433),
.B(n_1432),
.Y(n_5352)
);

INVx1_ASAP7_75t_L g5353 ( 
.A(n_5267),
.Y(n_5353)
);

INVx1_ASAP7_75t_L g5354 ( 
.A(n_5273),
.Y(n_5354)
);

INVx1_ASAP7_75t_L g5355 ( 
.A(n_5274),
.Y(n_5355)
);

BUFx3_ASAP7_75t_L g5356 ( 
.A(n_5300),
.Y(n_5356)
);

OR2x2_ASAP7_75t_L g5357 ( 
.A(n_5260),
.B(n_116),
.Y(n_5357)
);

OR2x2_ASAP7_75t_L g5358 ( 
.A(n_5184),
.B(n_117),
.Y(n_5358)
);

OR2x2_ASAP7_75t_L g5359 ( 
.A(n_5288),
.B(n_118),
.Y(n_5359)
);

INVx1_ASAP7_75t_L g5360 ( 
.A(n_5264),
.Y(n_5360)
);

INVx1_ASAP7_75t_L g5361 ( 
.A(n_5265),
.Y(n_5361)
);

INVx1_ASAP7_75t_L g5362 ( 
.A(n_5255),
.Y(n_5362)
);

INVx1_ASAP7_75t_L g5363 ( 
.A(n_5262),
.Y(n_5363)
);

INVx2_ASAP7_75t_L g5364 ( 
.A(n_5215),
.Y(n_5364)
);

HB1xp67_ASAP7_75t_L g5365 ( 
.A(n_5192),
.Y(n_5365)
);

INVx2_ASAP7_75t_SL g5366 ( 
.A(n_5292),
.Y(n_5366)
);

HB1xp67_ASAP7_75t_L g5367 ( 
.A(n_5188),
.Y(n_5367)
);

BUFx2_ASAP7_75t_L g5368 ( 
.A(n_5196),
.Y(n_5368)
);

INVx2_ASAP7_75t_L g5369 ( 
.A(n_5301),
.Y(n_5369)
);

AND2x2_ASAP7_75t_L g5370 ( 
.A(n_5172),
.B(n_119),
.Y(n_5370)
);

AO21x2_ASAP7_75t_L g5371 ( 
.A1(n_5295),
.A2(n_119),
.B(n_120),
.Y(n_5371)
);

BUFx3_ASAP7_75t_L g5372 ( 
.A(n_5300),
.Y(n_5372)
);

INVx1_ASAP7_75t_L g5373 ( 
.A(n_5237),
.Y(n_5373)
);

AOI22xp33_ASAP7_75t_SL g5374 ( 
.A1(n_5223),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.Y(n_5374)
);

AOI21x1_ASAP7_75t_L g5375 ( 
.A1(n_5226),
.A2(n_122),
.B(n_123),
.Y(n_5375)
);

INVx2_ASAP7_75t_L g5376 ( 
.A(n_5305),
.Y(n_5376)
);

BUFx2_ASAP7_75t_L g5377 ( 
.A(n_5175),
.Y(n_5377)
);

OR2x2_ASAP7_75t_L g5378 ( 
.A(n_5212),
.B(n_124),
.Y(n_5378)
);

INVx1_ASAP7_75t_L g5379 ( 
.A(n_5257),
.Y(n_5379)
);

OAI21x1_ASAP7_75t_L g5380 ( 
.A1(n_5191),
.A2(n_1438),
.B(n_1437),
.Y(n_5380)
);

AND2x4_ASAP7_75t_L g5381 ( 
.A(n_5224),
.B(n_1440),
.Y(n_5381)
);

INVx1_ASAP7_75t_L g5382 ( 
.A(n_5195),
.Y(n_5382)
);

INVx2_ASAP7_75t_SL g5383 ( 
.A(n_5317),
.Y(n_5383)
);

NAND2xp5_ASAP7_75t_L g5384 ( 
.A(n_5206),
.B(n_124),
.Y(n_5384)
);

HB1xp67_ASAP7_75t_L g5385 ( 
.A(n_5217),
.Y(n_5385)
);

INVx1_ASAP7_75t_L g5386 ( 
.A(n_5229),
.Y(n_5386)
);

AND2x2_ASAP7_75t_L g5387 ( 
.A(n_5187),
.B(n_126),
.Y(n_5387)
);

NOR2xp33_ASAP7_75t_L g5388 ( 
.A(n_5256),
.B(n_126),
.Y(n_5388)
);

INVx1_ASAP7_75t_L g5389 ( 
.A(n_5293),
.Y(n_5389)
);

INVx1_ASAP7_75t_L g5390 ( 
.A(n_5243),
.Y(n_5390)
);

NAND2xp5_ASAP7_75t_L g5391 ( 
.A(n_5247),
.B(n_127),
.Y(n_5391)
);

INVx1_ASAP7_75t_L g5392 ( 
.A(n_5242),
.Y(n_5392)
);

INVx4_ASAP7_75t_L g5393 ( 
.A(n_5269),
.Y(n_5393)
);

INVx3_ASAP7_75t_L g5394 ( 
.A(n_5297),
.Y(n_5394)
);

INVx1_ASAP7_75t_L g5395 ( 
.A(n_5261),
.Y(n_5395)
);

INVx2_ASAP7_75t_SL g5396 ( 
.A(n_5170),
.Y(n_5396)
);

INVx2_ASAP7_75t_L g5397 ( 
.A(n_5251),
.Y(n_5397)
);

INVx1_ASAP7_75t_L g5398 ( 
.A(n_5246),
.Y(n_5398)
);

INVx1_ASAP7_75t_L g5399 ( 
.A(n_5252),
.Y(n_5399)
);

INVx2_ASAP7_75t_L g5400 ( 
.A(n_5219),
.Y(n_5400)
);

INVx1_ASAP7_75t_L g5401 ( 
.A(n_5199),
.Y(n_5401)
);

INVx1_ASAP7_75t_L g5402 ( 
.A(n_5253),
.Y(n_5402)
);

INVx2_ASAP7_75t_L g5403 ( 
.A(n_5294),
.Y(n_5403)
);

BUFx2_ASAP7_75t_L g5404 ( 
.A(n_5176),
.Y(n_5404)
);

INVx1_ASAP7_75t_L g5405 ( 
.A(n_5190),
.Y(n_5405)
);

AOI21xp5_ASAP7_75t_L g5406 ( 
.A1(n_5178),
.A2(n_5222),
.B(n_5179),
.Y(n_5406)
);

INVx2_ASAP7_75t_L g5407 ( 
.A(n_5279),
.Y(n_5407)
);

INVx1_ASAP7_75t_L g5408 ( 
.A(n_5248),
.Y(n_5408)
);

INVx2_ASAP7_75t_L g5409 ( 
.A(n_5241),
.Y(n_5409)
);

HB1xp67_ASAP7_75t_L g5410 ( 
.A(n_5203),
.Y(n_5410)
);

INVx1_ASAP7_75t_L g5411 ( 
.A(n_5303),
.Y(n_5411)
);

INVx1_ASAP7_75t_L g5412 ( 
.A(n_5250),
.Y(n_5412)
);

OAI21xp5_ASAP7_75t_L g5413 ( 
.A1(n_5220),
.A2(n_128),
.B(n_129),
.Y(n_5413)
);

OAI21x1_ASAP7_75t_L g5414 ( 
.A1(n_5177),
.A2(n_1444),
.B(n_1443),
.Y(n_5414)
);

INVx1_ASAP7_75t_L g5415 ( 
.A(n_5296),
.Y(n_5415)
);

INVx1_ASAP7_75t_L g5416 ( 
.A(n_5290),
.Y(n_5416)
);

INVx2_ASAP7_75t_L g5417 ( 
.A(n_5203),
.Y(n_5417)
);

INVx1_ASAP7_75t_L g5418 ( 
.A(n_5231),
.Y(n_5418)
);

INVx1_ASAP7_75t_L g5419 ( 
.A(n_5233),
.Y(n_5419)
);

BUFx4f_ASAP7_75t_L g5420 ( 
.A(n_5299),
.Y(n_5420)
);

CKINVDCx6p67_ASAP7_75t_R g5421 ( 
.A(n_5309),
.Y(n_5421)
);

BUFx2_ASAP7_75t_L g5422 ( 
.A(n_5259),
.Y(n_5422)
);

INVx1_ASAP7_75t_L g5423 ( 
.A(n_5233),
.Y(n_5423)
);

AND2x2_ASAP7_75t_L g5424 ( 
.A(n_5302),
.B(n_5180),
.Y(n_5424)
);

AND2x4_ASAP7_75t_L g5425 ( 
.A(n_5311),
.B(n_1445),
.Y(n_5425)
);

INVx2_ASAP7_75t_L g5426 ( 
.A(n_5289),
.Y(n_5426)
);

HB1xp67_ASAP7_75t_L g5427 ( 
.A(n_5221),
.Y(n_5427)
);

AOI22xp33_ASAP7_75t_L g5428 ( 
.A1(n_5197),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_5428)
);

NOR2xp33_ASAP7_75t_L g5429 ( 
.A(n_5235),
.B(n_130),
.Y(n_5429)
);

INVx1_ASAP7_75t_L g5430 ( 
.A(n_5268),
.Y(n_5430)
);

INVx1_ASAP7_75t_L g5431 ( 
.A(n_5271),
.Y(n_5431)
);

INVx1_ASAP7_75t_L g5432 ( 
.A(n_5281),
.Y(n_5432)
);

BUFx2_ASAP7_75t_L g5433 ( 
.A(n_5312),
.Y(n_5433)
);

OAI21x1_ASAP7_75t_L g5434 ( 
.A1(n_5185),
.A2(n_1448),
.B(n_1446),
.Y(n_5434)
);

INVx2_ASAP7_75t_L g5435 ( 
.A(n_5315),
.Y(n_5435)
);

INVx2_ASAP7_75t_L g5436 ( 
.A(n_5276),
.Y(n_5436)
);

AND2x2_ASAP7_75t_L g5437 ( 
.A(n_5280),
.B(n_131),
.Y(n_5437)
);

INVx1_ASAP7_75t_L g5438 ( 
.A(n_5275),
.Y(n_5438)
);

INVx1_ASAP7_75t_L g5439 ( 
.A(n_5238),
.Y(n_5439)
);

INVx1_ASAP7_75t_L g5440 ( 
.A(n_5282),
.Y(n_5440)
);

AND2x4_ASAP7_75t_L g5441 ( 
.A(n_5287),
.B(n_5254),
.Y(n_5441)
);

NAND2x1p5_ASAP7_75t_L g5442 ( 
.A(n_5314),
.B(n_5298),
.Y(n_5442)
);

HB1xp67_ASAP7_75t_L g5443 ( 
.A(n_5304),
.Y(n_5443)
);

HB1xp67_ASAP7_75t_L g5444 ( 
.A(n_5277),
.Y(n_5444)
);

INVx3_ASAP7_75t_L g5445 ( 
.A(n_5316),
.Y(n_5445)
);

INVx2_ASAP7_75t_L g5446 ( 
.A(n_5313),
.Y(n_5446)
);

INVx1_ASAP7_75t_L g5447 ( 
.A(n_5263),
.Y(n_5447)
);

AND2x2_ASAP7_75t_L g5448 ( 
.A(n_5285),
.B(n_132),
.Y(n_5448)
);

AND2x2_ASAP7_75t_L g5449 ( 
.A(n_5310),
.B(n_133),
.Y(n_5449)
);

O2A1O1Ixp33_ASAP7_75t_L g5450 ( 
.A1(n_5258),
.A2(n_5284),
.B(n_5266),
.C(n_5227),
.Y(n_5450)
);

AND2x4_ASAP7_75t_L g5451 ( 
.A(n_5232),
.B(n_1453),
.Y(n_5451)
);

HB1xp67_ASAP7_75t_L g5452 ( 
.A(n_5307),
.Y(n_5452)
);

INVx1_ASAP7_75t_L g5453 ( 
.A(n_5286),
.Y(n_5453)
);

NOR2x1_ASAP7_75t_R g5454 ( 
.A(n_5218),
.B(n_133),
.Y(n_5454)
);

BUFx4_ASAP7_75t_SL g5455 ( 
.A(n_5240),
.Y(n_5455)
);

OAI21x1_ASAP7_75t_L g5456 ( 
.A1(n_5201),
.A2(n_1459),
.B(n_1454),
.Y(n_5456)
);

OR2x2_ASAP7_75t_L g5457 ( 
.A(n_5205),
.B(n_134),
.Y(n_5457)
);

INVx2_ASAP7_75t_SL g5458 ( 
.A(n_5270),
.Y(n_5458)
);

INVx1_ASAP7_75t_L g5459 ( 
.A(n_5308),
.Y(n_5459)
);

INVx1_ASAP7_75t_L g5460 ( 
.A(n_5306),
.Y(n_5460)
);

HB1xp67_ASAP7_75t_L g5461 ( 
.A(n_5194),
.Y(n_5461)
);

BUFx3_ASAP7_75t_L g5462 ( 
.A(n_5186),
.Y(n_5462)
);

INVx2_ASAP7_75t_L g5463 ( 
.A(n_5173),
.Y(n_5463)
);

INVx1_ASAP7_75t_L g5464 ( 
.A(n_5211),
.Y(n_5464)
);

OAI21xp5_ASAP7_75t_L g5465 ( 
.A1(n_5220),
.A2(n_134),
.B(n_135),
.Y(n_5465)
);

INVx1_ASAP7_75t_L g5466 ( 
.A(n_5211),
.Y(n_5466)
);

INVx2_ASAP7_75t_L g5467 ( 
.A(n_5173),
.Y(n_5467)
);

BUFx2_ASAP7_75t_L g5468 ( 
.A(n_5208),
.Y(n_5468)
);

BUFx2_ASAP7_75t_L g5469 ( 
.A(n_5208),
.Y(n_5469)
);

INVx2_ASAP7_75t_L g5470 ( 
.A(n_5173),
.Y(n_5470)
);

INVx1_ASAP7_75t_L g5471 ( 
.A(n_5211),
.Y(n_5471)
);

AND2x2_ASAP7_75t_L g5472 ( 
.A(n_5214),
.B(n_137),
.Y(n_5472)
);

OAI21x1_ASAP7_75t_L g5473 ( 
.A1(n_5225),
.A2(n_1461),
.B(n_1460),
.Y(n_5473)
);

INVx1_ASAP7_75t_L g5474 ( 
.A(n_5211),
.Y(n_5474)
);

OR2x2_ASAP7_75t_L g5475 ( 
.A(n_5194),
.B(n_138),
.Y(n_5475)
);

INVx2_ASAP7_75t_L g5476 ( 
.A(n_5173),
.Y(n_5476)
);

AND2x4_ASAP7_75t_L g5477 ( 
.A(n_5214),
.B(n_1462),
.Y(n_5477)
);

BUFx3_ASAP7_75t_L g5478 ( 
.A(n_5186),
.Y(n_5478)
);

AND2x2_ASAP7_75t_L g5479 ( 
.A(n_5214),
.B(n_138),
.Y(n_5479)
);

INVx1_ASAP7_75t_L g5480 ( 
.A(n_5211),
.Y(n_5480)
);

AOI22xp33_ASAP7_75t_L g5481 ( 
.A1(n_5406),
.A2(n_141),
.B1(n_139),
.B2(n_140),
.Y(n_5481)
);

INVx2_ASAP7_75t_L g5482 ( 
.A(n_5389),
.Y(n_5482)
);

INVx2_ASAP7_75t_L g5483 ( 
.A(n_5321),
.Y(n_5483)
);

INVx2_ASAP7_75t_L g5484 ( 
.A(n_5463),
.Y(n_5484)
);

INVx2_ASAP7_75t_L g5485 ( 
.A(n_5467),
.Y(n_5485)
);

HB1xp67_ASAP7_75t_L g5486 ( 
.A(n_5320),
.Y(n_5486)
);

INVx2_ASAP7_75t_L g5487 ( 
.A(n_5470),
.Y(n_5487)
);

AND2x2_ASAP7_75t_L g5488 ( 
.A(n_5367),
.B(n_139),
.Y(n_5488)
);

AO21x2_ASAP7_75t_L g5489 ( 
.A1(n_5401),
.A2(n_141),
.B(n_142),
.Y(n_5489)
);

AOI22xp33_ASAP7_75t_L g5490 ( 
.A1(n_5413),
.A2(n_145),
.B1(n_143),
.B2(n_144),
.Y(n_5490)
);

HB1xp67_ASAP7_75t_L g5491 ( 
.A(n_5461),
.Y(n_5491)
);

AOI22xp33_ASAP7_75t_SL g5492 ( 
.A1(n_5465),
.A2(n_145),
.B1(n_146),
.B2(n_144),
.Y(n_5492)
);

INVx1_ASAP7_75t_L g5493 ( 
.A(n_5329),
.Y(n_5493)
);

AND2x2_ASAP7_75t_L g5494 ( 
.A(n_5335),
.B(n_143),
.Y(n_5494)
);

INVx3_ASAP7_75t_L g5495 ( 
.A(n_5393),
.Y(n_5495)
);

AND2x2_ASAP7_75t_L g5496 ( 
.A(n_5377),
.B(n_147),
.Y(n_5496)
);

INVx2_ASAP7_75t_L g5497 ( 
.A(n_5476),
.Y(n_5497)
);

INVx4_ASAP7_75t_L g5498 ( 
.A(n_5326),
.Y(n_5498)
);

INVx2_ASAP7_75t_L g5499 ( 
.A(n_5369),
.Y(n_5499)
);

HB1xp67_ASAP7_75t_L g5500 ( 
.A(n_5333),
.Y(n_5500)
);

INVx1_ASAP7_75t_L g5501 ( 
.A(n_5331),
.Y(n_5501)
);

INVx1_ASAP7_75t_L g5502 ( 
.A(n_5338),
.Y(n_5502)
);

AO31x2_ASAP7_75t_L g5503 ( 
.A1(n_5402),
.A2(n_151),
.A3(n_148),
.B(n_149),
.Y(n_5503)
);

INVx2_ASAP7_75t_L g5504 ( 
.A(n_5376),
.Y(n_5504)
);

AND2x2_ASAP7_75t_L g5505 ( 
.A(n_5365),
.B(n_148),
.Y(n_5505)
);

INVx4_ASAP7_75t_L g5506 ( 
.A(n_5334),
.Y(n_5506)
);

INVx1_ASAP7_75t_L g5507 ( 
.A(n_5339),
.Y(n_5507)
);

INVx1_ASAP7_75t_L g5508 ( 
.A(n_5340),
.Y(n_5508)
);

AOI22xp5_ASAP7_75t_L g5509 ( 
.A1(n_5460),
.A2(n_156),
.B1(n_152),
.B2(n_155),
.Y(n_5509)
);

INVx2_ASAP7_75t_L g5510 ( 
.A(n_5322),
.Y(n_5510)
);

INVx2_ASAP7_75t_L g5511 ( 
.A(n_5464),
.Y(n_5511)
);

BUFx6f_ASAP7_75t_L g5512 ( 
.A(n_5342),
.Y(n_5512)
);

AND2x2_ASAP7_75t_L g5513 ( 
.A(n_5405),
.B(n_152),
.Y(n_5513)
);

INVx1_ASAP7_75t_L g5514 ( 
.A(n_5343),
.Y(n_5514)
);

NAND2xp5_ASAP7_75t_L g5515 ( 
.A(n_5418),
.B(n_156),
.Y(n_5515)
);

INVx3_ASAP7_75t_L g5516 ( 
.A(n_5336),
.Y(n_5516)
);

AND2x2_ASAP7_75t_L g5517 ( 
.A(n_5368),
.B(n_157),
.Y(n_5517)
);

HB1xp67_ASAP7_75t_L g5518 ( 
.A(n_5348),
.Y(n_5518)
);

AOI22xp33_ASAP7_75t_L g5519 ( 
.A1(n_5439),
.A2(n_159),
.B1(n_157),
.B2(n_158),
.Y(n_5519)
);

BUFx2_ASAP7_75t_L g5520 ( 
.A(n_5337),
.Y(n_5520)
);

INVx2_ASAP7_75t_L g5521 ( 
.A(n_5466),
.Y(n_5521)
);

HB1xp67_ASAP7_75t_L g5522 ( 
.A(n_5373),
.Y(n_5522)
);

BUFx2_ASAP7_75t_R g5523 ( 
.A(n_5404),
.Y(n_5523)
);

NAND2xp5_ASAP7_75t_L g5524 ( 
.A(n_5427),
.B(n_159),
.Y(n_5524)
);

NAND2xp5_ASAP7_75t_L g5525 ( 
.A(n_5390),
.B(n_160),
.Y(n_5525)
);

INVx1_ASAP7_75t_L g5526 ( 
.A(n_5471),
.Y(n_5526)
);

INVx2_ASAP7_75t_L g5527 ( 
.A(n_5474),
.Y(n_5527)
);

HB1xp67_ASAP7_75t_L g5528 ( 
.A(n_5386),
.Y(n_5528)
);

AND2x2_ASAP7_75t_L g5529 ( 
.A(n_5382),
.B(n_160),
.Y(n_5529)
);

BUFx2_ASAP7_75t_L g5530 ( 
.A(n_5468),
.Y(n_5530)
);

AND2x4_ASAP7_75t_L g5531 ( 
.A(n_5469),
.B(n_161),
.Y(n_5531)
);

INVx1_ASAP7_75t_L g5532 ( 
.A(n_5480),
.Y(n_5532)
);

INVx2_ASAP7_75t_L g5533 ( 
.A(n_5323),
.Y(n_5533)
);

AND2x4_ASAP7_75t_L g5534 ( 
.A(n_5417),
.B(n_161),
.Y(n_5534)
);

AND2x2_ASAP7_75t_L g5535 ( 
.A(n_5385),
.B(n_163),
.Y(n_5535)
);

BUFx2_ASAP7_75t_L g5536 ( 
.A(n_5346),
.Y(n_5536)
);

BUFx2_ASAP7_75t_L g5537 ( 
.A(n_5328),
.Y(n_5537)
);

AND2x2_ASAP7_75t_L g5538 ( 
.A(n_5395),
.B(n_163),
.Y(n_5538)
);

BUFx2_ASAP7_75t_L g5539 ( 
.A(n_5419),
.Y(n_5539)
);

INVx3_ASAP7_75t_L g5540 ( 
.A(n_5341),
.Y(n_5540)
);

BUFx3_ASAP7_75t_L g5541 ( 
.A(n_5422),
.Y(n_5541)
);

BUFx6f_ASAP7_75t_L g5542 ( 
.A(n_5342),
.Y(n_5542)
);

AND2x2_ASAP7_75t_L g5543 ( 
.A(n_5364),
.B(n_164),
.Y(n_5543)
);

BUFx6f_ASAP7_75t_L g5544 ( 
.A(n_5356),
.Y(n_5544)
);

INVxp67_ASAP7_75t_L g5545 ( 
.A(n_5399),
.Y(n_5545)
);

BUFx2_ASAP7_75t_L g5546 ( 
.A(n_5423),
.Y(n_5546)
);

AND2x4_ASAP7_75t_L g5547 ( 
.A(n_5407),
.B(n_165),
.Y(n_5547)
);

INVx2_ASAP7_75t_L g5548 ( 
.A(n_5324),
.Y(n_5548)
);

NAND2xp5_ASAP7_75t_L g5549 ( 
.A(n_5392),
.B(n_5379),
.Y(n_5549)
);

INVx2_ASAP7_75t_L g5550 ( 
.A(n_5347),
.Y(n_5550)
);

OR2x2_ASAP7_75t_L g5551 ( 
.A(n_5397),
.B(n_165),
.Y(n_5551)
);

INVx5_ASAP7_75t_L g5552 ( 
.A(n_5425),
.Y(n_5552)
);

INVx2_ASAP7_75t_L g5553 ( 
.A(n_5345),
.Y(n_5553)
);

OR2x2_ASAP7_75t_L g5554 ( 
.A(n_5398),
.B(n_166),
.Y(n_5554)
);

AND2x2_ASAP7_75t_L g5555 ( 
.A(n_5412),
.B(n_166),
.Y(n_5555)
);

NAND2xp5_ASAP7_75t_L g5556 ( 
.A(n_5403),
.B(n_167),
.Y(n_5556)
);

INVx1_ASAP7_75t_L g5557 ( 
.A(n_5350),
.Y(n_5557)
);

BUFx3_ASAP7_75t_L g5558 ( 
.A(n_5421),
.Y(n_5558)
);

INVx1_ASAP7_75t_L g5559 ( 
.A(n_5353),
.Y(n_5559)
);

INVx1_ASAP7_75t_L g5560 ( 
.A(n_5354),
.Y(n_5560)
);

INVx1_ASAP7_75t_L g5561 ( 
.A(n_5355),
.Y(n_5561)
);

AND2x2_ASAP7_75t_L g5562 ( 
.A(n_5424),
.B(n_168),
.Y(n_5562)
);

INVx3_ASAP7_75t_L g5563 ( 
.A(n_5372),
.Y(n_5563)
);

HB1xp67_ASAP7_75t_L g5564 ( 
.A(n_5411),
.Y(n_5564)
);

INVx1_ASAP7_75t_L g5565 ( 
.A(n_5360),
.Y(n_5565)
);

INVx2_ASAP7_75t_L g5566 ( 
.A(n_5366),
.Y(n_5566)
);

NAND2xp5_ASAP7_75t_L g5567 ( 
.A(n_5408),
.B(n_5415),
.Y(n_5567)
);

INVx2_ASAP7_75t_L g5568 ( 
.A(n_5383),
.Y(n_5568)
);

INVx2_ASAP7_75t_SL g5569 ( 
.A(n_5344),
.Y(n_5569)
);

BUFx3_ASAP7_75t_L g5570 ( 
.A(n_5318),
.Y(n_5570)
);

NOR2xp33_ASAP7_75t_L g5571 ( 
.A(n_5327),
.B(n_168),
.Y(n_5571)
);

AND2x2_ASAP7_75t_L g5572 ( 
.A(n_5426),
.B(n_169),
.Y(n_5572)
);

INVx2_ASAP7_75t_L g5573 ( 
.A(n_5361),
.Y(n_5573)
);

AND2x2_ASAP7_75t_L g5574 ( 
.A(n_5410),
.B(n_170),
.Y(n_5574)
);

INVx2_ASAP7_75t_SL g5575 ( 
.A(n_5396),
.Y(n_5575)
);

INVx2_ASAP7_75t_L g5576 ( 
.A(n_5362),
.Y(n_5576)
);

NAND2xp5_ASAP7_75t_L g5577 ( 
.A(n_5330),
.B(n_171),
.Y(n_5577)
);

AND2x2_ASAP7_75t_L g5578 ( 
.A(n_5319),
.B(n_171),
.Y(n_5578)
);

INVx1_ASAP7_75t_L g5579 ( 
.A(n_5363),
.Y(n_5579)
);

AND2x2_ASAP7_75t_L g5580 ( 
.A(n_5433),
.B(n_172),
.Y(n_5580)
);

AND2x2_ASAP7_75t_L g5581 ( 
.A(n_5431),
.B(n_173),
.Y(n_5581)
);

BUFx3_ASAP7_75t_L g5582 ( 
.A(n_5462),
.Y(n_5582)
);

NAND2xp5_ASAP7_75t_L g5583 ( 
.A(n_5438),
.B(n_174),
.Y(n_5583)
);

AND2x2_ASAP7_75t_L g5584 ( 
.A(n_5432),
.B(n_5325),
.Y(n_5584)
);

NAND2xp5_ASAP7_75t_L g5585 ( 
.A(n_5436),
.B(n_174),
.Y(n_5585)
);

AND2x2_ASAP7_75t_L g5586 ( 
.A(n_5441),
.B(n_5394),
.Y(n_5586)
);

INVx1_ASAP7_75t_L g5587 ( 
.A(n_5400),
.Y(n_5587)
);

INVxp67_ASAP7_75t_SL g5588 ( 
.A(n_5332),
.Y(n_5588)
);

INVx2_ASAP7_75t_L g5589 ( 
.A(n_5409),
.Y(n_5589)
);

OR2x2_ASAP7_75t_SL g5590 ( 
.A(n_5446),
.B(n_175),
.Y(n_5590)
);

INVx1_ASAP7_75t_L g5591 ( 
.A(n_5359),
.Y(n_5591)
);

AOI21x1_ASAP7_75t_L g5592 ( 
.A1(n_5391),
.A2(n_176),
.B(n_177),
.Y(n_5592)
);

AND2x2_ASAP7_75t_L g5593 ( 
.A(n_5435),
.B(n_176),
.Y(n_5593)
);

OR2x2_ASAP7_75t_L g5594 ( 
.A(n_5358),
.B(n_177),
.Y(n_5594)
);

INVx2_ASAP7_75t_SL g5595 ( 
.A(n_5478),
.Y(n_5595)
);

INVx2_ASAP7_75t_L g5596 ( 
.A(n_5416),
.Y(n_5596)
);

AOI22xp33_ASAP7_75t_L g5597 ( 
.A1(n_5440),
.A2(n_180),
.B1(n_178),
.B2(n_179),
.Y(n_5597)
);

INVx2_ASAP7_75t_R g5598 ( 
.A(n_5455),
.Y(n_5598)
);

INVx2_ASAP7_75t_L g5599 ( 
.A(n_5475),
.Y(n_5599)
);

OAI22xp5_ASAP7_75t_L g5600 ( 
.A1(n_5428),
.A2(n_182),
.B1(n_178),
.B2(n_181),
.Y(n_5600)
);

INVx1_ASAP7_75t_L g5601 ( 
.A(n_5357),
.Y(n_5601)
);

INVx3_ASAP7_75t_L g5602 ( 
.A(n_5445),
.Y(n_5602)
);

INVx1_ASAP7_75t_L g5603 ( 
.A(n_5430),
.Y(n_5603)
);

BUFx3_ASAP7_75t_L g5604 ( 
.A(n_5420),
.Y(n_5604)
);

AND2x2_ASAP7_75t_L g5605 ( 
.A(n_5472),
.B(n_182),
.Y(n_5605)
);

INVx2_ASAP7_75t_L g5606 ( 
.A(n_5378),
.Y(n_5606)
);

INVx2_ASAP7_75t_L g5607 ( 
.A(n_5453),
.Y(n_5607)
);

AND2x4_ASAP7_75t_L g5608 ( 
.A(n_5349),
.B(n_183),
.Y(n_5608)
);

AOI22xp33_ASAP7_75t_SL g5609 ( 
.A1(n_5443),
.A2(n_185),
.B1(n_186),
.B2(n_184),
.Y(n_5609)
);

BUFx3_ASAP7_75t_L g5610 ( 
.A(n_5437),
.Y(n_5610)
);

INVx1_ASAP7_75t_L g5611 ( 
.A(n_5371),
.Y(n_5611)
);

INVx1_ASAP7_75t_L g5612 ( 
.A(n_5384),
.Y(n_5612)
);

AOI22xp5_ASAP7_75t_L g5613 ( 
.A1(n_5447),
.A2(n_186),
.B1(n_183),
.B2(n_185),
.Y(n_5613)
);

AOI22xp5_ASAP7_75t_L g5614 ( 
.A1(n_5452),
.A2(n_5451),
.B1(n_5374),
.B2(n_5444),
.Y(n_5614)
);

NOR2xp33_ASAP7_75t_L g5615 ( 
.A(n_5429),
.B(n_5388),
.Y(n_5615)
);

AND2x2_ASAP7_75t_L g5616 ( 
.A(n_5479),
.B(n_187),
.Y(n_5616)
);

INVx2_ASAP7_75t_L g5617 ( 
.A(n_5457),
.Y(n_5617)
);

INVx2_ASAP7_75t_SL g5618 ( 
.A(n_5387),
.Y(n_5618)
);

HB1xp67_ASAP7_75t_L g5619 ( 
.A(n_5375),
.Y(n_5619)
);

AND2x2_ASAP7_75t_L g5620 ( 
.A(n_5370),
.B(n_187),
.Y(n_5620)
);

AND2x2_ASAP7_75t_L g5621 ( 
.A(n_5449),
.B(n_5381),
.Y(n_5621)
);

INVx1_ASAP7_75t_L g5622 ( 
.A(n_5414),
.Y(n_5622)
);

NAND2xp5_ASAP7_75t_L g5623 ( 
.A(n_5459),
.B(n_188),
.Y(n_5623)
);

INVx1_ASAP7_75t_L g5624 ( 
.A(n_5380),
.Y(n_5624)
);

NAND2xp5_ASAP7_75t_L g5625 ( 
.A(n_5458),
.B(n_188),
.Y(n_5625)
);

NAND2xp5_ASAP7_75t_L g5626 ( 
.A(n_5450),
.B(n_189),
.Y(n_5626)
);

INVx1_ASAP7_75t_L g5627 ( 
.A(n_5351),
.Y(n_5627)
);

OAI22xp5_ASAP7_75t_L g5628 ( 
.A1(n_5442),
.A2(n_191),
.B1(n_189),
.B2(n_190),
.Y(n_5628)
);

HB1xp67_ASAP7_75t_L g5629 ( 
.A(n_5473),
.Y(n_5629)
);

INVx1_ASAP7_75t_L g5630 ( 
.A(n_5352),
.Y(n_5630)
);

OR2x2_ASAP7_75t_L g5631 ( 
.A(n_5477),
.B(n_5448),
.Y(n_5631)
);

INVx3_ASAP7_75t_L g5632 ( 
.A(n_5456),
.Y(n_5632)
);

OR2x2_ASAP7_75t_L g5633 ( 
.A(n_5434),
.B(n_190),
.Y(n_5633)
);

INVx1_ASAP7_75t_L g5634 ( 
.A(n_5454),
.Y(n_5634)
);

INVx1_ASAP7_75t_L g5635 ( 
.A(n_5329),
.Y(n_5635)
);

INVx2_ASAP7_75t_L g5636 ( 
.A(n_5389),
.Y(n_5636)
);

INVxp67_ASAP7_75t_SL g5637 ( 
.A(n_5320),
.Y(n_5637)
);

INVx1_ASAP7_75t_L g5638 ( 
.A(n_5329),
.Y(n_5638)
);

HB1xp67_ASAP7_75t_L g5639 ( 
.A(n_5320),
.Y(n_5639)
);

INVx2_ASAP7_75t_L g5640 ( 
.A(n_5389),
.Y(n_5640)
);

INVx1_ASAP7_75t_L g5641 ( 
.A(n_5329),
.Y(n_5641)
);

AOI22xp33_ASAP7_75t_L g5642 ( 
.A1(n_5406),
.A2(n_193),
.B1(n_191),
.B2(n_192),
.Y(n_5642)
);

AOI22xp33_ASAP7_75t_L g5643 ( 
.A1(n_5406),
.A2(n_195),
.B1(n_193),
.B2(n_194),
.Y(n_5643)
);

BUFx6f_ASAP7_75t_L g5644 ( 
.A(n_5342),
.Y(n_5644)
);

BUFx2_ASAP7_75t_L g5645 ( 
.A(n_5337),
.Y(n_5645)
);

INVx1_ASAP7_75t_L g5646 ( 
.A(n_5329),
.Y(n_5646)
);

INVx2_ASAP7_75t_L g5647 ( 
.A(n_5389),
.Y(n_5647)
);

AOI22xp33_ASAP7_75t_L g5648 ( 
.A1(n_5406),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.Y(n_5648)
);

INVx3_ASAP7_75t_SL g5649 ( 
.A(n_5326),
.Y(n_5649)
);

OAI22xp5_ASAP7_75t_L g5650 ( 
.A1(n_5413),
.A2(n_200),
.B1(n_198),
.B2(n_199),
.Y(n_5650)
);

OR2x2_ASAP7_75t_L g5651 ( 
.A(n_5367),
.B(n_199),
.Y(n_5651)
);

INVx2_ASAP7_75t_SL g5652 ( 
.A(n_5422),
.Y(n_5652)
);

INVx2_ASAP7_75t_L g5653 ( 
.A(n_5389),
.Y(n_5653)
);

OR2x2_ASAP7_75t_L g5654 ( 
.A(n_5367),
.B(n_200),
.Y(n_5654)
);

OAI21xp5_ASAP7_75t_SL g5655 ( 
.A1(n_5406),
.A2(n_201),
.B(n_203),
.Y(n_5655)
);

BUFx2_ASAP7_75t_L g5656 ( 
.A(n_5337),
.Y(n_5656)
);

BUFx3_ASAP7_75t_L g5657 ( 
.A(n_5422),
.Y(n_5657)
);

OAI21xp33_ASAP7_75t_L g5658 ( 
.A1(n_5406),
.A2(n_204),
.B(n_205),
.Y(n_5658)
);

INVx2_ASAP7_75t_L g5659 ( 
.A(n_5389),
.Y(n_5659)
);

INVx1_ASAP7_75t_L g5660 ( 
.A(n_5329),
.Y(n_5660)
);

AOI22xp33_ASAP7_75t_SL g5661 ( 
.A1(n_5406),
.A2(n_206),
.B1(n_207),
.B2(n_205),
.Y(n_5661)
);

AND2x2_ASAP7_75t_L g5662 ( 
.A(n_5367),
.B(n_204),
.Y(n_5662)
);

INVx1_ASAP7_75t_L g5663 ( 
.A(n_5518),
.Y(n_5663)
);

AND2x2_ASAP7_75t_L g5664 ( 
.A(n_5520),
.B(n_206),
.Y(n_5664)
);

HB1xp67_ASAP7_75t_L g5665 ( 
.A(n_5564),
.Y(n_5665)
);

INVx1_ASAP7_75t_L g5666 ( 
.A(n_5522),
.Y(n_5666)
);

AND2x2_ASAP7_75t_L g5667 ( 
.A(n_5645),
.B(n_207),
.Y(n_5667)
);

AND2x2_ASAP7_75t_L g5668 ( 
.A(n_5656),
.B(n_208),
.Y(n_5668)
);

AND2x2_ASAP7_75t_L g5669 ( 
.A(n_5530),
.B(n_208),
.Y(n_5669)
);

INVx2_ASAP7_75t_L g5670 ( 
.A(n_5589),
.Y(n_5670)
);

INVx2_ASAP7_75t_L g5671 ( 
.A(n_5482),
.Y(n_5671)
);

INVx2_ASAP7_75t_L g5672 ( 
.A(n_5636),
.Y(n_5672)
);

INVx2_ASAP7_75t_L g5673 ( 
.A(n_5640),
.Y(n_5673)
);

INVx1_ASAP7_75t_L g5674 ( 
.A(n_5603),
.Y(n_5674)
);

BUFx3_ASAP7_75t_L g5675 ( 
.A(n_5558),
.Y(n_5675)
);

INVx2_ASAP7_75t_L g5676 ( 
.A(n_5647),
.Y(n_5676)
);

AOI22xp33_ASAP7_75t_SL g5677 ( 
.A1(n_5650),
.A2(n_211),
.B1(n_209),
.B2(n_210),
.Y(n_5677)
);

HB1xp67_ASAP7_75t_L g5678 ( 
.A(n_5486),
.Y(n_5678)
);

BUFx3_ASAP7_75t_L g5679 ( 
.A(n_5570),
.Y(n_5679)
);

INVx1_ASAP7_75t_L g5680 ( 
.A(n_5493),
.Y(n_5680)
);

INVx1_ASAP7_75t_SL g5681 ( 
.A(n_5523),
.Y(n_5681)
);

INVx2_ASAP7_75t_L g5682 ( 
.A(n_5653),
.Y(n_5682)
);

INVx2_ASAP7_75t_L g5683 ( 
.A(n_5659),
.Y(n_5683)
);

INVx1_ASAP7_75t_L g5684 ( 
.A(n_5501),
.Y(n_5684)
);

OR2x2_ASAP7_75t_L g5685 ( 
.A(n_5491),
.B(n_209),
.Y(n_5685)
);

NAND2xp5_ASAP7_75t_L g5686 ( 
.A(n_5617),
.B(n_211),
.Y(n_5686)
);

INVx2_ASAP7_75t_L g5687 ( 
.A(n_5539),
.Y(n_5687)
);

INVx2_ASAP7_75t_L g5688 ( 
.A(n_5546),
.Y(n_5688)
);

AND2x4_ASAP7_75t_L g5689 ( 
.A(n_5541),
.B(n_212),
.Y(n_5689)
);

CKINVDCx8_ASAP7_75t_R g5690 ( 
.A(n_5544),
.Y(n_5690)
);

INVx2_ASAP7_75t_SL g5691 ( 
.A(n_5657),
.Y(n_5691)
);

AOI222xp33_ASAP7_75t_L g5692 ( 
.A1(n_5626),
.A2(n_5658),
.B1(n_5655),
.B2(n_5490),
.C1(n_5600),
.C2(n_5597),
.Y(n_5692)
);

INVx2_ASAP7_75t_L g5693 ( 
.A(n_5587),
.Y(n_5693)
);

AND2x2_ASAP7_75t_L g5694 ( 
.A(n_5537),
.B(n_212),
.Y(n_5694)
);

INVx1_ASAP7_75t_L g5695 ( 
.A(n_5502),
.Y(n_5695)
);

NAND2xp5_ASAP7_75t_L g5696 ( 
.A(n_5639),
.B(n_213),
.Y(n_5696)
);

AOI222xp33_ASAP7_75t_SL g5697 ( 
.A1(n_5612),
.A2(n_215),
.B1(n_217),
.B2(n_213),
.C1(n_214),
.C2(n_216),
.Y(n_5697)
);

AO21x2_ASAP7_75t_L g5698 ( 
.A1(n_5611),
.A2(n_214),
.B(n_215),
.Y(n_5698)
);

INVx1_ASAP7_75t_L g5699 ( 
.A(n_5507),
.Y(n_5699)
);

AND2x2_ASAP7_75t_L g5700 ( 
.A(n_5652),
.B(n_216),
.Y(n_5700)
);

AND2x2_ASAP7_75t_L g5701 ( 
.A(n_5536),
.B(n_219),
.Y(n_5701)
);

INVx1_ASAP7_75t_L g5702 ( 
.A(n_5508),
.Y(n_5702)
);

INVx1_ASAP7_75t_L g5703 ( 
.A(n_5635),
.Y(n_5703)
);

HB1xp67_ASAP7_75t_L g5704 ( 
.A(n_5500),
.Y(n_5704)
);

AND2x4_ASAP7_75t_L g5705 ( 
.A(n_5495),
.B(n_219),
.Y(n_5705)
);

INVx1_ASAP7_75t_L g5706 ( 
.A(n_5638),
.Y(n_5706)
);

INVx2_ASAP7_75t_L g5707 ( 
.A(n_5607),
.Y(n_5707)
);

AND2x2_ASAP7_75t_L g5708 ( 
.A(n_5569),
.B(n_220),
.Y(n_5708)
);

AND2x2_ASAP7_75t_L g5709 ( 
.A(n_5584),
.B(n_220),
.Y(n_5709)
);

OR2x2_ASAP7_75t_L g5710 ( 
.A(n_5637),
.B(n_221),
.Y(n_5710)
);

AND2x2_ASAP7_75t_L g5711 ( 
.A(n_5586),
.B(n_221),
.Y(n_5711)
);

INVx2_ASAP7_75t_L g5712 ( 
.A(n_5573),
.Y(n_5712)
);

AO21x2_ASAP7_75t_L g5713 ( 
.A1(n_5619),
.A2(n_223),
.B(n_224),
.Y(n_5713)
);

AND2x2_ASAP7_75t_L g5714 ( 
.A(n_5606),
.B(n_223),
.Y(n_5714)
);

INVx2_ASAP7_75t_L g5715 ( 
.A(n_5553),
.Y(n_5715)
);

BUFx3_ASAP7_75t_L g5716 ( 
.A(n_5649),
.Y(n_5716)
);

INVx1_ASAP7_75t_L g5717 ( 
.A(n_5641),
.Y(n_5717)
);

NAND2xp5_ASAP7_75t_L g5718 ( 
.A(n_5588),
.B(n_224),
.Y(n_5718)
);

INVx1_ASAP7_75t_L g5719 ( 
.A(n_5646),
.Y(n_5719)
);

NAND2xp5_ASAP7_75t_L g5720 ( 
.A(n_5545),
.B(n_225),
.Y(n_5720)
);

INVx1_ASAP7_75t_L g5721 ( 
.A(n_5660),
.Y(n_5721)
);

OR2x2_ASAP7_75t_L g5722 ( 
.A(n_5599),
.B(n_225),
.Y(n_5722)
);

INVxp67_ASAP7_75t_L g5723 ( 
.A(n_5549),
.Y(n_5723)
);

AND2x2_ASAP7_75t_L g5724 ( 
.A(n_5516),
.B(n_226),
.Y(n_5724)
);

AND2x2_ASAP7_75t_L g5725 ( 
.A(n_5602),
.B(n_227),
.Y(n_5725)
);

INVx1_ASAP7_75t_L g5726 ( 
.A(n_5557),
.Y(n_5726)
);

AND2x2_ASAP7_75t_L g5727 ( 
.A(n_5601),
.B(n_227),
.Y(n_5727)
);

AND2x2_ASAP7_75t_L g5728 ( 
.A(n_5591),
.B(n_228),
.Y(n_5728)
);

AND2x2_ASAP7_75t_L g5729 ( 
.A(n_5566),
.B(n_229),
.Y(n_5729)
);

AND2x2_ASAP7_75t_L g5730 ( 
.A(n_5568),
.B(n_230),
.Y(n_5730)
);

AND2x2_ASAP7_75t_L g5731 ( 
.A(n_5540),
.B(n_233),
.Y(n_5731)
);

INVx1_ASAP7_75t_L g5732 ( 
.A(n_5559),
.Y(n_5732)
);

INVx1_ASAP7_75t_L g5733 ( 
.A(n_5560),
.Y(n_5733)
);

INVx2_ASAP7_75t_L g5734 ( 
.A(n_5576),
.Y(n_5734)
);

INVx2_ASAP7_75t_L g5735 ( 
.A(n_5596),
.Y(n_5735)
);

NAND2xp5_ASAP7_75t_L g5736 ( 
.A(n_5567),
.B(n_234),
.Y(n_5736)
);

INVx1_ASAP7_75t_L g5737 ( 
.A(n_5561),
.Y(n_5737)
);

AND2x2_ASAP7_75t_L g5738 ( 
.A(n_5563),
.B(n_5598),
.Y(n_5738)
);

INVx2_ASAP7_75t_L g5739 ( 
.A(n_5483),
.Y(n_5739)
);

INVx1_ASAP7_75t_L g5740 ( 
.A(n_5565),
.Y(n_5740)
);

INVx1_ASAP7_75t_L g5741 ( 
.A(n_5579),
.Y(n_5741)
);

A2O1A1Ixp33_ASAP7_75t_L g5742 ( 
.A1(n_5614),
.A2(n_242),
.B(n_250),
.C(n_234),
.Y(n_5742)
);

INVx1_ASAP7_75t_L g5743 ( 
.A(n_5514),
.Y(n_5743)
);

NAND2xp5_ASAP7_75t_L g5744 ( 
.A(n_5526),
.B(n_235),
.Y(n_5744)
);

AOI22xp33_ASAP7_75t_L g5745 ( 
.A1(n_5492),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.Y(n_5745)
);

NAND2xp5_ASAP7_75t_L g5746 ( 
.A(n_5532),
.B(n_236),
.Y(n_5746)
);

HB1xp67_ASAP7_75t_L g5747 ( 
.A(n_5528),
.Y(n_5747)
);

INVx1_ASAP7_75t_L g5748 ( 
.A(n_5510),
.Y(n_5748)
);

INVx3_ASAP7_75t_L g5749 ( 
.A(n_5506),
.Y(n_5749)
);

INVx2_ASAP7_75t_L g5750 ( 
.A(n_5484),
.Y(n_5750)
);

AOI221x1_ASAP7_75t_L g5751 ( 
.A1(n_5615),
.A2(n_240),
.B1(n_238),
.B2(n_239),
.C(n_241),
.Y(n_5751)
);

INVx3_ASAP7_75t_L g5752 ( 
.A(n_5544),
.Y(n_5752)
);

OR2x2_ASAP7_75t_L g5753 ( 
.A(n_5511),
.B(n_5521),
.Y(n_5753)
);

INVx2_ASAP7_75t_L g5754 ( 
.A(n_5485),
.Y(n_5754)
);

INVx1_ASAP7_75t_L g5755 ( 
.A(n_5527),
.Y(n_5755)
);

INVx2_ASAP7_75t_L g5756 ( 
.A(n_5487),
.Y(n_5756)
);

AND2x2_ASAP7_75t_L g5757 ( 
.A(n_5618),
.B(n_238),
.Y(n_5757)
);

AND2x2_ASAP7_75t_L g5758 ( 
.A(n_5575),
.B(n_240),
.Y(n_5758)
);

AND2x2_ASAP7_75t_L g5759 ( 
.A(n_5595),
.B(n_241),
.Y(n_5759)
);

HB1xp67_ASAP7_75t_L g5760 ( 
.A(n_5497),
.Y(n_5760)
);

INVx2_ASAP7_75t_L g5761 ( 
.A(n_5499),
.Y(n_5761)
);

BUFx3_ASAP7_75t_L g5762 ( 
.A(n_5582),
.Y(n_5762)
);

OA21x2_ASAP7_75t_L g5763 ( 
.A1(n_5504),
.A2(n_243),
.B(n_244),
.Y(n_5763)
);

NAND2xp5_ASAP7_75t_L g5764 ( 
.A(n_5533),
.B(n_244),
.Y(n_5764)
);

INVx1_ASAP7_75t_L g5765 ( 
.A(n_5548),
.Y(n_5765)
);

INVx3_ASAP7_75t_L g5766 ( 
.A(n_5512),
.Y(n_5766)
);

INVx2_ASAP7_75t_L g5767 ( 
.A(n_5550),
.Y(n_5767)
);

AND2x4_ASAP7_75t_SL g5768 ( 
.A(n_5498),
.B(n_245),
.Y(n_5768)
);

INVx2_ASAP7_75t_L g5769 ( 
.A(n_5554),
.Y(n_5769)
);

AOI22xp5_ASAP7_75t_L g5770 ( 
.A1(n_5661),
.A2(n_247),
.B1(n_245),
.B2(n_246),
.Y(n_5770)
);

NOR2x1_ASAP7_75t_SL g5771 ( 
.A(n_5651),
.B(n_247),
.Y(n_5771)
);

INVx1_ASAP7_75t_L g5772 ( 
.A(n_5551),
.Y(n_5772)
);

AND2x2_ASAP7_75t_L g5773 ( 
.A(n_5610),
.B(n_248),
.Y(n_5773)
);

INVx2_ASAP7_75t_L g5774 ( 
.A(n_5654),
.Y(n_5774)
);

OR2x2_ASAP7_75t_L g5775 ( 
.A(n_5524),
.B(n_248),
.Y(n_5775)
);

INVx2_ASAP7_75t_L g5776 ( 
.A(n_5574),
.Y(n_5776)
);

AOI221xp5_ASAP7_75t_L g5777 ( 
.A1(n_5609),
.A2(n_251),
.B1(n_249),
.B2(n_250),
.C(n_253),
.Y(n_5777)
);

OR2x2_ASAP7_75t_L g5778 ( 
.A(n_5577),
.B(n_249),
.Y(n_5778)
);

INVx1_ASAP7_75t_L g5779 ( 
.A(n_5525),
.Y(n_5779)
);

AND2x2_ASAP7_75t_L g5780 ( 
.A(n_5535),
.B(n_251),
.Y(n_5780)
);

INVx1_ASAP7_75t_L g5781 ( 
.A(n_5556),
.Y(n_5781)
);

AND2x2_ASAP7_75t_L g5782 ( 
.A(n_5621),
.B(n_254),
.Y(n_5782)
);

OR2x2_ASAP7_75t_L g5783 ( 
.A(n_5624),
.B(n_254),
.Y(n_5783)
);

INVx4_ASAP7_75t_L g5784 ( 
.A(n_5512),
.Y(n_5784)
);

INVx2_ASAP7_75t_L g5785 ( 
.A(n_5517),
.Y(n_5785)
);

INVxp67_ASAP7_75t_SL g5786 ( 
.A(n_5629),
.Y(n_5786)
);

NOR2x1_ASAP7_75t_L g5787 ( 
.A(n_5489),
.B(n_255),
.Y(n_5787)
);

AND2x2_ASAP7_75t_L g5788 ( 
.A(n_5555),
.B(n_256),
.Y(n_5788)
);

INVx2_ASAP7_75t_L g5789 ( 
.A(n_5572),
.Y(n_5789)
);

HB1xp67_ASAP7_75t_L g5790 ( 
.A(n_5488),
.Y(n_5790)
);

BUFx3_ASAP7_75t_L g5791 ( 
.A(n_5542),
.Y(n_5791)
);

HB1xp67_ASAP7_75t_L g5792 ( 
.A(n_5662),
.Y(n_5792)
);

INVx1_ASAP7_75t_L g5793 ( 
.A(n_5529),
.Y(n_5793)
);

INVx1_ASAP7_75t_L g5794 ( 
.A(n_5505),
.Y(n_5794)
);

INVx1_ASAP7_75t_L g5795 ( 
.A(n_5543),
.Y(n_5795)
);

INVx1_ASAP7_75t_L g5796 ( 
.A(n_5513),
.Y(n_5796)
);

AOI22xp33_ASAP7_75t_L g5797 ( 
.A1(n_5552),
.A2(n_259),
.B1(n_257),
.B2(n_258),
.Y(n_5797)
);

INVx1_ASAP7_75t_L g5798 ( 
.A(n_5627),
.Y(n_5798)
);

INVx2_ASAP7_75t_SL g5799 ( 
.A(n_5542),
.Y(n_5799)
);

INVx2_ASAP7_75t_L g5800 ( 
.A(n_5630),
.Y(n_5800)
);

INVx2_ASAP7_75t_L g5801 ( 
.A(n_5531),
.Y(n_5801)
);

INVx1_ASAP7_75t_L g5802 ( 
.A(n_5515),
.Y(n_5802)
);

NAND2xp5_ASAP7_75t_L g5803 ( 
.A(n_5538),
.B(n_5580),
.Y(n_5803)
);

INVx1_ASAP7_75t_L g5804 ( 
.A(n_5503),
.Y(n_5804)
);

BUFx2_ASAP7_75t_L g5805 ( 
.A(n_5608),
.Y(n_5805)
);

INVx1_ASAP7_75t_L g5806 ( 
.A(n_5503),
.Y(n_5806)
);

INVxp67_ASAP7_75t_SL g5807 ( 
.A(n_5585),
.Y(n_5807)
);

INVx2_ASAP7_75t_L g5808 ( 
.A(n_5496),
.Y(n_5808)
);

INVx1_ASAP7_75t_L g5809 ( 
.A(n_5581),
.Y(n_5809)
);

HB1xp67_ASAP7_75t_L g5810 ( 
.A(n_5622),
.Y(n_5810)
);

AOI33xp33_ASAP7_75t_L g5811 ( 
.A1(n_5519),
.A2(n_260),
.A3(n_262),
.B1(n_257),
.B2(n_259),
.B3(n_261),
.Y(n_5811)
);

AND2x2_ASAP7_75t_L g5812 ( 
.A(n_5494),
.B(n_261),
.Y(n_5812)
);

OR2x2_ASAP7_75t_L g5813 ( 
.A(n_5594),
.B(n_5562),
.Y(n_5813)
);

INVx2_ASAP7_75t_L g5814 ( 
.A(n_5644),
.Y(n_5814)
);

HB1xp67_ASAP7_75t_L g5815 ( 
.A(n_5632),
.Y(n_5815)
);

AND2x4_ASAP7_75t_L g5816 ( 
.A(n_5604),
.B(n_262),
.Y(n_5816)
);

OR2x2_ASAP7_75t_L g5817 ( 
.A(n_5625),
.B(n_263),
.Y(n_5817)
);

HB1xp67_ASAP7_75t_L g5818 ( 
.A(n_5593),
.Y(n_5818)
);

HB1xp67_ASAP7_75t_L g5819 ( 
.A(n_5592),
.Y(n_5819)
);

OAI21xp5_ASAP7_75t_L g5820 ( 
.A1(n_5509),
.A2(n_263),
.B(n_264),
.Y(n_5820)
);

INVx2_ASAP7_75t_L g5821 ( 
.A(n_5644),
.Y(n_5821)
);

INVx2_ASAP7_75t_L g5822 ( 
.A(n_5631),
.Y(n_5822)
);

INVx2_ASAP7_75t_L g5823 ( 
.A(n_5534),
.Y(n_5823)
);

INVx1_ASAP7_75t_L g5824 ( 
.A(n_5583),
.Y(n_5824)
);

INVx1_ASAP7_75t_L g5825 ( 
.A(n_5547),
.Y(n_5825)
);

INVx2_ASAP7_75t_L g5826 ( 
.A(n_5578),
.Y(n_5826)
);

BUFx6f_ASAP7_75t_L g5827 ( 
.A(n_5634),
.Y(n_5827)
);

INVx2_ASAP7_75t_L g5828 ( 
.A(n_5633),
.Y(n_5828)
);

NAND2xp5_ASAP7_75t_L g5829 ( 
.A(n_5571),
.B(n_264),
.Y(n_5829)
);

AND2x2_ASAP7_75t_L g5830 ( 
.A(n_5605),
.B(n_265),
.Y(n_5830)
);

AND2x2_ASAP7_75t_L g5831 ( 
.A(n_5616),
.B(n_5620),
.Y(n_5831)
);

INVx2_ASAP7_75t_L g5832 ( 
.A(n_5590),
.Y(n_5832)
);

NOR2xp33_ASAP7_75t_L g5833 ( 
.A(n_5623),
.B(n_266),
.Y(n_5833)
);

INVx1_ASAP7_75t_SL g5834 ( 
.A(n_5552),
.Y(n_5834)
);

BUFx3_ASAP7_75t_L g5835 ( 
.A(n_5613),
.Y(n_5835)
);

INVx2_ASAP7_75t_L g5836 ( 
.A(n_5628),
.Y(n_5836)
);

INVx1_ASAP7_75t_L g5837 ( 
.A(n_5481),
.Y(n_5837)
);

NAND2xp5_ASAP7_75t_SL g5838 ( 
.A(n_5648),
.B(n_267),
.Y(n_5838)
);

INVx3_ASAP7_75t_L g5839 ( 
.A(n_5642),
.Y(n_5839)
);

BUFx3_ASAP7_75t_L g5840 ( 
.A(n_5643),
.Y(n_5840)
);

INVx1_ASAP7_75t_L g5841 ( 
.A(n_5518),
.Y(n_5841)
);

BUFx2_ASAP7_75t_L g5842 ( 
.A(n_5541),
.Y(n_5842)
);

INVx2_ASAP7_75t_L g5843 ( 
.A(n_5589),
.Y(n_5843)
);

INVx2_ASAP7_75t_SL g5844 ( 
.A(n_5541),
.Y(n_5844)
);

NAND2xp5_ASAP7_75t_L g5845 ( 
.A(n_5617),
.B(n_267),
.Y(n_5845)
);

OR2x2_ASAP7_75t_L g5846 ( 
.A(n_5603),
.B(n_268),
.Y(n_5846)
);

AND2x2_ASAP7_75t_L g5847 ( 
.A(n_5520),
.B(n_268),
.Y(n_5847)
);

INVx2_ASAP7_75t_L g5848 ( 
.A(n_5589),
.Y(n_5848)
);

HB1xp67_ASAP7_75t_L g5849 ( 
.A(n_5564),
.Y(n_5849)
);

NAND2xp5_ASAP7_75t_L g5850 ( 
.A(n_5617),
.B(n_269),
.Y(n_5850)
);

AND2x2_ASAP7_75t_L g5851 ( 
.A(n_5520),
.B(n_269),
.Y(n_5851)
);

INVx1_ASAP7_75t_L g5852 ( 
.A(n_5518),
.Y(n_5852)
);

BUFx2_ASAP7_75t_L g5853 ( 
.A(n_5541),
.Y(n_5853)
);

AND2x2_ASAP7_75t_L g5854 ( 
.A(n_5520),
.B(n_270),
.Y(n_5854)
);

BUFx6f_ASAP7_75t_L g5855 ( 
.A(n_5570),
.Y(n_5855)
);

AND2x2_ASAP7_75t_L g5856 ( 
.A(n_5520),
.B(n_270),
.Y(n_5856)
);

INVx1_ASAP7_75t_L g5857 ( 
.A(n_5518),
.Y(n_5857)
);

AND2x2_ASAP7_75t_L g5858 ( 
.A(n_5520),
.B(n_271),
.Y(n_5858)
);

AND2x2_ASAP7_75t_L g5859 ( 
.A(n_5520),
.B(n_272),
.Y(n_5859)
);

INVx2_ASAP7_75t_SL g5860 ( 
.A(n_5541),
.Y(n_5860)
);

AOI21xp5_ASAP7_75t_L g5861 ( 
.A1(n_5655),
.A2(n_273),
.B(n_274),
.Y(n_5861)
);

INVx1_ASAP7_75t_L g5862 ( 
.A(n_5518),
.Y(n_5862)
);

AND2x2_ASAP7_75t_L g5863 ( 
.A(n_5520),
.B(n_273),
.Y(n_5863)
);

INVx1_ASAP7_75t_L g5864 ( 
.A(n_5518),
.Y(n_5864)
);

AND2x2_ASAP7_75t_L g5865 ( 
.A(n_5520),
.B(n_275),
.Y(n_5865)
);

INVx2_ASAP7_75t_SL g5866 ( 
.A(n_5541),
.Y(n_5866)
);

INVx1_ASAP7_75t_L g5867 ( 
.A(n_5674),
.Y(n_5867)
);

NOR2xp33_ASAP7_75t_L g5868 ( 
.A(n_5681),
.B(n_276),
.Y(n_5868)
);

AND2x2_ASAP7_75t_L g5869 ( 
.A(n_5738),
.B(n_277),
.Y(n_5869)
);

INVx2_ASAP7_75t_L g5870 ( 
.A(n_5827),
.Y(n_5870)
);

AND2x2_ASAP7_75t_L g5871 ( 
.A(n_5834),
.B(n_277),
.Y(n_5871)
);

NAND2xp5_ASAP7_75t_L g5872 ( 
.A(n_5807),
.B(n_278),
.Y(n_5872)
);

INVx1_ASAP7_75t_L g5873 ( 
.A(n_5741),
.Y(n_5873)
);

AND2x2_ASAP7_75t_L g5874 ( 
.A(n_5805),
.B(n_278),
.Y(n_5874)
);

INVx1_ASAP7_75t_L g5875 ( 
.A(n_5680),
.Y(n_5875)
);

INVx1_ASAP7_75t_L g5876 ( 
.A(n_5684),
.Y(n_5876)
);

AND2x2_ASAP7_75t_L g5877 ( 
.A(n_5842),
.B(n_279),
.Y(n_5877)
);

INVxp67_ASAP7_75t_SL g5878 ( 
.A(n_5819),
.Y(n_5878)
);

INVx2_ASAP7_75t_L g5879 ( 
.A(n_5827),
.Y(n_5879)
);

OR2x2_ASAP7_75t_L g5880 ( 
.A(n_5678),
.B(n_279),
.Y(n_5880)
);

INVx2_ASAP7_75t_L g5881 ( 
.A(n_5753),
.Y(n_5881)
);

AND2x4_ASAP7_75t_SL g5882 ( 
.A(n_5855),
.B(n_5749),
.Y(n_5882)
);

INVx2_ASAP7_75t_L g5883 ( 
.A(n_5670),
.Y(n_5883)
);

NAND2xp5_ASAP7_75t_L g5884 ( 
.A(n_5828),
.B(n_280),
.Y(n_5884)
);

OR2x2_ASAP7_75t_L g5885 ( 
.A(n_5704),
.B(n_281),
.Y(n_5885)
);

BUFx2_ASAP7_75t_L g5886 ( 
.A(n_5853),
.Y(n_5886)
);

AND2x2_ASAP7_75t_L g5887 ( 
.A(n_5822),
.B(n_5687),
.Y(n_5887)
);

AND2x2_ASAP7_75t_L g5888 ( 
.A(n_5688),
.B(n_282),
.Y(n_5888)
);

AND2x4_ASAP7_75t_L g5889 ( 
.A(n_5675),
.B(n_283),
.Y(n_5889)
);

INVx1_ASAP7_75t_L g5890 ( 
.A(n_5695),
.Y(n_5890)
);

HB1xp67_ASAP7_75t_L g5891 ( 
.A(n_5747),
.Y(n_5891)
);

AND2x4_ASAP7_75t_L g5892 ( 
.A(n_5691),
.B(n_283),
.Y(n_5892)
);

NAND2xp5_ASAP7_75t_L g5893 ( 
.A(n_5723),
.B(n_285),
.Y(n_5893)
);

AND2x2_ASAP7_75t_L g5894 ( 
.A(n_5790),
.B(n_286),
.Y(n_5894)
);

AND2x2_ASAP7_75t_L g5895 ( 
.A(n_5792),
.B(n_287),
.Y(n_5895)
);

INVx2_ASAP7_75t_L g5896 ( 
.A(n_5843),
.Y(n_5896)
);

INVx2_ASAP7_75t_L g5897 ( 
.A(n_5848),
.Y(n_5897)
);

AND2x2_ASAP7_75t_L g5898 ( 
.A(n_5818),
.B(n_288),
.Y(n_5898)
);

BUFx3_ASAP7_75t_L g5899 ( 
.A(n_5679),
.Y(n_5899)
);

INVx5_ASAP7_75t_L g5900 ( 
.A(n_5855),
.Y(n_5900)
);

AOI222xp33_ASAP7_75t_L g5901 ( 
.A1(n_5820),
.A2(n_291),
.B1(n_293),
.B2(n_289),
.C1(n_290),
.C2(n_292),
.Y(n_5901)
);

AND2x2_ASAP7_75t_L g5902 ( 
.A(n_5769),
.B(n_289),
.Y(n_5902)
);

INVx1_ASAP7_75t_L g5903 ( 
.A(n_5699),
.Y(n_5903)
);

AND2x4_ASAP7_75t_L g5904 ( 
.A(n_5844),
.B(n_291),
.Y(n_5904)
);

OR2x2_ASAP7_75t_L g5905 ( 
.A(n_5774),
.B(n_292),
.Y(n_5905)
);

AND2x2_ASAP7_75t_L g5906 ( 
.A(n_5814),
.B(n_293),
.Y(n_5906)
);

INVx1_ASAP7_75t_L g5907 ( 
.A(n_5702),
.Y(n_5907)
);

AND2x2_ASAP7_75t_L g5908 ( 
.A(n_5821),
.B(n_294),
.Y(n_5908)
);

INVx1_ASAP7_75t_SL g5909 ( 
.A(n_5716),
.Y(n_5909)
);

OR2x2_ASAP7_75t_L g5910 ( 
.A(n_5781),
.B(n_295),
.Y(n_5910)
);

INVx2_ASAP7_75t_L g5911 ( 
.A(n_5767),
.Y(n_5911)
);

INVx1_ASAP7_75t_L g5912 ( 
.A(n_5703),
.Y(n_5912)
);

AND2x2_ASAP7_75t_L g5913 ( 
.A(n_5860),
.B(n_295),
.Y(n_5913)
);

AND2x2_ASAP7_75t_L g5914 ( 
.A(n_5866),
.B(n_296),
.Y(n_5914)
);

HB1xp67_ASAP7_75t_L g5915 ( 
.A(n_5665),
.Y(n_5915)
);

INVx1_ASAP7_75t_L g5916 ( 
.A(n_5706),
.Y(n_5916)
);

INVx1_ASAP7_75t_L g5917 ( 
.A(n_5717),
.Y(n_5917)
);

AND2x4_ASAP7_75t_L g5918 ( 
.A(n_5762),
.B(n_296),
.Y(n_5918)
);

HB1xp67_ASAP7_75t_L g5919 ( 
.A(n_5849),
.Y(n_5919)
);

INVx2_ASAP7_75t_L g5920 ( 
.A(n_5739),
.Y(n_5920)
);

INVx1_ASAP7_75t_L g5921 ( 
.A(n_5719),
.Y(n_5921)
);

NAND2xp5_ASAP7_75t_L g5922 ( 
.A(n_5779),
.B(n_297),
.Y(n_5922)
);

INVx1_ASAP7_75t_L g5923 ( 
.A(n_5721),
.Y(n_5923)
);

AND2x2_ASAP7_75t_L g5924 ( 
.A(n_5776),
.B(n_297),
.Y(n_5924)
);

AND2x2_ASAP7_75t_L g5925 ( 
.A(n_5772),
.B(n_298),
.Y(n_5925)
);

INVx2_ASAP7_75t_L g5926 ( 
.A(n_5750),
.Y(n_5926)
);

INVx1_ASAP7_75t_L g5927 ( 
.A(n_5726),
.Y(n_5927)
);

OR2x2_ASAP7_75t_L g5928 ( 
.A(n_5802),
.B(n_298),
.Y(n_5928)
);

INVx1_ASAP7_75t_L g5929 ( 
.A(n_5732),
.Y(n_5929)
);

OR2x2_ASAP7_75t_L g5930 ( 
.A(n_5824),
.B(n_299),
.Y(n_5930)
);

HB1xp67_ASAP7_75t_L g5931 ( 
.A(n_5804),
.Y(n_5931)
);

AND2x4_ASAP7_75t_L g5932 ( 
.A(n_5752),
.B(n_300),
.Y(n_5932)
);

AND2x2_ASAP7_75t_L g5933 ( 
.A(n_5785),
.B(n_300),
.Y(n_5933)
);

AND2x2_ASAP7_75t_L g5934 ( 
.A(n_5808),
.B(n_301),
.Y(n_5934)
);

INVx2_ASAP7_75t_L g5935 ( 
.A(n_5754),
.Y(n_5935)
);

INVx2_ASAP7_75t_L g5936 ( 
.A(n_5756),
.Y(n_5936)
);

NAND2xp5_ASAP7_75t_L g5937 ( 
.A(n_5663),
.B(n_301),
.Y(n_5937)
);

AND2x2_ASAP7_75t_L g5938 ( 
.A(n_5789),
.B(n_5826),
.Y(n_5938)
);

NAND2xp5_ASAP7_75t_L g5939 ( 
.A(n_5666),
.B(n_302),
.Y(n_5939)
);

NAND2xp5_ASAP7_75t_L g5940 ( 
.A(n_5841),
.B(n_302),
.Y(n_5940)
);

AND2x4_ASAP7_75t_L g5941 ( 
.A(n_5791),
.B(n_303),
.Y(n_5941)
);

HB1xp67_ASAP7_75t_L g5942 ( 
.A(n_5806),
.Y(n_5942)
);

AND2x4_ASAP7_75t_L g5943 ( 
.A(n_5784),
.B(n_303),
.Y(n_5943)
);

INVx3_ASAP7_75t_L g5944 ( 
.A(n_5690),
.Y(n_5944)
);

INVx2_ASAP7_75t_L g5945 ( 
.A(n_5761),
.Y(n_5945)
);

INVx2_ASAP7_75t_L g5946 ( 
.A(n_5800),
.Y(n_5946)
);

INVx2_ASAP7_75t_L g5947 ( 
.A(n_5671),
.Y(n_5947)
);

HB1xp67_ASAP7_75t_L g5948 ( 
.A(n_5760),
.Y(n_5948)
);

AND2x2_ASAP7_75t_L g5949 ( 
.A(n_5794),
.B(n_5809),
.Y(n_5949)
);

INVx2_ASAP7_75t_L g5950 ( 
.A(n_5672),
.Y(n_5950)
);

NAND2xp5_ASAP7_75t_L g5951 ( 
.A(n_5852),
.B(n_304),
.Y(n_5951)
);

OR2x2_ASAP7_75t_L g5952 ( 
.A(n_5857),
.B(n_304),
.Y(n_5952)
);

INVx2_ASAP7_75t_L g5953 ( 
.A(n_5673),
.Y(n_5953)
);

INVx2_ASAP7_75t_L g5954 ( 
.A(n_5676),
.Y(n_5954)
);

AND2x2_ASAP7_75t_SL g5955 ( 
.A(n_5768),
.B(n_305),
.Y(n_5955)
);

AND2x4_ASAP7_75t_L g5956 ( 
.A(n_5799),
.B(n_305),
.Y(n_5956)
);

INVx1_ASAP7_75t_L g5957 ( 
.A(n_5733),
.Y(n_5957)
);

NAND2xp5_ASAP7_75t_L g5958 ( 
.A(n_5862),
.B(n_306),
.Y(n_5958)
);

INVx2_ASAP7_75t_L g5959 ( 
.A(n_5682),
.Y(n_5959)
);

NAND2xp5_ASAP7_75t_L g5960 ( 
.A(n_5864),
.B(n_306),
.Y(n_5960)
);

NAND2xp5_ASAP7_75t_L g5961 ( 
.A(n_5718),
.B(n_307),
.Y(n_5961)
);

INVx1_ASAP7_75t_L g5962 ( 
.A(n_5737),
.Y(n_5962)
);

INVx2_ASAP7_75t_L g5963 ( 
.A(n_5683),
.Y(n_5963)
);

OR2x6_ASAP7_75t_L g5964 ( 
.A(n_5861),
.B(n_307),
.Y(n_5964)
);

AND2x4_ASAP7_75t_L g5965 ( 
.A(n_5766),
.B(n_308),
.Y(n_5965)
);

OR2x2_ASAP7_75t_L g5966 ( 
.A(n_5793),
.B(n_308),
.Y(n_5966)
);

OR2x2_ASAP7_75t_L g5967 ( 
.A(n_5796),
.B(n_309),
.Y(n_5967)
);

INVx1_ASAP7_75t_L g5968 ( 
.A(n_5740),
.Y(n_5968)
);

OR2x2_ASAP7_75t_L g5969 ( 
.A(n_5813),
.B(n_309),
.Y(n_5969)
);

OAI22xp5_ASAP7_75t_L g5970 ( 
.A1(n_5835),
.A2(n_312),
.B1(n_310),
.B2(n_311),
.Y(n_5970)
);

BUFx3_ASAP7_75t_L g5971 ( 
.A(n_5689),
.Y(n_5971)
);

NAND2xp5_ASAP7_75t_L g5972 ( 
.A(n_5686),
.B(n_310),
.Y(n_5972)
);

AND2x2_ASAP7_75t_L g5973 ( 
.A(n_5825),
.B(n_313),
.Y(n_5973)
);

HB1xp67_ASAP7_75t_L g5974 ( 
.A(n_5798),
.Y(n_5974)
);

HB1xp67_ASAP7_75t_L g5975 ( 
.A(n_5810),
.Y(n_5975)
);

NOR2xp33_ASAP7_75t_L g5976 ( 
.A(n_5832),
.B(n_313),
.Y(n_5976)
);

AND2x4_ASAP7_75t_L g5977 ( 
.A(n_5801),
.B(n_314),
.Y(n_5977)
);

INVxp67_ASAP7_75t_L g5978 ( 
.A(n_5771),
.Y(n_5978)
);

AND2x2_ASAP7_75t_L g5979 ( 
.A(n_5795),
.B(n_315),
.Y(n_5979)
);

INVx2_ASAP7_75t_L g5980 ( 
.A(n_5712),
.Y(n_5980)
);

BUFx3_ASAP7_75t_L g5981 ( 
.A(n_5759),
.Y(n_5981)
);

AND2x2_ASAP7_75t_L g5982 ( 
.A(n_5707),
.B(n_315),
.Y(n_5982)
);

AND2x2_ASAP7_75t_L g5983 ( 
.A(n_5735),
.B(n_316),
.Y(n_5983)
);

AND2x2_ASAP7_75t_L g5984 ( 
.A(n_5715),
.B(n_316),
.Y(n_5984)
);

AND2x4_ASAP7_75t_L g5985 ( 
.A(n_5823),
.B(n_317),
.Y(n_5985)
);

BUFx2_ASAP7_75t_SL g5986 ( 
.A(n_5705),
.Y(n_5986)
);

NAND2xp5_ASAP7_75t_L g5987 ( 
.A(n_5845),
.B(n_317),
.Y(n_5987)
);

INVx1_ASAP7_75t_L g5988 ( 
.A(n_5743),
.Y(n_5988)
);

INVx2_ASAP7_75t_L g5989 ( 
.A(n_5734),
.Y(n_5989)
);

OR2x2_ASAP7_75t_L g5990 ( 
.A(n_5748),
.B(n_319),
.Y(n_5990)
);

NAND2xp5_ASAP7_75t_L g5991 ( 
.A(n_5850),
.B(n_319),
.Y(n_5991)
);

AND2x2_ASAP7_75t_L g5992 ( 
.A(n_5831),
.B(n_5786),
.Y(n_5992)
);

AND2x2_ASAP7_75t_L g5993 ( 
.A(n_5765),
.B(n_320),
.Y(n_5993)
);

INVx2_ASAP7_75t_L g5994 ( 
.A(n_5693),
.Y(n_5994)
);

OR2x2_ASAP7_75t_L g5995 ( 
.A(n_5755),
.B(n_321),
.Y(n_5995)
);

INVx1_ASAP7_75t_L g5996 ( 
.A(n_5764),
.Y(n_5996)
);

AND2x2_ASAP7_75t_L g5997 ( 
.A(n_5664),
.B(n_321),
.Y(n_5997)
);

INVx1_ASAP7_75t_L g5998 ( 
.A(n_5783),
.Y(n_5998)
);

AND2x2_ASAP7_75t_L g5999 ( 
.A(n_5667),
.B(n_322),
.Y(n_5999)
);

NAND2xp5_ASAP7_75t_L g6000 ( 
.A(n_5744),
.B(n_323),
.Y(n_6000)
);

AOI22xp33_ASAP7_75t_L g6001 ( 
.A1(n_5840),
.A2(n_326),
.B1(n_324),
.B2(n_325),
.Y(n_6001)
);

HB1xp67_ASAP7_75t_L g6002 ( 
.A(n_5763),
.Y(n_6002)
);

AND2x2_ASAP7_75t_L g6003 ( 
.A(n_5668),
.B(n_324),
.Y(n_6003)
);

AND2x2_ASAP7_75t_L g6004 ( 
.A(n_5847),
.B(n_5863),
.Y(n_6004)
);

INVx2_ASAP7_75t_L g6005 ( 
.A(n_5815),
.Y(n_6005)
);

INVx1_ASAP7_75t_L g6006 ( 
.A(n_5722),
.Y(n_6006)
);

HB1xp67_ASAP7_75t_L g6007 ( 
.A(n_5846),
.Y(n_6007)
);

INVx1_ASAP7_75t_L g6008 ( 
.A(n_5720),
.Y(n_6008)
);

INVx1_ASAP7_75t_L g6009 ( 
.A(n_5746),
.Y(n_6009)
);

INVxp67_ASAP7_75t_L g6010 ( 
.A(n_5787),
.Y(n_6010)
);

INVx2_ASAP7_75t_L g6011 ( 
.A(n_5725),
.Y(n_6011)
);

INVx1_ASAP7_75t_L g6012 ( 
.A(n_5710),
.Y(n_6012)
);

INVx1_ASAP7_75t_L g6013 ( 
.A(n_5685),
.Y(n_6013)
);

NAND2xp5_ASAP7_75t_SL g6014 ( 
.A(n_5836),
.B(n_326),
.Y(n_6014)
);

INVx2_ASAP7_75t_L g6015 ( 
.A(n_5724),
.Y(n_6015)
);

INVxp67_ASAP7_75t_L g6016 ( 
.A(n_5713),
.Y(n_6016)
);

NOR2xp67_ASAP7_75t_L g6017 ( 
.A(n_5694),
.B(n_327),
.Y(n_6017)
);

INVx2_ASAP7_75t_L g6018 ( 
.A(n_5729),
.Y(n_6018)
);

HB1xp67_ASAP7_75t_L g6019 ( 
.A(n_5698),
.Y(n_6019)
);

INVx1_ASAP7_75t_L g6020 ( 
.A(n_5714),
.Y(n_6020)
);

NAND2xp5_ASAP7_75t_L g6021 ( 
.A(n_5736),
.B(n_327),
.Y(n_6021)
);

NAND2xp5_ASAP7_75t_L g6022 ( 
.A(n_5701),
.B(n_328),
.Y(n_6022)
);

OR2x2_ASAP7_75t_L g6023 ( 
.A(n_5803),
.B(n_328),
.Y(n_6023)
);

INVx2_ASAP7_75t_L g6024 ( 
.A(n_5730),
.Y(n_6024)
);

INVx1_ASAP7_75t_L g6025 ( 
.A(n_5696),
.Y(n_6025)
);

AND2x2_ASAP7_75t_L g6026 ( 
.A(n_5851),
.B(n_329),
.Y(n_6026)
);

BUFx3_ASAP7_75t_L g6027 ( 
.A(n_5700),
.Y(n_6027)
);

AND2x2_ASAP7_75t_L g6028 ( 
.A(n_5854),
.B(n_5856),
.Y(n_6028)
);

INVx1_ASAP7_75t_L g6029 ( 
.A(n_5728),
.Y(n_6029)
);

INVx1_ASAP7_75t_L g6030 ( 
.A(n_5727),
.Y(n_6030)
);

AND2x4_ASAP7_75t_L g6031 ( 
.A(n_5858),
.B(n_330),
.Y(n_6031)
);

NAND2xp5_ASAP7_75t_L g6032 ( 
.A(n_5669),
.B(n_330),
.Y(n_6032)
);

AND2x4_ASAP7_75t_L g6033 ( 
.A(n_5859),
.B(n_331),
.Y(n_6033)
);

NAND2xp5_ASAP7_75t_L g6034 ( 
.A(n_5865),
.B(n_331),
.Y(n_6034)
);

INVx1_ASAP7_75t_L g6035 ( 
.A(n_5708),
.Y(n_6035)
);

NAND2xp5_ASAP7_75t_L g6036 ( 
.A(n_5709),
.B(n_332),
.Y(n_6036)
);

AND2x4_ASAP7_75t_SL g6037 ( 
.A(n_5816),
.B(n_5773),
.Y(n_6037)
);

AND2x2_ASAP7_75t_L g6038 ( 
.A(n_5711),
.B(n_332),
.Y(n_6038)
);

INVxp67_ASAP7_75t_SL g6039 ( 
.A(n_5817),
.Y(n_6039)
);

INVx2_ASAP7_75t_L g6040 ( 
.A(n_5731),
.Y(n_6040)
);

NOR2xp33_ASAP7_75t_SL g6041 ( 
.A(n_5742),
.B(n_334),
.Y(n_6041)
);

INVx2_ASAP7_75t_L g6042 ( 
.A(n_5758),
.Y(n_6042)
);

AND2x2_ASAP7_75t_L g6043 ( 
.A(n_5757),
.B(n_5782),
.Y(n_6043)
);

AND2x2_ASAP7_75t_L g6044 ( 
.A(n_5780),
.B(n_334),
.Y(n_6044)
);

INVx1_ASAP7_75t_L g6045 ( 
.A(n_5775),
.Y(n_6045)
);

AND2x2_ASAP7_75t_L g6046 ( 
.A(n_5788),
.B(n_335),
.Y(n_6046)
);

NAND2xp5_ASAP7_75t_L g6047 ( 
.A(n_5839),
.B(n_335),
.Y(n_6047)
);

AND2x2_ASAP7_75t_L g6048 ( 
.A(n_5812),
.B(n_336),
.Y(n_6048)
);

HB1xp67_ASAP7_75t_L g6049 ( 
.A(n_5778),
.Y(n_6049)
);

INVx2_ASAP7_75t_L g6050 ( 
.A(n_5830),
.Y(n_6050)
);

AND2x2_ASAP7_75t_L g6051 ( 
.A(n_5837),
.B(n_336),
.Y(n_6051)
);

NAND2xp5_ASAP7_75t_L g6052 ( 
.A(n_5833),
.B(n_5829),
.Y(n_6052)
);

INVx1_ASAP7_75t_L g6053 ( 
.A(n_5751),
.Y(n_6053)
);

INVx4_ASAP7_75t_L g6054 ( 
.A(n_5697),
.Y(n_6054)
);

HB1xp67_ASAP7_75t_L g6055 ( 
.A(n_5692),
.Y(n_6055)
);

AND2x2_ASAP7_75t_L g6056 ( 
.A(n_5797),
.B(n_337),
.Y(n_6056)
);

HB1xp67_ASAP7_75t_L g6057 ( 
.A(n_5838),
.Y(n_6057)
);

INVx1_ASAP7_75t_L g6058 ( 
.A(n_5811),
.Y(n_6058)
);

INVx1_ASAP7_75t_L g6059 ( 
.A(n_5770),
.Y(n_6059)
);

OR2x2_ASAP7_75t_L g6060 ( 
.A(n_5745),
.B(n_337),
.Y(n_6060)
);

OR2x2_ASAP7_75t_L g6061 ( 
.A(n_5677),
.B(n_338),
.Y(n_6061)
);

INVx1_ASAP7_75t_L g6062 ( 
.A(n_5777),
.Y(n_6062)
);

AND2x2_ASAP7_75t_L g6063 ( 
.A(n_5738),
.B(n_338),
.Y(n_6063)
);

INVx1_ASAP7_75t_L g6064 ( 
.A(n_5674),
.Y(n_6064)
);

INVx2_ASAP7_75t_L g6065 ( 
.A(n_5827),
.Y(n_6065)
);

OR2x2_ASAP7_75t_L g6066 ( 
.A(n_5678),
.B(n_339),
.Y(n_6066)
);

INVx2_ASAP7_75t_L g6067 ( 
.A(n_5827),
.Y(n_6067)
);

INVx1_ASAP7_75t_L g6068 ( 
.A(n_5674),
.Y(n_6068)
);

INVx4_ASAP7_75t_L g6069 ( 
.A(n_5855),
.Y(n_6069)
);

INVx2_ASAP7_75t_L g6070 ( 
.A(n_5827),
.Y(n_6070)
);

AND2x2_ASAP7_75t_L g6071 ( 
.A(n_5738),
.B(n_340),
.Y(n_6071)
);

AND2x4_ASAP7_75t_L g6072 ( 
.A(n_5738),
.B(n_341),
.Y(n_6072)
);

BUFx3_ASAP7_75t_L g6073 ( 
.A(n_5679),
.Y(n_6073)
);

BUFx3_ASAP7_75t_L g6074 ( 
.A(n_5679),
.Y(n_6074)
);

INVx1_ASAP7_75t_L g6075 ( 
.A(n_5674),
.Y(n_6075)
);

AND2x2_ASAP7_75t_L g6076 ( 
.A(n_5738),
.B(n_341),
.Y(n_6076)
);

NAND2xp5_ASAP7_75t_L g6077 ( 
.A(n_5807),
.B(n_342),
.Y(n_6077)
);

NAND2xp5_ASAP7_75t_L g6078 ( 
.A(n_5807),
.B(n_342),
.Y(n_6078)
);

NAND2xp5_ASAP7_75t_L g6079 ( 
.A(n_5807),
.B(n_344),
.Y(n_6079)
);

INVx1_ASAP7_75t_L g6080 ( 
.A(n_5674),
.Y(n_6080)
);

AND2x2_ASAP7_75t_L g6081 ( 
.A(n_5738),
.B(n_345),
.Y(n_6081)
);

NAND2xp5_ASAP7_75t_L g6082 ( 
.A(n_5807),
.B(n_345),
.Y(n_6082)
);

INVx1_ASAP7_75t_L g6083 ( 
.A(n_5674),
.Y(n_6083)
);

INVx3_ASAP7_75t_L g6084 ( 
.A(n_5690),
.Y(n_6084)
);

INVx2_ASAP7_75t_L g6085 ( 
.A(n_5827),
.Y(n_6085)
);

AND2x2_ASAP7_75t_L g6086 ( 
.A(n_5738),
.B(n_346),
.Y(n_6086)
);

AND2x4_ASAP7_75t_SL g6087 ( 
.A(n_5855),
.B(n_346),
.Y(n_6087)
);

AND2x4_ASAP7_75t_L g6088 ( 
.A(n_5738),
.B(n_347),
.Y(n_6088)
);

AND2x2_ASAP7_75t_L g6089 ( 
.A(n_5738),
.B(n_347),
.Y(n_6089)
);

AND2x2_ASAP7_75t_L g6090 ( 
.A(n_5738),
.B(n_348),
.Y(n_6090)
);

INVx1_ASAP7_75t_L g6091 ( 
.A(n_5674),
.Y(n_6091)
);

INVx2_ASAP7_75t_L g6092 ( 
.A(n_5827),
.Y(n_6092)
);

INVx2_ASAP7_75t_L g6093 ( 
.A(n_5827),
.Y(n_6093)
);

AND2x2_ASAP7_75t_L g6094 ( 
.A(n_5738),
.B(n_348),
.Y(n_6094)
);

AND2x2_ASAP7_75t_L g6095 ( 
.A(n_5738),
.B(n_350),
.Y(n_6095)
);

AND2x2_ASAP7_75t_L g6096 ( 
.A(n_5738),
.B(n_350),
.Y(n_6096)
);

AOI22xp33_ASAP7_75t_L g6097 ( 
.A1(n_5840),
.A2(n_353),
.B1(n_351),
.B2(n_352),
.Y(n_6097)
);

AOI22xp5_ASAP7_75t_L g6098 ( 
.A1(n_5697),
.A2(n_354),
.B1(n_352),
.B2(n_353),
.Y(n_6098)
);

AND2x2_ASAP7_75t_L g6099 ( 
.A(n_5738),
.B(n_355),
.Y(n_6099)
);

AND2x2_ASAP7_75t_L g6100 ( 
.A(n_5738),
.B(n_355),
.Y(n_6100)
);

AND2x2_ASAP7_75t_L g6101 ( 
.A(n_5738),
.B(n_356),
.Y(n_6101)
);

NAND2xp5_ASAP7_75t_L g6102 ( 
.A(n_5807),
.B(n_356),
.Y(n_6102)
);

INVx2_ASAP7_75t_L g6103 ( 
.A(n_5827),
.Y(n_6103)
);

INVx2_ASAP7_75t_SL g6104 ( 
.A(n_5675),
.Y(n_6104)
);

INVx1_ASAP7_75t_L g6105 ( 
.A(n_5674),
.Y(n_6105)
);

INVx1_ASAP7_75t_SL g6106 ( 
.A(n_5681),
.Y(n_6106)
);

INVxp67_ASAP7_75t_SL g6107 ( 
.A(n_5819),
.Y(n_6107)
);

NAND2xp5_ASAP7_75t_L g6108 ( 
.A(n_5807),
.B(n_357),
.Y(n_6108)
);

AND2x2_ASAP7_75t_L g6109 ( 
.A(n_5738),
.B(n_357),
.Y(n_6109)
);

INVx2_ASAP7_75t_L g6110 ( 
.A(n_5827),
.Y(n_6110)
);

INVx2_ASAP7_75t_SL g6111 ( 
.A(n_5675),
.Y(n_6111)
);

OR2x2_ASAP7_75t_L g6112 ( 
.A(n_5678),
.B(n_360),
.Y(n_6112)
);

INVx2_ASAP7_75t_L g6113 ( 
.A(n_5827),
.Y(n_6113)
);

AND2x2_ASAP7_75t_L g6114 ( 
.A(n_5738),
.B(n_360),
.Y(n_6114)
);

AND2x2_ASAP7_75t_L g6115 ( 
.A(n_5738),
.B(n_361),
.Y(n_6115)
);

AND2x2_ASAP7_75t_L g6116 ( 
.A(n_5738),
.B(n_362),
.Y(n_6116)
);

INVx1_ASAP7_75t_SL g6117 ( 
.A(n_5681),
.Y(n_6117)
);

INVx2_ASAP7_75t_L g6118 ( 
.A(n_5827),
.Y(n_6118)
);

INVx1_ASAP7_75t_L g6119 ( 
.A(n_5674),
.Y(n_6119)
);

INVx1_ASAP7_75t_L g6120 ( 
.A(n_5674),
.Y(n_6120)
);

INVx1_ASAP7_75t_L g6121 ( 
.A(n_5674),
.Y(n_6121)
);

INVx1_ASAP7_75t_L g6122 ( 
.A(n_5674),
.Y(n_6122)
);

INVx2_ASAP7_75t_L g6123 ( 
.A(n_5827),
.Y(n_6123)
);

INVx2_ASAP7_75t_L g6124 ( 
.A(n_5827),
.Y(n_6124)
);

BUFx2_ASAP7_75t_L g6125 ( 
.A(n_5738),
.Y(n_6125)
);

BUFx3_ASAP7_75t_L g6126 ( 
.A(n_5679),
.Y(n_6126)
);

AND2x2_ASAP7_75t_L g6127 ( 
.A(n_6125),
.B(n_363),
.Y(n_6127)
);

INVx1_ASAP7_75t_L g6128 ( 
.A(n_5931),
.Y(n_6128)
);

AND2x2_ASAP7_75t_L g6129 ( 
.A(n_5886),
.B(n_363),
.Y(n_6129)
);

INVx2_ASAP7_75t_L g6130 ( 
.A(n_5944),
.Y(n_6130)
);

INVx2_ASAP7_75t_L g6131 ( 
.A(n_6084),
.Y(n_6131)
);

OAI22xp5_ASAP7_75t_L g6132 ( 
.A1(n_6054),
.A2(n_366),
.B1(n_364),
.B2(n_365),
.Y(n_6132)
);

INVx4_ASAP7_75t_L g6133 ( 
.A(n_5900),
.Y(n_6133)
);

INVx2_ASAP7_75t_L g6134 ( 
.A(n_5900),
.Y(n_6134)
);

INVx2_ASAP7_75t_SL g6135 ( 
.A(n_5882),
.Y(n_6135)
);

INVx2_ASAP7_75t_L g6136 ( 
.A(n_6069),
.Y(n_6136)
);

OAI221xp5_ASAP7_75t_L g6137 ( 
.A1(n_6055),
.A2(n_366),
.B1(n_364),
.B2(n_365),
.C(n_367),
.Y(n_6137)
);

AND2x2_ASAP7_75t_L g6138 ( 
.A(n_5992),
.B(n_368),
.Y(n_6138)
);

INVx1_ASAP7_75t_L g6139 ( 
.A(n_5942),
.Y(n_6139)
);

INVx1_ASAP7_75t_L g6140 ( 
.A(n_5867),
.Y(n_6140)
);

INVx1_ASAP7_75t_L g6141 ( 
.A(n_5873),
.Y(n_6141)
);

AO21x2_ASAP7_75t_L g6142 ( 
.A1(n_5878),
.A2(n_368),
.B(n_369),
.Y(n_6142)
);

BUFx2_ASAP7_75t_L g6143 ( 
.A(n_5978),
.Y(n_6143)
);

OAI22xp5_ASAP7_75t_L g6144 ( 
.A1(n_6098),
.A2(n_374),
.B1(n_369),
.B2(n_373),
.Y(n_6144)
);

AO21x2_ASAP7_75t_L g6145 ( 
.A1(n_6107),
.A2(n_373),
.B(n_375),
.Y(n_6145)
);

AOI211xp5_ASAP7_75t_SL g6146 ( 
.A1(n_6041),
.A2(n_378),
.B(n_376),
.C(n_377),
.Y(n_6146)
);

AND2x4_ASAP7_75t_L g6147 ( 
.A(n_5870),
.B(n_5879),
.Y(n_6147)
);

BUFx2_ASAP7_75t_L g6148 ( 
.A(n_6010),
.Y(n_6148)
);

BUFx3_ASAP7_75t_L g6149 ( 
.A(n_5899),
.Y(n_6149)
);

AND2x2_ASAP7_75t_L g6150 ( 
.A(n_6049),
.B(n_376),
.Y(n_6150)
);

AO21x2_ASAP7_75t_L g6151 ( 
.A1(n_6019),
.A2(n_377),
.B(n_378),
.Y(n_6151)
);

INVx1_ASAP7_75t_L g6152 ( 
.A(n_5875),
.Y(n_6152)
);

INVxp67_ASAP7_75t_L g6153 ( 
.A(n_6057),
.Y(n_6153)
);

OAI31xp33_ASAP7_75t_L g6154 ( 
.A1(n_6053),
.A2(n_381),
.A3(n_379),
.B(n_380),
.Y(n_6154)
);

INVx2_ASAP7_75t_L g6155 ( 
.A(n_6065),
.Y(n_6155)
);

HB1xp67_ASAP7_75t_L g6156 ( 
.A(n_5891),
.Y(n_6156)
);

INVx2_ASAP7_75t_L g6157 ( 
.A(n_6067),
.Y(n_6157)
);

INVx1_ASAP7_75t_L g6158 ( 
.A(n_5876),
.Y(n_6158)
);

AOI22xp5_ASAP7_75t_L g6159 ( 
.A1(n_6062),
.A2(n_383),
.B1(n_380),
.B2(n_382),
.Y(n_6159)
);

INVx2_ASAP7_75t_L g6160 ( 
.A(n_6070),
.Y(n_6160)
);

AOI22xp33_ASAP7_75t_L g6161 ( 
.A1(n_6058),
.A2(n_385),
.B1(n_382),
.B2(n_384),
.Y(n_6161)
);

INVx1_ASAP7_75t_L g6162 ( 
.A(n_5890),
.Y(n_6162)
);

INVx2_ASAP7_75t_L g6163 ( 
.A(n_6085),
.Y(n_6163)
);

INVx2_ASAP7_75t_L g6164 ( 
.A(n_6092),
.Y(n_6164)
);

OA21x2_ASAP7_75t_L g6165 ( 
.A1(n_6016),
.A2(n_384),
.B(n_385),
.Y(n_6165)
);

INVx2_ASAP7_75t_L g6166 ( 
.A(n_6093),
.Y(n_6166)
);

INVx1_ASAP7_75t_L g6167 ( 
.A(n_5903),
.Y(n_6167)
);

OAI21x1_ASAP7_75t_L g6168 ( 
.A1(n_6005),
.A2(n_386),
.B(n_387),
.Y(n_6168)
);

INVx2_ASAP7_75t_SL g6169 ( 
.A(n_6073),
.Y(n_6169)
);

NOR2xp33_ASAP7_75t_SL g6170 ( 
.A(n_6106),
.B(n_386),
.Y(n_6170)
);

AOI22xp33_ASAP7_75t_L g6171 ( 
.A1(n_6059),
.A2(n_389),
.B1(n_387),
.B2(n_388),
.Y(n_6171)
);

INVx1_ASAP7_75t_L g6172 ( 
.A(n_5907),
.Y(n_6172)
);

NAND2xp5_ASAP7_75t_SL g6173 ( 
.A(n_5909),
.B(n_6117),
.Y(n_6173)
);

NAND2xp5_ASAP7_75t_L g6174 ( 
.A(n_6039),
.B(n_390),
.Y(n_6174)
);

AOI22xp33_ASAP7_75t_L g6175 ( 
.A1(n_5901),
.A2(n_393),
.B1(n_391),
.B2(n_392),
.Y(n_6175)
);

OAI21xp33_ASAP7_75t_L g6176 ( 
.A1(n_6001),
.A2(n_391),
.B(n_393),
.Y(n_6176)
);

INVx1_ASAP7_75t_L g6177 ( 
.A(n_5912),
.Y(n_6177)
);

INVx1_ASAP7_75t_L g6178 ( 
.A(n_5916),
.Y(n_6178)
);

INVx1_ASAP7_75t_L g6179 ( 
.A(n_5917),
.Y(n_6179)
);

INVx1_ASAP7_75t_L g6180 ( 
.A(n_5921),
.Y(n_6180)
);

INVxp67_ASAP7_75t_SL g6181 ( 
.A(n_6002),
.Y(n_6181)
);

NOR2xp33_ASAP7_75t_L g6182 ( 
.A(n_6104),
.B(n_394),
.Y(n_6182)
);

AND2x2_ASAP7_75t_L g6183 ( 
.A(n_5887),
.B(n_394),
.Y(n_6183)
);

AOI22xp33_ASAP7_75t_L g6184 ( 
.A1(n_5964),
.A2(n_397),
.B1(n_395),
.B2(n_396),
.Y(n_6184)
);

INVx1_ASAP7_75t_L g6185 ( 
.A(n_5923),
.Y(n_6185)
);

INVx2_ASAP7_75t_L g6186 ( 
.A(n_6103),
.Y(n_6186)
);

OAI22xp5_ASAP7_75t_L g6187 ( 
.A1(n_6110),
.A2(n_6113),
.B1(n_6123),
.B2(n_6118),
.Y(n_6187)
);

INVx1_ASAP7_75t_SL g6188 ( 
.A(n_5986),
.Y(n_6188)
);

INVx1_ASAP7_75t_L g6189 ( 
.A(n_5927),
.Y(n_6189)
);

INVx1_ASAP7_75t_L g6190 ( 
.A(n_5929),
.Y(n_6190)
);

INVx1_ASAP7_75t_L g6191 ( 
.A(n_5957),
.Y(n_6191)
);

INVx1_ASAP7_75t_L g6192 ( 
.A(n_5962),
.Y(n_6192)
);

HB1xp67_ASAP7_75t_L g6193 ( 
.A(n_5915),
.Y(n_6193)
);

AOI22xp33_ASAP7_75t_L g6194 ( 
.A1(n_5964),
.A2(n_398),
.B1(n_395),
.B2(n_397),
.Y(n_6194)
);

INVx2_ASAP7_75t_SL g6195 ( 
.A(n_6074),
.Y(n_6195)
);

INVx1_ASAP7_75t_L g6196 ( 
.A(n_5968),
.Y(n_6196)
);

INVx2_ASAP7_75t_L g6197 ( 
.A(n_6124),
.Y(n_6197)
);

OAI221xp5_ASAP7_75t_L g6198 ( 
.A1(n_6061),
.A2(n_401),
.B1(n_399),
.B2(n_400),
.C(n_402),
.Y(n_6198)
);

AOI221xp5_ASAP7_75t_L g6199 ( 
.A1(n_5970),
.A2(n_401),
.B1(n_399),
.B2(n_400),
.C(n_404),
.Y(n_6199)
);

OAI21x1_ASAP7_75t_L g6200 ( 
.A1(n_5946),
.A2(n_404),
.B(n_405),
.Y(n_6200)
);

OA21x2_ASAP7_75t_L g6201 ( 
.A1(n_5998),
.A2(n_406),
.B(n_407),
.Y(n_6201)
);

NAND2xp5_ASAP7_75t_L g6202 ( 
.A(n_6045),
.B(n_406),
.Y(n_6202)
);

AOI22xp5_ASAP7_75t_L g6203 ( 
.A1(n_6008),
.A2(n_409),
.B1(n_407),
.B2(n_408),
.Y(n_6203)
);

INVx2_ASAP7_75t_L g6204 ( 
.A(n_6111),
.Y(n_6204)
);

INVxp67_ASAP7_75t_SL g6205 ( 
.A(n_6017),
.Y(n_6205)
);

OA21x2_ASAP7_75t_L g6206 ( 
.A1(n_5975),
.A2(n_410),
.B(n_411),
.Y(n_6206)
);

OR2x2_ASAP7_75t_L g6207 ( 
.A(n_5881),
.B(n_410),
.Y(n_6207)
);

INVx1_ASAP7_75t_L g6208 ( 
.A(n_5988),
.Y(n_6208)
);

AOI211x1_ASAP7_75t_L g6209 ( 
.A1(n_6014),
.A2(n_414),
.B(n_412),
.C(n_413),
.Y(n_6209)
);

INVxp67_ASAP7_75t_SL g6210 ( 
.A(n_5919),
.Y(n_6210)
);

AND2x2_ASAP7_75t_L g6211 ( 
.A(n_5938),
.B(n_412),
.Y(n_6211)
);

NAND2xp5_ASAP7_75t_SL g6212 ( 
.A(n_6126),
.B(n_413),
.Y(n_6212)
);

INVx2_ASAP7_75t_L g6213 ( 
.A(n_5981),
.Y(n_6213)
);

INVx2_ASAP7_75t_SL g6214 ( 
.A(n_5971),
.Y(n_6214)
);

AOI22xp5_ASAP7_75t_L g6215 ( 
.A1(n_5949),
.A2(n_416),
.B1(n_414),
.B2(n_415),
.Y(n_6215)
);

AOI33xp33_ASAP7_75t_L g6216 ( 
.A1(n_6097),
.A2(n_418),
.A3(n_420),
.B1(n_415),
.B2(n_417),
.B3(n_419),
.Y(n_6216)
);

INVx1_ASAP7_75t_L g6217 ( 
.A(n_6064),
.Y(n_6217)
);

INVx2_ASAP7_75t_SL g6218 ( 
.A(n_6037),
.Y(n_6218)
);

OAI21xp5_ASAP7_75t_L g6219 ( 
.A1(n_6047),
.A2(n_417),
.B(n_418),
.Y(n_6219)
);

INVxp67_ASAP7_75t_SL g6220 ( 
.A(n_5948),
.Y(n_6220)
);

OAI21xp5_ASAP7_75t_L g6221 ( 
.A1(n_5976),
.A2(n_420),
.B(n_421),
.Y(n_6221)
);

INVxp67_ASAP7_75t_SL g6222 ( 
.A(n_6007),
.Y(n_6222)
);

INVx1_ASAP7_75t_L g6223 ( 
.A(n_6068),
.Y(n_6223)
);

OAI21x1_ASAP7_75t_L g6224 ( 
.A1(n_5994),
.A2(n_421),
.B(n_422),
.Y(n_6224)
);

INVx2_ASAP7_75t_L g6225 ( 
.A(n_6027),
.Y(n_6225)
);

AND2x2_ASAP7_75t_L g6226 ( 
.A(n_6006),
.B(n_423),
.Y(n_6226)
);

INVx1_ASAP7_75t_L g6227 ( 
.A(n_6075),
.Y(n_6227)
);

INVx2_ASAP7_75t_L g6228 ( 
.A(n_6040),
.Y(n_6228)
);

INVx2_ASAP7_75t_L g6229 ( 
.A(n_6011),
.Y(n_6229)
);

AND2x2_ASAP7_75t_L g6230 ( 
.A(n_6025),
.B(n_423),
.Y(n_6230)
);

INVx1_ASAP7_75t_L g6231 ( 
.A(n_6080),
.Y(n_6231)
);

NAND4xp25_ASAP7_75t_L g6232 ( 
.A(n_5868),
.B(n_426),
.C(n_427),
.D(n_425),
.Y(n_6232)
);

OR2x2_ASAP7_75t_L g6233 ( 
.A(n_6009),
.B(n_424),
.Y(n_6233)
);

NAND4xp25_ASAP7_75t_L g6234 ( 
.A(n_6012),
.B(n_429),
.C(n_430),
.D(n_425),
.Y(n_6234)
);

NAND3xp33_ASAP7_75t_L g6235 ( 
.A(n_5996),
.B(n_6077),
.C(n_5872),
.Y(n_6235)
);

OAI221xp5_ASAP7_75t_L g6236 ( 
.A1(n_6060),
.A2(n_430),
.B1(n_424),
.B2(n_429),
.C(n_431),
.Y(n_6236)
);

OR2x2_ASAP7_75t_L g6237 ( 
.A(n_6013),
.B(n_431),
.Y(n_6237)
);

NAND2xp5_ASAP7_75t_L g6238 ( 
.A(n_6042),
.B(n_6018),
.Y(n_6238)
);

INVx1_ASAP7_75t_L g6239 ( 
.A(n_6083),
.Y(n_6239)
);

AND2x4_ASAP7_75t_L g6240 ( 
.A(n_6072),
.B(n_432),
.Y(n_6240)
);

AO31x2_ASAP7_75t_L g6241 ( 
.A1(n_6078),
.A2(n_435),
.A3(n_433),
.B(n_434),
.Y(n_6241)
);

AO21x2_ASAP7_75t_L g6242 ( 
.A1(n_6079),
.A2(n_436),
.B(n_437),
.Y(n_6242)
);

BUFx3_ASAP7_75t_L g6243 ( 
.A(n_6088),
.Y(n_6243)
);

INVx3_ASAP7_75t_L g6244 ( 
.A(n_5943),
.Y(n_6244)
);

AO21x2_ASAP7_75t_L g6245 ( 
.A1(n_6082),
.A2(n_436),
.B(n_438),
.Y(n_6245)
);

INVx2_ASAP7_75t_L g6246 ( 
.A(n_6015),
.Y(n_6246)
);

AND2x2_ASAP7_75t_L g6247 ( 
.A(n_5869),
.B(n_439),
.Y(n_6247)
);

OAI22xp5_ASAP7_75t_L g6248 ( 
.A1(n_6029),
.A2(n_441),
.B1(n_439),
.B2(n_440),
.Y(n_6248)
);

AND2x2_ASAP7_75t_L g6249 ( 
.A(n_6063),
.B(n_442),
.Y(n_6249)
);

INVx2_ASAP7_75t_L g6250 ( 
.A(n_6050),
.Y(n_6250)
);

AND2x2_ASAP7_75t_L g6251 ( 
.A(n_6071),
.B(n_442),
.Y(n_6251)
);

INVxp67_ASAP7_75t_L g6252 ( 
.A(n_6076),
.Y(n_6252)
);

AOI221x1_ASAP7_75t_L g6253 ( 
.A1(n_6102),
.A2(n_445),
.B1(n_443),
.B2(n_444),
.C(n_446),
.Y(n_6253)
);

BUFx2_ASAP7_75t_L g6254 ( 
.A(n_6081),
.Y(n_6254)
);

INVx1_ASAP7_75t_L g6255 ( 
.A(n_6091),
.Y(n_6255)
);

AND2x2_ASAP7_75t_L g6256 ( 
.A(n_6086),
.B(n_445),
.Y(n_6256)
);

OR2x2_ASAP7_75t_L g6257 ( 
.A(n_5947),
.B(n_446),
.Y(n_6257)
);

INVx2_ASAP7_75t_SL g6258 ( 
.A(n_5871),
.Y(n_6258)
);

AND2x2_ASAP7_75t_L g6259 ( 
.A(n_6089),
.B(n_447),
.Y(n_6259)
);

AOI22xp33_ASAP7_75t_L g6260 ( 
.A1(n_6020),
.A2(n_6056),
.B1(n_6024),
.B2(n_6030),
.Y(n_6260)
);

INVx2_ASAP7_75t_L g6261 ( 
.A(n_5883),
.Y(n_6261)
);

BUFx2_ASAP7_75t_L g6262 ( 
.A(n_6090),
.Y(n_6262)
);

OA21x2_ASAP7_75t_L g6263 ( 
.A1(n_6105),
.A2(n_449),
.B(n_451),
.Y(n_6263)
);

INVx1_ASAP7_75t_L g6264 ( 
.A(n_6119),
.Y(n_6264)
);

AND2x2_ASAP7_75t_L g6265 ( 
.A(n_6094),
.B(n_6095),
.Y(n_6265)
);

AOI22xp33_ASAP7_75t_L g6266 ( 
.A1(n_6035),
.A2(n_453),
.B1(n_451),
.B2(n_452),
.Y(n_6266)
);

OAI33xp33_ASAP7_75t_L g6267 ( 
.A1(n_6108),
.A2(n_455),
.A3(n_457),
.B1(n_453),
.B2(n_454),
.B3(n_456),
.Y(n_6267)
);

NAND3xp33_ASAP7_75t_L g6268 ( 
.A(n_5893),
.B(n_454),
.C(n_455),
.Y(n_6268)
);

INVx1_ASAP7_75t_L g6269 ( 
.A(n_6120),
.Y(n_6269)
);

INVx2_ASAP7_75t_SL g6270 ( 
.A(n_5932),
.Y(n_6270)
);

BUFx3_ASAP7_75t_L g6271 ( 
.A(n_5892),
.Y(n_6271)
);

NAND4xp25_ASAP7_75t_L g6272 ( 
.A(n_6052),
.B(n_461),
.C(n_462),
.D(n_459),
.Y(n_6272)
);

INVx2_ASAP7_75t_L g6273 ( 
.A(n_5896),
.Y(n_6273)
);

AOI21xp5_ASAP7_75t_L g6274 ( 
.A1(n_5961),
.A2(n_458),
.B(n_459),
.Y(n_6274)
);

INVx2_ASAP7_75t_L g6275 ( 
.A(n_5897),
.Y(n_6275)
);

INVx1_ASAP7_75t_SL g6276 ( 
.A(n_6004),
.Y(n_6276)
);

BUFx2_ASAP7_75t_L g6277 ( 
.A(n_6096),
.Y(n_6277)
);

INVx2_ASAP7_75t_L g6278 ( 
.A(n_5911),
.Y(n_6278)
);

INVx1_ASAP7_75t_L g6279 ( 
.A(n_6121),
.Y(n_6279)
);

INVx2_ASAP7_75t_L g6280 ( 
.A(n_5920),
.Y(n_6280)
);

INVx1_ASAP7_75t_L g6281 ( 
.A(n_6122),
.Y(n_6281)
);

AND2x2_ASAP7_75t_L g6282 ( 
.A(n_6099),
.B(n_458),
.Y(n_6282)
);

INVx2_ASAP7_75t_L g6283 ( 
.A(n_5926),
.Y(n_6283)
);

OR2x6_ASAP7_75t_L g6284 ( 
.A(n_6100),
.B(n_6101),
.Y(n_6284)
);

AOI21xp33_ASAP7_75t_L g6285 ( 
.A1(n_6023),
.A2(n_462),
.B(n_463),
.Y(n_6285)
);

BUFx3_ASAP7_75t_L g6286 ( 
.A(n_5904),
.Y(n_6286)
);

INVx2_ASAP7_75t_L g6287 ( 
.A(n_5935),
.Y(n_6287)
);

INVx1_ASAP7_75t_L g6288 ( 
.A(n_5974),
.Y(n_6288)
);

INVx2_ASAP7_75t_L g6289 ( 
.A(n_5936),
.Y(n_6289)
);

INVx2_ASAP7_75t_L g6290 ( 
.A(n_5945),
.Y(n_6290)
);

OAI33xp33_ASAP7_75t_L g6291 ( 
.A1(n_5937),
.A2(n_465),
.A3(n_467),
.B1(n_463),
.B2(n_464),
.B3(n_466),
.Y(n_6291)
);

HB1xp67_ASAP7_75t_L g6292 ( 
.A(n_5950),
.Y(n_6292)
);

AOI21xp33_ASAP7_75t_L g6293 ( 
.A1(n_5884),
.A2(n_464),
.B(n_465),
.Y(n_6293)
);

INVx1_ASAP7_75t_L g6294 ( 
.A(n_5953),
.Y(n_6294)
);

INVx1_ASAP7_75t_L g6295 ( 
.A(n_5954),
.Y(n_6295)
);

NAND2xp5_ASAP7_75t_L g6296 ( 
.A(n_6109),
.B(n_468),
.Y(n_6296)
);

AOI22xp33_ASAP7_75t_L g6297 ( 
.A1(n_5959),
.A2(n_471),
.B1(n_469),
.B2(n_470),
.Y(n_6297)
);

OAI211xp5_ASAP7_75t_L g6298 ( 
.A1(n_5939),
.A2(n_473),
.B(n_470),
.C(n_472),
.Y(n_6298)
);

BUFx2_ASAP7_75t_L g6299 ( 
.A(n_6114),
.Y(n_6299)
);

INVx1_ASAP7_75t_L g6300 ( 
.A(n_5963),
.Y(n_6300)
);

OAI31xp33_ASAP7_75t_L g6301 ( 
.A1(n_6115),
.A2(n_475),
.A3(n_473),
.B(n_474),
.Y(n_6301)
);

INVx1_ASAP7_75t_SL g6302 ( 
.A(n_6028),
.Y(n_6302)
);

BUFx3_ASAP7_75t_L g6303 ( 
.A(n_5889),
.Y(n_6303)
);

INVx1_ASAP7_75t_SL g6304 ( 
.A(n_5955),
.Y(n_6304)
);

INVx1_ASAP7_75t_L g6305 ( 
.A(n_5980),
.Y(n_6305)
);

INVx1_ASAP7_75t_L g6306 ( 
.A(n_5989),
.Y(n_6306)
);

INVx2_ASAP7_75t_L g6307 ( 
.A(n_5905),
.Y(n_6307)
);

BUFx6f_ASAP7_75t_L g6308 ( 
.A(n_5941),
.Y(n_6308)
);

OAI33xp33_ASAP7_75t_L g6309 ( 
.A1(n_5940),
.A2(n_477),
.A3(n_480),
.B1(n_474),
.B2(n_476),
.B3(n_479),
.Y(n_6309)
);

AND2x2_ASAP7_75t_L g6310 ( 
.A(n_6116),
.B(n_476),
.Y(n_6310)
);

INVx1_ASAP7_75t_L g6311 ( 
.A(n_5990),
.Y(n_6311)
);

NOR2x1_ASAP7_75t_L g6312 ( 
.A(n_5880),
.B(n_477),
.Y(n_6312)
);

OAI222xp33_ASAP7_75t_L g6313 ( 
.A1(n_5969),
.A2(n_481),
.B1(n_483),
.B2(n_484),
.C1(n_480),
.C2(n_482),
.Y(n_6313)
);

INVx1_ASAP7_75t_L g6314 ( 
.A(n_6222),
.Y(n_6314)
);

INVx1_ASAP7_75t_L g6315 ( 
.A(n_6156),
.Y(n_6315)
);

AND2x2_ASAP7_75t_L g6316 ( 
.A(n_6188),
.B(n_6135),
.Y(n_6316)
);

INVx1_ASAP7_75t_L g6317 ( 
.A(n_6193),
.Y(n_6317)
);

AND2x2_ASAP7_75t_L g6318 ( 
.A(n_6130),
.B(n_6043),
.Y(n_6318)
);

AND2x4_ASAP7_75t_L g6319 ( 
.A(n_6133),
.B(n_6134),
.Y(n_6319)
);

AND2x2_ASAP7_75t_L g6320 ( 
.A(n_6131),
.B(n_6051),
.Y(n_6320)
);

INVxp67_ASAP7_75t_SL g6321 ( 
.A(n_6173),
.Y(n_6321)
);

OR2x2_ASAP7_75t_L g6322 ( 
.A(n_6276),
.B(n_5951),
.Y(n_6322)
);

AND2x4_ASAP7_75t_L g6323 ( 
.A(n_6169),
.B(n_5874),
.Y(n_6323)
);

NAND2xp5_ASAP7_75t_L g6324 ( 
.A(n_6205),
.B(n_5894),
.Y(n_6324)
);

OR2x2_ASAP7_75t_L g6325 ( 
.A(n_6302),
.B(n_5958),
.Y(n_6325)
);

NAND2xp5_ASAP7_75t_L g6326 ( 
.A(n_6148),
.B(n_5895),
.Y(n_6326)
);

INVx1_ASAP7_75t_L g6327 ( 
.A(n_6220),
.Y(n_6327)
);

INVx1_ASAP7_75t_L g6328 ( 
.A(n_6210),
.Y(n_6328)
);

INVx1_ASAP7_75t_L g6329 ( 
.A(n_6181),
.Y(n_6329)
);

INVx4_ASAP7_75t_L g6330 ( 
.A(n_6149),
.Y(n_6330)
);

BUFx2_ASAP7_75t_SL g6331 ( 
.A(n_6195),
.Y(n_6331)
);

NAND2xp5_ASAP7_75t_L g6332 ( 
.A(n_6258),
.B(n_5898),
.Y(n_6332)
);

INVx1_ASAP7_75t_L g6333 ( 
.A(n_6311),
.Y(n_6333)
);

AND2x2_ASAP7_75t_L g6334 ( 
.A(n_6143),
.B(n_5925),
.Y(n_6334)
);

OR2x2_ASAP7_75t_L g6335 ( 
.A(n_6307),
.B(n_5960),
.Y(n_6335)
);

INVx2_ASAP7_75t_L g6336 ( 
.A(n_6243),
.Y(n_6336)
);

INVx1_ASAP7_75t_L g6337 ( 
.A(n_6140),
.Y(n_6337)
);

INVx1_ASAP7_75t_L g6338 ( 
.A(n_6141),
.Y(n_6338)
);

INVx2_ASAP7_75t_L g6339 ( 
.A(n_6308),
.Y(n_6339)
);

INVx1_ASAP7_75t_L g6340 ( 
.A(n_6152),
.Y(n_6340)
);

INVx1_ASAP7_75t_L g6341 ( 
.A(n_6158),
.Y(n_6341)
);

INVx1_ASAP7_75t_L g6342 ( 
.A(n_6162),
.Y(n_6342)
);

AND2x4_ASAP7_75t_SL g6343 ( 
.A(n_6308),
.B(n_6244),
.Y(n_6343)
);

INVx1_ASAP7_75t_L g6344 ( 
.A(n_6167),
.Y(n_6344)
);

NAND2xp5_ASAP7_75t_L g6345 ( 
.A(n_6254),
.B(n_5993),
.Y(n_6345)
);

OR2x2_ASAP7_75t_L g6346 ( 
.A(n_6153),
.B(n_6238),
.Y(n_6346)
);

AND2x4_ASAP7_75t_SL g6347 ( 
.A(n_6136),
.B(n_5965),
.Y(n_6347)
);

INVx1_ASAP7_75t_L g6348 ( 
.A(n_6172),
.Y(n_6348)
);

INVx1_ASAP7_75t_L g6349 ( 
.A(n_6177),
.Y(n_6349)
);

INVx2_ASAP7_75t_SL g6350 ( 
.A(n_6271),
.Y(n_6350)
);

INVx1_ASAP7_75t_L g6351 ( 
.A(n_6178),
.Y(n_6351)
);

HB1xp67_ASAP7_75t_L g6352 ( 
.A(n_6262),
.Y(n_6352)
);

INVx1_ASAP7_75t_L g6353 ( 
.A(n_6179),
.Y(n_6353)
);

AND2x2_ASAP7_75t_L g6354 ( 
.A(n_6218),
.B(n_5979),
.Y(n_6354)
);

HB1xp67_ASAP7_75t_L g6355 ( 
.A(n_6277),
.Y(n_6355)
);

NAND4xp25_ASAP7_75t_L g6356 ( 
.A(n_6146),
.B(n_6175),
.C(n_6260),
.D(n_6154),
.Y(n_6356)
);

NOR2x1p5_ASAP7_75t_L g6357 ( 
.A(n_6213),
.B(n_6034),
.Y(n_6357)
);

INVx1_ASAP7_75t_L g6358 ( 
.A(n_6180),
.Y(n_6358)
);

INVx1_ASAP7_75t_L g6359 ( 
.A(n_6185),
.Y(n_6359)
);

AND2x4_ASAP7_75t_L g6360 ( 
.A(n_6214),
.B(n_5913),
.Y(n_6360)
);

NOR2xp67_ASAP7_75t_L g6361 ( 
.A(n_6204),
.B(n_5885),
.Y(n_6361)
);

INVx2_ASAP7_75t_SL g6362 ( 
.A(n_6286),
.Y(n_6362)
);

INVx2_ASAP7_75t_L g6363 ( 
.A(n_6303),
.Y(n_6363)
);

AND2x2_ASAP7_75t_L g6364 ( 
.A(n_6299),
.B(n_5973),
.Y(n_6364)
);

INVx1_ASAP7_75t_L g6365 ( 
.A(n_6189),
.Y(n_6365)
);

NOR2x1_ASAP7_75t_L g6366 ( 
.A(n_6151),
.B(n_6066),
.Y(n_6366)
);

INVx1_ASAP7_75t_L g6367 ( 
.A(n_6190),
.Y(n_6367)
);

AND2x2_ASAP7_75t_L g6368 ( 
.A(n_6265),
.B(n_5877),
.Y(n_6368)
);

HB1xp67_ASAP7_75t_L g6369 ( 
.A(n_6165),
.Y(n_6369)
);

HB1xp67_ASAP7_75t_L g6370 ( 
.A(n_6206),
.Y(n_6370)
);

AND2x2_ASAP7_75t_L g6371 ( 
.A(n_6225),
.B(n_5888),
.Y(n_6371)
);

INVx2_ASAP7_75t_L g6372 ( 
.A(n_6270),
.Y(n_6372)
);

INVx1_ASAP7_75t_L g6373 ( 
.A(n_6191),
.Y(n_6373)
);

OR2x2_ASAP7_75t_L g6374 ( 
.A(n_6250),
.B(n_5922),
.Y(n_6374)
);

INVx1_ASAP7_75t_L g6375 ( 
.A(n_6192),
.Y(n_6375)
);

INVx2_ASAP7_75t_SL g6376 ( 
.A(n_6240),
.Y(n_6376)
);

AND2x2_ASAP7_75t_L g6377 ( 
.A(n_6252),
.B(n_5902),
.Y(n_6377)
);

AND2x2_ASAP7_75t_L g6378 ( 
.A(n_6147),
.B(n_5914),
.Y(n_6378)
);

INVx1_ASAP7_75t_L g6379 ( 
.A(n_6196),
.Y(n_6379)
);

INVx2_ASAP7_75t_SL g6380 ( 
.A(n_6284),
.Y(n_6380)
);

INVx2_ASAP7_75t_L g6381 ( 
.A(n_6284),
.Y(n_6381)
);

OR2x2_ASAP7_75t_L g6382 ( 
.A(n_6228),
.B(n_5966),
.Y(n_6382)
);

OR2x2_ASAP7_75t_L g6383 ( 
.A(n_6229),
.B(n_5967),
.Y(n_6383)
);

NAND2xp33_ASAP7_75t_SL g6384 ( 
.A(n_6142),
.B(n_6112),
.Y(n_6384)
);

AND2x2_ASAP7_75t_L g6385 ( 
.A(n_6155),
.B(n_5906),
.Y(n_6385)
);

INVx1_ASAP7_75t_L g6386 ( 
.A(n_6208),
.Y(n_6386)
);

INVx1_ASAP7_75t_L g6387 ( 
.A(n_6217),
.Y(n_6387)
);

NAND2x1_ASAP7_75t_L g6388 ( 
.A(n_6288),
.B(n_6031),
.Y(n_6388)
);

NAND2xp5_ASAP7_75t_L g6389 ( 
.A(n_6304),
.B(n_5910),
.Y(n_6389)
);

AND2x2_ASAP7_75t_L g6390 ( 
.A(n_6157),
.B(n_5908),
.Y(n_6390)
);

OR2x2_ASAP7_75t_L g6391 ( 
.A(n_6246),
.B(n_5928),
.Y(n_6391)
);

INVx2_ASAP7_75t_L g6392 ( 
.A(n_6257),
.Y(n_6392)
);

INVxp67_ASAP7_75t_L g6393 ( 
.A(n_6145),
.Y(n_6393)
);

INVx1_ASAP7_75t_L g6394 ( 
.A(n_6223),
.Y(n_6394)
);

NAND3xp33_ASAP7_75t_L g6395 ( 
.A(n_6253),
.B(n_5930),
.C(n_5995),
.Y(n_6395)
);

INVx1_ASAP7_75t_L g6396 ( 
.A(n_6227),
.Y(n_6396)
);

INVxp67_ASAP7_75t_SL g6397 ( 
.A(n_6312),
.Y(n_6397)
);

AND2x2_ASAP7_75t_L g6398 ( 
.A(n_6160),
.B(n_5997),
.Y(n_6398)
);

INVx4_ASAP7_75t_L g6399 ( 
.A(n_6129),
.Y(n_6399)
);

INVx3_ASAP7_75t_L g6400 ( 
.A(n_6163),
.Y(n_6400)
);

AND2x2_ASAP7_75t_L g6401 ( 
.A(n_6164),
.B(n_5999),
.Y(n_6401)
);

OR2x2_ASAP7_75t_L g6402 ( 
.A(n_6235),
.B(n_5952),
.Y(n_6402)
);

INVx1_ASAP7_75t_L g6403 ( 
.A(n_6231),
.Y(n_6403)
);

INVx1_ASAP7_75t_SL g6404 ( 
.A(n_6127),
.Y(n_6404)
);

INVx1_ASAP7_75t_L g6405 ( 
.A(n_6239),
.Y(n_6405)
);

NAND2xp5_ASAP7_75t_L g6406 ( 
.A(n_6242),
.B(n_5933),
.Y(n_6406)
);

AND2x2_ASAP7_75t_L g6407 ( 
.A(n_6166),
.B(n_6003),
.Y(n_6407)
);

AND2x2_ASAP7_75t_L g6408 ( 
.A(n_6186),
.B(n_6026),
.Y(n_6408)
);

NAND2xp5_ASAP7_75t_L g6409 ( 
.A(n_6245),
.B(n_5934),
.Y(n_6409)
);

AND2x2_ASAP7_75t_L g6410 ( 
.A(n_6197),
.B(n_5924),
.Y(n_6410)
);

AND2x2_ASAP7_75t_L g6411 ( 
.A(n_6138),
.B(n_6046),
.Y(n_6411)
);

AND2x4_ASAP7_75t_L g6412 ( 
.A(n_6183),
.B(n_6226),
.Y(n_6412)
);

INVx1_ASAP7_75t_SL g6413 ( 
.A(n_6150),
.Y(n_6413)
);

INVx1_ASAP7_75t_L g6414 ( 
.A(n_6255),
.Y(n_6414)
);

INVx1_ASAP7_75t_L g6415 ( 
.A(n_6264),
.Y(n_6415)
);

OR2x2_ASAP7_75t_L g6416 ( 
.A(n_6261),
.B(n_6000),
.Y(n_6416)
);

NAND2xp5_ASAP7_75t_L g6417 ( 
.A(n_6274),
.B(n_5982),
.Y(n_6417)
);

NOR2x1_ASAP7_75t_L g6418 ( 
.A(n_6201),
.B(n_6263),
.Y(n_6418)
);

AND2x4_ASAP7_75t_L g6419 ( 
.A(n_6211),
.B(n_5956),
.Y(n_6419)
);

INVx1_ASAP7_75t_L g6420 ( 
.A(n_6269),
.Y(n_6420)
);

AND2x2_ASAP7_75t_L g6421 ( 
.A(n_6230),
.B(n_6044),
.Y(n_6421)
);

INVx1_ASAP7_75t_L g6422 ( 
.A(n_6279),
.Y(n_6422)
);

OAI21xp33_ASAP7_75t_L g6423 ( 
.A1(n_6216),
.A2(n_6021),
.B(n_5987),
.Y(n_6423)
);

INVx1_ASAP7_75t_L g6424 ( 
.A(n_6281),
.Y(n_6424)
);

AND2x2_ASAP7_75t_L g6425 ( 
.A(n_6292),
.B(n_6048),
.Y(n_6425)
);

NAND2x1_ASAP7_75t_L g6426 ( 
.A(n_6128),
.B(n_6033),
.Y(n_6426)
);

NAND2xp5_ASAP7_75t_L g6427 ( 
.A(n_6241),
.B(n_5983),
.Y(n_6427)
);

INVx1_ASAP7_75t_L g6428 ( 
.A(n_6139),
.Y(n_6428)
);

AND2x2_ASAP7_75t_L g6429 ( 
.A(n_6187),
.B(n_6038),
.Y(n_6429)
);

INVx2_ASAP7_75t_L g6430 ( 
.A(n_6207),
.Y(n_6430)
);

INVx1_ASAP7_75t_L g6431 ( 
.A(n_6294),
.Y(n_6431)
);

INVx1_ASAP7_75t_L g6432 ( 
.A(n_6295),
.Y(n_6432)
);

AND2x2_ASAP7_75t_L g6433 ( 
.A(n_6247),
.B(n_5985),
.Y(n_6433)
);

OR2x2_ASAP7_75t_L g6434 ( 
.A(n_6273),
.B(n_5972),
.Y(n_6434)
);

INVx1_ASAP7_75t_L g6435 ( 
.A(n_6300),
.Y(n_6435)
);

OR2x6_ASAP7_75t_L g6436 ( 
.A(n_6212),
.B(n_5918),
.Y(n_6436)
);

AND2x4_ASAP7_75t_L g6437 ( 
.A(n_6249),
.B(n_5977),
.Y(n_6437)
);

AND2x2_ASAP7_75t_L g6438 ( 
.A(n_6251),
.B(n_5984),
.Y(n_6438)
);

INVx1_ASAP7_75t_L g6439 ( 
.A(n_6305),
.Y(n_6439)
);

INVx1_ASAP7_75t_L g6440 ( 
.A(n_6306),
.Y(n_6440)
);

INVx2_ASAP7_75t_L g6441 ( 
.A(n_6275),
.Y(n_6441)
);

AND2x2_ASAP7_75t_L g6442 ( 
.A(n_6256),
.B(n_6022),
.Y(n_6442)
);

OR2x2_ASAP7_75t_L g6443 ( 
.A(n_6278),
.B(n_5991),
.Y(n_6443)
);

INVx2_ASAP7_75t_L g6444 ( 
.A(n_6280),
.Y(n_6444)
);

NAND2xp5_ASAP7_75t_L g6445 ( 
.A(n_6241),
.B(n_6032),
.Y(n_6445)
);

NAND2xp5_ASAP7_75t_L g6446 ( 
.A(n_6202),
.B(n_6036),
.Y(n_6446)
);

NAND2xp5_ASAP7_75t_L g6447 ( 
.A(n_6174),
.B(n_6233),
.Y(n_6447)
);

INVx1_ASAP7_75t_L g6448 ( 
.A(n_6283),
.Y(n_6448)
);

NOR4xp25_ASAP7_75t_L g6449 ( 
.A(n_6132),
.B(n_6087),
.C(n_483),
.D(n_479),
.Y(n_6449)
);

AND2x2_ASAP7_75t_L g6450 ( 
.A(n_6331),
.B(n_6287),
.Y(n_6450)
);

INVx2_ASAP7_75t_SL g6451 ( 
.A(n_6343),
.Y(n_6451)
);

AND2x2_ASAP7_75t_L g6452 ( 
.A(n_6316),
.B(n_6289),
.Y(n_6452)
);

INVx1_ASAP7_75t_L g6453 ( 
.A(n_6352),
.Y(n_6453)
);

INVx1_ASAP7_75t_L g6454 ( 
.A(n_6355),
.Y(n_6454)
);

NAND2xp5_ASAP7_75t_L g6455 ( 
.A(n_6397),
.B(n_6290),
.Y(n_6455)
);

HB1xp67_ASAP7_75t_L g6456 ( 
.A(n_6361),
.Y(n_6456)
);

AND2x2_ASAP7_75t_L g6457 ( 
.A(n_6319),
.B(n_6259),
.Y(n_6457)
);

OR2x2_ASAP7_75t_L g6458 ( 
.A(n_6404),
.B(n_6237),
.Y(n_6458)
);

HB1xp67_ASAP7_75t_L g6459 ( 
.A(n_6334),
.Y(n_6459)
);

AND2x2_ASAP7_75t_L g6460 ( 
.A(n_6330),
.B(n_6282),
.Y(n_6460)
);

AND2x2_ASAP7_75t_L g6461 ( 
.A(n_6368),
.B(n_6310),
.Y(n_6461)
);

INVxp33_ASAP7_75t_L g6462 ( 
.A(n_6388),
.Y(n_6462)
);

OR2x2_ASAP7_75t_L g6463 ( 
.A(n_6413),
.B(n_6268),
.Y(n_6463)
);

INVx1_ASAP7_75t_SL g6464 ( 
.A(n_6347),
.Y(n_6464)
);

INVx3_ASAP7_75t_L g6465 ( 
.A(n_6323),
.Y(n_6465)
);

AOI21xp5_ASAP7_75t_L g6466 ( 
.A1(n_6384),
.A2(n_6170),
.B(n_6221),
.Y(n_6466)
);

AND2x2_ASAP7_75t_L g6467 ( 
.A(n_6429),
.B(n_6182),
.Y(n_6467)
);

OAI32xp33_ASAP7_75t_L g6468 ( 
.A1(n_6370),
.A2(n_6144),
.A3(n_6272),
.B1(n_6234),
.B2(n_6232),
.Y(n_6468)
);

INVxp67_ASAP7_75t_L g6469 ( 
.A(n_6369),
.Y(n_6469)
);

AND2x2_ASAP7_75t_L g6470 ( 
.A(n_6378),
.B(n_6296),
.Y(n_6470)
);

AND2x2_ASAP7_75t_L g6471 ( 
.A(n_6364),
.B(n_6168),
.Y(n_6471)
);

INVx2_ASAP7_75t_L g6472 ( 
.A(n_6360),
.Y(n_6472)
);

INVx2_ASAP7_75t_L g6473 ( 
.A(n_6350),
.Y(n_6473)
);

INVx1_ASAP7_75t_L g6474 ( 
.A(n_6314),
.Y(n_6474)
);

AND2x2_ASAP7_75t_L g6475 ( 
.A(n_6354),
.B(n_6399),
.Y(n_6475)
);

NAND2xp5_ASAP7_75t_L g6476 ( 
.A(n_6321),
.B(n_6301),
.Y(n_6476)
);

INVx1_ASAP7_75t_L g6477 ( 
.A(n_6327),
.Y(n_6477)
);

INVxp67_ASAP7_75t_L g6478 ( 
.A(n_6366),
.Y(n_6478)
);

CKINVDCx20_ASAP7_75t_R g6479 ( 
.A(n_6433),
.Y(n_6479)
);

INVx2_ASAP7_75t_L g6480 ( 
.A(n_6362),
.Y(n_6480)
);

INVx1_ASAP7_75t_L g6481 ( 
.A(n_6328),
.Y(n_6481)
);

INVx2_ASAP7_75t_L g6482 ( 
.A(n_6380),
.Y(n_6482)
);

INVx1_ASAP7_75t_L g6483 ( 
.A(n_6329),
.Y(n_6483)
);

NOR2xp67_ASAP7_75t_SL g6484 ( 
.A(n_6363),
.B(n_6298),
.Y(n_6484)
);

NAND2xp5_ASAP7_75t_L g6485 ( 
.A(n_6449),
.B(n_6219),
.Y(n_6485)
);

AND2x2_ASAP7_75t_L g6486 ( 
.A(n_6339),
.B(n_6285),
.Y(n_6486)
);

OAI222xp33_ASAP7_75t_L g6487 ( 
.A1(n_6418),
.A2(n_6137),
.B1(n_6198),
.B2(n_6236),
.C1(n_6215),
.C2(n_6159),
.Y(n_6487)
);

INVx2_ASAP7_75t_L g6488 ( 
.A(n_6426),
.Y(n_6488)
);

INVx1_ASAP7_75t_L g6489 ( 
.A(n_6315),
.Y(n_6489)
);

INVx1_ASAP7_75t_L g6490 ( 
.A(n_6317),
.Y(n_6490)
);

INVx1_ASAP7_75t_SL g6491 ( 
.A(n_6436),
.Y(n_6491)
);

INVx3_ASAP7_75t_L g6492 ( 
.A(n_6437),
.Y(n_6492)
);

NAND2xp5_ASAP7_75t_L g6493 ( 
.A(n_6412),
.B(n_6293),
.Y(n_6493)
);

INVx1_ASAP7_75t_L g6494 ( 
.A(n_6430),
.Y(n_6494)
);

AND2x2_ASAP7_75t_L g6495 ( 
.A(n_6318),
.B(n_6200),
.Y(n_6495)
);

INVx1_ASAP7_75t_L g6496 ( 
.A(n_6392),
.Y(n_6496)
);

OR2x2_ASAP7_75t_L g6497 ( 
.A(n_6389),
.B(n_6248),
.Y(n_6497)
);

INVxp67_ASAP7_75t_SL g6498 ( 
.A(n_6393),
.Y(n_6498)
);

INVx1_ASAP7_75t_L g6499 ( 
.A(n_6337),
.Y(n_6499)
);

BUFx2_ASAP7_75t_L g6500 ( 
.A(n_6436),
.Y(n_6500)
);

INVx1_ASAP7_75t_L g6501 ( 
.A(n_6338),
.Y(n_6501)
);

OR2x2_ASAP7_75t_L g6502 ( 
.A(n_6324),
.B(n_6224),
.Y(n_6502)
);

INVx1_ASAP7_75t_L g6503 ( 
.A(n_6340),
.Y(n_6503)
);

AND2x2_ASAP7_75t_L g6504 ( 
.A(n_6381),
.B(n_6336),
.Y(n_6504)
);

NOR2xp33_ASAP7_75t_L g6505 ( 
.A(n_6376),
.B(n_6267),
.Y(n_6505)
);

INVx1_ASAP7_75t_L g6506 ( 
.A(n_6341),
.Y(n_6506)
);

AND2x2_ASAP7_75t_L g6507 ( 
.A(n_6320),
.B(n_6203),
.Y(n_6507)
);

AND2x2_ASAP7_75t_L g6508 ( 
.A(n_6425),
.B(n_6161),
.Y(n_6508)
);

NAND2xp33_ASAP7_75t_L g6509 ( 
.A(n_6395),
.B(n_6184),
.Y(n_6509)
);

BUFx2_ASAP7_75t_SL g6510 ( 
.A(n_6372),
.Y(n_6510)
);

INVx1_ASAP7_75t_L g6511 ( 
.A(n_6342),
.Y(n_6511)
);

OR2x2_ASAP7_75t_L g6512 ( 
.A(n_6326),
.B(n_6402),
.Y(n_6512)
);

INVx1_ASAP7_75t_L g6513 ( 
.A(n_6344),
.Y(n_6513)
);

OR2x2_ASAP7_75t_L g6514 ( 
.A(n_6332),
.B(n_6194),
.Y(n_6514)
);

INVx1_ASAP7_75t_L g6515 ( 
.A(n_6348),
.Y(n_6515)
);

INVx2_ASAP7_75t_L g6516 ( 
.A(n_6419),
.Y(n_6516)
);

OAI22xp33_ASAP7_75t_SL g6517 ( 
.A1(n_6445),
.A2(n_6291),
.B1(n_6309),
.B2(n_6313),
.Y(n_6517)
);

NAND2xp5_ASAP7_75t_L g6518 ( 
.A(n_6421),
.B(n_6209),
.Y(n_6518)
);

INVx1_ASAP7_75t_L g6519 ( 
.A(n_6349),
.Y(n_6519)
);

NOR2xp33_ASAP7_75t_L g6520 ( 
.A(n_6356),
.B(n_6176),
.Y(n_6520)
);

OAI21xp33_ASAP7_75t_L g6521 ( 
.A1(n_6346),
.A2(n_6199),
.B(n_6171),
.Y(n_6521)
);

AND2x2_ASAP7_75t_L g6522 ( 
.A(n_6442),
.B(n_6266),
.Y(n_6522)
);

AND2x2_ASAP7_75t_L g6523 ( 
.A(n_6371),
.B(n_6297),
.Y(n_6523)
);

INVx1_ASAP7_75t_L g6524 ( 
.A(n_6351),
.Y(n_6524)
);

INVxp67_ASAP7_75t_L g6525 ( 
.A(n_6411),
.Y(n_6525)
);

INVx1_ASAP7_75t_SL g6526 ( 
.A(n_6438),
.Y(n_6526)
);

INVx1_ASAP7_75t_L g6527 ( 
.A(n_6353),
.Y(n_6527)
);

INVx1_ASAP7_75t_L g6528 ( 
.A(n_6358),
.Y(n_6528)
);

INVx1_ASAP7_75t_L g6529 ( 
.A(n_6359),
.Y(n_6529)
);

AND2x2_ASAP7_75t_L g6530 ( 
.A(n_6398),
.B(n_482),
.Y(n_6530)
);

OAI22xp5_ASAP7_75t_L g6531 ( 
.A1(n_6406),
.A2(n_486),
.B1(n_487),
.B2(n_485),
.Y(n_6531)
);

AND2x2_ASAP7_75t_L g6532 ( 
.A(n_6401),
.B(n_484),
.Y(n_6532)
);

INVx2_ASAP7_75t_L g6533 ( 
.A(n_6407),
.Y(n_6533)
);

NOR2xp33_ASAP7_75t_L g6534 ( 
.A(n_6423),
.B(n_485),
.Y(n_6534)
);

OR2x2_ASAP7_75t_L g6535 ( 
.A(n_6345),
.B(n_486),
.Y(n_6535)
);

INVx2_ASAP7_75t_SL g6536 ( 
.A(n_6408),
.Y(n_6536)
);

INVx1_ASAP7_75t_L g6537 ( 
.A(n_6365),
.Y(n_6537)
);

INVx1_ASAP7_75t_L g6538 ( 
.A(n_6367),
.Y(n_6538)
);

AND2x4_ASAP7_75t_L g6539 ( 
.A(n_6385),
.B(n_488),
.Y(n_6539)
);

INVx1_ASAP7_75t_L g6540 ( 
.A(n_6373),
.Y(n_6540)
);

NAND2xp5_ASAP7_75t_L g6541 ( 
.A(n_6390),
.B(n_489),
.Y(n_6541)
);

AOI32xp33_ASAP7_75t_L g6542 ( 
.A1(n_6409),
.A2(n_491),
.A3(n_489),
.B1(n_490),
.B2(n_492),
.Y(n_6542)
);

NAND2xp5_ASAP7_75t_L g6543 ( 
.A(n_6410),
.B(n_490),
.Y(n_6543)
);

AND2x2_ASAP7_75t_L g6544 ( 
.A(n_6377),
.B(n_491),
.Y(n_6544)
);

NAND2xp5_ASAP7_75t_SL g6545 ( 
.A(n_6417),
.B(n_493),
.Y(n_6545)
);

NAND2xp5_ASAP7_75t_L g6546 ( 
.A(n_6357),
.B(n_493),
.Y(n_6546)
);

NAND2xp5_ASAP7_75t_L g6547 ( 
.A(n_6400),
.B(n_494),
.Y(n_6547)
);

NAND2xp5_ASAP7_75t_SL g6548 ( 
.A(n_6427),
.B(n_495),
.Y(n_6548)
);

AND2x2_ASAP7_75t_SL g6549 ( 
.A(n_6322),
.B(n_495),
.Y(n_6549)
);

AND2x2_ASAP7_75t_L g6550 ( 
.A(n_6335),
.B(n_496),
.Y(n_6550)
);

INVx2_ASAP7_75t_L g6551 ( 
.A(n_6391),
.Y(n_6551)
);

CKINVDCx8_ASAP7_75t_R g6552 ( 
.A(n_6447),
.Y(n_6552)
);

OR2x2_ASAP7_75t_L g6553 ( 
.A(n_6325),
.B(n_496),
.Y(n_6553)
);

NAND2xp5_ASAP7_75t_L g6554 ( 
.A(n_6441),
.B(n_497),
.Y(n_6554)
);

INVx1_ASAP7_75t_L g6555 ( 
.A(n_6375),
.Y(n_6555)
);

AND2x2_ASAP7_75t_L g6556 ( 
.A(n_6416),
.B(n_6434),
.Y(n_6556)
);

INVx1_ASAP7_75t_L g6557 ( 
.A(n_6379),
.Y(n_6557)
);

NAND2x1_ASAP7_75t_L g6558 ( 
.A(n_6444),
.B(n_497),
.Y(n_6558)
);

INVxp67_ASAP7_75t_SL g6559 ( 
.A(n_6382),
.Y(n_6559)
);

NAND2xp5_ASAP7_75t_L g6560 ( 
.A(n_6333),
.B(n_498),
.Y(n_6560)
);

INVx2_ASAP7_75t_SL g6561 ( 
.A(n_6383),
.Y(n_6561)
);

AOI21xp33_ASAP7_75t_SL g6562 ( 
.A1(n_6374),
.A2(n_498),
.B(n_499),
.Y(n_6562)
);

INVx1_ASAP7_75t_L g6563 ( 
.A(n_6386),
.Y(n_6563)
);

NAND2xp5_ASAP7_75t_L g6564 ( 
.A(n_6448),
.B(n_499),
.Y(n_6564)
);

INVx2_ASAP7_75t_L g6565 ( 
.A(n_6443),
.Y(n_6565)
);

OR2x2_ASAP7_75t_L g6566 ( 
.A(n_6446),
.B(n_500),
.Y(n_6566)
);

NOR2x1_ASAP7_75t_L g6567 ( 
.A(n_6428),
.B(n_501),
.Y(n_6567)
);

NAND2xp5_ASAP7_75t_L g6568 ( 
.A(n_6431),
.B(n_501),
.Y(n_6568)
);

NAND2xp5_ASAP7_75t_L g6569 ( 
.A(n_6432),
.B(n_502),
.Y(n_6569)
);

INVx3_ASAP7_75t_L g6570 ( 
.A(n_6435),
.Y(n_6570)
);

INVx1_ASAP7_75t_L g6571 ( 
.A(n_6387),
.Y(n_6571)
);

AND2x2_ASAP7_75t_L g6572 ( 
.A(n_6439),
.B(n_6440),
.Y(n_6572)
);

AND2x2_ASAP7_75t_L g6573 ( 
.A(n_6394),
.B(n_502),
.Y(n_6573)
);

INVx2_ASAP7_75t_L g6574 ( 
.A(n_6396),
.Y(n_6574)
);

INVx1_ASAP7_75t_L g6575 ( 
.A(n_6403),
.Y(n_6575)
);

INVx1_ASAP7_75t_L g6576 ( 
.A(n_6405),
.Y(n_6576)
);

INVx1_ASAP7_75t_L g6577 ( 
.A(n_6414),
.Y(n_6577)
);

INVx1_ASAP7_75t_L g6578 ( 
.A(n_6415),
.Y(n_6578)
);

INVx1_ASAP7_75t_L g6579 ( 
.A(n_6420),
.Y(n_6579)
);

INVx1_ASAP7_75t_L g6580 ( 
.A(n_6422),
.Y(n_6580)
);

NAND2xp5_ASAP7_75t_L g6581 ( 
.A(n_6424),
.B(n_503),
.Y(n_6581)
);

NOR2xp33_ASAP7_75t_L g6582 ( 
.A(n_6464),
.B(n_6451),
.Y(n_6582)
);

AND2x2_ASAP7_75t_L g6583 ( 
.A(n_6457),
.B(n_504),
.Y(n_6583)
);

NOR2xp33_ASAP7_75t_L g6584 ( 
.A(n_6479),
.B(n_504),
.Y(n_6584)
);

NOR2xp33_ASAP7_75t_L g6585 ( 
.A(n_6491),
.B(n_505),
.Y(n_6585)
);

NAND2xp5_ASAP7_75t_L g6586 ( 
.A(n_6459),
.B(n_505),
.Y(n_6586)
);

INVx1_ASAP7_75t_L g6587 ( 
.A(n_6453),
.Y(n_6587)
);

AND2x2_ASAP7_75t_L g6588 ( 
.A(n_6460),
.B(n_506),
.Y(n_6588)
);

NAND2xp5_ASAP7_75t_L g6589 ( 
.A(n_6456),
.B(n_508),
.Y(n_6589)
);

AND2x2_ASAP7_75t_L g6590 ( 
.A(n_6475),
.B(n_6500),
.Y(n_6590)
);

HB1xp67_ASAP7_75t_L g6591 ( 
.A(n_6558),
.Y(n_6591)
);

INVx2_ASAP7_75t_L g6592 ( 
.A(n_6465),
.Y(n_6592)
);

NAND2x1p5_ASAP7_75t_SL g6593 ( 
.A(n_6482),
.B(n_509),
.Y(n_6593)
);

INVx1_ASAP7_75t_L g6594 ( 
.A(n_6454),
.Y(n_6594)
);

NAND2xp5_ASAP7_75t_L g6595 ( 
.A(n_6549),
.B(n_509),
.Y(n_6595)
);

AND2x2_ASAP7_75t_L g6596 ( 
.A(n_6510),
.B(n_510),
.Y(n_6596)
);

INVx1_ASAP7_75t_SL g6597 ( 
.A(n_6450),
.Y(n_6597)
);

INVx3_ASAP7_75t_L g6598 ( 
.A(n_6492),
.Y(n_6598)
);

INVx1_ASAP7_75t_L g6599 ( 
.A(n_6559),
.Y(n_6599)
);

INVx1_ASAP7_75t_SL g6600 ( 
.A(n_6526),
.Y(n_6600)
);

AOI221xp5_ASAP7_75t_L g6601 ( 
.A1(n_6478),
.A2(n_513),
.B1(n_511),
.B2(n_512),
.C(n_514),
.Y(n_6601)
);

INVx1_ASAP7_75t_L g6602 ( 
.A(n_6573),
.Y(n_6602)
);

AND2x2_ASAP7_75t_L g6603 ( 
.A(n_6452),
.B(n_512),
.Y(n_6603)
);

NAND2xp5_ASAP7_75t_SL g6604 ( 
.A(n_6517),
.B(n_515),
.Y(n_6604)
);

HB1xp67_ASAP7_75t_L g6605 ( 
.A(n_6567),
.Y(n_6605)
);

AND2x2_ASAP7_75t_L g6606 ( 
.A(n_6461),
.B(n_516),
.Y(n_6606)
);

INVx1_ASAP7_75t_L g6607 ( 
.A(n_6544),
.Y(n_6607)
);

AND2x4_ASAP7_75t_L g6608 ( 
.A(n_6473),
.B(n_6480),
.Y(n_6608)
);

INVx1_ASAP7_75t_L g6609 ( 
.A(n_6458),
.Y(n_6609)
);

NOR3xp33_ASAP7_75t_L g6610 ( 
.A(n_6509),
.B(n_6520),
.C(n_6476),
.Y(n_6610)
);

NAND2xp33_ASAP7_75t_SL g6611 ( 
.A(n_6462),
.B(n_6484),
.Y(n_6611)
);

INVx1_ASAP7_75t_SL g6612 ( 
.A(n_6471),
.Y(n_6612)
);

NAND2xp5_ASAP7_75t_L g6613 ( 
.A(n_6472),
.B(n_516),
.Y(n_6613)
);

OR2x2_ASAP7_75t_L g6614 ( 
.A(n_6518),
.B(n_517),
.Y(n_6614)
);

OR2x2_ASAP7_75t_L g6615 ( 
.A(n_6497),
.B(n_517),
.Y(n_6615)
);

INVx1_ASAP7_75t_L g6616 ( 
.A(n_6554),
.Y(n_6616)
);

OR2x2_ASAP7_75t_L g6617 ( 
.A(n_6512),
.B(n_518),
.Y(n_6617)
);

AND2x2_ASAP7_75t_SL g6618 ( 
.A(n_6485),
.B(n_518),
.Y(n_6618)
);

OAI31xp33_ASAP7_75t_L g6619 ( 
.A1(n_6487),
.A2(n_521),
.A3(n_519),
.B(n_520),
.Y(n_6619)
);

NAND2xp5_ASAP7_75t_L g6620 ( 
.A(n_6504),
.B(n_522),
.Y(n_6620)
);

CKINVDCx16_ASAP7_75t_R g6621 ( 
.A(n_6463),
.Y(n_6621)
);

INVx1_ASAP7_75t_L g6622 ( 
.A(n_6561),
.Y(n_6622)
);

INVx2_ASAP7_75t_L g6623 ( 
.A(n_6488),
.Y(n_6623)
);

INVx2_ASAP7_75t_L g6624 ( 
.A(n_6516),
.Y(n_6624)
);

AND2x2_ASAP7_75t_L g6625 ( 
.A(n_6495),
.B(n_523),
.Y(n_6625)
);

AOI21xp5_ASAP7_75t_L g6626 ( 
.A1(n_6466),
.A2(n_524),
.B(n_525),
.Y(n_6626)
);

INVx1_ASAP7_75t_SL g6627 ( 
.A(n_6467),
.Y(n_6627)
);

OR2x2_ASAP7_75t_L g6628 ( 
.A(n_6525),
.B(n_524),
.Y(n_6628)
);

CKINVDCx20_ASAP7_75t_R g6629 ( 
.A(n_6552),
.Y(n_6629)
);

NAND4xp25_ASAP7_75t_L g6630 ( 
.A(n_6505),
.B(n_527),
.C(n_525),
.D(n_526),
.Y(n_6630)
);

INVx1_ASAP7_75t_L g6631 ( 
.A(n_6550),
.Y(n_6631)
);

NAND2xp5_ASAP7_75t_L g6632 ( 
.A(n_6508),
.B(n_526),
.Y(n_6632)
);

INVx1_ASAP7_75t_L g6633 ( 
.A(n_6551),
.Y(n_6633)
);

NOR2xp33_ASAP7_75t_L g6634 ( 
.A(n_6468),
.B(n_528),
.Y(n_6634)
);

AND2x2_ASAP7_75t_L g6635 ( 
.A(n_6470),
.B(n_528),
.Y(n_6635)
);

OR2x2_ASAP7_75t_L g6636 ( 
.A(n_6455),
.B(n_529),
.Y(n_6636)
);

AOI22xp33_ASAP7_75t_L g6637 ( 
.A1(n_6521),
.A2(n_6536),
.B1(n_6533),
.B2(n_6514),
.Y(n_6637)
);

AND2x2_ASAP7_75t_L g6638 ( 
.A(n_6486),
.B(n_529),
.Y(n_6638)
);

INVx1_ASAP7_75t_L g6639 ( 
.A(n_6530),
.Y(n_6639)
);

NAND2x1p5_ASAP7_75t_L g6640 ( 
.A(n_6539),
.B(n_530),
.Y(n_6640)
);

AOI33xp33_ASAP7_75t_L g6641 ( 
.A1(n_6489),
.A2(n_534),
.A3(n_537),
.B1(n_531),
.B2(n_533),
.B3(n_535),
.Y(n_6641)
);

NOR3xp33_ASAP7_75t_L g6642 ( 
.A(n_6494),
.B(n_531),
.C(n_534),
.Y(n_6642)
);

INVx1_ASAP7_75t_L g6643 ( 
.A(n_6532),
.Y(n_6643)
);

AND2x2_ASAP7_75t_L g6644 ( 
.A(n_6556),
.B(n_535),
.Y(n_6644)
);

AND2x2_ASAP7_75t_L g6645 ( 
.A(n_6507),
.B(n_537),
.Y(n_6645)
);

INVx1_ASAP7_75t_SL g6646 ( 
.A(n_6553),
.Y(n_6646)
);

INVx2_ASAP7_75t_L g6647 ( 
.A(n_6539),
.Y(n_6647)
);

HB1xp67_ASAP7_75t_L g6648 ( 
.A(n_6469),
.Y(n_6648)
);

AND2x4_ASAP7_75t_L g6649 ( 
.A(n_6496),
.B(n_6565),
.Y(n_6649)
);

NAND2xp5_ASAP7_75t_L g6650 ( 
.A(n_6542),
.B(n_538),
.Y(n_6650)
);

AND2x2_ASAP7_75t_L g6651 ( 
.A(n_6523),
.B(n_539),
.Y(n_6651)
);

INVx1_ASAP7_75t_L g6652 ( 
.A(n_6498),
.Y(n_6652)
);

OR2x2_ASAP7_75t_L g6653 ( 
.A(n_6493),
.B(n_539),
.Y(n_6653)
);

NAND2xp33_ASAP7_75t_SL g6654 ( 
.A(n_6545),
.B(n_540),
.Y(n_6654)
);

NAND2xp5_ASAP7_75t_L g6655 ( 
.A(n_6522),
.B(n_540),
.Y(n_6655)
);

NAND2xp33_ASAP7_75t_R g6656 ( 
.A(n_6562),
.B(n_541),
.Y(n_6656)
);

NAND2xp5_ASAP7_75t_L g6657 ( 
.A(n_6534),
.B(n_541),
.Y(n_6657)
);

NAND2xp5_ASAP7_75t_L g6658 ( 
.A(n_6531),
.B(n_542),
.Y(n_6658)
);

AND2x2_ASAP7_75t_L g6659 ( 
.A(n_6474),
.B(n_542),
.Y(n_6659)
);

INVx1_ASAP7_75t_L g6660 ( 
.A(n_6564),
.Y(n_6660)
);

INVx1_ASAP7_75t_L g6661 ( 
.A(n_6477),
.Y(n_6661)
);

NAND2xp5_ASAP7_75t_L g6662 ( 
.A(n_6548),
.B(n_544),
.Y(n_6662)
);

AND2x2_ASAP7_75t_L g6663 ( 
.A(n_6481),
.B(n_545),
.Y(n_6663)
);

NOR3xp33_ASAP7_75t_SL g6664 ( 
.A(n_6490),
.B(n_6483),
.C(n_6499),
.Y(n_6664)
);

INVx1_ASAP7_75t_SL g6665 ( 
.A(n_6502),
.Y(n_6665)
);

AND2x2_ASAP7_75t_L g6666 ( 
.A(n_6535),
.B(n_6566),
.Y(n_6666)
);

INVx2_ASAP7_75t_L g6667 ( 
.A(n_6570),
.Y(n_6667)
);

NOR2xp33_ASAP7_75t_L g6668 ( 
.A(n_6546),
.B(n_545),
.Y(n_6668)
);

INVx2_ASAP7_75t_L g6669 ( 
.A(n_6572),
.Y(n_6669)
);

NAND2xp5_ASAP7_75t_L g6670 ( 
.A(n_6541),
.B(n_6543),
.Y(n_6670)
);

AOI31xp33_ASAP7_75t_L g6671 ( 
.A1(n_6501),
.A2(n_550),
.A3(n_547),
.B(n_548),
.Y(n_6671)
);

INVx1_ASAP7_75t_L g6672 ( 
.A(n_6547),
.Y(n_6672)
);

INVx1_ASAP7_75t_L g6673 ( 
.A(n_6568),
.Y(n_6673)
);

NOR3xp33_ASAP7_75t_SL g6674 ( 
.A(n_6503),
.B(n_547),
.C(n_548),
.Y(n_6674)
);

INVx1_ASAP7_75t_L g6675 ( 
.A(n_6569),
.Y(n_6675)
);

INVx1_ASAP7_75t_L g6676 ( 
.A(n_6581),
.Y(n_6676)
);

OR2x2_ASAP7_75t_L g6677 ( 
.A(n_6560),
.B(n_550),
.Y(n_6677)
);

OAI31xp33_ASAP7_75t_L g6678 ( 
.A1(n_6506),
.A2(n_553),
.A3(n_551),
.B(n_552),
.Y(n_6678)
);

AND2x2_ASAP7_75t_L g6679 ( 
.A(n_6574),
.B(n_551),
.Y(n_6679)
);

AND2x2_ASAP7_75t_L g6680 ( 
.A(n_6511),
.B(n_552),
.Y(n_6680)
);

INVx1_ASAP7_75t_L g6681 ( 
.A(n_6513),
.Y(n_6681)
);

INVx1_ASAP7_75t_SL g6682 ( 
.A(n_6515),
.Y(n_6682)
);

AND2x2_ASAP7_75t_L g6683 ( 
.A(n_6519),
.B(n_553),
.Y(n_6683)
);

NAND2xp5_ASAP7_75t_L g6684 ( 
.A(n_6524),
.B(n_554),
.Y(n_6684)
);

INVx1_ASAP7_75t_SL g6685 ( 
.A(n_6527),
.Y(n_6685)
);

INVx1_ASAP7_75t_L g6686 ( 
.A(n_6528),
.Y(n_6686)
);

INVx1_ASAP7_75t_SL g6687 ( 
.A(n_6529),
.Y(n_6687)
);

INVx1_ASAP7_75t_L g6688 ( 
.A(n_6537),
.Y(n_6688)
);

AND2x2_ASAP7_75t_L g6689 ( 
.A(n_6538),
.B(n_554),
.Y(n_6689)
);

OR2x2_ASAP7_75t_L g6690 ( 
.A(n_6540),
.B(n_555),
.Y(n_6690)
);

AND2x2_ASAP7_75t_L g6691 ( 
.A(n_6555),
.B(n_556),
.Y(n_6691)
);

AND2x4_ASAP7_75t_L g6692 ( 
.A(n_6557),
.B(n_557),
.Y(n_6692)
);

AND2x2_ASAP7_75t_L g6693 ( 
.A(n_6563),
.B(n_557),
.Y(n_6693)
);

AOI33xp33_ASAP7_75t_L g6694 ( 
.A1(n_6571),
.A2(n_6578),
.A3(n_6576),
.B1(n_6579),
.B2(n_6577),
.B3(n_6575),
.Y(n_6694)
);

AND2x2_ASAP7_75t_L g6695 ( 
.A(n_6580),
.B(n_558),
.Y(n_6695)
);

NOR2xp67_ASAP7_75t_SL g6696 ( 
.A(n_6552),
.B(n_559),
.Y(n_6696)
);

AND2x2_ASAP7_75t_L g6697 ( 
.A(n_6464),
.B(n_559),
.Y(n_6697)
);

AND2x4_ASAP7_75t_L g6698 ( 
.A(n_6451),
.B(n_560),
.Y(n_6698)
);

INVx2_ASAP7_75t_L g6699 ( 
.A(n_6479),
.Y(n_6699)
);

INVx1_ASAP7_75t_L g6700 ( 
.A(n_6459),
.Y(n_6700)
);

AND2x2_ASAP7_75t_L g6701 ( 
.A(n_6464),
.B(n_561),
.Y(n_6701)
);

AND2x2_ASAP7_75t_L g6702 ( 
.A(n_6464),
.B(n_561),
.Y(n_6702)
);

INVx1_ASAP7_75t_L g6703 ( 
.A(n_6459),
.Y(n_6703)
);

NAND2xp5_ASAP7_75t_L g6704 ( 
.A(n_6491),
.B(n_562),
.Y(n_6704)
);

AND2x2_ASAP7_75t_L g6705 ( 
.A(n_6464),
.B(n_563),
.Y(n_6705)
);

INVx1_ASAP7_75t_L g6706 ( 
.A(n_6459),
.Y(n_6706)
);

INVx2_ASAP7_75t_L g6707 ( 
.A(n_6479),
.Y(n_6707)
);

AND2x2_ASAP7_75t_L g6708 ( 
.A(n_6464),
.B(n_563),
.Y(n_6708)
);

INVx3_ASAP7_75t_L g6709 ( 
.A(n_6465),
.Y(n_6709)
);

NOR2xp33_ASAP7_75t_L g6710 ( 
.A(n_6464),
.B(n_564),
.Y(n_6710)
);

NAND2xp5_ASAP7_75t_L g6711 ( 
.A(n_6491),
.B(n_565),
.Y(n_6711)
);

NAND2xp5_ASAP7_75t_L g6712 ( 
.A(n_6491),
.B(n_565),
.Y(n_6712)
);

NAND4xp25_ASAP7_75t_L g6713 ( 
.A(n_6491),
.B(n_568),
.C(n_566),
.D(n_567),
.Y(n_6713)
);

AND2x4_ASAP7_75t_L g6714 ( 
.A(n_6699),
.B(n_567),
.Y(n_6714)
);

INVx1_ASAP7_75t_SL g6715 ( 
.A(n_6629),
.Y(n_6715)
);

NAND2x1p5_ASAP7_75t_L g6716 ( 
.A(n_6696),
.B(n_568),
.Y(n_6716)
);

NAND2xp5_ASAP7_75t_L g6717 ( 
.A(n_6621),
.B(n_569),
.Y(n_6717)
);

INVx2_ASAP7_75t_L g6718 ( 
.A(n_6707),
.Y(n_6718)
);

NAND2xp5_ASAP7_75t_L g6719 ( 
.A(n_6597),
.B(n_6591),
.Y(n_6719)
);

INVx1_ASAP7_75t_L g6720 ( 
.A(n_6605),
.Y(n_6720)
);

NAND2xp5_ASAP7_75t_SL g6721 ( 
.A(n_6619),
.B(n_570),
.Y(n_6721)
);

INVx2_ASAP7_75t_L g6722 ( 
.A(n_6640),
.Y(n_6722)
);

HB1xp67_ASAP7_75t_L g6723 ( 
.A(n_6596),
.Y(n_6723)
);

OAI21xp33_ASAP7_75t_L g6724 ( 
.A1(n_6582),
.A2(n_570),
.B(n_571),
.Y(n_6724)
);

AND2x2_ASAP7_75t_L g6725 ( 
.A(n_6590),
.B(n_571),
.Y(n_6725)
);

INVx1_ASAP7_75t_L g6726 ( 
.A(n_6648),
.Y(n_6726)
);

INVx1_ASAP7_75t_L g6727 ( 
.A(n_6700),
.Y(n_6727)
);

INVx1_ASAP7_75t_L g6728 ( 
.A(n_6703),
.Y(n_6728)
);

INVx1_ASAP7_75t_L g6729 ( 
.A(n_6706),
.Y(n_6729)
);

INVx1_ASAP7_75t_L g6730 ( 
.A(n_6599),
.Y(n_6730)
);

NAND2xp5_ASAP7_75t_L g6731 ( 
.A(n_6627),
.B(n_573),
.Y(n_6731)
);

OR2x2_ASAP7_75t_L g6732 ( 
.A(n_6593),
.B(n_6600),
.Y(n_6732)
);

OR2x2_ASAP7_75t_L g6733 ( 
.A(n_6614),
.B(n_573),
.Y(n_6733)
);

AND2x2_ASAP7_75t_L g6734 ( 
.A(n_6598),
.B(n_574),
.Y(n_6734)
);

INVx1_ASAP7_75t_L g6735 ( 
.A(n_6644),
.Y(n_6735)
);

AND2x2_ASAP7_75t_L g6736 ( 
.A(n_6709),
.B(n_574),
.Y(n_6736)
);

INVxp67_ASAP7_75t_L g6737 ( 
.A(n_6656),
.Y(n_6737)
);

HB1xp67_ASAP7_75t_L g6738 ( 
.A(n_6698),
.Y(n_6738)
);

AND2x2_ASAP7_75t_L g6739 ( 
.A(n_6697),
.B(n_575),
.Y(n_6739)
);

NAND4xp25_ASAP7_75t_L g6740 ( 
.A(n_6610),
.B(n_578),
.C(n_576),
.D(n_577),
.Y(n_6740)
);

AOI21xp5_ASAP7_75t_L g6741 ( 
.A1(n_6604),
.A2(n_577),
.B(n_578),
.Y(n_6741)
);

OR2x2_ASAP7_75t_L g6742 ( 
.A(n_6622),
.B(n_580),
.Y(n_6742)
);

OR2x2_ASAP7_75t_L g6743 ( 
.A(n_6615),
.B(n_580),
.Y(n_6743)
);

AND2x2_ASAP7_75t_L g6744 ( 
.A(n_6701),
.B(n_581),
.Y(n_6744)
);

AND2x2_ASAP7_75t_L g6745 ( 
.A(n_6702),
.B(n_6705),
.Y(n_6745)
);

INVxp67_ASAP7_75t_L g6746 ( 
.A(n_6584),
.Y(n_6746)
);

INVxp67_ASAP7_75t_L g6747 ( 
.A(n_6611),
.Y(n_6747)
);

INVx2_ASAP7_75t_L g6748 ( 
.A(n_6608),
.Y(n_6748)
);

NAND2xp5_ASAP7_75t_L g6749 ( 
.A(n_6618),
.B(n_581),
.Y(n_6749)
);

INVx1_ASAP7_75t_L g6750 ( 
.A(n_6708),
.Y(n_6750)
);

AND2x2_ASAP7_75t_L g6751 ( 
.A(n_6592),
.B(n_582),
.Y(n_6751)
);

INVx1_ASAP7_75t_L g6752 ( 
.A(n_6606),
.Y(n_6752)
);

INVx1_ASAP7_75t_L g6753 ( 
.A(n_6609),
.Y(n_6753)
);

INVx1_ASAP7_75t_L g6754 ( 
.A(n_6704),
.Y(n_6754)
);

NAND2xp5_ASAP7_75t_L g6755 ( 
.A(n_6612),
.B(n_582),
.Y(n_6755)
);

AND2x2_ASAP7_75t_L g6756 ( 
.A(n_6645),
.B(n_583),
.Y(n_6756)
);

HB1xp67_ASAP7_75t_L g6757 ( 
.A(n_6647),
.Y(n_6757)
);

AND2x2_ASAP7_75t_L g6758 ( 
.A(n_6651),
.B(n_584),
.Y(n_6758)
);

NAND2xp5_ASAP7_75t_L g6759 ( 
.A(n_6710),
.B(n_6583),
.Y(n_6759)
);

XOR2x2_ASAP7_75t_L g6760 ( 
.A(n_6634),
.B(n_585),
.Y(n_6760)
);

NAND2xp5_ASAP7_75t_L g6761 ( 
.A(n_6588),
.B(n_585),
.Y(n_6761)
);

AND2x4_ASAP7_75t_L g6762 ( 
.A(n_6624),
.B(n_586),
.Y(n_6762)
);

INVx1_ASAP7_75t_L g6763 ( 
.A(n_6711),
.Y(n_6763)
);

INVx1_ASAP7_75t_SL g6764 ( 
.A(n_6654),
.Y(n_6764)
);

INVx1_ASAP7_75t_L g6765 ( 
.A(n_6712),
.Y(n_6765)
);

OR2x2_ASAP7_75t_L g6766 ( 
.A(n_6617),
.B(n_586),
.Y(n_6766)
);

HB1xp67_ASAP7_75t_L g6767 ( 
.A(n_6603),
.Y(n_6767)
);

NAND2xp5_ASAP7_75t_L g6768 ( 
.A(n_6623),
.B(n_588),
.Y(n_6768)
);

INVx1_ASAP7_75t_L g6769 ( 
.A(n_6607),
.Y(n_6769)
);

NAND2xp5_ASAP7_75t_L g6770 ( 
.A(n_6635),
.B(n_588),
.Y(n_6770)
);

OR2x2_ASAP7_75t_L g6771 ( 
.A(n_6646),
.B(n_589),
.Y(n_6771)
);

INVx1_ASAP7_75t_L g6772 ( 
.A(n_6628),
.Y(n_6772)
);

BUFx2_ASAP7_75t_L g6773 ( 
.A(n_6649),
.Y(n_6773)
);

AND2x2_ASAP7_75t_L g6774 ( 
.A(n_6639),
.B(n_589),
.Y(n_6774)
);

AND2x2_ASAP7_75t_L g6775 ( 
.A(n_6643),
.B(n_590),
.Y(n_6775)
);

NAND2xp5_ASAP7_75t_L g6776 ( 
.A(n_6625),
.B(n_590),
.Y(n_6776)
);

OR2x2_ASAP7_75t_L g6777 ( 
.A(n_6632),
.B(n_591),
.Y(n_6777)
);

OR2x2_ASAP7_75t_L g6778 ( 
.A(n_6665),
.B(n_591),
.Y(n_6778)
);

AND2x4_ASAP7_75t_L g6779 ( 
.A(n_6669),
.B(n_592),
.Y(n_6779)
);

NAND2xp5_ASAP7_75t_SL g6780 ( 
.A(n_6626),
.B(n_592),
.Y(n_6780)
);

HB1xp67_ASAP7_75t_L g6781 ( 
.A(n_6589),
.Y(n_6781)
);

INVx1_ASAP7_75t_L g6782 ( 
.A(n_6652),
.Y(n_6782)
);

NOR2xp67_ASAP7_75t_L g6783 ( 
.A(n_6667),
.B(n_594),
.Y(n_6783)
);

OR2x2_ASAP7_75t_L g6784 ( 
.A(n_6655),
.B(n_593),
.Y(n_6784)
);

INVx2_ASAP7_75t_L g6785 ( 
.A(n_6692),
.Y(n_6785)
);

INVx1_ASAP7_75t_L g6786 ( 
.A(n_6690),
.Y(n_6786)
);

BUFx2_ASAP7_75t_L g6787 ( 
.A(n_6664),
.Y(n_6787)
);

INVx1_ASAP7_75t_L g6788 ( 
.A(n_6620),
.Y(n_6788)
);

NAND2xp5_ASAP7_75t_L g6789 ( 
.A(n_6585),
.B(n_593),
.Y(n_6789)
);

INVx4_ASAP7_75t_L g6790 ( 
.A(n_6679),
.Y(n_6790)
);

INVx1_ASAP7_75t_L g6791 ( 
.A(n_6659),
.Y(n_6791)
);

INVx3_ASAP7_75t_L g6792 ( 
.A(n_6633),
.Y(n_6792)
);

AND2x4_ASAP7_75t_L g6793 ( 
.A(n_6631),
.B(n_594),
.Y(n_6793)
);

NOR2x1_ASAP7_75t_L g6794 ( 
.A(n_6630),
.B(n_595),
.Y(n_6794)
);

AND2x2_ASAP7_75t_L g6795 ( 
.A(n_6666),
.B(n_595),
.Y(n_6795)
);

AND2x2_ASAP7_75t_L g6796 ( 
.A(n_6638),
.B(n_6602),
.Y(n_6796)
);

NOR2xp33_ASAP7_75t_L g6797 ( 
.A(n_6713),
.B(n_597),
.Y(n_6797)
);

OR2x2_ASAP7_75t_L g6798 ( 
.A(n_6653),
.B(n_597),
.Y(n_6798)
);

INVx1_ASAP7_75t_L g6799 ( 
.A(n_6663),
.Y(n_6799)
);

AND2x2_ASAP7_75t_L g6800 ( 
.A(n_6637),
.B(n_6672),
.Y(n_6800)
);

INVx1_ASAP7_75t_L g6801 ( 
.A(n_6613),
.Y(n_6801)
);

INVx1_ASAP7_75t_L g6802 ( 
.A(n_6680),
.Y(n_6802)
);

HB1xp67_ASAP7_75t_L g6803 ( 
.A(n_6586),
.Y(n_6803)
);

AND2x4_ASAP7_75t_L g6804 ( 
.A(n_6587),
.B(n_598),
.Y(n_6804)
);

NOR2xp33_ASAP7_75t_L g6805 ( 
.A(n_6650),
.B(n_598),
.Y(n_6805)
);

NAND2xp5_ASAP7_75t_L g6806 ( 
.A(n_6668),
.B(n_599),
.Y(n_6806)
);

INVx2_ASAP7_75t_L g6807 ( 
.A(n_6683),
.Y(n_6807)
);

NAND2xp5_ASAP7_75t_L g6808 ( 
.A(n_6594),
.B(n_599),
.Y(n_6808)
);

OR2x2_ASAP7_75t_L g6809 ( 
.A(n_6636),
.B(n_600),
.Y(n_6809)
);

NAND3xp33_ASAP7_75t_L g6810 ( 
.A(n_6642),
.B(n_601),
.C(n_602),
.Y(n_6810)
);

NAND2xp5_ASAP7_75t_L g6811 ( 
.A(n_6689),
.B(n_602),
.Y(n_6811)
);

INVx1_ASAP7_75t_L g6812 ( 
.A(n_6691),
.Y(n_6812)
);

INVx1_ASAP7_75t_L g6813 ( 
.A(n_6693),
.Y(n_6813)
);

OR2x2_ASAP7_75t_L g6814 ( 
.A(n_6670),
.B(n_6682),
.Y(n_6814)
);

INVx2_ASAP7_75t_SL g6815 ( 
.A(n_6695),
.Y(n_6815)
);

INVx2_ASAP7_75t_L g6816 ( 
.A(n_6677),
.Y(n_6816)
);

INVx3_ASAP7_75t_L g6817 ( 
.A(n_6685),
.Y(n_6817)
);

INVx1_ASAP7_75t_L g6818 ( 
.A(n_6684),
.Y(n_6818)
);

NAND2xp5_ASAP7_75t_L g6819 ( 
.A(n_6678),
.B(n_603),
.Y(n_6819)
);

NAND2xp5_ASAP7_75t_L g6820 ( 
.A(n_6674),
.B(n_603),
.Y(n_6820)
);

O2A1O1Ixp33_ASAP7_75t_L g6821 ( 
.A1(n_6671),
.A2(n_607),
.B(n_604),
.C(n_606),
.Y(n_6821)
);

NAND2xp5_ASAP7_75t_L g6822 ( 
.A(n_6687),
.B(n_604),
.Y(n_6822)
);

INVx2_ASAP7_75t_L g6823 ( 
.A(n_6661),
.Y(n_6823)
);

CKINVDCx16_ASAP7_75t_R g6824 ( 
.A(n_6595),
.Y(n_6824)
);

AND2x2_ASAP7_75t_L g6825 ( 
.A(n_6660),
.B(n_607),
.Y(n_6825)
);

AOI211xp5_ASAP7_75t_L g6826 ( 
.A1(n_6601),
.A2(n_610),
.B(n_608),
.C(n_609),
.Y(n_6826)
);

OR2x2_ASAP7_75t_L g6827 ( 
.A(n_6673),
.B(n_610),
.Y(n_6827)
);

INVx2_ASAP7_75t_L g6828 ( 
.A(n_6616),
.Y(n_6828)
);

INVx1_ASAP7_75t_L g6829 ( 
.A(n_6694),
.Y(n_6829)
);

AND2x2_ASAP7_75t_L g6830 ( 
.A(n_6675),
.B(n_6676),
.Y(n_6830)
);

NAND2xp5_ASAP7_75t_L g6831 ( 
.A(n_6641),
.B(n_611),
.Y(n_6831)
);

INVx1_ASAP7_75t_SL g6832 ( 
.A(n_6662),
.Y(n_6832)
);

NOR2xp33_ASAP7_75t_L g6833 ( 
.A(n_6657),
.B(n_6658),
.Y(n_6833)
);

AND2x2_ASAP7_75t_L g6834 ( 
.A(n_6681),
.B(n_612),
.Y(n_6834)
);

INVx2_ASAP7_75t_L g6835 ( 
.A(n_6686),
.Y(n_6835)
);

INVx2_ASAP7_75t_L g6836 ( 
.A(n_6688),
.Y(n_6836)
);

NAND2xp5_ASAP7_75t_L g6837 ( 
.A(n_6621),
.B(n_613),
.Y(n_6837)
);

NAND2xp5_ASAP7_75t_L g6838 ( 
.A(n_6621),
.B(n_613),
.Y(n_6838)
);

AND2x2_ASAP7_75t_L g6839 ( 
.A(n_6590),
.B(n_614),
.Y(n_6839)
);

INVx2_ASAP7_75t_L g6840 ( 
.A(n_6699),
.Y(n_6840)
);

NOR2x1_ASAP7_75t_L g6841 ( 
.A(n_6629),
.B(n_615),
.Y(n_6841)
);

INVx2_ASAP7_75t_L g6842 ( 
.A(n_6699),
.Y(n_6842)
);

AND2x2_ASAP7_75t_L g6843 ( 
.A(n_6590),
.B(n_615),
.Y(n_6843)
);

INVx1_ASAP7_75t_L g6844 ( 
.A(n_6605),
.Y(n_6844)
);

INVx1_ASAP7_75t_L g6845 ( 
.A(n_6605),
.Y(n_6845)
);

INVx1_ASAP7_75t_L g6846 ( 
.A(n_6605),
.Y(n_6846)
);

OR2x2_ASAP7_75t_L g6847 ( 
.A(n_6593),
.B(n_616),
.Y(n_6847)
);

NOR2xp33_ASAP7_75t_L g6848 ( 
.A(n_6629),
.B(n_617),
.Y(n_6848)
);

NAND2xp5_ASAP7_75t_L g6849 ( 
.A(n_6621),
.B(n_617),
.Y(n_6849)
);

NAND2xp5_ASAP7_75t_L g6850 ( 
.A(n_6621),
.B(n_618),
.Y(n_6850)
);

AND2x4_ASAP7_75t_L g6851 ( 
.A(n_6699),
.B(n_618),
.Y(n_6851)
);

BUFx2_ASAP7_75t_L g6852 ( 
.A(n_6629),
.Y(n_6852)
);

INVx1_ASAP7_75t_L g6853 ( 
.A(n_6605),
.Y(n_6853)
);

AND2x4_ASAP7_75t_L g6854 ( 
.A(n_6699),
.B(n_619),
.Y(n_6854)
);

INVx1_ASAP7_75t_L g6855 ( 
.A(n_6605),
.Y(n_6855)
);

NOR2xp33_ASAP7_75t_L g6856 ( 
.A(n_6629),
.B(n_619),
.Y(n_6856)
);

AND2x2_ASAP7_75t_L g6857 ( 
.A(n_6590),
.B(n_620),
.Y(n_6857)
);

AND2x2_ASAP7_75t_L g6858 ( 
.A(n_6590),
.B(n_620),
.Y(n_6858)
);

AND2x2_ASAP7_75t_L g6859 ( 
.A(n_6590),
.B(n_621),
.Y(n_6859)
);

INVxp67_ASAP7_75t_SL g6860 ( 
.A(n_6605),
.Y(n_6860)
);

NAND2xp5_ASAP7_75t_L g6861 ( 
.A(n_6621),
.B(n_621),
.Y(n_6861)
);

INVx1_ASAP7_75t_L g6862 ( 
.A(n_6605),
.Y(n_6862)
);

AND2x2_ASAP7_75t_L g6863 ( 
.A(n_6590),
.B(n_622),
.Y(n_6863)
);

INVx1_ASAP7_75t_L g6864 ( 
.A(n_6605),
.Y(n_6864)
);

AOI22xp5_ASAP7_75t_L g6865 ( 
.A1(n_6610),
.A2(n_624),
.B1(n_622),
.B2(n_623),
.Y(n_6865)
);

INVx2_ASAP7_75t_SL g6866 ( 
.A(n_6596),
.Y(n_6866)
);

INVx2_ASAP7_75t_L g6867 ( 
.A(n_6699),
.Y(n_6867)
);

INVx1_ASAP7_75t_L g6868 ( 
.A(n_6605),
.Y(n_6868)
);

NAND2xp5_ASAP7_75t_SL g6869 ( 
.A(n_6621),
.B(n_625),
.Y(n_6869)
);

INVxp67_ASAP7_75t_L g6870 ( 
.A(n_6605),
.Y(n_6870)
);

NOR2xp33_ASAP7_75t_L g6871 ( 
.A(n_6629),
.B(n_625),
.Y(n_6871)
);

INVx1_ASAP7_75t_SL g6872 ( 
.A(n_6629),
.Y(n_6872)
);

AND2x4_ASAP7_75t_L g6873 ( 
.A(n_6699),
.B(n_626),
.Y(n_6873)
);

NAND2xp5_ASAP7_75t_L g6874 ( 
.A(n_6621),
.B(n_626),
.Y(n_6874)
);

AND2x2_ASAP7_75t_L g6875 ( 
.A(n_6590),
.B(n_628),
.Y(n_6875)
);

AND2x2_ASAP7_75t_L g6876 ( 
.A(n_6590),
.B(n_629),
.Y(n_6876)
);

OR2x2_ASAP7_75t_L g6877 ( 
.A(n_6593),
.B(n_630),
.Y(n_6877)
);

INVx1_ASAP7_75t_L g6878 ( 
.A(n_6605),
.Y(n_6878)
);

INVx1_ASAP7_75t_SL g6879 ( 
.A(n_6629),
.Y(n_6879)
);

NAND2x1_ASAP7_75t_L g6880 ( 
.A(n_6598),
.B(n_630),
.Y(n_6880)
);

INVx1_ASAP7_75t_L g6881 ( 
.A(n_6605),
.Y(n_6881)
);

CKINVDCx5p33_ASAP7_75t_R g6882 ( 
.A(n_6629),
.Y(n_6882)
);

INVxp67_ASAP7_75t_L g6883 ( 
.A(n_6605),
.Y(n_6883)
);

OR2x2_ASAP7_75t_L g6884 ( 
.A(n_6593),
.B(n_631),
.Y(n_6884)
);

NAND2xp5_ASAP7_75t_L g6885 ( 
.A(n_6621),
.B(n_631),
.Y(n_6885)
);

AND2x2_ASAP7_75t_L g6886 ( 
.A(n_6590),
.B(n_632),
.Y(n_6886)
);

INVxp67_ASAP7_75t_L g6887 ( 
.A(n_6605),
.Y(n_6887)
);

INVx1_ASAP7_75t_L g6888 ( 
.A(n_6605),
.Y(n_6888)
);

AND2x2_ASAP7_75t_L g6889 ( 
.A(n_6590),
.B(n_632),
.Y(n_6889)
);

INVx1_ASAP7_75t_L g6890 ( 
.A(n_6605),
.Y(n_6890)
);

NOR3xp33_ASAP7_75t_L g6891 ( 
.A(n_6604),
.B(n_634),
.C(n_636),
.Y(n_6891)
);

NAND2xp5_ASAP7_75t_L g6892 ( 
.A(n_6621),
.B(n_634),
.Y(n_6892)
);

AND2x4_ASAP7_75t_L g6893 ( 
.A(n_6699),
.B(n_636),
.Y(n_6893)
);

OR2x2_ASAP7_75t_L g6894 ( 
.A(n_6593),
.B(n_637),
.Y(n_6894)
);

OR2x2_ASAP7_75t_L g6895 ( 
.A(n_6593),
.B(n_638),
.Y(n_6895)
);

NAND2xp5_ASAP7_75t_L g6896 ( 
.A(n_6621),
.B(n_638),
.Y(n_6896)
);

INVx1_ASAP7_75t_L g6897 ( 
.A(n_6605),
.Y(n_6897)
);

NAND2x1p5_ASAP7_75t_L g6898 ( 
.A(n_6696),
.B(n_639),
.Y(n_6898)
);

INVx1_ASAP7_75t_L g6899 ( 
.A(n_6605),
.Y(n_6899)
);

AND2x2_ASAP7_75t_L g6900 ( 
.A(n_6590),
.B(n_639),
.Y(n_6900)
);

AND2x2_ASAP7_75t_L g6901 ( 
.A(n_6590),
.B(n_640),
.Y(n_6901)
);

AND2x2_ASAP7_75t_L g6902 ( 
.A(n_6590),
.B(n_640),
.Y(n_6902)
);

INVx1_ASAP7_75t_L g6903 ( 
.A(n_6605),
.Y(n_6903)
);

INVx1_ASAP7_75t_L g6904 ( 
.A(n_6605),
.Y(n_6904)
);

NAND4xp25_ASAP7_75t_SL g6905 ( 
.A(n_6619),
.B(n_643),
.C(n_641),
.D(n_642),
.Y(n_6905)
);

NAND2xp5_ASAP7_75t_L g6906 ( 
.A(n_6715),
.B(n_641),
.Y(n_6906)
);

INVxp67_ASAP7_75t_SL g6907 ( 
.A(n_6841),
.Y(n_6907)
);

AOI22xp5_ASAP7_75t_L g6908 ( 
.A1(n_6882),
.A2(n_646),
.B1(n_644),
.B2(n_645),
.Y(n_6908)
);

OAI22xp5_ASAP7_75t_L g6909 ( 
.A1(n_6787),
.A2(n_6747),
.B1(n_6737),
.B2(n_6829),
.Y(n_6909)
);

HB1xp67_ASAP7_75t_L g6910 ( 
.A(n_6783),
.Y(n_6910)
);

AOI21xp5_ASAP7_75t_L g6911 ( 
.A1(n_6869),
.A2(n_644),
.B(n_647),
.Y(n_6911)
);

NOR2xp33_ASAP7_75t_L g6912 ( 
.A(n_6872),
.B(n_648),
.Y(n_6912)
);

OR2x2_ASAP7_75t_L g6913 ( 
.A(n_6732),
.B(n_648),
.Y(n_6913)
);

INVx1_ASAP7_75t_L g6914 ( 
.A(n_6738),
.Y(n_6914)
);

INVx2_ASAP7_75t_L g6915 ( 
.A(n_6852),
.Y(n_6915)
);

NAND3xp33_ASAP7_75t_SL g6916 ( 
.A(n_6891),
.B(n_649),
.C(n_650),
.Y(n_6916)
);

INVx2_ASAP7_75t_L g6917 ( 
.A(n_6773),
.Y(n_6917)
);

OR2x2_ASAP7_75t_L g6918 ( 
.A(n_6719),
.B(n_651),
.Y(n_6918)
);

NAND2xp5_ASAP7_75t_L g6919 ( 
.A(n_6879),
.B(n_651),
.Y(n_6919)
);

INVx2_ASAP7_75t_L g6920 ( 
.A(n_6880),
.Y(n_6920)
);

INVx1_ASAP7_75t_SL g6921 ( 
.A(n_6745),
.Y(n_6921)
);

AND2x2_ASAP7_75t_L g6922 ( 
.A(n_6723),
.B(n_6866),
.Y(n_6922)
);

INVxp67_ASAP7_75t_L g6923 ( 
.A(n_6757),
.Y(n_6923)
);

NAND2xp5_ASAP7_75t_L g6924 ( 
.A(n_6860),
.B(n_652),
.Y(n_6924)
);

NOR2xp67_ASAP7_75t_L g6925 ( 
.A(n_6817),
.B(n_652),
.Y(n_6925)
);

OAI221xp5_ASAP7_75t_SL g6926 ( 
.A1(n_6870),
.A2(n_655),
.B1(n_653),
.B2(n_654),
.C(n_656),
.Y(n_6926)
);

OAI221xp5_ASAP7_75t_L g6927 ( 
.A1(n_6883),
.A2(n_655),
.B1(n_653),
.B2(n_654),
.C(n_656),
.Y(n_6927)
);

INVxp67_ASAP7_75t_L g6928 ( 
.A(n_6848),
.Y(n_6928)
);

NAND2xp5_ASAP7_75t_SL g6929 ( 
.A(n_6824),
.B(n_657),
.Y(n_6929)
);

AOI22xp33_ASAP7_75t_SL g6930 ( 
.A1(n_6800),
.A2(n_659),
.B1(n_657),
.B2(n_658),
.Y(n_6930)
);

INVxp67_ASAP7_75t_L g6931 ( 
.A(n_6856),
.Y(n_6931)
);

INVx2_ASAP7_75t_L g6932 ( 
.A(n_6748),
.Y(n_6932)
);

BUFx2_ASAP7_75t_L g6933 ( 
.A(n_6767),
.Y(n_6933)
);

OAI22xp33_ASAP7_75t_L g6934 ( 
.A1(n_6847),
.A2(n_661),
.B1(n_659),
.B2(n_660),
.Y(n_6934)
);

AND2x2_ASAP7_75t_L g6935 ( 
.A(n_6796),
.B(n_660),
.Y(n_6935)
);

OAI22xp33_ASAP7_75t_L g6936 ( 
.A1(n_6877),
.A2(n_664),
.B1(n_662),
.B2(n_663),
.Y(n_6936)
);

NOR2x1_ASAP7_75t_L g6937 ( 
.A(n_6740),
.B(n_662),
.Y(n_6937)
);

OAI21xp5_ASAP7_75t_SL g6938 ( 
.A1(n_6764),
.A2(n_663),
.B(n_665),
.Y(n_6938)
);

AOI22xp5_ASAP7_75t_L g6939 ( 
.A1(n_6905),
.A2(n_668),
.B1(n_665),
.B2(n_667),
.Y(n_6939)
);

OAI21xp5_ASAP7_75t_L g6940 ( 
.A1(n_6741),
.A2(n_672),
.B(n_671),
.Y(n_6940)
);

AOI21xp33_ASAP7_75t_L g6941 ( 
.A1(n_6887),
.A2(n_669),
.B(n_671),
.Y(n_6941)
);

AND2x2_ASAP7_75t_L g6942 ( 
.A(n_6725),
.B(n_6839),
.Y(n_6942)
);

NAND2xp5_ASAP7_75t_SL g6943 ( 
.A(n_6884),
.B(n_669),
.Y(n_6943)
);

NOR3xp33_ASAP7_75t_L g6944 ( 
.A(n_6746),
.B(n_672),
.C(n_673),
.Y(n_6944)
);

INVx1_ASAP7_75t_L g6945 ( 
.A(n_6739),
.Y(n_6945)
);

OR2x2_ASAP7_75t_L g6946 ( 
.A(n_6717),
.B(n_6837),
.Y(n_6946)
);

OAI22xp5_ASAP7_75t_SL g6947 ( 
.A1(n_6894),
.A2(n_675),
.B1(n_673),
.B2(n_674),
.Y(n_6947)
);

NAND2xp5_ASAP7_75t_L g6948 ( 
.A(n_6843),
.B(n_6857),
.Y(n_6948)
);

INVx1_ASAP7_75t_L g6949 ( 
.A(n_6744),
.Y(n_6949)
);

INVx1_ASAP7_75t_L g6950 ( 
.A(n_6858),
.Y(n_6950)
);

INVx1_ASAP7_75t_L g6951 ( 
.A(n_6859),
.Y(n_6951)
);

AND2x2_ASAP7_75t_L g6952 ( 
.A(n_6863),
.B(n_675),
.Y(n_6952)
);

NAND2xp33_ASAP7_75t_SL g6953 ( 
.A(n_6895),
.B(n_6838),
.Y(n_6953)
);

INVx1_ASAP7_75t_L g6954 ( 
.A(n_6875),
.Y(n_6954)
);

XOR2x2_ASAP7_75t_L g6955 ( 
.A(n_6760),
.B(n_6794),
.Y(n_6955)
);

AOI22xp5_ASAP7_75t_L g6956 ( 
.A1(n_6721),
.A2(n_678),
.B1(n_676),
.B2(n_677),
.Y(n_6956)
);

NAND2xp5_ASAP7_75t_L g6957 ( 
.A(n_6876),
.B(n_676),
.Y(n_6957)
);

OAI221xp5_ASAP7_75t_L g6958 ( 
.A1(n_6849),
.A2(n_681),
.B1(n_679),
.B2(n_680),
.C(n_682),
.Y(n_6958)
);

INVx1_ASAP7_75t_L g6959 ( 
.A(n_6886),
.Y(n_6959)
);

INVx2_ASAP7_75t_SL g6960 ( 
.A(n_6734),
.Y(n_6960)
);

INVx1_ASAP7_75t_L g6961 ( 
.A(n_6889),
.Y(n_6961)
);

INVxp67_ASAP7_75t_L g6962 ( 
.A(n_6871),
.Y(n_6962)
);

AOI22xp5_ASAP7_75t_L g6963 ( 
.A1(n_6718),
.A2(n_685),
.B1(n_683),
.B2(n_684),
.Y(n_6963)
);

AND2x2_ASAP7_75t_L g6964 ( 
.A(n_6900),
.B(n_683),
.Y(n_6964)
);

OAI22xp5_ASAP7_75t_L g6965 ( 
.A1(n_6865),
.A2(n_688),
.B1(n_686),
.B2(n_687),
.Y(n_6965)
);

AOI22xp33_ASAP7_75t_SL g6966 ( 
.A1(n_6726),
.A2(n_6844),
.B1(n_6845),
.B2(n_6720),
.Y(n_6966)
);

INVx1_ASAP7_75t_L g6967 ( 
.A(n_6901),
.Y(n_6967)
);

OAI22xp5_ASAP7_75t_L g6968 ( 
.A1(n_6850),
.A2(n_689),
.B1(n_686),
.B2(n_687),
.Y(n_6968)
);

OR2x2_ASAP7_75t_L g6969 ( 
.A(n_6861),
.B(n_690),
.Y(n_6969)
);

OAI22xp5_ASAP7_75t_L g6970 ( 
.A1(n_6874),
.A2(n_693),
.B1(n_690),
.B2(n_691),
.Y(n_6970)
);

INVxp67_ASAP7_75t_SL g6971 ( 
.A(n_6716),
.Y(n_6971)
);

INVx1_ASAP7_75t_L g6972 ( 
.A(n_6902),
.Y(n_6972)
);

NAND2xp5_ASAP7_75t_L g6973 ( 
.A(n_6750),
.B(n_691),
.Y(n_6973)
);

AOI22xp33_ASAP7_75t_L g6974 ( 
.A1(n_6840),
.A2(n_696),
.B1(n_694),
.B2(n_695),
.Y(n_6974)
);

INVx1_ASAP7_75t_L g6975 ( 
.A(n_6758),
.Y(n_6975)
);

NOR2xp33_ASAP7_75t_L g6976 ( 
.A(n_6790),
.B(n_694),
.Y(n_6976)
);

OAI21xp33_ASAP7_75t_L g6977 ( 
.A1(n_6842),
.A2(n_695),
.B(n_696),
.Y(n_6977)
);

INVx1_ASAP7_75t_SL g6978 ( 
.A(n_6885),
.Y(n_6978)
);

NAND2xp5_ASAP7_75t_L g6979 ( 
.A(n_6722),
.B(n_697),
.Y(n_6979)
);

NOR2xp33_ASAP7_75t_L g6980 ( 
.A(n_6892),
.B(n_698),
.Y(n_6980)
);

NAND2xp5_ASAP7_75t_L g6981 ( 
.A(n_6736),
.B(n_698),
.Y(n_6981)
);

INVxp67_ASAP7_75t_SL g6982 ( 
.A(n_6898),
.Y(n_6982)
);

OAI31xp33_ASAP7_75t_L g6983 ( 
.A1(n_6896),
.A2(n_701),
.A3(n_699),
.B(n_700),
.Y(n_6983)
);

AND2x2_ASAP7_75t_L g6984 ( 
.A(n_6785),
.B(n_701),
.Y(n_6984)
);

INVx1_ASAP7_75t_L g6985 ( 
.A(n_6795),
.Y(n_6985)
);

AOI22xp5_ASAP7_75t_L g6986 ( 
.A1(n_6867),
.A2(n_705),
.B1(n_703),
.B2(n_704),
.Y(n_6986)
);

OAI21xp33_ASAP7_75t_SL g6987 ( 
.A1(n_6846),
.A2(n_704),
.B(n_706),
.Y(n_6987)
);

NAND2xp5_ASAP7_75t_L g6988 ( 
.A(n_6815),
.B(n_707),
.Y(n_6988)
);

AOI222xp33_ASAP7_75t_L g6989 ( 
.A1(n_6853),
.A2(n_709),
.B1(n_711),
.B2(n_707),
.C1(n_708),
.C2(n_710),
.Y(n_6989)
);

AND2x2_ASAP7_75t_L g6990 ( 
.A(n_6735),
.B(n_709),
.Y(n_6990)
);

AOI322xp5_ASAP7_75t_L g6991 ( 
.A1(n_6855),
.A2(n_717),
.A3(n_716),
.B1(n_713),
.B2(n_710),
.C1(n_711),
.C2(n_714),
.Y(n_6991)
);

INVx1_ASAP7_75t_SL g6992 ( 
.A(n_6771),
.Y(n_6992)
);

OAI221xp5_ASAP7_75t_L g6993 ( 
.A1(n_6862),
.A2(n_716),
.B1(n_713),
.B2(n_714),
.C(n_718),
.Y(n_6993)
);

NAND2xp5_ASAP7_75t_L g6994 ( 
.A(n_6864),
.B(n_718),
.Y(n_6994)
);

INVx1_ASAP7_75t_L g6995 ( 
.A(n_6756),
.Y(n_6995)
);

OAI211xp5_ASAP7_75t_L g6996 ( 
.A1(n_6868),
.A2(n_721),
.B(n_719),
.C(n_720),
.Y(n_6996)
);

INVx1_ASAP7_75t_L g6997 ( 
.A(n_6743),
.Y(n_6997)
);

AOI22xp33_ASAP7_75t_SL g6998 ( 
.A1(n_6878),
.A2(n_725),
.B1(n_722),
.B2(n_723),
.Y(n_6998)
);

OAI22xp5_ASAP7_75t_L g6999 ( 
.A1(n_6810),
.A2(n_725),
.B1(n_722),
.B2(n_723),
.Y(n_6999)
);

OAI22xp5_ASAP7_75t_L g7000 ( 
.A1(n_6826),
.A2(n_728),
.B1(n_726),
.B2(n_727),
.Y(n_7000)
);

AND2x2_ASAP7_75t_L g7001 ( 
.A(n_6752),
.B(n_727),
.Y(n_7001)
);

OAI21xp5_ASAP7_75t_L g7002 ( 
.A1(n_6780),
.A2(n_6821),
.B(n_6881),
.Y(n_7002)
);

A2O1A1Ixp33_ASAP7_75t_L g7003 ( 
.A1(n_6805),
.A2(n_731),
.B(n_728),
.C(n_730),
.Y(n_7003)
);

AOI22xp5_ASAP7_75t_L g7004 ( 
.A1(n_6888),
.A2(n_733),
.B1(n_731),
.B2(n_732),
.Y(n_7004)
);

OAI22xp33_ASAP7_75t_SL g7005 ( 
.A1(n_6890),
.A2(n_734),
.B1(n_732),
.B2(n_733),
.Y(n_7005)
);

OAI221xp5_ASAP7_75t_L g7006 ( 
.A1(n_6897),
.A2(n_736),
.B1(n_734),
.B2(n_735),
.C(n_737),
.Y(n_7006)
);

INVx2_ASAP7_75t_L g7007 ( 
.A(n_6714),
.Y(n_7007)
);

INVx1_ASAP7_75t_L g7008 ( 
.A(n_6899),
.Y(n_7008)
);

NOR2xp33_ASAP7_75t_L g7009 ( 
.A(n_6724),
.B(n_6903),
.Y(n_7009)
);

AOI21xp33_ASAP7_75t_L g7010 ( 
.A1(n_6814),
.A2(n_735),
.B(n_736),
.Y(n_7010)
);

NAND2xp5_ASAP7_75t_L g7011 ( 
.A(n_6904),
.B(n_738),
.Y(n_7011)
);

INVx1_ASAP7_75t_L g7012 ( 
.A(n_6766),
.Y(n_7012)
);

OAI22xp33_ASAP7_75t_L g7013 ( 
.A1(n_6819),
.A2(n_740),
.B1(n_738),
.B2(n_739),
.Y(n_7013)
);

NAND3xp33_ASAP7_75t_L g7014 ( 
.A(n_6727),
.B(n_6729),
.C(n_6728),
.Y(n_7014)
);

AO22x1_ASAP7_75t_L g7015 ( 
.A1(n_6753),
.A2(n_748),
.B1(n_756),
.B2(n_739),
.Y(n_7015)
);

AOI22xp33_ASAP7_75t_L g7016 ( 
.A1(n_6807),
.A2(n_6833),
.B1(n_6791),
.B2(n_6802),
.Y(n_7016)
);

NAND2xp5_ASAP7_75t_L g7017 ( 
.A(n_6762),
.B(n_741),
.Y(n_7017)
);

INVx1_ASAP7_75t_L g7018 ( 
.A(n_6751),
.Y(n_7018)
);

OAI21xp33_ASAP7_75t_L g7019 ( 
.A1(n_6759),
.A2(n_741),
.B(n_742),
.Y(n_7019)
);

OAI22xp33_ASAP7_75t_L g7020 ( 
.A1(n_6831),
.A2(n_745),
.B1(n_743),
.B2(n_744),
.Y(n_7020)
);

AOI22xp5_ASAP7_75t_L g7021 ( 
.A1(n_6799),
.A2(n_746),
.B1(n_744),
.B2(n_745),
.Y(n_7021)
);

OAI21xp5_ASAP7_75t_SL g7022 ( 
.A1(n_6832),
.A2(n_747),
.B(n_748),
.Y(n_7022)
);

NAND2xp5_ASAP7_75t_L g7023 ( 
.A(n_6812),
.B(n_747),
.Y(n_7023)
);

INVx1_ASAP7_75t_SL g7024 ( 
.A(n_6778),
.Y(n_7024)
);

NAND2x1_ASAP7_75t_L g7025 ( 
.A(n_6792),
.B(n_749),
.Y(n_7025)
);

OAI22xp5_ASAP7_75t_L g7026 ( 
.A1(n_6813),
.A2(n_6820),
.B1(n_6763),
.B2(n_6765),
.Y(n_7026)
);

INVx2_ASAP7_75t_L g7027 ( 
.A(n_6851),
.Y(n_7027)
);

OAI21xp5_ASAP7_75t_SL g7028 ( 
.A1(n_6782),
.A2(n_750),
.B(n_751),
.Y(n_7028)
);

INVx1_ASAP7_75t_SL g7029 ( 
.A(n_6749),
.Y(n_7029)
);

AND2x2_ASAP7_75t_L g7030 ( 
.A(n_6816),
.B(n_750),
.Y(n_7030)
);

NOR2xp33_ASAP7_75t_L g7031 ( 
.A(n_6731),
.B(n_751),
.Y(n_7031)
);

INVx1_ASAP7_75t_L g7032 ( 
.A(n_6742),
.Y(n_7032)
);

INVx1_ASAP7_75t_L g7033 ( 
.A(n_6798),
.Y(n_7033)
);

INVx1_ASAP7_75t_L g7034 ( 
.A(n_6774),
.Y(n_7034)
);

AND2x4_ASAP7_75t_L g7035 ( 
.A(n_6786),
.B(n_752),
.Y(n_7035)
);

OAI21xp5_ASAP7_75t_L g7036 ( 
.A1(n_6755),
.A2(n_754),
.B(n_753),
.Y(n_7036)
);

OAI221xp5_ASAP7_75t_L g7037 ( 
.A1(n_6769),
.A2(n_757),
.B1(n_752),
.B2(n_755),
.C(n_758),
.Y(n_7037)
);

INVx1_ASAP7_75t_L g7038 ( 
.A(n_6775),
.Y(n_7038)
);

AND2x2_ASAP7_75t_L g7039 ( 
.A(n_6754),
.B(n_755),
.Y(n_7039)
);

AND2x4_ASAP7_75t_L g7040 ( 
.A(n_6730),
.B(n_759),
.Y(n_7040)
);

NAND2xp5_ASAP7_75t_SL g7041 ( 
.A(n_6772),
.B(n_759),
.Y(n_7041)
);

NAND2xp5_ASAP7_75t_SL g7042 ( 
.A(n_6733),
.B(n_760),
.Y(n_7042)
);

OAI21xp33_ASAP7_75t_L g7043 ( 
.A1(n_6788),
.A2(n_761),
.B(n_762),
.Y(n_7043)
);

OAI21xp5_ASAP7_75t_L g7044 ( 
.A1(n_6822),
.A2(n_764),
.B(n_763),
.Y(n_7044)
);

INVx1_ASAP7_75t_L g7045 ( 
.A(n_6761),
.Y(n_7045)
);

OR2x2_ASAP7_75t_L g7046 ( 
.A(n_6768),
.B(n_761),
.Y(n_7046)
);

O2A1O1Ixp33_ASAP7_75t_L g7047 ( 
.A1(n_6808),
.A2(n_765),
.B(n_763),
.C(n_764),
.Y(n_7047)
);

INVx1_ASAP7_75t_L g7048 ( 
.A(n_6776),
.Y(n_7048)
);

A2O1A1Ixp33_ASAP7_75t_L g7049 ( 
.A1(n_6797),
.A2(n_6835),
.B(n_6836),
.C(n_6823),
.Y(n_7049)
);

AOI21xp5_ASAP7_75t_L g7050 ( 
.A1(n_6806),
.A2(n_765),
.B(n_766),
.Y(n_7050)
);

OAI322xp33_ASAP7_75t_L g7051 ( 
.A1(n_6828),
.A2(n_771),
.A3(n_770),
.B1(n_768),
.B2(n_766),
.C1(n_767),
.C2(n_769),
.Y(n_7051)
);

INVx1_ASAP7_75t_SL g7052 ( 
.A(n_6933),
.Y(n_7052)
);

INVx1_ASAP7_75t_L g7053 ( 
.A(n_6910),
.Y(n_7053)
);

NAND2xp5_ASAP7_75t_L g7054 ( 
.A(n_6907),
.B(n_6825),
.Y(n_7054)
);

INVx1_ASAP7_75t_L g7055 ( 
.A(n_6925),
.Y(n_7055)
);

XOR2xp5_ASAP7_75t_L g7056 ( 
.A(n_6955),
.B(n_6781),
.Y(n_7056)
);

INVx1_ASAP7_75t_L g7057 ( 
.A(n_6922),
.Y(n_7057)
);

NAND2xp33_ASAP7_75t_SL g7058 ( 
.A(n_7025),
.B(n_6920),
.Y(n_7058)
);

NAND2xp5_ASAP7_75t_L g7059 ( 
.A(n_6921),
.B(n_6834),
.Y(n_7059)
);

AND2x2_ASAP7_75t_L g7060 ( 
.A(n_6917),
.B(n_6803),
.Y(n_7060)
);

INVx1_ASAP7_75t_SL g7061 ( 
.A(n_6913),
.Y(n_7061)
);

NAND2xp5_ASAP7_75t_L g7062 ( 
.A(n_6915),
.B(n_6914),
.Y(n_7062)
);

AOI21xp33_ASAP7_75t_SL g7063 ( 
.A1(n_6923),
.A2(n_6809),
.B(n_6827),
.Y(n_7063)
);

INVx2_ASAP7_75t_L g7064 ( 
.A(n_6942),
.Y(n_7064)
);

NOR2xp33_ASAP7_75t_L g7065 ( 
.A(n_6938),
.B(n_6777),
.Y(n_7065)
);

NAND2xp5_ASAP7_75t_L g7066 ( 
.A(n_7015),
.B(n_6779),
.Y(n_7066)
);

INVx1_ASAP7_75t_L g7067 ( 
.A(n_6935),
.Y(n_7067)
);

INVx2_ASAP7_75t_L g7068 ( 
.A(n_6952),
.Y(n_7068)
);

INVx1_ASAP7_75t_L g7069 ( 
.A(n_6964),
.Y(n_7069)
);

INVx1_ASAP7_75t_L g7070 ( 
.A(n_6984),
.Y(n_7070)
);

AND2x2_ASAP7_75t_L g7071 ( 
.A(n_6971),
.B(n_6830),
.Y(n_7071)
);

INVxp33_ASAP7_75t_L g7072 ( 
.A(n_6912),
.Y(n_7072)
);

INVx2_ASAP7_75t_L g7073 ( 
.A(n_7035),
.Y(n_7073)
);

NAND2x1p5_ASAP7_75t_L g7074 ( 
.A(n_6992),
.B(n_7024),
.Y(n_7074)
);

INVx1_ASAP7_75t_L g7075 ( 
.A(n_6906),
.Y(n_7075)
);

INVxp67_ASAP7_75t_SL g7076 ( 
.A(n_6929),
.Y(n_7076)
);

INVx1_ASAP7_75t_L g7077 ( 
.A(n_6919),
.Y(n_7077)
);

INVx1_ASAP7_75t_L g7078 ( 
.A(n_6948),
.Y(n_7078)
);

NAND2xp5_ASAP7_75t_L g7079 ( 
.A(n_6982),
.B(n_6804),
.Y(n_7079)
);

INVx1_ASAP7_75t_L g7080 ( 
.A(n_6918),
.Y(n_7080)
);

NAND2xp5_ASAP7_75t_L g7081 ( 
.A(n_6960),
.B(n_6801),
.Y(n_7081)
);

NAND2xp5_ASAP7_75t_L g7082 ( 
.A(n_6939),
.B(n_6793),
.Y(n_7082)
);

INVx1_ASAP7_75t_L g7083 ( 
.A(n_6990),
.Y(n_7083)
);

INVx1_ASAP7_75t_L g7084 ( 
.A(n_7001),
.Y(n_7084)
);

NOR2xp33_ASAP7_75t_L g7085 ( 
.A(n_6950),
.B(n_6784),
.Y(n_7085)
);

OR2x2_ASAP7_75t_L g7086 ( 
.A(n_6951),
.B(n_6818),
.Y(n_7086)
);

INVx2_ASAP7_75t_L g7087 ( 
.A(n_7035),
.Y(n_7087)
);

AND2x2_ASAP7_75t_L g7088 ( 
.A(n_7007),
.B(n_6854),
.Y(n_7088)
);

NAND2xp5_ASAP7_75t_L g7089 ( 
.A(n_6930),
.B(n_6873),
.Y(n_7089)
);

INVx1_ASAP7_75t_L g7090 ( 
.A(n_6924),
.Y(n_7090)
);

NAND2xp5_ASAP7_75t_L g7091 ( 
.A(n_6954),
.B(n_6959),
.Y(n_7091)
);

NAND2xp5_ASAP7_75t_L g7092 ( 
.A(n_6961),
.B(n_6893),
.Y(n_7092)
);

INVx2_ASAP7_75t_L g7093 ( 
.A(n_7027),
.Y(n_7093)
);

INVx1_ASAP7_75t_L g7094 ( 
.A(n_6967),
.Y(n_7094)
);

AND2x2_ASAP7_75t_L g7095 ( 
.A(n_6932),
.B(n_6770),
.Y(n_7095)
);

NAND3xp33_ASAP7_75t_L g7096 ( 
.A(n_6966),
.B(n_6811),
.C(n_6789),
.Y(n_7096)
);

OAI21xp5_ASAP7_75t_L g7097 ( 
.A1(n_6909),
.A2(n_767),
.B(n_769),
.Y(n_7097)
);

NAND2xp5_ASAP7_75t_L g7098 ( 
.A(n_6972),
.B(n_771),
.Y(n_7098)
);

OR2x2_ASAP7_75t_L g7099 ( 
.A(n_6985),
.B(n_6945),
.Y(n_7099)
);

AND2x2_ASAP7_75t_L g7100 ( 
.A(n_6949),
.B(n_772),
.Y(n_7100)
);

INVxp67_ASAP7_75t_SL g7101 ( 
.A(n_6947),
.Y(n_7101)
);

NAND2xp5_ASAP7_75t_L g7102 ( 
.A(n_6998),
.B(n_6975),
.Y(n_7102)
);

AND2x2_ASAP7_75t_L g7103 ( 
.A(n_6995),
.B(n_773),
.Y(n_7103)
);

AOI21xp33_ASAP7_75t_L g7104 ( 
.A1(n_7009),
.A2(n_774),
.B(n_775),
.Y(n_7104)
);

NAND2xp5_ASAP7_75t_L g7105 ( 
.A(n_7034),
.B(n_774),
.Y(n_7105)
);

NOR2xp33_ASAP7_75t_L g7106 ( 
.A(n_6928),
.B(n_775),
.Y(n_7106)
);

NAND2x1p5_ASAP7_75t_L g7107 ( 
.A(n_7032),
.B(n_776),
.Y(n_7107)
);

INVx1_ASAP7_75t_L g7108 ( 
.A(n_6957),
.Y(n_7108)
);

INVx1_ASAP7_75t_L g7109 ( 
.A(n_7040),
.Y(n_7109)
);

INVx1_ASAP7_75t_L g7110 ( 
.A(n_7040),
.Y(n_7110)
);

INVx1_ASAP7_75t_L g7111 ( 
.A(n_6981),
.Y(n_7111)
);

NAND2xp5_ASAP7_75t_L g7112 ( 
.A(n_7038),
.B(n_776),
.Y(n_7112)
);

INVx1_ASAP7_75t_L g7113 ( 
.A(n_7030),
.Y(n_7113)
);

INVx1_ASAP7_75t_L g7114 ( 
.A(n_6969),
.Y(n_7114)
);

AND2x2_ASAP7_75t_L g7115 ( 
.A(n_7002),
.B(n_777),
.Y(n_7115)
);

NAND3xp33_ASAP7_75t_L g7116 ( 
.A(n_6987),
.B(n_778),
.C(n_779),
.Y(n_7116)
);

INVx1_ASAP7_75t_L g7117 ( 
.A(n_6988),
.Y(n_7117)
);

INVx2_ASAP7_75t_SL g7118 ( 
.A(n_7039),
.Y(n_7118)
);

NAND2xp5_ASAP7_75t_L g7119 ( 
.A(n_6989),
.B(n_780),
.Y(n_7119)
);

NOR2xp33_ASAP7_75t_L g7120 ( 
.A(n_6931),
.B(n_781),
.Y(n_7120)
);

INVx1_ASAP7_75t_L g7121 ( 
.A(n_7017),
.Y(n_7121)
);

NAND2xp5_ASAP7_75t_L g7122 ( 
.A(n_7018),
.B(n_782),
.Y(n_7122)
);

NOR2xp33_ASAP7_75t_L g7123 ( 
.A(n_6962),
.B(n_783),
.Y(n_7123)
);

INVx1_ASAP7_75t_L g7124 ( 
.A(n_6946),
.Y(n_7124)
);

OR2x2_ASAP7_75t_L g7125 ( 
.A(n_6978),
.B(n_784),
.Y(n_7125)
);

NAND2xp5_ASAP7_75t_L g7126 ( 
.A(n_6934),
.B(n_784),
.Y(n_7126)
);

INVx1_ASAP7_75t_L g7127 ( 
.A(n_6979),
.Y(n_7127)
);

INVx1_ASAP7_75t_L g7128 ( 
.A(n_6976),
.Y(n_7128)
);

AND2x2_ASAP7_75t_L g7129 ( 
.A(n_6937),
.B(n_785),
.Y(n_7129)
);

NAND2xp33_ASAP7_75t_L g7130 ( 
.A(n_6944),
.B(n_785),
.Y(n_7130)
);

NAND2xp5_ASAP7_75t_L g7131 ( 
.A(n_6936),
.B(n_786),
.Y(n_7131)
);

INVx1_ASAP7_75t_L g7132 ( 
.A(n_7046),
.Y(n_7132)
);

NAND2x1p5_ASAP7_75t_L g7133 ( 
.A(n_6997),
.B(n_786),
.Y(n_7133)
);

OAI21xp5_ASAP7_75t_SL g7134 ( 
.A1(n_7016),
.A2(n_787),
.B(n_788),
.Y(n_7134)
);

NAND2xp5_ASAP7_75t_L g7135 ( 
.A(n_7012),
.B(n_788),
.Y(n_7135)
);

INVx2_ASAP7_75t_L g7136 ( 
.A(n_7033),
.Y(n_7136)
);

INVxp67_ASAP7_75t_L g7137 ( 
.A(n_6980),
.Y(n_7137)
);

INVx3_ASAP7_75t_L g7138 ( 
.A(n_7008),
.Y(n_7138)
);

INVx1_ASAP7_75t_SL g7139 ( 
.A(n_6953),
.Y(n_7139)
);

NOR2x1_ASAP7_75t_L g7140 ( 
.A(n_7022),
.B(n_789),
.Y(n_7140)
);

NOR2xp33_ASAP7_75t_L g7141 ( 
.A(n_6943),
.B(n_789),
.Y(n_7141)
);

NAND3xp33_ASAP7_75t_L g7142 ( 
.A(n_7014),
.B(n_792),
.C(n_793),
.Y(n_7142)
);

INVx1_ASAP7_75t_L g7143 ( 
.A(n_6994),
.Y(n_7143)
);

INVx1_ASAP7_75t_L g7144 ( 
.A(n_7011),
.Y(n_7144)
);

NAND2x1p5_ASAP7_75t_L g7145 ( 
.A(n_7042),
.B(n_794),
.Y(n_7145)
);

INVx1_ASAP7_75t_L g7146 ( 
.A(n_6973),
.Y(n_7146)
);

NAND2xp33_ASAP7_75t_L g7147 ( 
.A(n_7019),
.B(n_795),
.Y(n_7147)
);

CKINVDCx14_ASAP7_75t_R g7148 ( 
.A(n_7026),
.Y(n_7148)
);

NAND2xp5_ASAP7_75t_L g7149 ( 
.A(n_6956),
.B(n_7050),
.Y(n_7149)
);

AND2x2_ASAP7_75t_L g7150 ( 
.A(n_7029),
.B(n_795),
.Y(n_7150)
);

INVx1_ASAP7_75t_L g7151 ( 
.A(n_7023),
.Y(n_7151)
);

OR2x2_ASAP7_75t_L g7152 ( 
.A(n_6916),
.B(n_797),
.Y(n_7152)
);

INVx1_ASAP7_75t_L g7153 ( 
.A(n_7041),
.Y(n_7153)
);

AND2x2_ASAP7_75t_L g7154 ( 
.A(n_6940),
.B(n_797),
.Y(n_7154)
);

OR2x2_ASAP7_75t_L g7155 ( 
.A(n_7000),
.B(n_798),
.Y(n_7155)
);

INVx1_ASAP7_75t_SL g7156 ( 
.A(n_6911),
.Y(n_7156)
);

NAND2xp5_ASAP7_75t_L g7157 ( 
.A(n_7031),
.B(n_799),
.Y(n_7157)
);

AOI22xp33_ASAP7_75t_L g7158 ( 
.A1(n_7045),
.A2(n_802),
.B1(n_800),
.B2(n_801),
.Y(n_7158)
);

INVx1_ASAP7_75t_L g7159 ( 
.A(n_7005),
.Y(n_7159)
);

INVx2_ASAP7_75t_L g7160 ( 
.A(n_7048),
.Y(n_7160)
);

NAND2xp5_ASAP7_75t_SL g7161 ( 
.A(n_6983),
.B(n_800),
.Y(n_7161)
);

INVx1_ASAP7_75t_L g7162 ( 
.A(n_6977),
.Y(n_7162)
);

INVx1_ASAP7_75t_L g7163 ( 
.A(n_7004),
.Y(n_7163)
);

AND2x2_ASAP7_75t_L g7164 ( 
.A(n_7036),
.B(n_801),
.Y(n_7164)
);

NAND2x1p5_ASAP7_75t_L g7165 ( 
.A(n_6908),
.B(n_802),
.Y(n_7165)
);

OR2x2_ASAP7_75t_L g7166 ( 
.A(n_7049),
.B(n_804),
.Y(n_7166)
);

OR2x2_ASAP7_75t_L g7167 ( 
.A(n_7028),
.B(n_806),
.Y(n_7167)
);

INVx1_ASAP7_75t_L g7168 ( 
.A(n_6968),
.Y(n_7168)
);

INVx1_ASAP7_75t_L g7169 ( 
.A(n_6970),
.Y(n_7169)
);

NAND2xp5_ASAP7_75t_L g7170 ( 
.A(n_7003),
.B(n_7013),
.Y(n_7170)
);

AOI22xp33_ASAP7_75t_L g7171 ( 
.A1(n_7020),
.A2(n_809),
.B1(n_806),
.B2(n_807),
.Y(n_7171)
);

INVx1_ASAP7_75t_SL g7172 ( 
.A(n_7010),
.Y(n_7172)
);

INVx1_ASAP7_75t_L g7173 ( 
.A(n_6963),
.Y(n_7173)
);

INVx1_ASAP7_75t_L g7174 ( 
.A(n_6986),
.Y(n_7174)
);

HB1xp67_ASAP7_75t_L g7175 ( 
.A(n_7044),
.Y(n_7175)
);

INVx1_ASAP7_75t_L g7176 ( 
.A(n_7021),
.Y(n_7176)
);

INVx2_ASAP7_75t_L g7177 ( 
.A(n_6993),
.Y(n_7177)
);

NAND2xp5_ASAP7_75t_L g7178 ( 
.A(n_7043),
.B(n_807),
.Y(n_7178)
);

INVx1_ASAP7_75t_L g7179 ( 
.A(n_6996),
.Y(n_7179)
);

NAND2xp5_ASAP7_75t_L g7180 ( 
.A(n_6991),
.B(n_810),
.Y(n_7180)
);

INVx1_ASAP7_75t_L g7181 ( 
.A(n_6999),
.Y(n_7181)
);

OR2x2_ASAP7_75t_L g7182 ( 
.A(n_6926),
.B(n_810),
.Y(n_7182)
);

NAND2xp5_ASAP7_75t_L g7183 ( 
.A(n_6965),
.B(n_811),
.Y(n_7183)
);

NAND2xp5_ASAP7_75t_L g7184 ( 
.A(n_6974),
.B(n_811),
.Y(n_7184)
);

INVx1_ASAP7_75t_L g7185 ( 
.A(n_7051),
.Y(n_7185)
);

BUFx2_ASAP7_75t_L g7186 ( 
.A(n_6941),
.Y(n_7186)
);

OAI22xp33_ASAP7_75t_L g7187 ( 
.A1(n_6958),
.A2(n_814),
.B1(n_812),
.B2(n_813),
.Y(n_7187)
);

OR2x2_ASAP7_75t_L g7188 ( 
.A(n_6927),
.B(n_812),
.Y(n_7188)
);

NOR2x1_ASAP7_75t_L g7189 ( 
.A(n_7047),
.B(n_813),
.Y(n_7189)
);

INVx1_ASAP7_75t_SL g7190 ( 
.A(n_7006),
.Y(n_7190)
);

INVx1_ASAP7_75t_L g7191 ( 
.A(n_7037),
.Y(n_7191)
);

NOR2xp67_ASAP7_75t_L g7192 ( 
.A(n_6910),
.B(n_814),
.Y(n_7192)
);

INVx2_ASAP7_75t_L g7193 ( 
.A(n_6933),
.Y(n_7193)
);

NOR2xp33_ASAP7_75t_L g7194 ( 
.A(n_6910),
.B(n_815),
.Y(n_7194)
);

AND2x2_ASAP7_75t_L g7195 ( 
.A(n_6922),
.B(n_816),
.Y(n_7195)
);

INVx1_ASAP7_75t_L g7196 ( 
.A(n_6910),
.Y(n_7196)
);

NAND2xp5_ASAP7_75t_L g7197 ( 
.A(n_6907),
.B(n_817),
.Y(n_7197)
);

INVx1_ASAP7_75t_L g7198 ( 
.A(n_6910),
.Y(n_7198)
);

NOR2x1_ASAP7_75t_L g7199 ( 
.A(n_6925),
.B(n_817),
.Y(n_7199)
);

NAND2xp5_ASAP7_75t_L g7200 ( 
.A(n_6907),
.B(n_818),
.Y(n_7200)
);

NAND2xp5_ASAP7_75t_L g7201 ( 
.A(n_6907),
.B(n_818),
.Y(n_7201)
);

INVx1_ASAP7_75t_L g7202 ( 
.A(n_6910),
.Y(n_7202)
);

AOI22xp5_ASAP7_75t_L g7203 ( 
.A1(n_6909),
.A2(n_821),
.B1(n_819),
.B2(n_820),
.Y(n_7203)
);

INVx1_ASAP7_75t_L g7204 ( 
.A(n_6910),
.Y(n_7204)
);

INVx1_ASAP7_75t_L g7205 ( 
.A(n_6910),
.Y(n_7205)
);

NAND2xp5_ASAP7_75t_L g7206 ( 
.A(n_6907),
.B(n_821),
.Y(n_7206)
);

INVx1_ASAP7_75t_L g7207 ( 
.A(n_6910),
.Y(n_7207)
);

INVx1_ASAP7_75t_L g7208 ( 
.A(n_6910),
.Y(n_7208)
);

NAND2xp5_ASAP7_75t_L g7209 ( 
.A(n_6907),
.B(n_822),
.Y(n_7209)
);

NAND2xp5_ASAP7_75t_L g7210 ( 
.A(n_6907),
.B(n_822),
.Y(n_7210)
);

NAND2x1p5_ASAP7_75t_L g7211 ( 
.A(n_7025),
.B(n_823),
.Y(n_7211)
);

INVx1_ASAP7_75t_L g7212 ( 
.A(n_6910),
.Y(n_7212)
);

INVx1_ASAP7_75t_L g7213 ( 
.A(n_6910),
.Y(n_7213)
);

INVx1_ASAP7_75t_L g7214 ( 
.A(n_6910),
.Y(n_7214)
);

INVx1_ASAP7_75t_L g7215 ( 
.A(n_6910),
.Y(n_7215)
);

INVx2_ASAP7_75t_L g7216 ( 
.A(n_7211),
.Y(n_7216)
);

INVx1_ASAP7_75t_L g7217 ( 
.A(n_7199),
.Y(n_7217)
);

OR2x2_ASAP7_75t_L g7218 ( 
.A(n_7074),
.B(n_823),
.Y(n_7218)
);

INVx1_ASAP7_75t_L g7219 ( 
.A(n_7192),
.Y(n_7219)
);

INVx1_ASAP7_75t_L g7220 ( 
.A(n_7066),
.Y(n_7220)
);

AOI21xp33_ASAP7_75t_SL g7221 ( 
.A1(n_7055),
.A2(n_827),
.B(n_826),
.Y(n_7221)
);

XNOR2xp5_ASAP7_75t_L g7222 ( 
.A(n_7056),
.B(n_826),
.Y(n_7222)
);

INVx1_ASAP7_75t_L g7223 ( 
.A(n_7195),
.Y(n_7223)
);

A2O1A1Ixp33_ASAP7_75t_L g7224 ( 
.A1(n_7148),
.A2(n_828),
.B(n_830),
.C(n_827),
.Y(n_7224)
);

INVx1_ASAP7_75t_L g7225 ( 
.A(n_7133),
.Y(n_7225)
);

XNOR2xp5_ASAP7_75t_L g7226 ( 
.A(n_7096),
.B(n_828),
.Y(n_7226)
);

NOR3xp33_ASAP7_75t_SL g7227 ( 
.A(n_7058),
.B(n_825),
.C(n_831),
.Y(n_7227)
);

NAND2xp5_ASAP7_75t_L g7228 ( 
.A(n_7052),
.B(n_831),
.Y(n_7228)
);

NAND2xp5_ASAP7_75t_L g7229 ( 
.A(n_7073),
.B(n_832),
.Y(n_7229)
);

INVx1_ASAP7_75t_L g7230 ( 
.A(n_7107),
.Y(n_7230)
);

INVx1_ASAP7_75t_L g7231 ( 
.A(n_7087),
.Y(n_7231)
);

NAND2xp5_ASAP7_75t_L g7232 ( 
.A(n_7109),
.B(n_832),
.Y(n_7232)
);

NAND2xp5_ASAP7_75t_SL g7233 ( 
.A(n_7193),
.B(n_833),
.Y(n_7233)
);

INVx1_ASAP7_75t_L g7234 ( 
.A(n_7110),
.Y(n_7234)
);

INVx1_ASAP7_75t_L g7235 ( 
.A(n_7071),
.Y(n_7235)
);

NAND2xp5_ASAP7_75t_L g7236 ( 
.A(n_7101),
.B(n_833),
.Y(n_7236)
);

INVx2_ASAP7_75t_L g7237 ( 
.A(n_7064),
.Y(n_7237)
);

AOI221xp5_ASAP7_75t_L g7238 ( 
.A1(n_7185),
.A2(n_7159),
.B1(n_7179),
.B2(n_7115),
.C(n_7097),
.Y(n_7238)
);

AND2x2_ASAP7_75t_L g7239 ( 
.A(n_7088),
.B(n_834),
.Y(n_7239)
);

INVx1_ASAP7_75t_L g7240 ( 
.A(n_7057),
.Y(n_7240)
);

NAND2xp5_ASAP7_75t_L g7241 ( 
.A(n_7053),
.B(n_834),
.Y(n_7241)
);

NAND2xp5_ASAP7_75t_L g7242 ( 
.A(n_7196),
.B(n_835),
.Y(n_7242)
);

NAND3xp33_ASAP7_75t_L g7243 ( 
.A(n_7116),
.B(n_836),
.C(n_837),
.Y(n_7243)
);

INVx1_ASAP7_75t_L g7244 ( 
.A(n_7059),
.Y(n_7244)
);

INVx3_ASAP7_75t_L g7245 ( 
.A(n_7138),
.Y(n_7245)
);

XNOR2x2_ASAP7_75t_L g7246 ( 
.A(n_7142),
.B(n_836),
.Y(n_7246)
);

AND2x2_ASAP7_75t_L g7247 ( 
.A(n_7060),
.B(n_837),
.Y(n_7247)
);

NAND2xp33_ASAP7_75t_L g7248 ( 
.A(n_7140),
.B(n_839),
.Y(n_7248)
);

NOR3xp33_ASAP7_75t_SL g7249 ( 
.A(n_7062),
.B(n_840),
.C(n_841),
.Y(n_7249)
);

NAND2xp33_ASAP7_75t_R g7250 ( 
.A(n_7138),
.B(n_840),
.Y(n_7250)
);

INVx2_ASAP7_75t_L g7251 ( 
.A(n_7145),
.Y(n_7251)
);

NAND2xp5_ASAP7_75t_L g7252 ( 
.A(n_7198),
.B(n_841),
.Y(n_7252)
);

AOI31xp33_ASAP7_75t_L g7253 ( 
.A1(n_7072),
.A2(n_844),
.A3(n_845),
.B(n_843),
.Y(n_7253)
);

CKINVDCx14_ASAP7_75t_R g7254 ( 
.A(n_7186),
.Y(n_7254)
);

INVx2_ASAP7_75t_L g7255 ( 
.A(n_7099),
.Y(n_7255)
);

NOR4xp25_ASAP7_75t_SL g7256 ( 
.A(n_7161),
.B(n_845),
.C(n_842),
.D(n_843),
.Y(n_7256)
);

NAND2xp5_ASAP7_75t_SL g7257 ( 
.A(n_7063),
.B(n_846),
.Y(n_7257)
);

NOR2xp33_ASAP7_75t_L g7258 ( 
.A(n_7061),
.B(n_848),
.Y(n_7258)
);

OR2x2_ASAP7_75t_L g7259 ( 
.A(n_7089),
.B(n_848),
.Y(n_7259)
);

INVx1_ASAP7_75t_L g7260 ( 
.A(n_7202),
.Y(n_7260)
);

NAND2xp5_ASAP7_75t_L g7261 ( 
.A(n_7204),
.B(n_849),
.Y(n_7261)
);

INVx2_ASAP7_75t_L g7262 ( 
.A(n_7205),
.Y(n_7262)
);

NAND2x1p5_ASAP7_75t_SL g7263 ( 
.A(n_7118),
.B(n_850),
.Y(n_7263)
);

NAND2xp5_ASAP7_75t_SL g7264 ( 
.A(n_7139),
.B(n_851),
.Y(n_7264)
);

INVx2_ASAP7_75t_L g7265 ( 
.A(n_7207),
.Y(n_7265)
);

INVx1_ASAP7_75t_L g7266 ( 
.A(n_7208),
.Y(n_7266)
);

OR2x2_ASAP7_75t_L g7267 ( 
.A(n_7212),
.B(n_851),
.Y(n_7267)
);

XNOR2xp5_ASAP7_75t_L g7268 ( 
.A(n_7190),
.B(n_853),
.Y(n_7268)
);

INVx1_ASAP7_75t_L g7269 ( 
.A(n_7213),
.Y(n_7269)
);

AND2x2_ASAP7_75t_L g7270 ( 
.A(n_7093),
.B(n_852),
.Y(n_7270)
);

CKINVDCx20_ASAP7_75t_R g7271 ( 
.A(n_7082),
.Y(n_7271)
);

INVx1_ASAP7_75t_L g7272 ( 
.A(n_7214),
.Y(n_7272)
);

NOR2xp33_ASAP7_75t_L g7273 ( 
.A(n_7215),
.B(n_852),
.Y(n_7273)
);

INVx1_ASAP7_75t_L g7274 ( 
.A(n_7100),
.Y(n_7274)
);

INVxp67_ASAP7_75t_L g7275 ( 
.A(n_7194),
.Y(n_7275)
);

INVx1_ASAP7_75t_L g7276 ( 
.A(n_7103),
.Y(n_7276)
);

INVx1_ASAP7_75t_SL g7277 ( 
.A(n_7129),
.Y(n_7277)
);

INVx1_ASAP7_75t_L g7278 ( 
.A(n_7054),
.Y(n_7278)
);

INVx1_ASAP7_75t_L g7279 ( 
.A(n_7092),
.Y(n_7279)
);

XOR2x2_ASAP7_75t_L g7280 ( 
.A(n_7189),
.B(n_854),
.Y(n_7280)
);

NAND2xp5_ASAP7_75t_L g7281 ( 
.A(n_7067),
.B(n_854),
.Y(n_7281)
);

AOI21xp5_ASAP7_75t_L g7282 ( 
.A1(n_7079),
.A2(n_855),
.B(n_856),
.Y(n_7282)
);

INVx1_ASAP7_75t_L g7283 ( 
.A(n_7197),
.Y(n_7283)
);

INVx1_ASAP7_75t_L g7284 ( 
.A(n_7200),
.Y(n_7284)
);

NAND2xp5_ASAP7_75t_L g7285 ( 
.A(n_7069),
.B(n_855),
.Y(n_7285)
);

NAND2xp5_ASAP7_75t_SL g7286 ( 
.A(n_7136),
.B(n_857),
.Y(n_7286)
);

CKINVDCx5p33_ASAP7_75t_R g7287 ( 
.A(n_7172),
.Y(n_7287)
);

NOR3xp33_ASAP7_75t_L g7288 ( 
.A(n_7091),
.B(n_868),
.C(n_857),
.Y(n_7288)
);

AND2x2_ASAP7_75t_L g7289 ( 
.A(n_7068),
.B(n_7076),
.Y(n_7289)
);

INVx1_ASAP7_75t_L g7290 ( 
.A(n_7201),
.Y(n_7290)
);

AND2x2_ASAP7_75t_L g7291 ( 
.A(n_7095),
.B(n_858),
.Y(n_7291)
);

AND2x2_ASAP7_75t_L g7292 ( 
.A(n_7083),
.B(n_860),
.Y(n_7292)
);

INVx2_ASAP7_75t_L g7293 ( 
.A(n_7125),
.Y(n_7293)
);

INVx1_ASAP7_75t_L g7294 ( 
.A(n_7206),
.Y(n_7294)
);

INVx1_ASAP7_75t_L g7295 ( 
.A(n_7209),
.Y(n_7295)
);

OAI21xp5_ASAP7_75t_SL g7296 ( 
.A1(n_7134),
.A2(n_860),
.B(n_861),
.Y(n_7296)
);

NAND2xp5_ASAP7_75t_SL g7297 ( 
.A(n_7065),
.B(n_861),
.Y(n_7297)
);

AND2x2_ASAP7_75t_L g7298 ( 
.A(n_7084),
.B(n_863),
.Y(n_7298)
);

NAND2xp5_ASAP7_75t_L g7299 ( 
.A(n_7070),
.B(n_863),
.Y(n_7299)
);

OR2x2_ASAP7_75t_L g7300 ( 
.A(n_7182),
.B(n_864),
.Y(n_7300)
);

NAND2xp5_ASAP7_75t_L g7301 ( 
.A(n_7150),
.B(n_864),
.Y(n_7301)
);

INVx1_ASAP7_75t_L g7302 ( 
.A(n_7210),
.Y(n_7302)
);

NAND2xp5_ASAP7_75t_L g7303 ( 
.A(n_7113),
.B(n_866),
.Y(n_7303)
);

AND2x2_ASAP7_75t_L g7304 ( 
.A(n_7154),
.B(n_867),
.Y(n_7304)
);

INVx1_ASAP7_75t_L g7305 ( 
.A(n_7166),
.Y(n_7305)
);

NAND2xp5_ASAP7_75t_L g7306 ( 
.A(n_7094),
.B(n_867),
.Y(n_7306)
);

NAND2xp5_ASAP7_75t_L g7307 ( 
.A(n_7164),
.B(n_868),
.Y(n_7307)
);

INVx1_ASAP7_75t_L g7308 ( 
.A(n_7098),
.Y(n_7308)
);

NOR3xp33_ASAP7_75t_SL g7309 ( 
.A(n_7102),
.B(n_869),
.C(n_870),
.Y(n_7309)
);

HB1xp67_ASAP7_75t_L g7310 ( 
.A(n_7175),
.Y(n_7310)
);

AND2x2_ASAP7_75t_L g7311 ( 
.A(n_7165),
.B(n_7124),
.Y(n_7311)
);

NAND2xp5_ASAP7_75t_SL g7312 ( 
.A(n_7217),
.B(n_7187),
.Y(n_7312)
);

INVx2_ASAP7_75t_L g7313 ( 
.A(n_7245),
.Y(n_7313)
);

OAI321xp33_ASAP7_75t_L g7314 ( 
.A1(n_7220),
.A2(n_7081),
.A3(n_7169),
.B1(n_7168),
.B2(n_7078),
.C(n_7137),
.Y(n_7314)
);

INVx1_ASAP7_75t_L g7315 ( 
.A(n_7218),
.Y(n_7315)
);

NOR4xp25_ASAP7_75t_L g7316 ( 
.A(n_7219),
.B(n_7156),
.C(n_7191),
.D(n_7181),
.Y(n_7316)
);

INVx1_ASAP7_75t_L g7317 ( 
.A(n_7239),
.Y(n_7317)
);

NOR3xp33_ASAP7_75t_L g7318 ( 
.A(n_7238),
.B(n_7085),
.C(n_7080),
.Y(n_7318)
);

OAI31xp33_ASAP7_75t_SL g7319 ( 
.A1(n_7222),
.A2(n_7153),
.A3(n_7163),
.B(n_7176),
.Y(n_7319)
);

NAND2xp5_ASAP7_75t_SL g7320 ( 
.A(n_7216),
.B(n_7203),
.Y(n_7320)
);

NAND4xp75_ASAP7_75t_L g7321 ( 
.A(n_7257),
.B(n_7077),
.C(n_7075),
.D(n_7128),
.Y(n_7321)
);

OAI21xp5_ASAP7_75t_SL g7322 ( 
.A1(n_7226),
.A2(n_7162),
.B(n_7173),
.Y(n_7322)
);

AOI22xp5_ASAP7_75t_L g7323 ( 
.A1(n_7271),
.A2(n_7254),
.B1(n_7287),
.B2(n_7235),
.Y(n_7323)
);

AOI21xp33_ASAP7_75t_L g7324 ( 
.A1(n_7248),
.A2(n_7086),
.B(n_7170),
.Y(n_7324)
);

AND4x1_ASAP7_75t_L g7325 ( 
.A(n_7227),
.B(n_7106),
.C(n_7123),
.D(n_7120),
.Y(n_7325)
);

AOI321xp33_ASAP7_75t_L g7326 ( 
.A1(n_7231),
.A2(n_7114),
.A3(n_7132),
.B1(n_7160),
.B2(n_7090),
.C(n_7144),
.Y(n_7326)
);

AOI21xp5_ASAP7_75t_L g7327 ( 
.A1(n_7310),
.A2(n_7130),
.B(n_7147),
.Y(n_7327)
);

NAND4xp25_ASAP7_75t_L g7328 ( 
.A(n_7289),
.B(n_7174),
.C(n_7149),
.D(n_7177),
.Y(n_7328)
);

NOR2xp67_ASAP7_75t_L g7329 ( 
.A(n_7221),
.B(n_7152),
.Y(n_7329)
);

OAI22xp5_ASAP7_75t_L g7330 ( 
.A1(n_7237),
.A2(n_7171),
.B1(n_7180),
.B2(n_7119),
.Y(n_7330)
);

NOR3x1_ASAP7_75t_SL g7331 ( 
.A(n_7268),
.B(n_7104),
.C(n_7105),
.Y(n_7331)
);

O2A1O1Ixp33_ASAP7_75t_L g7332 ( 
.A1(n_7224),
.A2(n_7253),
.B(n_7236),
.C(n_7264),
.Y(n_7332)
);

AND2x2_ASAP7_75t_L g7333 ( 
.A(n_7311),
.B(n_7223),
.Y(n_7333)
);

INVx2_ASAP7_75t_L g7334 ( 
.A(n_7247),
.Y(n_7334)
);

NAND2xp5_ASAP7_75t_L g7335 ( 
.A(n_7234),
.B(n_7141),
.Y(n_7335)
);

OR2x2_ASAP7_75t_L g7336 ( 
.A(n_7263),
.B(n_7135),
.Y(n_7336)
);

NAND2xp5_ASAP7_75t_L g7337 ( 
.A(n_7277),
.B(n_7108),
.Y(n_7337)
);

INVx1_ASAP7_75t_L g7338 ( 
.A(n_7291),
.Y(n_7338)
);

NAND2xp5_ASAP7_75t_L g7339 ( 
.A(n_7255),
.B(n_7111),
.Y(n_7339)
);

INVx1_ASAP7_75t_L g7340 ( 
.A(n_7270),
.Y(n_7340)
);

NAND2xp5_ASAP7_75t_L g7341 ( 
.A(n_7292),
.B(n_7121),
.Y(n_7341)
);

NOR2x1_ASAP7_75t_L g7342 ( 
.A(n_7225),
.B(n_7126),
.Y(n_7342)
);

NAND3xp33_ASAP7_75t_L g7343 ( 
.A(n_7309),
.B(n_7117),
.C(n_7127),
.Y(n_7343)
);

AOI21xp5_ASAP7_75t_L g7344 ( 
.A1(n_7297),
.A2(n_7131),
.B(n_7112),
.Y(n_7344)
);

NAND2xp5_ASAP7_75t_L g7345 ( 
.A(n_7298),
.B(n_7146),
.Y(n_7345)
);

AOI22xp5_ASAP7_75t_L g7346 ( 
.A1(n_7244),
.A2(n_7143),
.B1(n_7151),
.B2(n_7122),
.Y(n_7346)
);

INVx1_ASAP7_75t_L g7347 ( 
.A(n_7267),
.Y(n_7347)
);

AOI21xp5_ASAP7_75t_L g7348 ( 
.A1(n_7233),
.A2(n_7157),
.B(n_7183),
.Y(n_7348)
);

AOI221xp5_ASAP7_75t_L g7349 ( 
.A1(n_7260),
.A2(n_7184),
.B1(n_7158),
.B2(n_7178),
.C(n_7155),
.Y(n_7349)
);

NOR2xp33_ASAP7_75t_SL g7350 ( 
.A(n_7230),
.B(n_7167),
.Y(n_7350)
);

NOR4xp25_ASAP7_75t_L g7351 ( 
.A(n_7266),
.B(n_7188),
.C(n_875),
.D(n_871),
.Y(n_7351)
);

NAND3xp33_ASAP7_75t_L g7352 ( 
.A(n_7249),
.B(n_871),
.C(n_872),
.Y(n_7352)
);

NAND2xp5_ASAP7_75t_L g7353 ( 
.A(n_7304),
.B(n_7240),
.Y(n_7353)
);

INVxp67_ASAP7_75t_SL g7354 ( 
.A(n_7250),
.Y(n_7354)
);

AOI221xp5_ASAP7_75t_L g7355 ( 
.A1(n_7269),
.A2(n_877),
.B1(n_872),
.B2(n_876),
.C(n_878),
.Y(n_7355)
);

NAND2xp5_ASAP7_75t_L g7356 ( 
.A(n_7274),
.B(n_877),
.Y(n_7356)
);

NAND2xp5_ASAP7_75t_L g7357 ( 
.A(n_7276),
.B(n_879),
.Y(n_7357)
);

INVx1_ASAP7_75t_L g7358 ( 
.A(n_7259),
.Y(n_7358)
);

AOI21xp5_ASAP7_75t_L g7359 ( 
.A1(n_7280),
.A2(n_879),
.B(n_880),
.Y(n_7359)
);

NAND2xp5_ASAP7_75t_SL g7360 ( 
.A(n_7251),
.B(n_880),
.Y(n_7360)
);

INVx1_ASAP7_75t_L g7361 ( 
.A(n_7228),
.Y(n_7361)
);

NAND3xp33_ASAP7_75t_SL g7362 ( 
.A(n_7256),
.B(n_881),
.C(n_882),
.Y(n_7362)
);

NAND2xp5_ASAP7_75t_L g7363 ( 
.A(n_7262),
.B(n_881),
.Y(n_7363)
);

AOI21xp5_ASAP7_75t_L g7364 ( 
.A1(n_7282),
.A2(n_883),
.B(n_884),
.Y(n_7364)
);

AO22x2_ASAP7_75t_SL g7365 ( 
.A1(n_7265),
.A2(n_887),
.B1(n_885),
.B2(n_886),
.Y(n_7365)
);

NAND2xp5_ASAP7_75t_SL g7366 ( 
.A(n_7293),
.B(n_886),
.Y(n_7366)
);

OAI21xp5_ASAP7_75t_L g7367 ( 
.A1(n_7243),
.A2(n_887),
.B(n_888),
.Y(n_7367)
);

NOR3xp33_ASAP7_75t_L g7368 ( 
.A(n_7278),
.B(n_889),
.C(n_890),
.Y(n_7368)
);

NAND2xp5_ASAP7_75t_L g7369 ( 
.A(n_7258),
.B(n_7273),
.Y(n_7369)
);

NAND3xp33_ASAP7_75t_SL g7370 ( 
.A(n_7296),
.B(n_890),
.C(n_892),
.Y(n_7370)
);

NOR3xp33_ASAP7_75t_SL g7371 ( 
.A(n_7272),
.B(n_892),
.C(n_893),
.Y(n_7371)
);

A2O1A1Ixp33_ASAP7_75t_L g7372 ( 
.A1(n_7288),
.A2(n_895),
.B(n_893),
.C(n_894),
.Y(n_7372)
);

NOR3xp33_ASAP7_75t_L g7373 ( 
.A(n_7279),
.B(n_894),
.C(n_897),
.Y(n_7373)
);

INVx1_ASAP7_75t_L g7374 ( 
.A(n_7232),
.Y(n_7374)
);

NAND2xp5_ASAP7_75t_L g7375 ( 
.A(n_7365),
.B(n_7305),
.Y(n_7375)
);

NOR2xp67_ASAP7_75t_L g7376 ( 
.A(n_7362),
.B(n_7275),
.Y(n_7376)
);

NAND5xp2_ASAP7_75t_L g7377 ( 
.A(n_7319),
.B(n_7290),
.C(n_7294),
.D(n_7284),
.E(n_7283),
.Y(n_7377)
);

AOI21xp5_ASAP7_75t_L g7378 ( 
.A1(n_7354),
.A2(n_7327),
.B(n_7312),
.Y(n_7378)
);

NAND3xp33_ASAP7_75t_L g7379 ( 
.A(n_7318),
.B(n_7242),
.C(n_7241),
.Y(n_7379)
);

NAND2xp5_ASAP7_75t_SL g7380 ( 
.A(n_7323),
.B(n_7229),
.Y(n_7380)
);

OAI222xp33_ASAP7_75t_L g7381 ( 
.A1(n_7342),
.A2(n_7302),
.B1(n_7295),
.B2(n_7308),
.C1(n_7252),
.C2(n_7261),
.Y(n_7381)
);

AND2x2_ASAP7_75t_L g7382 ( 
.A(n_7333),
.B(n_7300),
.Y(n_7382)
);

NOR3x1_ASAP7_75t_SL g7383 ( 
.A(n_7331),
.B(n_7246),
.C(n_7281),
.Y(n_7383)
);

BUFx2_ASAP7_75t_L g7384 ( 
.A(n_7371),
.Y(n_7384)
);

NAND4xp75_ASAP7_75t_L g7385 ( 
.A(n_7329),
.B(n_7306),
.C(n_7285),
.D(n_7303),
.Y(n_7385)
);

NAND2xp5_ASAP7_75t_L g7386 ( 
.A(n_7317),
.B(n_7301),
.Y(n_7386)
);

NOR2x1_ASAP7_75t_L g7387 ( 
.A(n_7343),
.B(n_7286),
.Y(n_7387)
);

A2O1A1O1Ixp25_ASAP7_75t_L g7388 ( 
.A1(n_7324),
.A2(n_7299),
.B(n_7307),
.C(n_900),
.D(n_898),
.Y(n_7388)
);

NOR3xp33_ASAP7_75t_L g7389 ( 
.A(n_7314),
.B(n_900),
.C(n_899),
.Y(n_7389)
);

NAND3xp33_ASAP7_75t_SL g7390 ( 
.A(n_7351),
.B(n_898),
.C(n_899),
.Y(n_7390)
);

OAI221xp5_ASAP7_75t_L g7391 ( 
.A1(n_7322),
.A2(n_903),
.B1(n_901),
.B2(n_902),
.C(n_904),
.Y(n_7391)
);

AOI221xp5_ASAP7_75t_SL g7392 ( 
.A1(n_7328),
.A2(n_904),
.B1(n_902),
.B2(n_903),
.C(n_905),
.Y(n_7392)
);

NAND4xp25_ASAP7_75t_L g7393 ( 
.A(n_7326),
.B(n_908),
.C(n_905),
.D(n_906),
.Y(n_7393)
);

NOR2xp33_ASAP7_75t_L g7394 ( 
.A(n_7350),
.B(n_7334),
.Y(n_7394)
);

OAI211xp5_ASAP7_75t_L g7395 ( 
.A1(n_7316),
.A2(n_909),
.B(n_906),
.C(n_908),
.Y(n_7395)
);

OA211x2_ASAP7_75t_L g7396 ( 
.A1(n_7370),
.A2(n_911),
.B(n_909),
.C(n_910),
.Y(n_7396)
);

OR3x1_ASAP7_75t_L g7397 ( 
.A(n_7338),
.B(n_910),
.C(n_912),
.Y(n_7397)
);

NAND4xp75_ASAP7_75t_L g7398 ( 
.A(n_7359),
.B(n_914),
.C(n_912),
.D(n_913),
.Y(n_7398)
);

NOR2xp33_ASAP7_75t_L g7399 ( 
.A(n_7352),
.B(n_913),
.Y(n_7399)
);

NAND3xp33_ASAP7_75t_L g7400 ( 
.A(n_7349),
.B(n_915),
.C(n_916),
.Y(n_7400)
);

NAND5xp2_ASAP7_75t_L g7401 ( 
.A(n_7332),
.B(n_917),
.C(n_915),
.D(n_916),
.E(n_918),
.Y(n_7401)
);

NOR3xp33_ASAP7_75t_L g7402 ( 
.A(n_7330),
.B(n_920),
.C(n_919),
.Y(n_7402)
);

NOR2xp33_ASAP7_75t_SL g7403 ( 
.A(n_7336),
.B(n_917),
.Y(n_7403)
);

AOI222xp33_ASAP7_75t_L g7404 ( 
.A1(n_7320),
.A2(n_922),
.B1(n_924),
.B2(n_919),
.C1(n_920),
.C2(n_923),
.Y(n_7404)
);

AND2x4_ASAP7_75t_L g7405 ( 
.A(n_7313),
.B(n_7315),
.Y(n_7405)
);

NOR2x1_ASAP7_75t_L g7406 ( 
.A(n_7321),
.B(n_923),
.Y(n_7406)
);

NAND2xp5_ASAP7_75t_SL g7407 ( 
.A(n_7364),
.B(n_925),
.Y(n_7407)
);

AOI211xp5_ASAP7_75t_L g7408 ( 
.A1(n_7367),
.A2(n_927),
.B(n_925),
.C(n_926),
.Y(n_7408)
);

AND2x2_ASAP7_75t_L g7409 ( 
.A(n_7340),
.B(n_927),
.Y(n_7409)
);

NOR3xp33_ASAP7_75t_L g7410 ( 
.A(n_7339),
.B(n_930),
.C(n_929),
.Y(n_7410)
);

INVx1_ASAP7_75t_L g7411 ( 
.A(n_7353),
.Y(n_7411)
);

OAI221xp5_ASAP7_75t_L g7412 ( 
.A1(n_7346),
.A2(n_930),
.B1(n_928),
.B2(n_929),
.C(n_932),
.Y(n_7412)
);

NOR2xp67_ASAP7_75t_L g7413 ( 
.A(n_7347),
.B(n_933),
.Y(n_7413)
);

NOR3xp33_ASAP7_75t_L g7414 ( 
.A(n_7337),
.B(n_934),
.C(n_933),
.Y(n_7414)
);

BUFx6f_ASAP7_75t_L g7415 ( 
.A(n_7405),
.Y(n_7415)
);

HB1xp67_ASAP7_75t_L g7416 ( 
.A(n_7413),
.Y(n_7416)
);

OAI22xp33_ASAP7_75t_L g7417 ( 
.A1(n_7403),
.A2(n_7363),
.B1(n_7357),
.B2(n_7356),
.Y(n_7417)
);

NOR2x1_ASAP7_75t_L g7418 ( 
.A(n_7397),
.B(n_7366),
.Y(n_7418)
);

INVx1_ASAP7_75t_L g7419 ( 
.A(n_7383),
.Y(n_7419)
);

NOR2xp33_ASAP7_75t_L g7420 ( 
.A(n_7393),
.B(n_7401),
.Y(n_7420)
);

OAI31xp33_ASAP7_75t_L g7421 ( 
.A1(n_7395),
.A2(n_7372),
.A3(n_7358),
.B(n_7361),
.Y(n_7421)
);

INVx1_ASAP7_75t_L g7422 ( 
.A(n_7382),
.Y(n_7422)
);

NAND4xp75_ASAP7_75t_L g7423 ( 
.A(n_7406),
.B(n_7335),
.C(n_7341),
.D(n_7345),
.Y(n_7423)
);

INVx2_ASAP7_75t_L g7424 ( 
.A(n_7405),
.Y(n_7424)
);

AOI21xp5_ASAP7_75t_L g7425 ( 
.A1(n_7378),
.A2(n_7360),
.B(n_7344),
.Y(n_7425)
);

NAND2xp5_ASAP7_75t_L g7426 ( 
.A(n_7409),
.B(n_7373),
.Y(n_7426)
);

NOR2xp67_ASAP7_75t_L g7427 ( 
.A(n_7390),
.B(n_7348),
.Y(n_7427)
);

AOI311xp33_ASAP7_75t_L g7428 ( 
.A1(n_7389),
.A2(n_7374),
.A3(n_7369),
.B(n_7368),
.C(n_7355),
.Y(n_7428)
);

OAI21xp5_ASAP7_75t_L g7429 ( 
.A1(n_7394),
.A2(n_7325),
.B(n_932),
.Y(n_7429)
);

NAND2xp5_ASAP7_75t_L g7430 ( 
.A(n_7376),
.B(n_934),
.Y(n_7430)
);

NOR2x1_ASAP7_75t_L g7431 ( 
.A(n_7398),
.B(n_935),
.Y(n_7431)
);

INVx1_ASAP7_75t_L g7432 ( 
.A(n_7375),
.Y(n_7432)
);

AOI22xp5_ASAP7_75t_L g7433 ( 
.A1(n_7384),
.A2(n_937),
.B1(n_935),
.B2(n_936),
.Y(n_7433)
);

OAI211xp5_ASAP7_75t_L g7434 ( 
.A1(n_7388),
.A2(n_939),
.B(n_937),
.C(n_938),
.Y(n_7434)
);

OAI22xp33_ASAP7_75t_L g7435 ( 
.A1(n_7391),
.A2(n_942),
.B1(n_938),
.B2(n_941),
.Y(n_7435)
);

OAI21xp5_ASAP7_75t_L g7436 ( 
.A1(n_7400),
.A2(n_942),
.B(n_943),
.Y(n_7436)
);

INVx1_ASAP7_75t_L g7437 ( 
.A(n_7396),
.Y(n_7437)
);

INVx1_ASAP7_75t_L g7438 ( 
.A(n_7387),
.Y(n_7438)
);

INVx1_ASAP7_75t_L g7439 ( 
.A(n_7415),
.Y(n_7439)
);

NOR3xp33_ASAP7_75t_SL g7440 ( 
.A(n_7434),
.B(n_7377),
.C(n_7381),
.Y(n_7440)
);

NOR2xp33_ASAP7_75t_L g7441 ( 
.A(n_7415),
.B(n_7407),
.Y(n_7441)
);

NOR3xp33_ASAP7_75t_L g7442 ( 
.A(n_7419),
.B(n_7379),
.C(n_7380),
.Y(n_7442)
);

NOR2x1p5_ASAP7_75t_L g7443 ( 
.A(n_7423),
.B(n_7385),
.Y(n_7443)
);

INVx2_ASAP7_75t_L g7444 ( 
.A(n_7424),
.Y(n_7444)
);

AND3x4_ASAP7_75t_L g7445 ( 
.A(n_7418),
.B(n_7402),
.C(n_7414),
.Y(n_7445)
);

OR2x2_ASAP7_75t_L g7446 ( 
.A(n_7430),
.B(n_7386),
.Y(n_7446)
);

AOI21xp5_ASAP7_75t_L g7447 ( 
.A1(n_7425),
.A2(n_7399),
.B(n_7411),
.Y(n_7447)
);

NOR2xp33_ASAP7_75t_L g7448 ( 
.A(n_7422),
.B(n_7412),
.Y(n_7448)
);

NAND4xp75_ASAP7_75t_L g7449 ( 
.A(n_7427),
.B(n_7392),
.C(n_7404),
.D(n_7410),
.Y(n_7449)
);

AND3x4_ASAP7_75t_L g7450 ( 
.A(n_7431),
.B(n_7408),
.C(n_943),
.Y(n_7450)
);

AND2x4_ASAP7_75t_L g7451 ( 
.A(n_7438),
.B(n_7437),
.Y(n_7451)
);

AND2x4_ASAP7_75t_L g7452 ( 
.A(n_7432),
.B(n_944),
.Y(n_7452)
);

AND2x2_ASAP7_75t_L g7453 ( 
.A(n_7420),
.B(n_945),
.Y(n_7453)
);

INVx2_ASAP7_75t_L g7454 ( 
.A(n_7416),
.Y(n_7454)
);

NOR2xp33_ASAP7_75t_L g7455 ( 
.A(n_7435),
.B(n_945),
.Y(n_7455)
);

OR2x2_ASAP7_75t_L g7456 ( 
.A(n_7426),
.B(n_946),
.Y(n_7456)
);

NOR3x1_ASAP7_75t_L g7457 ( 
.A(n_7436),
.B(n_947),
.C(n_948),
.Y(n_7457)
);

AOI221xp5_ASAP7_75t_L g7458 ( 
.A1(n_7442),
.A2(n_7417),
.B1(n_7429),
.B2(n_7421),
.C(n_7433),
.Y(n_7458)
);

HB1xp67_ASAP7_75t_L g7459 ( 
.A(n_7452),
.Y(n_7459)
);

INVx1_ASAP7_75t_L g7460 ( 
.A(n_7453),
.Y(n_7460)
);

INVx1_ASAP7_75t_L g7461 ( 
.A(n_7456),
.Y(n_7461)
);

BUFx2_ASAP7_75t_L g7462 ( 
.A(n_7444),
.Y(n_7462)
);

OR2x2_ASAP7_75t_L g7463 ( 
.A(n_7439),
.B(n_7428),
.Y(n_7463)
);

BUFx2_ASAP7_75t_L g7464 ( 
.A(n_7451),
.Y(n_7464)
);

HB1xp67_ASAP7_75t_L g7465 ( 
.A(n_7450),
.Y(n_7465)
);

NAND4xp75_ASAP7_75t_L g7466 ( 
.A(n_7440),
.B(n_951),
.C(n_949),
.D(n_950),
.Y(n_7466)
);

NAND3xp33_ASAP7_75t_SL g7467 ( 
.A(n_7445),
.B(n_950),
.C(n_951),
.Y(n_7467)
);

NOR2xp33_ASAP7_75t_L g7468 ( 
.A(n_7454),
.B(n_952),
.Y(n_7468)
);

NOR3x1_ASAP7_75t_L g7469 ( 
.A(n_7449),
.B(n_952),
.C(n_953),
.Y(n_7469)
);

NAND3xp33_ASAP7_75t_L g7470 ( 
.A(n_7455),
.B(n_953),
.C(n_955),
.Y(n_7470)
);

NAND2xp5_ASAP7_75t_L g7471 ( 
.A(n_7441),
.B(n_957),
.Y(n_7471)
);

XOR2xp5_ASAP7_75t_L g7472 ( 
.A(n_7466),
.B(n_7446),
.Y(n_7472)
);

AOI22xp5_ASAP7_75t_L g7473 ( 
.A1(n_7464),
.A2(n_7448),
.B1(n_7462),
.B2(n_7443),
.Y(n_7473)
);

AO22x2_ASAP7_75t_L g7474 ( 
.A1(n_7467),
.A2(n_7447),
.B1(n_7457),
.B2(n_958),
.Y(n_7474)
);

INVx1_ASAP7_75t_L g7475 ( 
.A(n_7459),
.Y(n_7475)
);

NAND2xp33_ASAP7_75t_L g7476 ( 
.A(n_7465),
.B(n_956),
.Y(n_7476)
);

NAND5xp2_ASAP7_75t_L g7477 ( 
.A(n_7473),
.B(n_7458),
.C(n_7460),
.D(n_7461),
.E(n_7471),
.Y(n_7477)
);

INVx1_ASAP7_75t_SL g7478 ( 
.A(n_7476),
.Y(n_7478)
);

OAI222xp33_ASAP7_75t_L g7479 ( 
.A1(n_7475),
.A2(n_7463),
.B1(n_7469),
.B2(n_7468),
.C1(n_7470),
.C2(n_958),
.Y(n_7479)
);

NOR2xp33_ASAP7_75t_L g7480 ( 
.A(n_7472),
.B(n_956),
.Y(n_7480)
);

AOI21xp5_ASAP7_75t_L g7481 ( 
.A1(n_7480),
.A2(n_7474),
.B(n_957),
.Y(n_7481)
);

AOI322xp5_ASAP7_75t_L g7482 ( 
.A1(n_7478),
.A2(n_964),
.A3(n_963),
.B1(n_961),
.B2(n_959),
.C1(n_960),
.C2(n_962),
.Y(n_7482)
);

INVx2_ASAP7_75t_L g7483 ( 
.A(n_7482),
.Y(n_7483)
);

BUFx12f_ASAP7_75t_L g7484 ( 
.A(n_7481),
.Y(n_7484)
);

AOI21xp5_ASAP7_75t_L g7485 ( 
.A1(n_7483),
.A2(n_7477),
.B(n_7479),
.Y(n_7485)
);

OAI21xp5_ASAP7_75t_L g7486 ( 
.A1(n_7484),
.A2(n_959),
.B(n_960),
.Y(n_7486)
);

INVx1_ASAP7_75t_L g7487 ( 
.A(n_7486),
.Y(n_7487)
);

AND2x4_ASAP7_75t_L g7488 ( 
.A(n_7485),
.B(n_962),
.Y(n_7488)
);

AOI221xp5_ASAP7_75t_SL g7489 ( 
.A1(n_7487),
.A2(n_966),
.B1(n_963),
.B2(n_965),
.C(n_967),
.Y(n_7489)
);

AOI22xp5_ASAP7_75t_L g7490 ( 
.A1(n_7489),
.A2(n_7488),
.B1(n_968),
.B2(n_966),
.Y(n_7490)
);

AOI221xp5_ASAP7_75t_L g7491 ( 
.A1(n_7489),
.A2(n_969),
.B1(n_967),
.B2(n_968),
.C(n_970),
.Y(n_7491)
);

AOI21x1_ASAP7_75t_L g7492 ( 
.A1(n_7491),
.A2(n_971),
.B(n_970),
.Y(n_7492)
);

OAI21xp33_ASAP7_75t_SL g7493 ( 
.A1(n_7490),
.A2(n_969),
.B(n_971),
.Y(n_7493)
);

INVx1_ASAP7_75t_L g7494 ( 
.A(n_7492),
.Y(n_7494)
);

INVx4_ASAP7_75t_L g7495 ( 
.A(n_7493),
.Y(n_7495)
);

AOI221xp5_ASAP7_75t_L g7496 ( 
.A1(n_7494),
.A2(n_974),
.B1(n_972),
.B2(n_973),
.C(n_975),
.Y(n_7496)
);

OR2x6_ASAP7_75t_L g7497 ( 
.A(n_7495),
.B(n_973),
.Y(n_7497)
);

AOI21xp5_ASAP7_75t_L g7498 ( 
.A1(n_7497),
.A2(n_974),
.B(n_975),
.Y(n_7498)
);

AOI211xp5_ASAP7_75t_L g7499 ( 
.A1(n_7498),
.A2(n_7496),
.B(n_978),
.C(n_977),
.Y(n_7499)
);


endmodule