module real_aes_6480_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_241;
wire n_168;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_0), .B(n_87), .C(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g124 ( .A(n_0), .Y(n_124) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_1), .A2(n_145), .B(n_148), .C(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g211 ( .A(n_2), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_3), .A2(n_140), .B(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_4), .B(n_221), .Y(n_535) );
AOI21xp33_ASAP7_75t_L g222 ( .A1(n_5), .A2(n_140), .B(n_223), .Y(n_222) );
AND2x6_ASAP7_75t_L g145 ( .A(n_6), .B(n_146), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_7), .A2(n_191), .B(n_192), .Y(n_190) );
INVx1_ASAP7_75t_L g108 ( .A(n_8), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_8), .B(n_41), .Y(n_125) );
OAI22xp5_ASAP7_75t_L g128 ( .A1(n_9), .A2(n_31), .B1(n_129), .B2(n_130), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_9), .Y(n_130) );
INVx1_ASAP7_75t_L g470 ( .A(n_10), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_11), .B(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g228 ( .A(n_12), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_13), .B(n_181), .Y(n_491) );
INVx1_ASAP7_75t_L g166 ( .A(n_14), .Y(n_166) );
INVx1_ASAP7_75t_L g199 ( .A(n_15), .Y(n_199) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_16), .A2(n_154), .B(n_200), .C(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_17), .B(n_221), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_18), .B(n_156), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g139 ( .A(n_19), .B(n_140), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_20), .B(n_571), .Y(n_570) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_21), .A2(n_180), .B(n_214), .C(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_22), .B(n_221), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_23), .B(n_181), .Y(n_524) );
A2O1A1Ixp33_ASAP7_75t_L g195 ( .A1(n_24), .A2(n_196), .B(n_198), .C(n_200), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_25), .B(n_181), .Y(n_510) );
CKINVDCx16_ASAP7_75t_R g520 ( .A(n_26), .Y(n_520) );
INVx1_ASAP7_75t_L g509 ( .A(n_27), .Y(n_509) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_28), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_29), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_30), .B(n_181), .Y(n_212) );
INVx1_ASAP7_75t_L g129 ( .A(n_31), .Y(n_129) );
INVx1_ASAP7_75t_L g567 ( .A(n_32), .Y(n_567) );
INVx1_ASAP7_75t_L g238 ( .A(n_33), .Y(n_238) );
INVx2_ASAP7_75t_L g143 ( .A(n_34), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_35), .Y(n_493) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_36), .A2(n_180), .B(n_229), .C(n_533), .Y(n_532) );
INVxp67_ASAP7_75t_L g568 ( .A(n_37), .Y(n_568) );
A2O1A1Ixp33_ASAP7_75t_L g147 ( .A1(n_38), .A2(n_145), .B(n_148), .C(n_151), .Y(n_147) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_39), .A2(n_148), .B(n_508), .C(n_513), .Y(n_507) );
CKINVDCx14_ASAP7_75t_R g531 ( .A(n_40), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_41), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g236 ( .A(n_42), .Y(n_236) );
A2O1A1Ixp33_ASAP7_75t_L g468 ( .A1(n_43), .A2(n_158), .B(n_226), .C(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_44), .B(n_181), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_45), .A2(n_102), .B1(n_113), .B2(n_743), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_46), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g564 ( .A(n_47), .Y(n_564) );
INVx1_ASAP7_75t_L g498 ( .A(n_48), .Y(n_498) );
CKINVDCx16_ASAP7_75t_R g239 ( .A(n_49), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_50), .B(n_140), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_51), .Y(n_126) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_52), .A2(n_148), .B1(n_214), .B2(n_235), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_53), .Y(n_168) );
CKINVDCx16_ASAP7_75t_R g207 ( .A(n_54), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_55), .A2(n_226), .B(n_227), .C(n_229), .Y(n_225) );
CKINVDCx14_ASAP7_75t_R g467 ( .A(n_56), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g276 ( .A(n_57), .Y(n_276) );
INVx1_ASAP7_75t_L g224 ( .A(n_58), .Y(n_224) );
INVx1_ASAP7_75t_L g146 ( .A(n_59), .Y(n_146) );
INVx1_ASAP7_75t_L g165 ( .A(n_60), .Y(n_165) );
INVx1_ASAP7_75t_SL g534 ( .A(n_61), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_62), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_63), .B(n_221), .Y(n_502) );
INVx1_ASAP7_75t_L g523 ( .A(n_64), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_SL g246 ( .A1(n_65), .A2(n_156), .B(n_229), .C(n_247), .Y(n_246) );
INVxp67_ASAP7_75t_L g248 ( .A(n_66), .Y(n_248) );
INVx1_ASAP7_75t_L g112 ( .A(n_67), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_68), .A2(n_140), .B(n_466), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_69), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g241 ( .A(n_70), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_71), .A2(n_140), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g269 ( .A(n_72), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_73), .A2(n_191), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g477 ( .A(n_74), .Y(n_477) );
CKINVDCx16_ASAP7_75t_R g506 ( .A(n_75), .Y(n_506) );
OAI22xp5_ASAP7_75t_SL g739 ( .A1(n_76), .A2(n_77), .B1(n_740), .B2(n_741), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_76), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_77), .Y(n_740) );
A2O1A1Ixp33_ASAP7_75t_L g270 ( .A1(n_78), .A2(n_145), .B(n_148), .C(n_271), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_79), .A2(n_140), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g480 ( .A(n_80), .Y(n_480) );
AOI222xp33_ASAP7_75t_SL g127 ( .A1(n_81), .A2(n_128), .B1(n_131), .B2(n_728), .C1(n_729), .C2(n_733), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_82), .B(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g163 ( .A(n_83), .Y(n_163) );
INVx1_ASAP7_75t_L g489 ( .A(n_84), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_85), .B(n_156), .Y(n_155) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_86), .A2(n_145), .B(n_148), .C(n_210), .Y(n_209) );
OR2x2_ASAP7_75t_L g121 ( .A(n_87), .B(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g457 ( .A(n_87), .Y(n_457) );
OR2x2_ASAP7_75t_L g727 ( .A(n_87), .B(n_123), .Y(n_727) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_88), .A2(n_148), .B(n_522), .C(n_525), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_89), .B(n_174), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g217 ( .A(n_90), .Y(n_217) );
A2O1A1Ixp33_ASAP7_75t_L g176 ( .A1(n_91), .A2(n_145), .B(n_148), .C(n_177), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_92), .Y(n_186) );
INVx1_ASAP7_75t_L g245 ( .A(n_93), .Y(n_245) );
CKINVDCx16_ASAP7_75t_R g193 ( .A(n_94), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_95), .B(n_153), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_96), .B(n_170), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_97), .B(n_170), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_98), .B(n_112), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_99), .A2(n_140), .B(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g501 ( .A(n_100), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
CKINVDCx6p67_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_105), .Y(n_744) );
CKINVDCx9p33_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g106 ( .A(n_107), .B(n_109), .Y(n_106) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
AOI22x1_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_127), .B1(n_736), .B2(n_737), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_119), .Y(n_114) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_SL g736 ( .A(n_116), .Y(n_736) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g737 ( .A1(n_119), .A2(n_738), .B(n_742), .Y(n_737) );
NOR2xp33_ASAP7_75t_SL g119 ( .A(n_120), .B(n_126), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_121), .Y(n_742) );
NOR2x2_ASAP7_75t_L g735 ( .A(n_122), .B(n_457), .Y(n_735) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OR2x2_ASAP7_75t_L g456 ( .A(n_123), .B(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
INVx1_ASAP7_75t_L g728 ( .A(n_128), .Y(n_728) );
OAI22xp5_ASAP7_75t_SL g131 ( .A1(n_132), .A2(n_456), .B1(n_458), .B2(n_727), .Y(n_131) );
INVx2_ASAP7_75t_L g730 ( .A(n_132), .Y(n_730) );
AND2x2_ASAP7_75t_SL g132 ( .A(n_133), .B(n_425), .Y(n_132) );
NOR3xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_318), .C(n_391), .Y(n_133) );
OAI211xp5_ASAP7_75t_SL g134 ( .A1(n_135), .A2(n_203), .B(n_250), .C(n_302), .Y(n_134) );
INVxp67_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_171), .Y(n_136) );
AND2x2_ASAP7_75t_L g266 ( .A(n_137), .B(n_267), .Y(n_266) );
INVx3_ASAP7_75t_L g285 ( .A(n_137), .Y(n_285) );
INVx2_ASAP7_75t_L g300 ( .A(n_137), .Y(n_300) );
INVx1_ASAP7_75t_L g330 ( .A(n_137), .Y(n_330) );
AND2x2_ASAP7_75t_L g380 ( .A(n_137), .B(n_301), .Y(n_380) );
AOI32xp33_ASAP7_75t_L g407 ( .A1(n_137), .A2(n_335), .A3(n_408), .B1(n_410), .B2(n_411), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_137), .B(n_256), .Y(n_413) );
AND2x2_ASAP7_75t_L g440 ( .A(n_137), .B(n_283), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_137), .B(n_449), .Y(n_448) );
OR2x6_ASAP7_75t_L g137 ( .A(n_138), .B(n_167), .Y(n_137) );
AOI21xp5_ASAP7_75t_SL g138 ( .A1(n_139), .A2(n_147), .B(n_160), .Y(n_138) );
BUFx2_ASAP7_75t_L g191 ( .A(n_140), .Y(n_191) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_145), .Y(n_140) );
NAND2x1p5_ASAP7_75t_L g208 ( .A(n_141), .B(n_145), .Y(n_208) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
INVx1_ASAP7_75t_L g512 ( .A(n_142), .Y(n_512) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g149 ( .A(n_143), .Y(n_149) );
INVx1_ASAP7_75t_L g215 ( .A(n_143), .Y(n_215) );
INVx1_ASAP7_75t_L g150 ( .A(n_144), .Y(n_150) );
INVx3_ASAP7_75t_L g154 ( .A(n_144), .Y(n_154) );
INVx1_ASAP7_75t_L g156 ( .A(n_144), .Y(n_156) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_144), .Y(n_181) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_144), .Y(n_197) );
INVx4_ASAP7_75t_SL g201 ( .A(n_145), .Y(n_201) );
BUFx3_ASAP7_75t_L g513 ( .A(n_145), .Y(n_513) );
INVx5_ASAP7_75t_L g194 ( .A(n_148), .Y(n_194) );
AND2x6_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
BUFx3_ASAP7_75t_L g159 ( .A(n_149), .Y(n_159) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_149), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_155), .B(n_157), .Y(n_151) );
O2A1O1Ixp33_ASAP7_75t_L g210 ( .A1(n_153), .A2(n_211), .B(n_212), .C(n_213), .Y(n_210) );
O2A1O1Ixp33_ASAP7_75t_L g508 ( .A1(n_153), .A2(n_509), .B(n_510), .C(n_511), .Y(n_508) );
OAI22xp33_ASAP7_75t_L g566 ( .A1(n_153), .A2(n_196), .B1(n_567), .B2(n_568), .Y(n_566) );
INVx5_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_154), .B(n_228), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_154), .B(n_248), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_154), .B(n_470), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_157), .A2(n_272), .B(n_273), .Y(n_271) );
O2A1O1Ixp5_ASAP7_75t_L g488 ( .A1(n_157), .A2(n_489), .B(n_490), .C(n_491), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_L g522 ( .A1(n_157), .A2(n_490), .B(n_523), .C(n_524), .Y(n_522) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g200 ( .A(n_159), .Y(n_200) );
INVx1_ASAP7_75t_L g274 ( .A(n_160), .Y(n_274) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AO21x2_ASAP7_75t_L g205 ( .A1(n_161), .A2(n_206), .B(n_216), .Y(n_205) );
AO21x2_ASAP7_75t_L g232 ( .A1(n_161), .A2(n_233), .B(n_240), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_161), .B(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_162), .Y(n_170) );
AND2x2_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
AND2x2_ASAP7_75t_SL g174 ( .A(n_163), .B(n_164), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_165), .B(n_166), .Y(n_164) );
NOR2xp33_ASAP7_75t_SL g167 ( .A(n_168), .B(n_169), .Y(n_167) );
INVx3_ASAP7_75t_L g221 ( .A(n_169), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_169), .B(n_493), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_169), .B(n_515), .Y(n_514) );
AO21x2_ASAP7_75t_L g518 ( .A1(n_169), .A2(n_519), .B(n_526), .Y(n_518) );
INVx4_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
OA21x2_ASAP7_75t_L g242 ( .A1(n_170), .A2(n_243), .B(n_249), .Y(n_242) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_170), .Y(n_474) );
AND2x2_ASAP7_75t_L g329 ( .A(n_171), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g351 ( .A(n_171), .Y(n_351) );
AND2x2_ASAP7_75t_L g436 ( .A(n_171), .B(n_266), .Y(n_436) );
AND2x2_ASAP7_75t_L g439 ( .A(n_171), .B(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_188), .Y(n_171) );
INVx2_ASAP7_75t_L g258 ( .A(n_172), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_172), .B(n_283), .Y(n_289) );
AND2x2_ASAP7_75t_L g299 ( .A(n_172), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g335 ( .A(n_172), .Y(n_335) );
AO21x2_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_175), .B(n_185), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_173), .B(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g571 ( .A(n_173), .Y(n_571) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g187 ( .A(n_174), .Y(n_187) );
OA21x2_ASAP7_75t_L g189 ( .A1(n_174), .A2(n_190), .B(n_202), .Y(n_189) );
OA21x2_ASAP7_75t_L g464 ( .A1(n_174), .A2(n_465), .B(n_471), .Y(n_464) );
O2A1O1Ixp33_ASAP7_75t_L g505 ( .A1(n_174), .A2(n_208), .B(n_506), .C(n_507), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_176), .B(n_184), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_182), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_180), .B(n_534), .Y(n_533) );
INVx4_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g226 ( .A(n_181), .Y(n_226) );
HB1xp67_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx3_ASAP7_75t_L g229 ( .A(n_183), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_186), .B(n_187), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_187), .B(n_217), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_187), .B(n_276), .Y(n_275) );
AO21x2_ASAP7_75t_L g484 ( .A1(n_187), .A2(n_485), .B(n_492), .Y(n_484) );
AND2x2_ASAP7_75t_L g277 ( .A(n_188), .B(n_258), .Y(n_277) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g259 ( .A(n_189), .Y(n_259) );
AND2x2_ASAP7_75t_L g301 ( .A(n_189), .B(n_283), .Y(n_301) );
AND2x2_ASAP7_75t_L g370 ( .A(n_189), .B(n_267), .Y(n_370) );
O2A1O1Ixp33_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_195), .C(n_201), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g223 ( .A1(n_194), .A2(n_201), .B(n_224), .C(n_225), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_L g244 ( .A1(n_194), .A2(n_201), .B(n_245), .C(n_246), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_SL g466 ( .A1(n_194), .A2(n_201), .B(n_467), .C(n_468), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_SL g476 ( .A1(n_194), .A2(n_201), .B(n_477), .C(n_478), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_SL g497 ( .A1(n_194), .A2(n_201), .B(n_498), .C(n_499), .Y(n_497) );
O2A1O1Ixp33_ASAP7_75t_L g530 ( .A1(n_194), .A2(n_201), .B(n_531), .C(n_532), .Y(n_530) );
O2A1O1Ixp33_ASAP7_75t_SL g563 ( .A1(n_194), .A2(n_201), .B(n_564), .C(n_565), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_196), .B(n_199), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_196), .B(n_480), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_196), .B(n_501), .Y(n_500) );
INVx4_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
OAI22xp5_ASAP7_75t_SL g235 ( .A1(n_197), .A2(n_236), .B1(n_237), .B2(n_238), .Y(n_235) );
INVx2_ASAP7_75t_L g237 ( .A(n_197), .Y(n_237) );
OAI22xp33_ASAP7_75t_L g233 ( .A1(n_201), .A2(n_208), .B1(n_234), .B2(n_239), .Y(n_233) );
INVx1_ASAP7_75t_L g525 ( .A(n_201), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_204), .B(n_218), .Y(n_203) );
OR2x2_ASAP7_75t_L g264 ( .A(n_204), .B(n_232), .Y(n_264) );
INVx1_ASAP7_75t_L g343 ( .A(n_204), .Y(n_343) );
AND2x2_ASAP7_75t_L g357 ( .A(n_204), .B(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_204), .B(n_231), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_204), .B(n_355), .Y(n_409) );
AND2x2_ASAP7_75t_L g417 ( .A(n_204), .B(n_418), .Y(n_417) );
INVx3_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx3_ASAP7_75t_L g254 ( .A(n_205), .Y(n_254) );
AND2x2_ASAP7_75t_L g324 ( .A(n_205), .B(n_232), .Y(n_324) );
OAI21xp5_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_208), .B(n_209), .Y(n_206) );
OAI21xp5_ASAP7_75t_L g268 ( .A1(n_208), .A2(n_269), .B(n_270), .Y(n_268) );
OAI21xp5_ASAP7_75t_L g485 ( .A1(n_208), .A2(n_486), .B(n_487), .Y(n_485) );
OAI21xp5_ASAP7_75t_L g519 ( .A1(n_208), .A2(n_520), .B(n_521), .Y(n_519) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx3_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_218), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g451 ( .A(n_218), .Y(n_451) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_231), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_219), .B(n_295), .Y(n_317) );
OR2x2_ASAP7_75t_L g346 ( .A(n_219), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g378 ( .A(n_219), .B(n_358), .Y(n_378) );
INVx1_ASAP7_75t_SL g398 ( .A(n_219), .Y(n_398) );
AND2x2_ASAP7_75t_L g402 ( .A(n_219), .B(n_263), .Y(n_402) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_SL g255 ( .A(n_220), .B(n_231), .Y(n_255) );
AND2x2_ASAP7_75t_L g262 ( .A(n_220), .B(n_242), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_220), .B(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g305 ( .A(n_220), .B(n_287), .Y(n_305) );
INVx1_ASAP7_75t_SL g312 ( .A(n_220), .Y(n_312) );
BUFx2_ASAP7_75t_L g323 ( .A(n_220), .Y(n_323) );
AND2x2_ASAP7_75t_L g339 ( .A(n_220), .B(n_254), .Y(n_339) );
AND2x2_ASAP7_75t_L g354 ( .A(n_220), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g418 ( .A(n_220), .B(n_232), .Y(n_418) );
OA21x2_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_230), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_231), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g342 ( .A(n_231), .B(n_343), .Y(n_342) );
AOI221xp5_ASAP7_75t_L g359 ( .A1(n_231), .A2(n_360), .B1(n_363), .B2(n_366), .C(n_371), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_231), .B(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_242), .Y(n_231) );
INVx3_ASAP7_75t_L g287 ( .A(n_232), .Y(n_287) );
INVx2_ASAP7_75t_L g490 ( .A(n_237), .Y(n_490) );
BUFx2_ASAP7_75t_L g297 ( .A(n_242), .Y(n_297) );
AND2x2_ASAP7_75t_L g311 ( .A(n_242), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g328 ( .A(n_242), .Y(n_328) );
OR2x2_ASAP7_75t_L g347 ( .A(n_242), .B(n_287), .Y(n_347) );
INVx3_ASAP7_75t_L g355 ( .A(n_242), .Y(n_355) );
AND2x2_ASAP7_75t_L g358 ( .A(n_242), .B(n_287), .Y(n_358) );
AOI221xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_256), .B1(n_260), .B2(n_265), .C(n_278), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_255), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_253), .B(n_327), .Y(n_452) );
OR2x2_ASAP7_75t_L g455 ( .A(n_253), .B(n_286), .Y(n_455) );
INVx1_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
OAI221xp5_ASAP7_75t_SL g278 ( .A1(n_254), .A2(n_279), .B1(n_286), .B2(n_288), .C(n_291), .Y(n_278) );
AND2x2_ASAP7_75t_L g295 ( .A(n_254), .B(n_287), .Y(n_295) );
AND2x2_ASAP7_75t_L g303 ( .A(n_254), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_254), .B(n_311), .Y(n_310) );
NAND2x1_ASAP7_75t_L g353 ( .A(n_254), .B(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g405 ( .A(n_254), .B(n_347), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_256), .A2(n_365), .B1(n_394), .B2(n_396), .Y(n_393) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AOI322xp5_ASAP7_75t_L g302 ( .A1(n_257), .A2(n_266), .A3(n_303), .B1(n_306), .B2(n_309), .C1(n_313), .C2(n_316), .Y(n_302) );
OR2x2_ASAP7_75t_L g314 ( .A(n_257), .B(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_258), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g293 ( .A(n_258), .B(n_267), .Y(n_293) );
INVx1_ASAP7_75t_L g308 ( .A(n_258), .Y(n_308) );
AND2x2_ASAP7_75t_L g374 ( .A(n_258), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g284 ( .A(n_259), .B(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g375 ( .A(n_259), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_259), .B(n_283), .Y(n_449) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_263), .B(n_398), .Y(n_397) );
INVx3_ASAP7_75t_SL g263 ( .A(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g349 ( .A(n_264), .B(n_296), .Y(n_349) );
OR2x2_ASAP7_75t_L g446 ( .A(n_264), .B(n_297), .Y(n_446) );
INVx1_ASAP7_75t_L g427 ( .A(n_265), .Y(n_427) );
AND2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_277), .Y(n_265) );
INVx4_ASAP7_75t_L g315 ( .A(n_266), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_266), .B(n_334), .Y(n_340) );
INVx2_ASAP7_75t_L g283 ( .A(n_267), .Y(n_283) );
AO21x2_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_274), .B(n_275), .Y(n_267) );
AO21x2_ASAP7_75t_L g560 ( .A1(n_274), .A2(n_561), .B(n_569), .Y(n_560) );
INVx1_ASAP7_75t_L g578 ( .A(n_274), .Y(n_578) );
INVx1_ASAP7_75t_L g365 ( .A(n_277), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_277), .B(n_337), .Y(n_406) );
AOI21xp33_ASAP7_75t_L g352 ( .A1(n_279), .A2(n_353), .B(n_356), .Y(n_352) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_284), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g337 ( .A(n_283), .Y(n_337) );
INVx1_ASAP7_75t_L g364 ( .A(n_283), .Y(n_364) );
INVx1_ASAP7_75t_L g290 ( .A(n_284), .Y(n_290) );
AND2x2_ASAP7_75t_L g292 ( .A(n_284), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g388 ( .A(n_285), .B(n_374), .Y(n_388) );
AND2x2_ASAP7_75t_L g410 ( .A(n_285), .B(n_370), .Y(n_410) );
BUFx2_ASAP7_75t_L g362 ( .A(n_287), .Y(n_362) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
AOI32xp33_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_294), .A3(n_295), .B1(n_296), .B2(n_298), .Y(n_291) );
INVx1_ASAP7_75t_L g372 ( .A(n_292), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_292), .A2(n_420), .B1(n_421), .B2(n_423), .Y(n_419) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_295), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_295), .B(n_354), .Y(n_395) );
AND2x2_ASAP7_75t_L g442 ( .A(n_295), .B(n_327), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_296), .B(n_343), .Y(n_390) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g443 ( .A(n_298), .Y(n_443) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
INVx1_ASAP7_75t_L g368 ( .A(n_299), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_301), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g415 ( .A(n_301), .B(n_335), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_301), .B(n_330), .Y(n_422) );
INVx1_ASAP7_75t_SL g404 ( .A(n_303), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_304), .B(n_355), .Y(n_382) );
NOR4xp25_ASAP7_75t_L g428 ( .A(n_304), .B(n_327), .C(n_429), .D(n_432), .Y(n_428) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_305), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVxp67_ASAP7_75t_L g385 ( .A(n_308), .Y(n_385) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OAI21xp33_ASAP7_75t_L g435 ( .A1(n_311), .A2(n_402), .B(n_436), .Y(n_435) );
AND2x4_ASAP7_75t_L g327 ( .A(n_312), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g376 ( .A(n_315), .Y(n_376) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND4xp25_ASAP7_75t_SL g318 ( .A(n_319), .B(n_344), .C(n_359), .D(n_379), .Y(n_318) );
O2A1O1Ixp33_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_325), .B(n_329), .C(n_331), .Y(n_319) );
INVx1_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_322), .B(n_324), .Y(n_321) );
INVx1_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g411 ( .A(n_324), .B(n_354), .Y(n_411) );
AND2x2_ASAP7_75t_L g420 ( .A(n_324), .B(n_398), .Y(n_420) );
INVx3_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_327), .B(n_362), .Y(n_424) );
AND2x2_ASAP7_75t_L g336 ( .A(n_330), .B(n_337), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_338), .B1(n_340), .B2(n_341), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_336), .Y(n_333) );
AND2x2_ASAP7_75t_L g434 ( .A(n_334), .B(n_380), .Y(n_434) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_336), .B(n_385), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_337), .B(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
O2A1O1Ixp33_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_348), .B(n_350), .C(n_352), .Y(n_344) );
AOI221xp5_ASAP7_75t_L g379 ( .A1(n_345), .A2(n_380), .B1(n_381), .B2(n_383), .C(n_386), .Y(n_379) );
INVx1_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OAI221xp5_ASAP7_75t_L g437 ( .A1(n_353), .A2(n_438), .B1(n_441), .B2(n_443), .C(n_444), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_354), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_362), .B(n_431), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
INVx1_ASAP7_75t_L g392 ( .A(n_364), .Y(n_392) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_367), .A2(n_387), .B1(n_389), .B2(n_390), .Y(n_386) );
OR2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AOI21xp33_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_373), .B(n_377), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_376), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_376), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OAI221xp5_ASAP7_75t_L g450 ( .A1(n_387), .A2(n_413), .B1(n_451), .B2(n_452), .C(n_453), .Y(n_450) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g432 ( .A(n_389), .Y(n_432) );
OAI211xp5_ASAP7_75t_SL g391 ( .A1(n_392), .A2(n_393), .B(n_399), .C(n_419), .Y(n_391) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AOI211xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_402), .B(n_403), .C(n_412), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
A2O1A1Ixp33_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_405), .B(n_406), .C(n_407), .Y(n_403) );
INVx1_ASAP7_75t_L g431 ( .A(n_409), .Y(n_431) );
OAI21xp5_ASAP7_75t_SL g453 ( .A1(n_410), .A2(n_436), .B(n_454), .Y(n_453) );
AOI21xp33_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_414), .B(n_416), .Y(n_412) );
INVx1_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
INVxp67_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OAI21xp5_ASAP7_75t_SL g445 ( .A1(n_422), .A2(n_446), .B(n_447), .Y(n_445) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
NOR3xp33_ASAP7_75t_L g425 ( .A(n_426), .B(n_437), .C(n_450), .Y(n_425) );
OAI211xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_428), .B(n_433), .C(n_435), .Y(n_426) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
CKINVDCx14_ASAP7_75t_R g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g732 ( .A(n_456), .Y(n_732) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OAI22xp5_ASAP7_75t_SL g729 ( .A1(n_459), .A2(n_727), .B1(n_730), .B2(n_731), .Y(n_729) );
XOR2xp5_ASAP7_75t_L g738 ( .A(n_459), .B(n_739), .Y(n_738) );
OR2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_657), .Y(n_459) );
NAND5xp2_ASAP7_75t_L g460 ( .A(n_461), .B(n_572), .C(n_604), .D(n_621), .E(n_644), .Y(n_460) );
AOI221xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_503), .B1(n_536), .B2(n_540), .C(n_544), .Y(n_461) );
INVx1_ASAP7_75t_L g684 ( .A(n_462), .Y(n_684) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_482), .Y(n_462) );
AND3x2_ASAP7_75t_L g659 ( .A(n_463), .B(n_484), .C(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_472), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_464), .B(n_542), .Y(n_541) );
BUFx3_ASAP7_75t_L g551 ( .A(n_464), .Y(n_551) );
AND2x2_ASAP7_75t_L g555 ( .A(n_464), .B(n_494), .Y(n_555) );
INVx2_ASAP7_75t_L g581 ( .A(n_464), .Y(n_581) );
OR2x2_ASAP7_75t_L g592 ( .A(n_464), .B(n_495), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_464), .B(n_483), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_464), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g671 ( .A(n_464), .B(n_495), .Y(n_671) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_472), .Y(n_554) );
AND2x2_ASAP7_75t_L g612 ( .A(n_472), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_472), .B(n_483), .Y(n_631) );
INVx1_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
OR2x2_ASAP7_75t_L g543 ( .A(n_473), .B(n_483), .Y(n_543) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_473), .Y(n_550) );
AND2x2_ASAP7_75t_L g598 ( .A(n_473), .B(n_495), .Y(n_598) );
NAND3xp33_ASAP7_75t_L g623 ( .A(n_473), .B(n_482), .C(n_581), .Y(n_623) );
AND2x2_ASAP7_75t_L g688 ( .A(n_473), .B(n_484), .Y(n_688) );
AND2x2_ASAP7_75t_L g722 ( .A(n_473), .B(n_483), .Y(n_722) );
OA21x2_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_475), .B(n_481), .Y(n_473) );
OA21x2_ASAP7_75t_L g495 ( .A1(n_474), .A2(n_496), .B(n_502), .Y(n_495) );
OA21x2_ASAP7_75t_L g528 ( .A1(n_474), .A2(n_529), .B(n_535), .Y(n_528) );
INVxp67_ASAP7_75t_L g552 ( .A(n_482), .Y(n_552) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_494), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_483), .B(n_581), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_483), .B(n_612), .Y(n_620) );
AND2x2_ASAP7_75t_L g670 ( .A(n_483), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g698 ( .A(n_483), .Y(n_698) );
INVx4_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g605 ( .A(n_484), .B(n_598), .Y(n_605) );
BUFx3_ASAP7_75t_L g637 ( .A(n_484), .Y(n_637) );
INVx2_ASAP7_75t_L g613 ( .A(n_494), .Y(n_613) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_495), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_503), .A2(n_673), .B1(n_675), .B2(n_676), .Y(n_672) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_516), .Y(n_503) );
AND2x2_ASAP7_75t_L g536 ( .A(n_504), .B(n_537), .Y(n_536) );
INVx3_ASAP7_75t_SL g547 ( .A(n_504), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_504), .B(n_576), .Y(n_608) );
OR2x2_ASAP7_75t_L g627 ( .A(n_504), .B(n_517), .Y(n_627) );
AND2x2_ASAP7_75t_L g632 ( .A(n_504), .B(n_584), .Y(n_632) );
AND2x2_ASAP7_75t_L g635 ( .A(n_504), .B(n_577), .Y(n_635) );
AND2x2_ASAP7_75t_L g647 ( .A(n_504), .B(n_528), .Y(n_647) );
AND2x2_ASAP7_75t_L g663 ( .A(n_504), .B(n_518), .Y(n_663) );
AND2x4_ASAP7_75t_L g666 ( .A(n_504), .B(n_538), .Y(n_666) );
OR2x2_ASAP7_75t_L g683 ( .A(n_504), .B(n_619), .Y(n_683) );
OR2x2_ASAP7_75t_L g714 ( .A(n_504), .B(n_560), .Y(n_714) );
NAND2xp5_ASAP7_75t_SL g716 ( .A(n_504), .B(n_642), .Y(n_716) );
OR2x6_ASAP7_75t_L g504 ( .A(n_505), .B(n_514), .Y(n_504) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_512), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g590 ( .A(n_516), .B(n_558), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_516), .B(n_577), .Y(n_709) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_528), .Y(n_516) );
AND2x2_ASAP7_75t_L g546 ( .A(n_517), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g576 ( .A(n_517), .B(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g584 ( .A(n_517), .B(n_560), .Y(n_584) );
AND2x2_ASAP7_75t_L g602 ( .A(n_517), .B(n_538), .Y(n_602) );
OR2x2_ASAP7_75t_L g619 ( .A(n_517), .B(n_577), .Y(n_619) );
INVx2_ASAP7_75t_SL g517 ( .A(n_518), .Y(n_517) );
BUFx2_ASAP7_75t_L g539 ( .A(n_518), .Y(n_539) );
AND2x2_ASAP7_75t_L g642 ( .A(n_518), .B(n_528), .Y(n_642) );
INVx2_ASAP7_75t_L g538 ( .A(n_528), .Y(n_538) );
INVx1_ASAP7_75t_L g654 ( .A(n_528), .Y(n_654) );
AND2x2_ASAP7_75t_L g704 ( .A(n_528), .B(n_547), .Y(n_704) );
AND2x2_ASAP7_75t_L g557 ( .A(n_537), .B(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g588 ( .A(n_537), .B(n_547), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_537), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
AND2x2_ASAP7_75t_L g575 ( .A(n_538), .B(n_547), .Y(n_575) );
OR2x2_ASAP7_75t_L g691 ( .A(n_539), .B(n_665), .Y(n_691) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_542), .B(n_671), .Y(n_677) );
INVx2_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
OAI32xp33_ASAP7_75t_L g633 ( .A1(n_543), .A2(n_634), .A3(n_636), .B1(n_638), .B2(n_639), .Y(n_633) );
OR2x2_ASAP7_75t_L g650 ( .A(n_543), .B(n_592), .Y(n_650) );
OAI21xp33_ASAP7_75t_SL g675 ( .A1(n_543), .A2(n_553), .B(n_580), .Y(n_675) );
OAI22xp33_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_548), .B1(n_553), .B2(n_556), .Y(n_544) );
INVxp33_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_546), .B(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_547), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g601 ( .A(n_547), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g701 ( .A(n_547), .B(n_642), .Y(n_701) );
OR2x2_ASAP7_75t_L g725 ( .A(n_547), .B(n_619), .Y(n_725) );
AOI21xp33_ASAP7_75t_L g708 ( .A1(n_548), .A2(n_607), .B(n_709), .Y(n_708) );
OR2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_552), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
INVx1_ASAP7_75t_L g585 ( .A(n_550), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_550), .B(n_555), .Y(n_603) );
AND2x2_ASAP7_75t_L g625 ( .A(n_551), .B(n_598), .Y(n_625) );
INVx1_ASAP7_75t_L g638 ( .A(n_551), .Y(n_638) );
OR2x2_ASAP7_75t_L g643 ( .A(n_551), .B(n_577), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_554), .B(n_592), .Y(n_591) );
OAI22xp33_ASAP7_75t_L g573 ( .A1(n_555), .A2(n_574), .B1(n_579), .B2(n_583), .Y(n_573) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_558), .A2(n_616), .B1(n_623), .B2(n_624), .Y(n_622) );
AND2x2_ASAP7_75t_L g700 ( .A(n_558), .B(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_SL g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_560), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g719 ( .A(n_560), .B(n_602), .Y(n_719) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
OA21x2_ASAP7_75t_L g577 ( .A1(n_562), .A2(n_570), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AOI221xp5_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_585), .B1(n_586), .B2(n_591), .C(n_593), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_575), .B(n_577), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_575), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g594 ( .A(n_576), .Y(n_594) );
O2A1O1Ixp33_ASAP7_75t_L g681 ( .A1(n_576), .A2(n_682), .B(n_683), .C(n_684), .Y(n_681) );
AND2x2_ASAP7_75t_L g686 ( .A(n_576), .B(n_666), .Y(n_686) );
O2A1O1Ixp33_ASAP7_75t_SL g724 ( .A1(n_576), .A2(n_665), .B(n_725), .C(n_726), .Y(n_724) );
BUFx3_ASAP7_75t_L g616 ( .A(n_577), .Y(n_616) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_580), .B(n_637), .Y(n_680) );
AOI211xp5_ASAP7_75t_L g699 ( .A1(n_580), .A2(n_700), .B(n_702), .C(n_708), .Y(n_699) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
INVxp67_ASAP7_75t_L g660 ( .A(n_582), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_584), .B(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_587), .B(n_589), .Y(n_586) );
INVx1_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
AOI211xp5_ASAP7_75t_L g604 ( .A1(n_588), .A2(n_605), .B(n_606), .C(n_614), .Y(n_604) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g689 ( .A(n_592), .Y(n_689) );
OR2x2_ASAP7_75t_L g706 ( .A(n_592), .B(n_636), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_595), .B1(n_600), .B2(n_603), .Y(n_593) );
OAI22xp33_ASAP7_75t_L g606 ( .A1(n_595), .A2(n_607), .B1(n_608), .B2(n_609), .Y(n_606) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_599), .Y(n_596) );
OR2x2_ASAP7_75t_L g693 ( .A(n_597), .B(n_637), .Y(n_693) );
INVx1_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g648 ( .A(n_598), .B(n_638), .Y(n_648) );
INVx1_ASAP7_75t_L g656 ( .A(n_599), .Y(n_656) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_602), .B(n_616), .Y(n_664) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
NAND2xp5_ASAP7_75t_SL g655 ( .A(n_612), .B(n_656), .Y(n_655) );
INVx2_ASAP7_75t_L g721 ( .A(n_613), .Y(n_721) );
AOI21xp33_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_617), .B(n_620), .Y(n_614) );
INVx1_ASAP7_75t_L g651 ( .A(n_615), .Y(n_651) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_616), .B(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_616), .B(n_647), .Y(n_646) );
NAND2x1p5_ASAP7_75t_L g667 ( .A(n_616), .B(n_642), .Y(n_667) );
NAND2xp5_ASAP7_75t_SL g674 ( .A(n_616), .B(n_663), .Y(n_674) );
OAI211xp5_ASAP7_75t_L g678 ( .A1(n_616), .A2(n_626), .B(n_666), .C(n_679), .Y(n_678) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
AOI221xp5_ASAP7_75t_SL g621 ( .A1(n_622), .A2(n_626), .B1(n_628), .B2(n_632), .C(n_633), .Y(n_621) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVxp67_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_630), .B(n_638), .Y(n_712) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
O2A1O1Ixp33_ASAP7_75t_L g723 ( .A1(n_632), .A2(n_647), .B(n_649), .C(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_635), .B(n_642), .Y(n_707) );
NAND2xp5_ASAP7_75t_SL g726 ( .A(n_636), .B(n_689), .Y(n_726) );
CKINVDCx16_ASAP7_75t_R g636 ( .A(n_637), .Y(n_636) );
INVxp33_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .Y(n_640) );
AOI21xp33_ASAP7_75t_SL g652 ( .A1(n_641), .A2(n_653), .B(n_655), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_641), .B(n_714), .Y(n_713) );
INVx2_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_642), .B(n_696), .Y(n_695) );
AOI221xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_648), .B1(n_649), .B2(n_651), .C(n_652), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_648), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g682 ( .A(n_654), .Y(n_682) );
NAND5xp2_ASAP7_75t_L g657 ( .A(n_658), .B(n_685), .C(n_699), .D(n_710), .E(n_723), .Y(n_657) );
AOI211xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_661), .B(n_668), .C(n_681), .Y(n_658) );
INVx2_ASAP7_75t_SL g705 ( .A(n_659), .Y(n_705) );
NAND4xp25_ASAP7_75t_SL g661 ( .A(n_662), .B(n_664), .C(n_665), .D(n_667), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx3_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OAI211xp5_ASAP7_75t_SL g668 ( .A1(n_667), .A2(n_669), .B(n_672), .C(n_678), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g669 ( .A(n_670), .Y(n_669) );
AOI221xp5_ASAP7_75t_L g710 ( .A1(n_670), .A2(n_711), .B1(n_713), .B2(n_715), .C(n_717), .Y(n_710) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AOI221xp5_ASAP7_75t_SL g685 ( .A1(n_686), .A2(n_687), .B1(n_690), .B2(n_692), .C(n_694), .Y(n_685) );
AND2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_693), .A2(n_716), .B1(n_718), .B2(n_720), .Y(n_717) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_705), .B1(n_706), .B2(n_707), .Y(n_702) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
INVx3_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_744), .Y(n_743) );
endmodule