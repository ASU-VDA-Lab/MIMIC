module fake_netlist_1_8082_n_35 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_35);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_35;
wire n_20;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_13;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_0), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_8), .Y(n_12) );
AOI21x1_ASAP7_75t_L g13 ( .A1(n_1), .A2(n_3), .B(n_6), .Y(n_13) );
AND2x2_ASAP7_75t_L g14 ( .A(n_5), .B(n_1), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_2), .Y(n_15) );
NOR2xp33_ASAP7_75t_R g16 ( .A(n_11), .B(n_0), .Y(n_16) );
O2A1O1Ixp33_ASAP7_75t_L g17 ( .A1(n_14), .A2(n_0), .B(n_1), .C(n_2), .Y(n_17) );
A2O1A1Ixp33_ASAP7_75t_L g18 ( .A1(n_14), .A2(n_3), .B(n_4), .C(n_6), .Y(n_18) );
AND2x4_ASAP7_75t_L g19 ( .A(n_14), .B(n_11), .Y(n_19) );
NAND2xp5_ASAP7_75t_SL g20 ( .A(n_12), .B(n_4), .Y(n_20) );
CKINVDCx5p33_ASAP7_75t_R g21 ( .A(n_16), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_19), .B(n_12), .Y(n_22) );
NAND2xp33_ASAP7_75t_L g23 ( .A(n_18), .B(n_15), .Y(n_23) );
CKINVDCx5p33_ASAP7_75t_R g24 ( .A(n_16), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_22), .Y(n_25) );
AND2x4_ASAP7_75t_SL g26 ( .A(n_22), .B(n_19), .Y(n_26) );
OR2x2_ASAP7_75t_L g27 ( .A(n_22), .B(n_20), .Y(n_27) );
INVxp67_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
NAND3xp33_ASAP7_75t_L g29 ( .A(n_27), .B(n_24), .C(n_21), .Y(n_29) );
NAND4xp25_ASAP7_75t_L g30 ( .A(n_28), .B(n_17), .C(n_29), .D(n_26), .Y(n_30) );
NAND3xp33_ASAP7_75t_L g31 ( .A(n_29), .B(n_23), .C(n_24), .Y(n_31) );
INVx2_ASAP7_75t_L g32 ( .A(n_31), .Y(n_32) );
NOR2x1_ASAP7_75t_L g33 ( .A(n_30), .B(n_23), .Y(n_33) );
NAND2x1_ASAP7_75t_L g34 ( .A(n_32), .B(n_13), .Y(n_34) );
AOI322xp5_ASAP7_75t_L g35 ( .A1(n_34), .A2(n_33), .A3(n_13), .B1(n_9), .B2(n_10), .C1(n_8), .C2(n_7), .Y(n_35) );
endmodule