module fake_ariane_514_n_1592 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_332, n_294, n_197, n_176, n_34, n_172, n_347, n_183, n_373, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_349, n_346, n_214, n_348, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_327, n_77, n_372, n_377, n_15, n_23, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_267, n_335, n_350, n_291, n_344, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_333, n_376, n_221, n_321, n_86, n_361, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_343, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_366, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_378, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_159, n_358, n_105, n_30, n_131, n_263, n_360, n_229, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_364, n_258, n_118, n_121, n_353, n_22, n_241, n_29, n_357, n_191, n_80, n_211, n_97, n_322, n_251, n_116, n_351, n_39, n_359, n_155, n_127, n_1592);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_347;
input n_183;
input n_373;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_267;
input n_335;
input n_350;
input n_291;
input n_344;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_333;
input n_376;
input n_221;
input n_321;
input n_86;
input n_361;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_343;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_378;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_360;
input n_229;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_118;
input n_121;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_191;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_351;
input n_39;
input n_359;
input n_155;
input n_127;

output n_1592;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_995;
wire n_1184;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_559;
wire n_495;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_611;
wire n_1295;
wire n_1013;
wire n_1495;
wire n_661;
wire n_533;
wire n_438;
wire n_1560;
wire n_1548;
wire n_440;
wire n_1396;
wire n_1230;
wire n_612;
wire n_512;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_380;
wire n_1585;
wire n_1432;
wire n_1108;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_762;
wire n_1253;
wire n_1468;
wire n_555;
wire n_804;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_436;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_698;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_404;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_706;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_1467;
wire n_1304;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1489;
wire n_1218;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_551;
wire n_417;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_1352;
wire n_643;
wire n_1492;
wire n_1441;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_1521;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1444;
wire n_820;
wire n_872;
wire n_1157;
wire n_1584;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_1552;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1587;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1482;
wire n_1361;
wire n_1057;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1458;
wire n_679;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_1479;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1571;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1591;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_946;
wire n_757;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1474;
wire n_1583;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_1129;
wire n_1252;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_1434;
wire n_1569;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

BUFx3_ASAP7_75t_L g379 ( 
.A(n_278),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_202),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_330),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_21),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_264),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_132),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_271),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_261),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_218),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_295),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_182),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_353),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_68),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_126),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_354),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_52),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_374),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_83),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_260),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_336),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_193),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_294),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_177),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_165),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_65),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_204),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_82),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_314),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_109),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_34),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_87),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_365),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_174),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_17),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_27),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_311),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_175),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_26),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_363),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_302),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_340),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_122),
.Y(n_420)
);

BUFx10_ASAP7_75t_L g421 ( 
.A(n_241),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_89),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_364),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_53),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_307),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_22),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_373),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_155),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_237),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_181),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_90),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_9),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_283),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_229),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_250),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_22),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_96),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_301),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_55),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_228),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_350),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_221),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_227),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_323),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_274),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_169),
.Y(n_446)
);

BUFx10_ASAP7_75t_L g447 ( 
.A(n_209),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_85),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_15),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_246),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_152),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_179),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_28),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_377),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_94),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_5),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_116),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g458 ( 
.A(n_326),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_316),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_62),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_52),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_304),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_105),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_259),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_240),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_258),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_200),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_92),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_226),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_21),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_308),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_113),
.Y(n_472)
);

BUFx5_ASAP7_75t_L g473 ( 
.A(n_223),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_78),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_168),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_366),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_134),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_254),
.Y(n_478)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_232),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_28),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g481 ( 
.A(n_355),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_189),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_49),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_103),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_245),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_59),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_63),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_173),
.Y(n_488)
);

BUFx10_ASAP7_75t_L g489 ( 
.A(n_266),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_262),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_101),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_3),
.Y(n_492)
);

CKINVDCx14_ASAP7_75t_R g493 ( 
.A(n_220),
.Y(n_493)
);

INVx2_ASAP7_75t_SL g494 ( 
.A(n_203),
.Y(n_494)
);

BUFx8_ASAP7_75t_SL g495 ( 
.A(n_357),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_71),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_312),
.Y(n_497)
);

INVxp33_ASAP7_75t_L g498 ( 
.A(n_170),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_305),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_137),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_178),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_325),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_293),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_372),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_320),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_239),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_248),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_12),
.Y(n_508)
);

INVxp67_ASAP7_75t_SL g509 ( 
.A(n_34),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_345),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_318),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_17),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_91),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_216),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_147),
.Y(n_515)
);

CKINVDCx16_ASAP7_75t_R g516 ( 
.A(n_371),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_184),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_75),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_104),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_171),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_131),
.Y(n_521)
);

BUFx10_ASAP7_75t_L g522 ( 
.A(n_121),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_327),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_44),
.Y(n_524)
);

INVxp67_ASAP7_75t_SL g525 ( 
.A(n_13),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_199),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_157),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_102),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_125),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_166),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_110),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_289),
.Y(n_532)
);

BUFx8_ASAP7_75t_SL g533 ( 
.A(n_67),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_107),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_40),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_257),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_244),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_129),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_160),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_196),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_58),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_303),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_344),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_284),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_55),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g546 ( 
.A(n_356),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_315),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_32),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_253),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_328),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_154),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_12),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_29),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_251),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_298),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_144),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_279),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_339),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_93),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_243),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_111),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_201),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_367),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_321),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_225),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_58),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_288),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_1),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_79),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_164),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_42),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_382),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_495),
.Y(n_573)
);

BUFx2_ASAP7_75t_L g574 ( 
.A(n_545),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_394),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_410),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_408),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_379),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_391),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_495),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_456),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_490),
.B(n_0),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_533),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_533),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_461),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_483),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_469),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_492),
.Y(n_588)
);

INVxp67_ASAP7_75t_SL g589 ( 
.A(n_456),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_412),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_524),
.Y(n_591)
);

INVxp67_ASAP7_75t_SL g592 ( 
.A(n_460),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_534),
.B(n_0),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_553),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_568),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_510),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_527),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_528),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_571),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_542),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_460),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_498),
.B(n_1),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_413),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_530),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_489),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_489),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_391),
.Y(n_607)
);

INVxp67_ASAP7_75t_SL g608 ( 
.A(n_509),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g609 ( 
.A(n_416),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_426),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_493),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_522),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_522),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_432),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_421),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_421),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_436),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_421),
.Y(n_618)
);

INVxp67_ASAP7_75t_SL g619 ( 
.A(n_498),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_381),
.B(n_390),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_447),
.Y(n_621)
);

INVxp67_ASAP7_75t_SL g622 ( 
.A(n_525),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_447),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_439),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_447),
.Y(n_625)
);

INVxp67_ASAP7_75t_L g626 ( 
.A(n_449),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g627 ( 
.A(n_493),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_391),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_453),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_415),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_395),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_470),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_396),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_397),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_402),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_480),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_404),
.Y(n_637)
);

NOR2xp67_ASAP7_75t_L g638 ( 
.A(n_486),
.B(n_2),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_407),
.Y(n_639)
);

BUFx2_ASAP7_75t_SL g640 ( 
.A(n_379),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_487),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_475),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_481),
.Y(n_643)
);

CKINVDCx20_ASAP7_75t_R g644 ( 
.A(n_516),
.Y(n_644)
);

CKINVDCx20_ASAP7_75t_R g645 ( 
.A(n_475),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_417),
.Y(n_646)
);

CKINVDCx20_ASAP7_75t_R g647 ( 
.A(n_502),
.Y(n_647)
);

CKINVDCx20_ASAP7_75t_R g648 ( 
.A(n_502),
.Y(n_648)
);

CKINVDCx16_ASAP7_75t_R g649 ( 
.A(n_424),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_508),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_512),
.Y(n_651)
);

CKINVDCx16_ASAP7_75t_R g652 ( 
.A(n_391),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_419),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_535),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_422),
.Y(n_655)
);

CKINVDCx20_ASAP7_75t_R g656 ( 
.A(n_541),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_548),
.B(n_2),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_433),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_552),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_566),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_437),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_380),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_570),
.Y(n_663)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_383),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_438),
.B(n_3),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_443),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_446),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_384),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_385),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_448),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_386),
.Y(n_671)
);

BUFx2_ASAP7_75t_L g672 ( 
.A(n_451),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_452),
.Y(n_673)
);

CKINVDCx16_ASAP7_75t_R g674 ( 
.A(n_472),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_472),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_455),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_387),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_464),
.Y(n_678)
);

CKINVDCx20_ASAP7_75t_R g679 ( 
.A(n_569),
.Y(n_679)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_388),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_468),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_474),
.Y(n_682)
);

CKINVDCx20_ASAP7_75t_R g683 ( 
.A(n_567),
.Y(n_683)
);

NOR2xp67_ASAP7_75t_L g684 ( 
.A(n_476),
.B(n_4),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_482),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_488),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_491),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_L g688 ( 
.A1(n_619),
.A2(n_501),
.B1(n_505),
.B2(n_499),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_621),
.B(n_431),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_596),
.Y(n_690)
);

HB1xp67_ASAP7_75t_L g691 ( 
.A(n_574),
.Y(n_691)
);

AND2x4_ASAP7_75t_L g692 ( 
.A(n_605),
.B(n_458),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_572),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_579),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_579),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_579),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_579),
.Y(n_697)
);

CKINVDCx20_ASAP7_75t_R g698 ( 
.A(n_603),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_649),
.B(n_485),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_575),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_597),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_577),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_598),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_600),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_573),
.Y(n_705)
);

CKINVDCx20_ASAP7_75t_R g706 ( 
.A(n_576),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_585),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_586),
.Y(n_708)
);

XNOR2xp5_ASAP7_75t_L g709 ( 
.A(n_587),
.B(n_546),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_580),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_588),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_591),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_594),
.Y(n_713)
);

INVx3_ASAP7_75t_L g714 ( 
.A(n_652),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_611),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_583),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_595),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_599),
.Y(n_718)
);

CKINVDCx20_ASAP7_75t_R g719 ( 
.A(n_627),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_589),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_630),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_589),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_592),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_592),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_674),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_626),
.B(n_479),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_607),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_615),
.B(n_511),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_607),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_R g730 ( 
.A(n_584),
.B(n_389),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_578),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_607),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_SL g733 ( 
.A1(n_643),
.A2(n_520),
.B1(n_523),
.B2(n_521),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_607),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_642),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_687),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_668),
.Y(n_737)
);

HB1xp67_ASAP7_75t_L g738 ( 
.A(n_610),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_628),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_644),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_669),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_628),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_606),
.B(n_494),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_616),
.B(n_526),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_628),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_671),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_686),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_677),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_685),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_631),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_662),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_633),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_593),
.A2(n_531),
.B1(n_536),
.B2(n_529),
.Y(n_753)
);

CKINVDCx16_ASAP7_75t_R g754 ( 
.A(n_650),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_663),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_R g756 ( 
.A(n_664),
.B(n_392),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_634),
.Y(n_757)
);

NAND2xp33_ASAP7_75t_SL g758 ( 
.A(n_582),
.B(n_537),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_590),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_618),
.B(n_543),
.Y(n_760)
);

AND2x4_ASAP7_75t_L g761 ( 
.A(n_612),
.B(n_544),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_679),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_628),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_675),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_623),
.B(n_549),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_675),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_675),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_625),
.B(n_559),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_613),
.B(n_560),
.Y(n_769)
);

HB1xp67_ASAP7_75t_L g770 ( 
.A(n_614),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_656),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_680),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_675),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_635),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_637),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_683),
.Y(n_776)
);

NAND2xp33_ASAP7_75t_SL g777 ( 
.A(n_657),
.B(n_562),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_617),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_731),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_735),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_693),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_714),
.B(n_629),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_699),
.B(n_632),
.Y(n_783)
);

NAND2xp33_ASAP7_75t_L g784 ( 
.A(n_737),
.B(n_636),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_700),
.Y(n_785)
);

NOR2x1p5_ASAP7_75t_L g786 ( 
.A(n_741),
.B(n_746),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_734),
.Y(n_787)
);

BUFx10_ASAP7_75t_L g788 ( 
.A(n_778),
.Y(n_788)
);

NAND3xp33_ASAP7_75t_L g789 ( 
.A(n_777),
.B(n_620),
.C(n_602),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_702),
.Y(n_790)
);

OR2x2_ASAP7_75t_L g791 ( 
.A(n_691),
.B(n_609),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_707),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_714),
.B(n_641),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_736),
.B(n_639),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_695),
.Y(n_795)
);

OR2x2_ASAP7_75t_L g796 ( 
.A(n_691),
.B(n_624),
.Y(n_796)
);

INVx5_ASAP7_75t_L g797 ( 
.A(n_725),
.Y(n_797)
);

NOR3xp33_ASAP7_75t_L g798 ( 
.A(n_777),
.B(n_665),
.C(n_622),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_708),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_725),
.B(n_608),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_739),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_742),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_695),
.Y(n_803)
);

OAI22xp33_ASAP7_75t_L g804 ( 
.A1(n_753),
.A2(n_622),
.B1(n_608),
.B2(n_672),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_688),
.A2(n_604),
.B1(n_684),
.B2(n_653),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_720),
.B(n_651),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_745),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_695),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_722),
.B(n_626),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_747),
.B(n_646),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_749),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_748),
.B(n_645),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_723),
.B(n_647),
.Y(n_813)
);

INVx4_ASAP7_75t_SL g814 ( 
.A(n_733),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_L g815 ( 
.A1(n_758),
.A2(n_655),
.B1(n_661),
.B2(n_658),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_689),
.B(n_648),
.Y(n_816)
);

INVx3_ASAP7_75t_L g817 ( 
.A(n_750),
.Y(n_817)
);

OR2x2_ASAP7_75t_L g818 ( 
.A(n_759),
.B(n_654),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_758),
.A2(n_761),
.B1(n_757),
.B2(n_752),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_724),
.B(n_640),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_764),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_730),
.B(n_659),
.Y(n_822)
);

OAI22xp33_ASAP7_75t_L g823 ( 
.A1(n_759),
.A2(n_581),
.B1(n_638),
.B2(n_660),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_738),
.B(n_581),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_711),
.A2(n_666),
.B1(n_670),
.B2(n_667),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_751),
.Y(n_826)
);

OR2x2_ASAP7_75t_L g827 ( 
.A(n_754),
.B(n_682),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_738),
.B(n_673),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_695),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_730),
.B(n_676),
.Y(n_830)
);

OAI22xp5_ASAP7_75t_L g831 ( 
.A1(n_769),
.A2(n_678),
.B1(n_681),
.B2(n_601),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_729),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_766),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_773),
.Y(n_834)
);

INVx2_ASAP7_75t_SL g835 ( 
.A(n_756),
.Y(n_835)
);

NAND2x1_ASAP7_75t_L g836 ( 
.A(n_774),
.B(n_775),
.Y(n_836)
);

BUFx4f_ASAP7_75t_L g837 ( 
.A(n_761),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_726),
.B(n_393),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_712),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_756),
.B(n_398),
.Y(n_840)
);

INVx5_ASAP7_75t_L g841 ( 
.A(n_729),
.Y(n_841)
);

INVx4_ASAP7_75t_L g842 ( 
.A(n_692),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_694),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_694),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_713),
.Y(n_845)
);

INVx2_ASAP7_75t_SL g846 ( 
.A(n_770),
.Y(n_846)
);

OR2x6_ASAP7_75t_L g847 ( 
.A(n_770),
.B(n_472),
.Y(n_847)
);

CKINVDCx20_ASAP7_75t_R g848 ( 
.A(n_706),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_692),
.B(n_399),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_728),
.B(n_473),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_743),
.B(n_769),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_743),
.B(n_400),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_696),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_744),
.B(n_401),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_760),
.B(n_403),
.Y(n_855)
);

INVx5_ASAP7_75t_L g856 ( 
.A(n_729),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_696),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_705),
.B(n_405),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_710),
.B(n_406),
.Y(n_859)
);

INVx3_ASAP7_75t_L g860 ( 
.A(n_697),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_765),
.B(n_473),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_717),
.A2(n_718),
.B1(n_768),
.B2(n_507),
.Y(n_862)
);

AND2x4_ASAP7_75t_L g863 ( 
.A(n_690),
.B(n_472),
.Y(n_863)
);

INVx5_ASAP7_75t_L g864 ( 
.A(n_729),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_697),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_727),
.Y(n_866)
);

AO22x2_ASAP7_75t_L g867 ( 
.A1(n_709),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_781),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_813),
.Y(n_869)
);

NOR2x1p5_ASAP7_75t_L g870 ( 
.A(n_818),
.B(n_716),
.Y(n_870)
);

BUFx2_ASAP7_75t_L g871 ( 
.A(n_848),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_837),
.B(n_701),
.Y(n_872)
);

AND2x4_ASAP7_75t_L g873 ( 
.A(n_797),
.B(n_703),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_826),
.Y(n_874)
);

INVx5_ASAP7_75t_L g875 ( 
.A(n_847),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_779),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_820),
.B(n_854),
.Y(n_877)
);

A2O1A1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_789),
.A2(n_809),
.B(n_798),
.C(n_806),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_855),
.B(n_704),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_838),
.B(n_409),
.Y(n_880)
);

AOI22xp5_ASAP7_75t_L g881 ( 
.A1(n_798),
.A2(n_762),
.B1(n_772),
.B2(n_755),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_811),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_811),
.B(n_411),
.Y(n_883)
);

INVxp67_ASAP7_75t_L g884 ( 
.A(n_783),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_837),
.B(n_776),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_780),
.Y(n_886)
);

BUFx8_ASAP7_75t_L g887 ( 
.A(n_846),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_843),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_782),
.B(n_771),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_785),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_844),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_817),
.B(n_800),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_790),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_816),
.B(n_721),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_792),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_817),
.B(n_414),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_799),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_793),
.B(n_418),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_800),
.B(n_420),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_824),
.B(n_423),
.Y(n_900)
);

CKINVDCx20_ASAP7_75t_R g901 ( 
.A(n_788),
.Y(n_901)
);

INVx2_ASAP7_75t_SL g902 ( 
.A(n_847),
.Y(n_902)
);

NAND3xp33_ASAP7_75t_L g903 ( 
.A(n_784),
.B(n_789),
.C(n_828),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_797),
.B(n_425),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_863),
.B(n_427),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_795),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_839),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_863),
.B(n_845),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_819),
.B(n_428),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_794),
.Y(n_910)
);

A2O1A1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_850),
.A2(n_861),
.B(n_851),
.C(n_810),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_794),
.Y(n_912)
);

AND2x2_ASAP7_75t_SL g913 ( 
.A(n_827),
.B(n_740),
.Y(n_913)
);

INVx5_ASAP7_75t_L g914 ( 
.A(n_847),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_SL g915 ( 
.A1(n_805),
.A2(n_698),
.B1(n_719),
.B2(n_715),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_835),
.B(n_429),
.Y(n_916)
);

INVx2_ASAP7_75t_SL g917 ( 
.A(n_797),
.Y(n_917)
);

INVx2_ASAP7_75t_SL g918 ( 
.A(n_791),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_788),
.B(n_6),
.Y(n_919)
);

NAND3xp33_ASAP7_75t_L g920 ( 
.A(n_850),
.B(n_763),
.C(n_727),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_853),
.Y(n_921)
);

NAND2xp33_ASAP7_75t_SL g922 ( 
.A(n_786),
.B(n_430),
.Y(n_922)
);

NAND3xp33_ASAP7_75t_L g923 ( 
.A(n_858),
.B(n_859),
.C(n_815),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_810),
.B(n_434),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_796),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_857),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_823),
.B(n_435),
.Y(n_927)
);

NAND2xp33_ASAP7_75t_L g928 ( 
.A(n_861),
.B(n_852),
.Y(n_928)
);

INVxp67_ASAP7_75t_L g929 ( 
.A(n_812),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_836),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_842),
.B(n_440),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_823),
.B(n_441),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_815),
.B(n_442),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_842),
.B(n_444),
.Y(n_934)
);

OR2x2_ASAP7_75t_L g935 ( 
.A(n_822),
.B(n_7),
.Y(n_935)
);

NAND3xp33_ASAP7_75t_L g936 ( 
.A(n_831),
.B(n_763),
.C(n_767),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_830),
.B(n_840),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_849),
.B(n_445),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_804),
.A2(n_454),
.B1(n_457),
.B2(n_450),
.Y(n_939)
);

O2A1O1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_831),
.A2(n_804),
.B(n_825),
.C(n_865),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_795),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_862),
.B(n_459),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_860),
.B(n_462),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_825),
.A2(n_465),
.B1(n_466),
.B2(n_463),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_814),
.B(n_7),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_866),
.Y(n_946)
);

NAND2x1_ASAP7_75t_L g947 ( 
.A(n_860),
.B(n_767),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_787),
.B(n_467),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_814),
.B(n_8),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_867),
.B(n_8),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_801),
.B(n_471),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_802),
.B(n_477),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_807),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_SL g954 ( 
.A(n_867),
.B(n_478),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_821),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_833),
.B(n_484),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_834),
.B(n_496),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_841),
.A2(n_500),
.B1(n_503),
.B2(n_497),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_795),
.B(n_504),
.Y(n_959)
);

AO22x1_ASAP7_75t_L g960 ( 
.A1(n_841),
.A2(n_513),
.B1(n_514),
.B2(n_506),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_803),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_803),
.B(n_515),
.Y(n_962)
);

NOR3x1_ASAP7_75t_L g963 ( 
.A(n_864),
.B(n_9),
.C(n_10),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_803),
.B(n_517),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_868),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_877),
.A2(n_829),
.B(n_808),
.Y(n_966)
);

OAI21xp5_ASAP7_75t_L g967 ( 
.A1(n_911),
.A2(n_856),
.B(n_841),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_869),
.A2(n_518),
.B1(n_532),
.B2(n_519),
.Y(n_968)
);

OAI21xp5_ASAP7_75t_L g969 ( 
.A1(n_920),
.A2(n_864),
.B(n_856),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_890),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_928),
.A2(n_829),
.B(n_808),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_R g972 ( 
.A(n_901),
.B(n_808),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_910),
.B(n_829),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_893),
.Y(n_974)
);

OAI22xp5_ASAP7_75t_L g975 ( 
.A1(n_878),
.A2(n_832),
.B1(n_538),
.B2(n_540),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_912),
.B(n_832),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_879),
.B(n_832),
.Y(n_977)
);

O2A1O1Ixp33_ASAP7_75t_SL g978 ( 
.A1(n_898),
.A2(n_880),
.B(n_896),
.C(n_883),
.Y(n_978)
);

HB1xp67_ASAP7_75t_L g979 ( 
.A(n_918),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_L g980 ( 
.A1(n_920),
.A2(n_864),
.B(n_856),
.Y(n_980)
);

AOI22xp5_ASAP7_75t_L g981 ( 
.A1(n_923),
.A2(n_539),
.B1(n_550),
.B2(n_547),
.Y(n_981)
);

NAND2xp33_ASAP7_75t_L g982 ( 
.A(n_882),
.B(n_473),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_892),
.B(n_551),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_924),
.A2(n_555),
.B(n_554),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_934),
.A2(n_557),
.B(n_556),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_930),
.A2(n_561),
.B(n_558),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_882),
.B(n_563),
.Y(n_987)
);

BUFx2_ASAP7_75t_L g988 ( 
.A(n_871),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_903),
.A2(n_564),
.B1(n_565),
.B2(n_507),
.Y(n_989)
);

HB1xp67_ASAP7_75t_L g990 ( 
.A(n_925),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_884),
.B(n_10),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_931),
.A2(n_507),
.B(n_732),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_876),
.Y(n_993)
);

OR2x2_ASAP7_75t_L g994 ( 
.A(n_889),
.B(n_11),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_937),
.A2(n_507),
.B(n_732),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_L g996 ( 
.A1(n_908),
.A2(n_473),
.B1(n_732),
.B2(n_14),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_947),
.A2(n_732),
.B(n_473),
.Y(n_997)
);

BUFx3_ASAP7_75t_L g998 ( 
.A(n_874),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_875),
.B(n_473),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_895),
.A2(n_66),
.B(n_64),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_897),
.A2(n_70),
.B(n_69),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_907),
.B(n_11),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_886),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_887),
.Y(n_1004)
);

INVx2_ASAP7_75t_SL g1005 ( 
.A(n_887),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_936),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_936),
.A2(n_73),
.B(n_72),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_900),
.A2(n_961),
.B(n_905),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_953),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_888),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_940),
.A2(n_15),
.B(n_13),
.C(n_14),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_916),
.B(n_16),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_959),
.A2(n_964),
.B(n_943),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_929),
.B(n_16),
.Y(n_1014)
);

AOI21xp33_ASAP7_75t_L g1015 ( 
.A1(n_939),
.A2(n_18),
.B(n_19),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_875),
.B(n_18),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_872),
.A2(n_23),
.B(n_19),
.C(n_20),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_913),
.B(n_20),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_875),
.B(n_23),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_914),
.B(n_899),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_914),
.B(n_24),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_881),
.B(n_914),
.Y(n_1022)
);

O2A1O1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_885),
.A2(n_927),
.B(n_932),
.C(n_904),
.Y(n_1023)
);

BUFx12f_ASAP7_75t_L g1024 ( 
.A(n_873),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_906),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_902),
.B(n_24),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_881),
.B(n_25),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_891),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_917),
.A2(n_76),
.B(n_74),
.Y(n_1029)
);

HB1xp67_ASAP7_75t_L g1030 ( 
.A(n_873),
.Y(n_1030)
);

O2A1O1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_933),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_948),
.A2(n_80),
.B(n_77),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_870),
.B(n_894),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_915),
.B(n_29),
.Y(n_1034)
);

AND2x2_ASAP7_75t_SL g1035 ( 
.A(n_954),
.B(n_30),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_909),
.B(n_30),
.Y(n_1036)
);

NOR2xp67_ASAP7_75t_L g1037 ( 
.A(n_938),
.B(n_81),
.Y(n_1037)
);

AND2x6_ASAP7_75t_L g1038 ( 
.A(n_949),
.B(n_84),
.Y(n_1038)
);

BUFx4f_ASAP7_75t_L g1039 ( 
.A(n_949),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_906),
.Y(n_1040)
);

INVxp67_ASAP7_75t_L g1041 ( 
.A(n_915),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_951),
.A2(n_956),
.B(n_952),
.Y(n_1042)
);

AOI22xp33_ASAP7_75t_L g1043 ( 
.A1(n_950),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_978),
.A2(n_960),
.B(n_962),
.Y(n_1044)
);

INVx2_ASAP7_75t_SL g1045 ( 
.A(n_1039),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_1013),
.A2(n_941),
.B(n_906),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_965),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_982),
.A2(n_941),
.B(n_957),
.Y(n_1048)
);

BUFx8_ASAP7_75t_L g1049 ( 
.A(n_1024),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_977),
.A2(n_941),
.B(n_922),
.Y(n_1050)
);

OAI21x1_ASAP7_75t_L g1051 ( 
.A1(n_967),
.A2(n_926),
.B(n_921),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_1027),
.A2(n_935),
.B(n_919),
.C(n_945),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_998),
.B(n_1030),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_1039),
.B(n_944),
.Y(n_1054)
);

AOI211x1_ASAP7_75t_L g1055 ( 
.A1(n_1015),
.A2(n_963),
.B(n_958),
.C(n_942),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_966),
.A2(n_946),
.B(n_955),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_970),
.Y(n_1057)
);

INVx2_ASAP7_75t_SL g1058 ( 
.A(n_972),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_974),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_1033),
.B(n_31),
.Y(n_1060)
);

AO31x2_ASAP7_75t_L g1061 ( 
.A1(n_1006),
.A2(n_206),
.A3(n_376),
.B(n_375),
.Y(n_1061)
);

OAI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_1008),
.A2(n_33),
.B(n_35),
.Y(n_1062)
);

AOI21x1_ASAP7_75t_L g1063 ( 
.A1(n_971),
.A2(n_88),
.B(n_86),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_1022),
.B(n_35),
.Y(n_1064)
);

INVx5_ASAP7_75t_L g1065 ( 
.A(n_1038),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_979),
.B(n_36),
.Y(n_1066)
);

OAI21x1_ASAP7_75t_L g1067 ( 
.A1(n_969),
.A2(n_97),
.B(n_95),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_1020),
.B(n_36),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1009),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_1025),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_991),
.A2(n_37),
.B(n_38),
.C(n_39),
.Y(n_1071)
);

OAI21xp33_ASAP7_75t_SL g1072 ( 
.A1(n_1012),
.A2(n_37),
.B(n_38),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_990),
.B(n_39),
.Y(n_1073)
);

AND3x4_ASAP7_75t_L g1074 ( 
.A(n_1004),
.B(n_40),
.C(n_41),
.Y(n_1074)
);

O2A1O1Ixp5_ASAP7_75t_L g1075 ( 
.A1(n_1036),
.A2(n_41),
.B(n_42),
.C(n_43),
.Y(n_1075)
);

CKINVDCx14_ASAP7_75t_R g1076 ( 
.A(n_988),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_1042),
.A2(n_99),
.B(n_98),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_980),
.A2(n_106),
.B(n_100),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1014),
.B(n_43),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_995),
.A2(n_112),
.B(n_108),
.Y(n_1080)
);

OAI22x1_ASAP7_75t_L g1081 ( 
.A1(n_1034),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_1081)
);

OAI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_973),
.A2(n_45),
.B(n_46),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1041),
.B(n_1003),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_1007),
.A2(n_115),
.B(n_114),
.Y(n_1084)
);

OAI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_976),
.A2(n_47),
.B(n_48),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_992),
.A2(n_118),
.B(n_117),
.Y(n_1086)
);

OAI21x1_ASAP7_75t_L g1087 ( 
.A1(n_997),
.A2(n_1032),
.B(n_1001),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_1025),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1035),
.B(n_47),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_984),
.A2(n_120),
.B(n_119),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_987),
.A2(n_124),
.B(n_123),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_SL g1092 ( 
.A1(n_1023),
.A2(n_48),
.B(n_49),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_1000),
.A2(n_128),
.B(n_127),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_1018),
.B(n_50),
.Y(n_1094)
);

NAND2x1p5_ASAP7_75t_L g1095 ( 
.A(n_1005),
.B(n_130),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_985),
.A2(n_135),
.B(n_133),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_1043),
.A2(n_50),
.B1(n_51),
.B2(n_53),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_993),
.B(n_983),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1010),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_994),
.B(n_51),
.Y(n_1100)
);

NAND2xp33_ASAP7_75t_L g1101 ( 
.A(n_1025),
.B(n_54),
.Y(n_1101)
);

A2O1A1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_1037),
.A2(n_54),
.B(n_56),
.C(n_57),
.Y(n_1102)
);

BUFx8_ASAP7_75t_SL g1103 ( 
.A(n_1016),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1028),
.B(n_56),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_1011),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_1105)
);

AOI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_968),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_1106)
);

HAxp5_ASAP7_75t_L g1107 ( 
.A(n_1031),
.B(n_61),
.CON(n_1107),
.SN(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1002),
.B(n_63),
.Y(n_1108)
);

INVxp67_ASAP7_75t_L g1109 ( 
.A(n_1026),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1038),
.B(n_1040),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_986),
.A2(n_136),
.B(n_138),
.Y(n_1111)
);

OAI22x1_ASAP7_75t_L g1112 ( 
.A1(n_981),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_1112)
);

AOI21x1_ASAP7_75t_L g1113 ( 
.A1(n_999),
.A2(n_142),
.B(n_143),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1083),
.B(n_1038),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_1049),
.Y(n_1115)
);

NAND2x1p5_ASAP7_75t_L g1116 ( 
.A(n_1058),
.B(n_1040),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1099),
.Y(n_1117)
);

BUFx2_ASAP7_75t_L g1118 ( 
.A(n_1076),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1052),
.B(n_1038),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1047),
.Y(n_1120)
);

NAND3xp33_ASAP7_75t_L g1121 ( 
.A(n_1079),
.B(n_1017),
.C(n_975),
.Y(n_1121)
);

BUFx8_ASAP7_75t_L g1122 ( 
.A(n_1053),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_1064),
.B(n_1019),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_1088),
.Y(n_1124)
);

NAND2x1p5_ASAP7_75t_L g1125 ( 
.A(n_1045),
.B(n_1040),
.Y(n_1125)
);

INVx1_ASAP7_75t_SL g1126 ( 
.A(n_1053),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1051),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_1065),
.B(n_1021),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_1094),
.A2(n_989),
.B1(n_996),
.B2(n_1029),
.Y(n_1129)
);

OR2x6_ASAP7_75t_L g1130 ( 
.A(n_1095),
.B(n_378),
.Y(n_1130)
);

HB1xp67_ASAP7_75t_L g1131 ( 
.A(n_1057),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1108),
.A2(n_145),
.B1(n_146),
.B2(n_148),
.Y(n_1132)
);

OA21x2_ASAP7_75t_L g1133 ( 
.A1(n_1062),
.A2(n_1087),
.B(n_1056),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1069),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_1060),
.B(n_370),
.Y(n_1135)
);

INVx3_ASAP7_75t_L g1136 ( 
.A(n_1065),
.Y(n_1136)
);

INVx2_ASAP7_75t_SL g1137 ( 
.A(n_1049),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_SL g1138 ( 
.A1(n_1082),
.A2(n_149),
.B(n_150),
.C(n_151),
.Y(n_1138)
);

OR2x2_ASAP7_75t_L g1139 ( 
.A(n_1059),
.B(n_153),
.Y(n_1139)
);

INVx2_ASAP7_75t_SL g1140 ( 
.A(n_1088),
.Y(n_1140)
);

AND2x2_ASAP7_75t_SL g1141 ( 
.A(n_1101),
.B(n_156),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1104),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1061),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1061),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1061),
.Y(n_1145)
);

INVx1_ASAP7_75t_SL g1146 ( 
.A(n_1103),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1100),
.B(n_369),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1098),
.Y(n_1148)
);

OR2x2_ASAP7_75t_L g1149 ( 
.A(n_1073),
.B(n_158),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1046),
.A2(n_159),
.B(n_161),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1109),
.B(n_368),
.Y(n_1151)
);

BUFx4_ASAP7_75t_SL g1152 ( 
.A(n_1074),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1081),
.B(n_162),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1068),
.B(n_362),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1068),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1089),
.B(n_163),
.Y(n_1156)
);

BUFx2_ASAP7_75t_L g1157 ( 
.A(n_1088),
.Y(n_1157)
);

OAI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1106),
.A2(n_1054),
.B1(n_1071),
.B2(n_1055),
.Y(n_1158)
);

BUFx3_ASAP7_75t_L g1159 ( 
.A(n_1070),
.Y(n_1159)
);

HB1xp67_ASAP7_75t_L g1160 ( 
.A(n_1070),
.Y(n_1160)
);

OR2x2_ASAP7_75t_L g1161 ( 
.A(n_1066),
.B(n_167),
.Y(n_1161)
);

BUFx3_ASAP7_75t_L g1162 ( 
.A(n_1110),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_1065),
.B(n_1050),
.Y(n_1163)
);

BUFx8_ASAP7_75t_SL g1164 ( 
.A(n_1113),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1075),
.Y(n_1165)
);

NAND2x1p5_ASAP7_75t_L g1166 ( 
.A(n_1067),
.B(n_172),
.Y(n_1166)
);

INVx5_ASAP7_75t_L g1167 ( 
.A(n_1107),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_L g1168 ( 
.A1(n_1097),
.A2(n_176),
.B1(n_180),
.B2(n_183),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1085),
.B(n_185),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1078),
.Y(n_1170)
);

A2O1A1Ixp33_ASAP7_75t_SL g1171 ( 
.A1(n_1090),
.A2(n_1096),
.B(n_1044),
.C(n_1111),
.Y(n_1171)
);

OR2x2_ASAP7_75t_L g1172 ( 
.A(n_1105),
.B(n_186),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1063),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_1048),
.B(n_187),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1077),
.A2(n_188),
.B(n_190),
.Y(n_1175)
);

BUFx3_ASAP7_75t_L g1176 ( 
.A(n_1092),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_1112),
.A2(n_191),
.B1(n_192),
.B2(n_194),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1102),
.B(n_1072),
.Y(n_1178)
);

BUFx3_ASAP7_75t_L g1179 ( 
.A(n_1080),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_1086),
.B(n_195),
.Y(n_1180)
);

INVx5_ASAP7_75t_L g1181 ( 
.A(n_1093),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_1084),
.B(n_361),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_1091),
.Y(n_1183)
);

OR2x6_ASAP7_75t_L g1184 ( 
.A(n_1058),
.B(n_197),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_1045),
.B(n_360),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1099),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1046),
.A2(n_198),
.B(n_205),
.Y(n_1187)
);

BUFx3_ASAP7_75t_L g1188 ( 
.A(n_1049),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_1088),
.Y(n_1189)
);

HB1xp67_ASAP7_75t_L g1190 ( 
.A(n_1131),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1173),
.A2(n_207),
.B(n_208),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1123),
.A2(n_1121),
.B(n_1169),
.Y(n_1192)
);

BUFx3_ASAP7_75t_L g1193 ( 
.A(n_1122),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_SL g1194 ( 
.A1(n_1167),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_1194)
);

BUFx3_ASAP7_75t_L g1195 ( 
.A(n_1122),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1117),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1186),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1127),
.A2(n_213),
.B(n_214),
.Y(n_1198)
);

BUFx2_ASAP7_75t_SL g1199 ( 
.A(n_1115),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1134),
.B(n_215),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1120),
.Y(n_1201)
);

INVx2_ASAP7_75t_SL g1202 ( 
.A(n_1124),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1134),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_1160),
.Y(n_1204)
);

OA21x2_ASAP7_75t_L g1205 ( 
.A1(n_1143),
.A2(n_1145),
.B(n_1144),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1148),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_1136),
.Y(n_1207)
);

CKINVDCx11_ASAP7_75t_R g1208 ( 
.A(n_1188),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1142),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1167),
.B(n_217),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1171),
.A2(n_359),
.B(n_222),
.Y(n_1211)
);

HB1xp67_ASAP7_75t_L g1212 ( 
.A(n_1155),
.Y(n_1212)
);

OAI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1167),
.A2(n_219),
.B1(n_224),
.B2(n_230),
.Y(n_1213)
);

INVx3_ASAP7_75t_L g1214 ( 
.A(n_1136),
.Y(n_1214)
);

CKINVDCx11_ASAP7_75t_R g1215 ( 
.A(n_1146),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1143),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_1152),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1144),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1127),
.Y(n_1219)
);

BUFx12f_ASAP7_75t_L g1220 ( 
.A(n_1137),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1170),
.Y(n_1221)
);

OR2x2_ASAP7_75t_L g1222 ( 
.A(n_1126),
.B(n_231),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_1118),
.Y(n_1223)
);

AOI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1163),
.A2(n_233),
.B(n_234),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1170),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1133),
.Y(n_1226)
);

INVx5_ASAP7_75t_L g1227 ( 
.A(n_1164),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1139),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1133),
.A2(n_235),
.B(n_236),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1179),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_1159),
.Y(n_1231)
);

AO21x2_ASAP7_75t_L g1232 ( 
.A1(n_1119),
.A2(n_238),
.B(n_242),
.Y(n_1232)
);

NAND2x1p5_ASAP7_75t_L g1233 ( 
.A(n_1162),
.B(n_247),
.Y(n_1233)
);

CKINVDCx16_ASAP7_75t_R g1234 ( 
.A(n_1184),
.Y(n_1234)
);

AO21x1_ASAP7_75t_L g1235 ( 
.A1(n_1158),
.A2(n_249),
.B(n_252),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1165),
.Y(n_1236)
);

AO21x2_ASAP7_75t_L g1237 ( 
.A1(n_1114),
.A2(n_255),
.B(n_256),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_SL g1238 ( 
.A1(n_1153),
.A2(n_1141),
.B1(n_1172),
.B2(n_1156),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1166),
.A2(n_263),
.B(n_265),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1157),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1184),
.B(n_267),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1124),
.B(n_268),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1124),
.Y(n_1243)
);

AOI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1178),
.A2(n_269),
.B(n_270),
.Y(n_1244)
);

NOR2x1_ASAP7_75t_R g1245 ( 
.A(n_1185),
.B(n_272),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1189),
.B(n_273),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1129),
.A2(n_275),
.B1(n_276),
.B2(n_277),
.Y(n_1247)
);

BUFx2_ASAP7_75t_L g1248 ( 
.A(n_1189),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1181),
.Y(n_1249)
);

HB1xp67_ASAP7_75t_L g1250 ( 
.A(n_1189),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1140),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_SL g1252 ( 
.A1(n_1135),
.A2(n_280),
.B1(n_281),
.B2(n_282),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1128),
.B(n_1185),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1177),
.A2(n_285),
.B1(n_286),
.B2(n_287),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_1128),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1154),
.B(n_290),
.Y(n_1256)
);

AOI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1130),
.A2(n_291),
.B1(n_292),
.B2(n_296),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1149),
.B(n_358),
.Y(n_1258)
);

CKINVDCx11_ASAP7_75t_R g1259 ( 
.A(n_1130),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1181),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1203),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1216),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1216),
.Y(n_1263)
);

BUFx2_ASAP7_75t_SL g1264 ( 
.A(n_1227),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1203),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1218),
.Y(n_1266)
);

INVxp67_ASAP7_75t_L g1267 ( 
.A(n_1240),
.Y(n_1267)
);

OA21x2_ASAP7_75t_L g1268 ( 
.A1(n_1226),
.A2(n_1187),
.B(n_1150),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1219),
.Y(n_1269)
);

INVx3_ASAP7_75t_L g1270 ( 
.A(n_1230),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1219),
.Y(n_1271)
);

OA21x2_ASAP7_75t_L g1272 ( 
.A1(n_1226),
.A2(n_1175),
.B(n_1182),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1229),
.A2(n_1191),
.B(n_1198),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1201),
.B(n_1182),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1221),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1190),
.B(n_1151),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1229),
.A2(n_1132),
.B(n_1168),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1221),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1225),
.Y(n_1279)
);

CKINVDCx11_ASAP7_75t_R g1280 ( 
.A(n_1208),
.Y(n_1280)
);

AO21x2_ASAP7_75t_L g1281 ( 
.A1(n_1236),
.A2(n_1138),
.B(n_1180),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1205),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1205),
.Y(n_1283)
);

INVx3_ASAP7_75t_L g1284 ( 
.A(n_1230),
.Y(n_1284)
);

CKINVDCx6p67_ASAP7_75t_R g1285 ( 
.A(n_1193),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1205),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1236),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1191),
.A2(n_1147),
.B(n_1181),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1249),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1249),
.Y(n_1290)
);

INVx3_ASAP7_75t_L g1291 ( 
.A(n_1260),
.Y(n_1291)
);

HB1xp67_ASAP7_75t_L g1292 ( 
.A(n_1204),
.Y(n_1292)
);

HB1xp67_ASAP7_75t_L g1293 ( 
.A(n_1212),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1200),
.B(n_1176),
.Y(n_1294)
);

AOI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1235),
.A2(n_1174),
.B(n_1180),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1260),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1200),
.B(n_1174),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1196),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1197),
.B(n_1161),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1209),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1206),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1232),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1228),
.B(n_1116),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1232),
.Y(n_1304)
);

OR2x6_ASAP7_75t_L g1305 ( 
.A(n_1233),
.B(n_1183),
.Y(n_1305)
);

AO21x2_ASAP7_75t_L g1306 ( 
.A1(n_1192),
.A2(n_1183),
.B(n_1125),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1232),
.Y(n_1307)
);

OR2x6_ASAP7_75t_L g1308 ( 
.A(n_1233),
.B(n_1183),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_SL g1309 ( 
.A1(n_1227),
.A2(n_1234),
.B1(n_1241),
.B2(n_1238),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1253),
.B(n_297),
.Y(n_1310)
);

INVx3_ASAP7_75t_L g1311 ( 
.A(n_1207),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1237),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1237),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1253),
.B(n_299),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1207),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1237),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1250),
.B(n_300),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1210),
.A2(n_306),
.B(n_309),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1198),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1207),
.B(n_310),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1214),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1223),
.B(n_313),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1214),
.Y(n_1323)
);

CKINVDCx11_ASAP7_75t_R g1324 ( 
.A(n_1208),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1214),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1244),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1243),
.B(n_317),
.Y(n_1327)
);

AO21x2_ASAP7_75t_L g1328 ( 
.A1(n_1235),
.A2(n_319),
.B(n_322),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1224),
.Y(n_1329)
);

INVx2_ASAP7_75t_SL g1330 ( 
.A(n_1227),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1239),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1248),
.B(n_324),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1291),
.B(n_1227),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_L g1334 ( 
.A(n_1285),
.B(n_1215),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1300),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1300),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1292),
.B(n_1227),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1278),
.Y(n_1338)
);

OR2x2_ASAP7_75t_L g1339 ( 
.A(n_1293),
.B(n_1269),
.Y(n_1339)
);

HB1xp67_ASAP7_75t_L g1340 ( 
.A(n_1267),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1311),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_1285),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1301),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_1330),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1301),
.Y(n_1345)
);

INVxp67_ASAP7_75t_SL g1346 ( 
.A(n_1276),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1274),
.B(n_1315),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1298),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1274),
.B(n_1251),
.Y(n_1349)
);

NAND2x1_ASAP7_75t_L g1350 ( 
.A(n_1315),
.B(n_1202),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1298),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1321),
.B(n_1255),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1261),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1291),
.B(n_1255),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1321),
.B(n_1255),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1261),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1309),
.A2(n_1259),
.B1(n_1256),
.B2(n_1254),
.Y(n_1357)
);

AND2x4_ASAP7_75t_L g1358 ( 
.A(n_1291),
.B(n_1255),
.Y(n_1358)
);

INVx3_ASAP7_75t_L g1359 ( 
.A(n_1311),
.Y(n_1359)
);

NAND3xp33_ASAP7_75t_L g1360 ( 
.A(n_1323),
.B(n_1257),
.C(n_1252),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1280),
.B(n_1215),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1323),
.B(n_1202),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1265),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1269),
.B(n_1193),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1279),
.Y(n_1365)
);

AND2x4_ASAP7_75t_L g1366 ( 
.A(n_1330),
.B(n_1195),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_1324),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1265),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_L g1369 ( 
.A(n_1322),
.B(n_1231),
.Y(n_1369)
);

OR2x2_ASAP7_75t_L g1370 ( 
.A(n_1271),
.B(n_1195),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1271),
.B(n_1275),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1325),
.B(n_1246),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_L g1373 ( 
.A(n_1322),
.B(n_1231),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1299),
.B(n_1294),
.Y(n_1374)
);

OR2x2_ASAP7_75t_L g1375 ( 
.A(n_1275),
.B(n_1199),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1325),
.B(n_1242),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1299),
.B(n_1259),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1294),
.B(n_1210),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1289),
.B(n_1242),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1289),
.B(n_1246),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1262),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1262),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1263),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1303),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1290),
.B(n_1256),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1263),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1266),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1266),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1346),
.B(n_1311),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1347),
.B(n_1297),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1340),
.B(n_1306),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1339),
.Y(n_1392)
);

NAND3xp33_ASAP7_75t_L g1393 ( 
.A(n_1375),
.B(n_1360),
.C(n_1339),
.Y(n_1393)
);

NAND3xp33_ASAP7_75t_L g1394 ( 
.A(n_1375),
.B(n_1296),
.C(n_1290),
.Y(n_1394)
);

NAND3xp33_ASAP7_75t_L g1395 ( 
.A(n_1378),
.B(n_1296),
.C(n_1303),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1349),
.B(n_1306),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_R g1397 ( 
.A(n_1367),
.B(n_1295),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1349),
.B(n_1306),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1374),
.B(n_1297),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1347),
.B(n_1384),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1352),
.B(n_1270),
.Y(n_1401)
);

NAND4xp25_ASAP7_75t_L g1402 ( 
.A(n_1369),
.B(n_1319),
.C(n_1326),
.D(n_1318),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1352),
.B(n_1270),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1355),
.B(n_1270),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1384),
.B(n_1264),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1385),
.B(n_1284),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1385),
.B(n_1335),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1344),
.B(n_1264),
.Y(n_1408)
);

AOI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1357),
.A2(n_1328),
.B1(n_1308),
.B2(n_1305),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1355),
.B(n_1284),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1377),
.B(n_1284),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1373),
.A2(n_1328),
.B1(n_1258),
.B2(n_1312),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1336),
.B(n_1326),
.Y(n_1413)
);

AOI221xp5_ASAP7_75t_L g1414 ( 
.A1(n_1343),
.A2(n_1312),
.B1(n_1328),
.B2(n_1213),
.C(n_1247),
.Y(n_1414)
);

OAI21xp5_ASAP7_75t_SL g1415 ( 
.A1(n_1361),
.A2(n_1295),
.B(n_1194),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1345),
.B(n_1272),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1337),
.A2(n_1314),
.B1(n_1310),
.B2(n_1308),
.Y(n_1417)
);

OAI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1364),
.A2(n_1305),
.B1(n_1308),
.B2(n_1272),
.Y(n_1418)
);

OAI221xp5_ASAP7_75t_L g1419 ( 
.A1(n_1364),
.A2(n_1317),
.B1(n_1332),
.B2(n_1329),
.C(n_1222),
.Y(n_1419)
);

NAND2x1_ASAP7_75t_L g1420 ( 
.A(n_1333),
.B(n_1305),
.Y(n_1420)
);

NAND2xp33_ASAP7_75t_L g1421 ( 
.A(n_1367),
.B(n_1217),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1372),
.B(n_1376),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1370),
.B(n_1272),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1338),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1413),
.Y(n_1425)
);

OAI21xp33_ASAP7_75t_L g1426 ( 
.A1(n_1402),
.A2(n_1362),
.B(n_1372),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1392),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1400),
.B(n_1341),
.Y(n_1428)
);

AND4x1_ASAP7_75t_L g1429 ( 
.A(n_1393),
.B(n_1334),
.C(n_1217),
.D(n_1220),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1391),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1416),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1389),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_1406),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1424),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1422),
.B(n_1341),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1407),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1390),
.B(n_1341),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1396),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1424),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1411),
.B(n_1359),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1398),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1401),
.B(n_1359),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1401),
.B(n_1359),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1403),
.Y(n_1444)
);

INVx1_ASAP7_75t_SL g1445 ( 
.A(n_1421),
.Y(n_1445)
);

INVx1_ASAP7_75t_SL g1446 ( 
.A(n_1421),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1423),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1399),
.B(n_1403),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1404),
.B(n_1376),
.Y(n_1449)
);

AND2x4_ASAP7_75t_L g1450 ( 
.A(n_1449),
.B(n_1366),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1425),
.B(n_1412),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1432),
.B(n_1370),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1427),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1427),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1449),
.B(n_1404),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1435),
.B(n_1437),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1425),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1436),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1431),
.B(n_1412),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1436),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1434),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1434),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1433),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_SL g1464 ( 
.A(n_1445),
.B(n_1397),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1431),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1463),
.B(n_1448),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1458),
.B(n_1426),
.Y(n_1467)
);

NAND2xp33_ASAP7_75t_SL g1468 ( 
.A(n_1450),
.B(n_1397),
.Y(n_1468)
);

AOI211xp5_ASAP7_75t_L g1469 ( 
.A1(n_1464),
.A2(n_1415),
.B(n_1419),
.C(n_1446),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1451),
.B(n_1447),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1453),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1450),
.B(n_1440),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1454),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1460),
.B(n_1447),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1457),
.Y(n_1475)
);

NAND2x1_ASAP7_75t_L g1476 ( 
.A(n_1456),
.B(n_1437),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1459),
.B(n_1438),
.Y(n_1477)
);

OAI21xp33_ASAP7_75t_L g1478 ( 
.A1(n_1459),
.A2(n_1429),
.B(n_1409),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1451),
.B(n_1438),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1465),
.B(n_1444),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1452),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1461),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1455),
.B(n_1441),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1456),
.B(n_1440),
.Y(n_1484)
);

NAND2x1_ASAP7_75t_SL g1485 ( 
.A(n_1481),
.B(n_1430),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1475),
.B(n_1462),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1471),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1484),
.B(n_1435),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1466),
.B(n_1428),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1473),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1469),
.A2(n_1342),
.B1(n_1414),
.B2(n_1395),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1478),
.B(n_1220),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1472),
.B(n_1428),
.Y(n_1493)
);

NOR2xp67_ASAP7_75t_L g1494 ( 
.A(n_1483),
.B(n_1394),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1482),
.Y(n_1495)
);

NAND2x1_ASAP7_75t_SL g1496 ( 
.A(n_1494),
.B(n_1469),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_L g1497 ( 
.A(n_1492),
.B(n_1478),
.Y(n_1497)
);

AOI32xp33_ASAP7_75t_L g1498 ( 
.A1(n_1491),
.A2(n_1468),
.A3(n_1467),
.B1(n_1477),
.B2(n_1479),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1485),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1487),
.Y(n_1500)
);

INVx3_ASAP7_75t_L g1501 ( 
.A(n_1489),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1490),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1495),
.Y(n_1503)
);

AOI21xp33_ASAP7_75t_L g1504 ( 
.A1(n_1491),
.A2(n_1486),
.B(n_1470),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1486),
.Y(n_1505)
);

NAND3xp33_ASAP7_75t_SL g1506 ( 
.A(n_1498),
.B(n_1476),
.C(n_1493),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1502),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1501),
.B(n_1488),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_SL g1509 ( 
.A(n_1499),
.B(n_1474),
.Y(n_1509)
);

BUFx2_ASAP7_75t_L g1510 ( 
.A(n_1501),
.Y(n_1510)
);

INVx1_ASAP7_75t_SL g1511 ( 
.A(n_1496),
.Y(n_1511)
);

NAND2xp33_ASAP7_75t_R g1512 ( 
.A(n_1497),
.B(n_1366),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1510),
.B(n_1503),
.Y(n_1513)
);

INVxp67_ASAP7_75t_L g1514 ( 
.A(n_1511),
.Y(n_1514)
);

NAND4xp25_ASAP7_75t_L g1515 ( 
.A(n_1506),
.B(n_1505),
.C(n_1500),
.D(n_1504),
.Y(n_1515)
);

AOI322xp5_ASAP7_75t_L g1516 ( 
.A1(n_1509),
.A2(n_1504),
.A3(n_1480),
.B1(n_1418),
.B2(n_1329),
.C1(n_1313),
.C2(n_1316),
.Y(n_1516)
);

NAND4xp25_ASAP7_75t_L g1517 ( 
.A(n_1507),
.B(n_1366),
.C(n_1408),
.D(n_1443),
.Y(n_1517)
);

NOR4xp25_ASAP7_75t_L g1518 ( 
.A(n_1508),
.B(n_1320),
.C(n_1327),
.D(n_1417),
.Y(n_1518)
);

OAI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1512),
.A2(n_1277),
.B(n_1320),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1512),
.A2(n_1418),
.B1(n_1313),
.B2(n_1316),
.Y(n_1520)
);

AOI321xp33_ASAP7_75t_L g1521 ( 
.A1(n_1509),
.A2(n_1380),
.A3(n_1379),
.B1(n_1327),
.B2(n_1245),
.C(n_1302),
.Y(n_1521)
);

NOR3xp33_ASAP7_75t_L g1522 ( 
.A(n_1514),
.B(n_1222),
.C(n_1239),
.Y(n_1522)
);

AOI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1515),
.A2(n_1350),
.B(n_1211),
.Y(n_1523)
);

NAND4xp75_ASAP7_75t_L g1524 ( 
.A(n_1513),
.B(n_1405),
.C(n_1379),
.D(n_1380),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_L g1525 ( 
.A(n_1517),
.B(n_1442),
.Y(n_1525)
);

OAI211xp5_ASAP7_75t_L g1526 ( 
.A1(n_1518),
.A2(n_1443),
.B(n_1442),
.C(n_1362),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1519),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1520),
.Y(n_1528)
);

AND3x4_ASAP7_75t_L g1529 ( 
.A(n_1521),
.B(n_1333),
.C(n_1358),
.Y(n_1529)
);

NOR3xp33_ASAP7_75t_L g1530 ( 
.A(n_1516),
.B(n_1420),
.C(n_1331),
.Y(n_1530)
);

AOI211xp5_ASAP7_75t_L g1531 ( 
.A1(n_1523),
.A2(n_1277),
.B(n_1333),
.C(n_1319),
.Y(n_1531)
);

NAND4xp25_ASAP7_75t_L g1532 ( 
.A(n_1525),
.B(n_1410),
.C(n_1331),
.D(n_1354),
.Y(n_1532)
);

NOR3xp33_ASAP7_75t_L g1533 ( 
.A(n_1527),
.B(n_1288),
.C(n_1439),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1522),
.B(n_1439),
.Y(n_1534)
);

NAND4xp25_ASAP7_75t_SL g1535 ( 
.A(n_1526),
.B(n_1353),
.C(n_1356),
.D(n_1363),
.Y(n_1535)
);

NAND3xp33_ASAP7_75t_SL g1536 ( 
.A(n_1529),
.B(n_1368),
.C(n_1302),
.Y(n_1536)
);

NOR3xp33_ASAP7_75t_L g1537 ( 
.A(n_1528),
.B(n_1288),
.C(n_1273),
.Y(n_1537)
);

OAI21xp5_ASAP7_75t_SL g1538 ( 
.A1(n_1530),
.A2(n_1358),
.B(n_1354),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1531),
.B(n_1524),
.Y(n_1539)
);

INVxp67_ASAP7_75t_L g1540 ( 
.A(n_1534),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1537),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1535),
.Y(n_1542)
);

AOI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1536),
.A2(n_1281),
.B1(n_1305),
.B2(n_1308),
.Y(n_1543)
);

INVxp67_ASAP7_75t_SL g1544 ( 
.A(n_1533),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1532),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1538),
.Y(n_1546)
);

AOI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1537),
.A2(n_1281),
.B1(n_1304),
.B2(n_1307),
.Y(n_1547)
);

NOR2x1_ASAP7_75t_L g1548 ( 
.A(n_1535),
.B(n_1281),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1544),
.Y(n_1549)
);

NOR3xp33_ASAP7_75t_L g1550 ( 
.A(n_1540),
.B(n_1541),
.C(n_1546),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1542),
.Y(n_1551)
);

INVx4_ASAP7_75t_L g1552 ( 
.A(n_1545),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1548),
.Y(n_1553)
);

NAND2xp33_ASAP7_75t_SL g1554 ( 
.A(n_1539),
.B(n_1354),
.Y(n_1554)
);

NOR4xp25_ASAP7_75t_L g1555 ( 
.A(n_1547),
.B(n_1348),
.C(n_1351),
.D(n_1371),
.Y(n_1555)
);

OAI22xp5_ASAP7_75t_SL g1556 ( 
.A1(n_1543),
.A2(n_1272),
.B1(n_1358),
.B2(n_1268),
.Y(n_1556)
);

NOR3xp33_ASAP7_75t_L g1557 ( 
.A(n_1540),
.B(n_1273),
.C(n_1304),
.Y(n_1557)
);

NOR4xp25_ASAP7_75t_L g1558 ( 
.A(n_1540),
.B(n_1371),
.C(n_1282),
.D(n_1307),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1539),
.B(n_1282),
.Y(n_1559)
);

NOR4xp75_ASAP7_75t_L g1560 ( 
.A(n_1539),
.B(n_329),
.C(n_331),
.D(n_332),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1546),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1542),
.B(n_1383),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1561),
.B(n_1387),
.Y(n_1563)
);

NOR2x1_ASAP7_75t_L g1564 ( 
.A(n_1552),
.B(n_333),
.Y(n_1564)
);

INVxp67_ASAP7_75t_L g1565 ( 
.A(n_1549),
.Y(n_1565)
);

NAND3xp33_ASAP7_75t_SL g1566 ( 
.A(n_1550),
.B(n_1283),
.C(n_1286),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1562),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1553),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1551),
.B(n_1268),
.Y(n_1569)
);

XOR2x2_ASAP7_75t_L g1570 ( 
.A(n_1560),
.B(n_334),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1564),
.B(n_1559),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1563),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1565),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1568),
.A2(n_1556),
.B1(n_1557),
.B2(n_1554),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1567),
.B(n_1555),
.Y(n_1575)
);

OAI211xp5_ASAP7_75t_SL g1576 ( 
.A1(n_1573),
.A2(n_1575),
.B(n_1571),
.C(n_1572),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1574),
.B(n_1570),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1572),
.B(n_1569),
.Y(n_1578)
);

OAI322xp33_ASAP7_75t_L g1579 ( 
.A1(n_1573),
.A2(n_1566),
.A3(n_1558),
.B1(n_1283),
.B2(n_1286),
.C1(n_1287),
.C2(n_1381),
.Y(n_1579)
);

NOR2x1_ASAP7_75t_L g1580 ( 
.A(n_1576),
.B(n_335),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1578),
.Y(n_1581)
);

OAI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1577),
.A2(n_1268),
.B(n_1388),
.Y(n_1582)
);

AOI21xp5_ASAP7_75t_L g1583 ( 
.A1(n_1581),
.A2(n_1579),
.B(n_1268),
.Y(n_1583)
);

AOI21xp33_ASAP7_75t_L g1584 ( 
.A1(n_1580),
.A2(n_337),
.B(n_338),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1582),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1584),
.A2(n_341),
.B(n_342),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1585),
.B(n_343),
.Y(n_1587)
);

OAI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1586),
.A2(n_1583),
.B(n_1287),
.Y(n_1588)
);

OAI222xp33_ASAP7_75t_L g1589 ( 
.A1(n_1587),
.A2(n_1388),
.B1(n_1386),
.B2(n_1382),
.C1(n_1381),
.C2(n_1365),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1588),
.A2(n_1386),
.B1(n_1382),
.B2(n_1365),
.Y(n_1590)
);

OAI221xp5_ASAP7_75t_R g1591 ( 
.A1(n_1590),
.A2(n_1589),
.B1(n_347),
.B2(n_348),
.C(n_349),
.Y(n_1591)
);

AOI211xp5_ASAP7_75t_L g1592 ( 
.A1(n_1591),
.A2(n_346),
.B(n_351),
.C(n_352),
.Y(n_1592)
);


endmodule