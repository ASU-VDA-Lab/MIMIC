module real_jpeg_1102_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_1),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_61)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_64),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_1),
.A2(n_35),
.B1(n_36),
.B2(n_64),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_1),
.A2(n_51),
.B1(n_53),
.B2(n_64),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_2),
.A2(n_62),
.B1(n_63),
.B2(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_2),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_162),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_2),
.A2(n_35),
.B1(n_36),
.B2(n_162),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_2),
.A2(n_51),
.B1(n_53),
.B2(n_162),
.Y(n_273)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_3),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_4),
.A2(n_62),
.B1(n_63),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_4),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_100),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_4),
.A2(n_35),
.B1(n_36),
.B2(n_100),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_4),
.A2(n_51),
.B1(n_53),
.B2(n_100),
.Y(n_217)
);

O2A1O1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_5),
.A2(n_29),
.B(n_33),
.C(n_34),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_5),
.B(n_29),
.Y(n_33)
);

AO22x2_ASAP7_75t_L g34 ( 
.A1(n_5),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_34)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_5),
.A2(n_11),
.B(n_29),
.C(n_212),
.Y(n_211)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_9),
.A2(n_35),
.B1(n_36),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_9),
.A2(n_51),
.B1(n_53),
.B2(n_57),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_57),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_9),
.A2(n_57),
.B1(n_62),
.B2(n_63),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_10),
.A2(n_62),
.B1(n_63),
.B2(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_10),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_122),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_122),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_10),
.A2(n_51),
.B1(n_53),
.B2(n_122),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_11),
.B(n_62),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_11),
.B(n_163),
.Y(n_200)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_11),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_11),
.B(n_34),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_213),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_11),
.B(n_48),
.C(n_51),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_11),
.A2(n_35),
.B1(n_36),
.B2(n_213),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_11),
.B(n_90),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_11),
.B(n_79),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_12),
.A2(n_35),
.B1(n_36),
.B2(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_55),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_12),
.A2(n_51),
.B1(n_53),
.B2(n_55),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_12),
.A2(n_55),
.B1(n_62),
.B2(n_63),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_13),
.A2(n_35),
.B1(n_36),
.B2(n_43),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_13),
.A2(n_43),
.B1(n_62),
.B2(n_63),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_13),
.A2(n_43),
.B1(n_51),
.B2(n_53),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_14),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_15),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_15),
.A2(n_40),
.B1(n_62),
.B2(n_63),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_15),
.A2(n_35),
.B1(n_36),
.B2(n_40),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_15),
.A2(n_40),
.B1(n_51),
.B2(n_53),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_326),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_313),
.B(n_325),
.Y(n_19)
);

AO21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_138),
.B(n_310),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_125),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_101),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_23),
.B(n_101),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_82),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_58),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_25),
.A2(n_26),
.B(n_44),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_25),
.B(n_58),
.C(n_82),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_44),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_27),
.A2(n_41),
.B1(n_42),
.B2(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_27),
.A2(n_39),
.B1(n_41),
.B2(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_27),
.A2(n_41),
.B1(n_76),
.B2(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_27),
.A2(n_179),
.B(n_181),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_27),
.A2(n_181),
.B(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_28),
.B(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_28),
.A2(n_34),
.B1(n_180),
.B2(n_197),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_28),
.A2(n_34),
.B(n_317),
.Y(n_316)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_29),
.A2(n_30),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

AOI32xp33_ASAP7_75t_L g183 ( 
.A1(n_29),
.A2(n_63),
.A3(n_68),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp33_ASAP7_75t_SL g185 ( 
.A(n_30),
.B(n_69),
.Y(n_185)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_34),
.B(n_159),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_36),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

OAI21xp33_ASAP7_75t_L g212 ( 
.A1(n_35),
.A2(n_38),
.B(n_213),
.Y(n_212)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_36),
.B(n_258),
.Y(n_257)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_41),
.A2(n_118),
.B(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_41),
.A2(n_158),
.B(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_50),
.B1(n_54),
.B2(n_56),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_45),
.A2(n_50),
.B1(n_54),
.B2(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_45),
.A2(n_50),
.B1(n_206),
.B2(n_240),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_45),
.A2(n_208),
.B(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_79),
.B(n_80),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_46),
.A2(n_79),
.B1(n_95),
.B2(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_46),
.A2(n_79),
.B1(n_116),
.B2(n_153),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_46),
.A2(n_205),
.B(n_207),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_46),
.B(n_209),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_48),
.A2(n_49),
.B1(n_51),
.B2(n_53),
.Y(n_50)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_50),
.A2(n_228),
.B(n_229),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_50),
.A2(n_229),
.B(n_240),
.Y(n_239)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_51),
.B(n_269),
.Y(n_268)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_73),
.B2(n_81),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_59),
.A2(n_60),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_SL g136 ( 
.A(n_60),
.B(n_74),
.C(n_78),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_60),
.B(n_129),
.C(n_136),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_65),
.B1(n_67),
.B2(n_72),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_61),
.A2(n_67),
.B(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_62),
.A2(n_63),
.B1(n_68),
.B2(n_69),
.Y(n_71)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

O2A1O1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_63),
.A2(n_65),
.B(n_213),
.C(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_65),
.A2(n_120),
.B(n_123),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_65),
.A2(n_67),
.B1(n_72),
.B2(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_66),
.A2(n_121),
.B1(n_161),
.B2(n_163),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_66),
.A2(n_163),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_66),
.A2(n_163),
.B1(n_320),
.B2(n_329),
.Y(n_328)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_71),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_67),
.B(n_99),
.Y(n_124)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_67),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_67),
.A2(n_97),
.B(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_77),
.B2(n_78),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_77),
.A2(n_78),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_78),
.B(n_130),
.C(n_134),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_79),
.B(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_86),
.B(n_96),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_83),
.A2(n_84),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_93),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_86),
.B1(n_96),
.B2(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_85),
.A2(n_86),
.B1(n_93),
.B2(n_148),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_90),
.B(n_91),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_87),
.A2(n_90),
.B1(n_113),
.B2(n_155),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_87),
.A2(n_213),
.B(n_246),
.Y(n_270)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_88),
.A2(n_89),
.B1(n_92),
.B2(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_88),
.A2(n_89),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_88),
.A2(n_89),
.B1(n_188),
.B2(n_203),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_88),
.B(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_88),
.A2(n_244),
.B(n_245),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_88),
.A2(n_89),
.B1(n_244),
.B2(n_278),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_89),
.A2(n_203),
.B(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_89),
.B(n_217),
.Y(n_246)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_90),
.A2(n_216),
.B(n_273),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_93),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_107),
.C(n_108),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_102),
.A2(n_103),
.B1(n_107),
.B2(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_141),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_117),
.C(n_119),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_109),
.A2(n_110),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_114),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_111),
.A2(n_114),
.B1(n_115),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_111),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_117),
.B(n_119),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_124),
.B(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_125),
.A2(n_311),
.B(n_312),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_137),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_126),
.B(n_137),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_136),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_131),
.Y(n_319)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_135),
.Y(n_317)
);

AO21x1_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_164),
.B(n_309),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_143),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_140),
.B(n_143),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.C(n_149),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_147),
.Y(n_167)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_167),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_156),
.C(n_160),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_150),
.A2(n_151),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_152),
.B(n_154),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_153),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_155),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_156),
.A2(n_157),
.B1(n_160),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_161),
.Y(n_177)
);

OAI21x1_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_190),
.B(n_308),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_166),
.B(n_168),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_173),
.C(n_175),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_169),
.B(n_173),
.Y(n_293)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_170),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_175),
.B(n_293),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.C(n_182),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_176),
.B(n_178),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_182),
.B(n_296),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_183),
.A2(n_186),
.B1(n_187),
.B2(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_183),
.Y(n_232)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_184),
.Y(n_222)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

AOI31xp33_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_290),
.A3(n_300),
.B(n_305),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_234),
.B(n_289),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_218),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_193),
.B(n_218),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_204),
.C(n_210),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_194),
.B(n_286),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_198),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_195),
.B(n_199),
.C(n_202),
.Y(n_233)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_204),
.B(n_210),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_211),
.B(n_214),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_230),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_219),
.B(n_231),
.C(n_233),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_223),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_220),
.B(n_225),
.C(n_226),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_284),
.B(n_288),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_253),
.B(n_283),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_247),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_237),
.B(n_247),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_241),
.C(n_242),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_238),
.A2(n_239),
.B1(n_241),
.B2(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_241),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_242),
.A2(n_243),
.B1(n_262),
.B2(n_264),
.Y(n_261)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_252),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_249),
.B(n_251),
.C(n_252),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_265),
.B(n_282),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_261),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_261),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_259),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_256),
.A2(n_257),
.B1(n_259),
.B2(n_280),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_259),
.Y(n_280)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_262),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_276),
.B(n_281),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_271),
.B(n_275),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_270),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_272),
.B(n_274),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_273),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_279),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_279),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_287),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_285),
.B(n_287),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

OAI21xp33_ASAP7_75t_L g305 ( 
.A1(n_291),
.A2(n_306),
.B(n_307),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_294),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_294),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_297),
.C(n_298),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_302),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_297),
.A2(n_298),
.B1(n_299),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_297),
.Y(n_303)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_304),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_304),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_324),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_324),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_323),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_318),
.B1(n_321),
.B2(n_322),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_316),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_318),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_321),
.C(n_323),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_331),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_330),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_328),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_330),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);


endmodule