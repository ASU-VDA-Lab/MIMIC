module fake_netlist_1_12390_n_732 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_93, n_51, n_39, n_732);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_93;
input n_51;
input n_39;
output n_732;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_659;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_666;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
NAND2xp5_ASAP7_75t_L g95 ( .A(n_89), .B(n_42), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_92), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_58), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_83), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_2), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_19), .Y(n_100) );
INVxp67_ASAP7_75t_SL g101 ( .A(n_27), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_76), .Y(n_102) );
BUFx3_ASAP7_75t_L g103 ( .A(n_88), .Y(n_103) );
BUFx3_ASAP7_75t_L g104 ( .A(n_61), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_47), .Y(n_105) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_74), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_62), .Y(n_107) );
INVx3_ASAP7_75t_L g108 ( .A(n_44), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_30), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_73), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_78), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_29), .Y(n_112) );
BUFx10_ASAP7_75t_L g113 ( .A(n_4), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_28), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_3), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_41), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_80), .Y(n_117) );
BUFx3_ASAP7_75t_L g118 ( .A(n_6), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_71), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_67), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_34), .Y(n_121) );
OR2x2_ASAP7_75t_L g122 ( .A(n_0), .B(n_81), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_15), .Y(n_123) );
BUFx2_ASAP7_75t_L g124 ( .A(n_37), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_69), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_11), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_46), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_4), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_0), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_54), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_26), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_25), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_39), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_3), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_96), .Y(n_135) );
OA21x2_ASAP7_75t_L g136 ( .A1(n_96), .A2(n_45), .B(n_93), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_124), .B(n_1), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_97), .Y(n_138) );
AND2x6_ASAP7_75t_L g139 ( .A(n_108), .B(n_22), .Y(n_139) );
AND2x2_ASAP7_75t_SL g140 ( .A(n_124), .B(n_94), .Y(n_140) );
AND2x2_ASAP7_75t_L g141 ( .A(n_113), .B(n_1), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g142 ( .A(n_128), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_100), .B(n_2), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_108), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_100), .B(n_5), .Y(n_145) );
INVx6_ASAP7_75t_L g146 ( .A(n_103), .Y(n_146) );
CKINVDCx8_ASAP7_75t_R g147 ( .A(n_109), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_106), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_108), .Y(n_149) );
OAI22xp5_ASAP7_75t_SL g150 ( .A1(n_123), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_97), .Y(n_151) );
AND2x2_ASAP7_75t_L g152 ( .A(n_113), .B(n_7), .Y(n_152) );
OA21x2_ASAP7_75t_L g153 ( .A1(n_98), .A2(n_49), .B(n_90), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_123), .B(n_8), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_137), .B(n_111), .Y(n_155) );
INVx2_ASAP7_75t_SL g156 ( .A(n_137), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_144), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_144), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_148), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_144), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_149), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_137), .B(n_112), .Y(n_162) );
NAND2xp33_ASAP7_75t_L g163 ( .A(n_139), .B(n_133), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_149), .Y(n_164) );
AND2x6_ASAP7_75t_L g165 ( .A(n_137), .B(n_98), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_141), .B(n_113), .Y(n_166) );
INVx2_ASAP7_75t_SL g167 ( .A(n_137), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_149), .Y(n_168) );
INVx4_ASAP7_75t_L g169 ( .A(n_139), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_135), .B(n_125), .Y(n_170) );
INVxp33_ASAP7_75t_L g171 ( .A(n_141), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_135), .B(n_103), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_138), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_148), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_138), .B(n_99), .Y(n_175) );
OAI22xp33_ASAP7_75t_L g176 ( .A1(n_143), .A2(n_134), .B1(n_115), .B2(n_126), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_151), .B(n_113), .Y(n_177) );
INVx3_ASAP7_75t_L g178 ( .A(n_139), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_141), .B(n_118), .Y(n_179) );
NAND2xp33_ASAP7_75t_L g180 ( .A(n_139), .B(n_122), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_148), .Y(n_181) );
OR2x2_ASAP7_75t_L g182 ( .A(n_152), .B(n_118), .Y(n_182) );
OR2x6_ASAP7_75t_L g183 ( .A(n_152), .B(n_122), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_151), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_166), .B(n_152), .Y(n_185) );
INVxp67_ASAP7_75t_SL g186 ( .A(n_182), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_157), .Y(n_187) );
AOI22xp33_ASAP7_75t_L g188 ( .A1(n_165), .A2(n_140), .B1(n_139), .B2(n_154), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_169), .B(n_147), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_157), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_158), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_166), .B(n_140), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_158), .Y(n_193) );
BUFx3_ASAP7_75t_L g194 ( .A(n_169), .Y(n_194) );
INVx8_ASAP7_75t_L g195 ( .A(n_165), .Y(n_195) );
AOI22xp5_ASAP7_75t_L g196 ( .A1(n_165), .A2(n_140), .B1(n_150), .B2(n_139), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_169), .B(n_147), .Y(n_197) );
NAND2xp33_ASAP7_75t_L g198 ( .A(n_165), .B(n_139), .Y(n_198) );
NOR2xp33_ASAP7_75t_SL g199 ( .A(n_169), .B(n_139), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_179), .B(n_147), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_160), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_176), .B(n_143), .Y(n_202) );
OAI21xp5_ASAP7_75t_L g203 ( .A1(n_178), .A2(n_153), .B(n_136), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_183), .Y(n_204) );
INVxp67_ASAP7_75t_L g205 ( .A(n_182), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_160), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_163), .A2(n_153), .B(n_136), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_161), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_161), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_156), .B(n_145), .Y(n_210) );
AND2x6_ASAP7_75t_SL g211 ( .A(n_183), .B(n_145), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_179), .B(n_154), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g213 ( .A1(n_165), .A2(n_150), .B1(n_139), .B2(n_134), .Y(n_213) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_165), .A2(n_146), .B1(n_129), .B2(n_102), .Y(n_214) );
INVx2_ASAP7_75t_SL g215 ( .A(n_165), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_177), .B(n_146), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_164), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_164), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_156), .B(n_129), .Y(n_219) );
HB1xp67_ASAP7_75t_L g220 ( .A(n_183), .Y(n_220) );
INVx2_ASAP7_75t_SL g221 ( .A(n_165), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_167), .B(n_129), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_167), .B(n_129), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_173), .B(n_101), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_186), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_185), .B(n_171), .Y(n_226) );
OAI21xp5_ASAP7_75t_L g227 ( .A1(n_207), .A2(n_178), .B(n_180), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_199), .A2(n_178), .B(n_155), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_212), .B(n_183), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_187), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_205), .B(n_183), .Y(n_231) );
BUFx3_ASAP7_75t_L g232 ( .A(n_195), .Y(n_232) );
NOR2xp67_ASAP7_75t_SL g233 ( .A(n_194), .B(n_178), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_192), .B(n_175), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_187), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_199), .A2(n_162), .B(n_184), .Y(n_236) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_220), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_196), .A2(n_213), .B(n_188), .C(n_191), .Y(n_238) );
O2A1O1Ixp5_ASAP7_75t_L g239 ( .A1(n_202), .A2(n_172), .B(n_170), .C(n_173), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_198), .A2(n_184), .B(n_170), .Y(n_240) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_195), .Y(n_241) );
OAI22xp5_ASAP7_75t_L g242 ( .A1(n_196), .A2(n_107), .B1(n_168), .B2(n_142), .Y(n_242) );
O2A1O1Ixp5_ASAP7_75t_L g243 ( .A1(n_203), .A2(n_168), .B(n_125), .C(n_131), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_204), .B(n_146), .Y(n_244) );
OAI22xp5_ASAP7_75t_L g245 ( .A1(n_195), .A2(n_146), .B1(n_102), .B2(n_114), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_203), .A2(n_210), .B(n_216), .Y(n_246) );
OR2x6_ASAP7_75t_L g247 ( .A(n_195), .B(n_129), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_211), .Y(n_248) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_195), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_200), .B(n_146), .Y(n_250) );
NOR2xp67_ASAP7_75t_L g251 ( .A(n_213), .B(n_8), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_187), .B(n_105), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_190), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_211), .B(n_105), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_194), .B(n_95), .Y(n_255) );
INVx3_ASAP7_75t_SL g256 ( .A(n_190), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_224), .Y(n_257) );
AOI21xp5_ASAP7_75t_SL g258 ( .A1(n_247), .A2(n_215), .B(n_221), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_246), .A2(n_189), .B(n_197), .Y(n_259) );
AOI221xp5_ASAP7_75t_L g260 ( .A1(n_226), .A2(n_224), .B1(n_191), .B2(n_206), .C(n_218), .Y(n_260) );
OAI21xp5_ASAP7_75t_L g261 ( .A1(n_243), .A2(n_201), .B(n_206), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_225), .Y(n_262) );
AO32x2_ASAP7_75t_L g263 ( .A1(n_245), .A2(n_221), .A3(n_215), .B1(n_153), .B2(n_136), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_L g264 ( .A1(n_238), .A2(n_201), .B(n_218), .C(n_190), .Y(n_264) );
AOI21x1_ASAP7_75t_L g265 ( .A1(n_227), .A2(n_136), .B(n_153), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_256), .B(n_194), .Y(n_266) );
AND2x4_ASAP7_75t_L g267 ( .A(n_232), .B(n_193), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_SL g268 ( .A1(n_238), .A2(n_235), .B(n_230), .C(n_253), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_234), .A2(n_223), .B(n_222), .Y(n_269) );
A2O1A1Ixp33_ASAP7_75t_L g270 ( .A1(n_239), .A2(n_217), .B(n_209), .C(n_208), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_252), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_237), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_240), .A2(n_219), .B(n_217), .Y(n_273) );
BUFx6f_ASAP7_75t_L g274 ( .A(n_256), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_229), .B(n_193), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_236), .A2(n_217), .B(n_209), .Y(n_276) );
AOI22xp5_ASAP7_75t_L g277 ( .A1(n_257), .A2(n_209), .B1(n_208), .B2(n_193), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_255), .A2(n_208), .B(n_214), .Y(n_278) );
AO31x2_ASAP7_75t_L g279 ( .A1(n_230), .A2(n_127), .A3(n_110), .B(n_114), .Y(n_279) );
BUFx10_ASAP7_75t_L g280 ( .A(n_254), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_260), .B(n_253), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_262), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_271), .B(n_231), .Y(n_283) );
OA21x2_ASAP7_75t_L g284 ( .A1(n_261), .A2(n_251), .B(n_250), .Y(n_284) );
OR2x2_ASAP7_75t_SL g285 ( .A(n_274), .B(n_136), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_275), .B(n_257), .Y(n_286) );
OA21x2_ASAP7_75t_L g287 ( .A1(n_265), .A2(n_228), .B(n_110), .Y(n_287) );
AO21x2_ASAP7_75t_L g288 ( .A1(n_268), .A2(n_255), .B(n_132), .Y(n_288) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_274), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_264), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_263), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_263), .Y(n_292) );
OAI21x1_ASAP7_75t_L g293 ( .A1(n_276), .A2(n_153), .B(n_120), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_263), .Y(n_294) );
OAI21x1_ASAP7_75t_L g295 ( .A1(n_259), .A2(n_132), .B(n_120), .Y(n_295) );
OAI21x1_ASAP7_75t_L g296 ( .A1(n_273), .A2(n_119), .B(n_121), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_277), .B(n_242), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_270), .Y(n_298) );
AND2x4_ASAP7_75t_SL g299 ( .A(n_274), .B(n_241), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_279), .Y(n_300) );
OAI21x1_ASAP7_75t_L g301 ( .A1(n_278), .A2(n_119), .B(n_121), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_269), .A2(n_247), .B(n_244), .Y(n_302) );
OAI21xp5_ASAP7_75t_L g303 ( .A1(n_281), .A2(n_258), .B(n_267), .Y(n_303) );
OAI22xp5_ASAP7_75t_L g304 ( .A1(n_297), .A2(n_248), .B1(n_247), .B2(n_267), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_290), .B(n_279), .Y(n_305) );
INVx3_ASAP7_75t_L g306 ( .A(n_299), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_300), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_300), .Y(n_308) );
OR2x6_ASAP7_75t_L g309 ( .A(n_284), .B(n_247), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_291), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_300), .B(n_279), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_290), .B(n_272), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_291), .Y(n_313) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_289), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_282), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_290), .B(n_116), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_282), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_291), .Y(n_318) );
INVxp67_ASAP7_75t_L g319 ( .A(n_289), .Y(n_319) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_284), .Y(n_320) );
OAI21xp5_ASAP7_75t_L g321 ( .A1(n_281), .A2(n_266), .B(n_116), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_296), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_286), .A2(n_248), .B1(n_280), .B2(n_104), .Y(n_323) );
AO21x2_ASAP7_75t_L g324 ( .A1(n_298), .A2(n_130), .B(n_127), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_286), .B(n_117), .Y(n_325) );
INVx1_ASAP7_75t_SL g326 ( .A(n_299), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_286), .B(n_117), .Y(n_327) );
OR2x2_ASAP7_75t_L g328 ( .A(n_297), .B(n_9), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_283), .B(n_9), .Y(n_329) );
NAND2x1p5_ASAP7_75t_L g330 ( .A(n_284), .B(n_241), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_296), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_291), .B(n_130), .Y(n_332) );
AO21x2_ASAP7_75t_L g333 ( .A1(n_298), .A2(n_292), .B(n_294), .Y(n_333) );
INVx2_ASAP7_75t_SL g334 ( .A(n_299), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_311), .B(n_292), .Y(n_335) );
NOR2x1_ASAP7_75t_L g336 ( .A(n_306), .B(n_288), .Y(n_336) );
BUFx2_ASAP7_75t_L g337 ( .A(n_309), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_311), .B(n_292), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_307), .B(n_292), .Y(n_339) );
AND2x2_ASAP7_75t_SL g340 ( .A(n_320), .B(n_284), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_311), .B(n_294), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_310), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_307), .B(n_294), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_308), .Y(n_344) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_314), .Y(n_345) );
AND2x4_ASAP7_75t_SL g346 ( .A(n_306), .B(n_298), .Y(n_346) );
INVx4_ASAP7_75t_L g347 ( .A(n_309), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_308), .B(n_294), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_310), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_310), .B(n_301), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_313), .B(n_301), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_313), .B(n_301), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_313), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_318), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_315), .B(n_283), .Y(n_355) );
AOI22xp33_ASAP7_75t_SL g356 ( .A1(n_304), .A2(n_284), .B1(n_288), .B2(n_299), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_318), .B(n_284), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_305), .B(n_295), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_318), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_333), .B(n_288), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_333), .Y(n_361) );
BUFx3_ASAP7_75t_L g362 ( .A(n_334), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_322), .B(n_288), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_315), .Y(n_364) );
BUFx3_ASAP7_75t_L g365 ( .A(n_334), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_317), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_317), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_322), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_333), .B(n_288), .Y(n_369) );
BUFx2_ASAP7_75t_L g370 ( .A(n_309), .Y(n_370) );
NOR2x1_ASAP7_75t_L g371 ( .A(n_306), .B(n_287), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_333), .B(n_296), .Y(n_372) );
BUFx2_ASAP7_75t_L g373 ( .A(n_309), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_331), .Y(n_374) );
BUFx3_ASAP7_75t_L g375 ( .A(n_334), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_332), .B(n_295), .Y(n_376) );
NAND2x1_ASAP7_75t_L g377 ( .A(n_309), .B(n_287), .Y(n_377) );
INVxp67_ASAP7_75t_L g378 ( .A(n_314), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_331), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_332), .Y(n_380) );
BUFx2_ASAP7_75t_L g381 ( .A(n_309), .Y(n_381) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_319), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_332), .B(n_295), .Y(n_383) );
INVx3_ASAP7_75t_L g384 ( .A(n_330), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_316), .B(n_287), .Y(n_385) );
AND2x4_ASAP7_75t_L g386 ( .A(n_320), .B(n_293), .Y(n_386) );
BUFx3_ASAP7_75t_L g387 ( .A(n_306), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_305), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_364), .B(n_325), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_335), .B(n_330), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_366), .B(n_325), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_345), .B(n_312), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_342), .Y(n_393) );
AND2x4_ASAP7_75t_L g394 ( .A(n_347), .B(n_326), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_335), .B(n_330), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_366), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_342), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_367), .B(n_327), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_342), .Y(n_399) );
NOR2x1_ASAP7_75t_L g400 ( .A(n_336), .B(n_329), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_349), .Y(n_401) );
AND2x4_ASAP7_75t_L g402 ( .A(n_347), .B(n_326), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_335), .B(n_330), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_338), .B(n_316), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_338), .B(n_316), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_345), .B(n_312), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_355), .B(n_327), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_338), .B(n_341), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_341), .B(n_324), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_367), .Y(n_410) );
INVxp67_ASAP7_75t_SL g411 ( .A(n_378), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_355), .B(n_327), .Y(n_412) );
AND2x4_ASAP7_75t_L g413 ( .A(n_347), .B(n_303), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_344), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_344), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_382), .Y(n_416) );
INVx2_ASAP7_75t_SL g417 ( .A(n_362), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_382), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_341), .B(n_319), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_343), .B(n_324), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_343), .B(n_324), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_343), .B(n_324), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_348), .B(n_303), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_348), .B(n_106), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_348), .B(n_388), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_388), .B(n_106), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_378), .B(n_328), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_339), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_388), .B(n_106), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_339), .Y(n_430) );
AND2x4_ASAP7_75t_L g431 ( .A(n_347), .B(n_106), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_380), .B(n_328), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_339), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_358), .B(n_329), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_358), .B(n_304), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_376), .A2(n_323), .B1(n_321), .B2(n_131), .Y(n_436) );
INVx3_ASAP7_75t_L g437 ( .A(n_347), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_376), .B(n_287), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_380), .B(n_321), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_376), .B(n_383), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_368), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_358), .B(n_285), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_383), .B(n_287), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_383), .B(n_287), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_356), .A2(n_302), .B1(n_104), .B2(n_293), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_380), .B(n_10), .Y(n_446) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_362), .Y(n_447) );
AND2x4_ASAP7_75t_L g448 ( .A(n_337), .B(n_302), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_385), .B(n_10), .Y(n_449) );
AND2x2_ASAP7_75t_SL g450 ( .A(n_337), .B(n_285), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_357), .B(n_148), .Y(n_451) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_362), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_365), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_368), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_365), .Y(n_455) );
AOI22xp33_ASAP7_75t_SL g456 ( .A1(n_337), .A2(n_293), .B1(n_285), .B2(n_232), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_357), .B(n_372), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_349), .Y(n_458) );
NAND2x1p5_ASAP7_75t_L g459 ( .A(n_387), .B(n_249), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_385), .B(n_11), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_357), .B(n_148), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_374), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_374), .B(n_12), .Y(n_463) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_365), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_353), .B(n_12), .Y(n_465) );
INVxp67_ASAP7_75t_L g466 ( .A(n_375), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_372), .B(n_148), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_416), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_408), .B(n_370), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_440), .B(n_353), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_418), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_440), .B(n_360), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_396), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_410), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_428), .B(n_360), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_408), .B(n_370), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_457), .B(n_354), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_414), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_430), .B(n_360), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_451), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_433), .B(n_369), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_457), .B(n_354), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_415), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_404), .B(n_359), .Y(n_484) );
NAND2x1p5_ASAP7_75t_L g485 ( .A(n_431), .B(n_375), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_411), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_392), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_404), .B(n_370), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_405), .B(n_373), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_405), .B(n_359), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_392), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_390), .B(n_373), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_424), .B(n_369), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_434), .B(n_373), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_390), .B(n_381), .Y(n_495) );
INVx1_ASAP7_75t_SL g496 ( .A(n_447), .Y(n_496) );
AND2x2_ASAP7_75t_SL g497 ( .A(n_450), .B(n_381), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_395), .B(n_375), .Y(n_498) );
INVx1_ASAP7_75t_SL g499 ( .A(n_452), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_406), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_395), .B(n_384), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_424), .B(n_369), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_406), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_407), .A2(n_356), .B1(n_340), .B2(n_363), .Y(n_504) );
INVx3_ASAP7_75t_L g505 ( .A(n_431), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_409), .B(n_372), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_441), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_454), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_393), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_409), .B(n_379), .Y(n_510) );
INVx1_ASAP7_75t_SL g511 ( .A(n_453), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_462), .Y(n_512) );
INVx3_ASAP7_75t_L g513 ( .A(n_431), .Y(n_513) );
NOR2xp67_ASAP7_75t_L g514 ( .A(n_437), .B(n_384), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_425), .B(n_379), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_419), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_425), .B(n_379), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_403), .B(n_384), .Y(n_518) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_467), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_420), .B(n_361), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_403), .B(n_384), .Y(n_521) );
INVx2_ASAP7_75t_SL g522 ( .A(n_417), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_420), .B(n_361), .Y(n_523) );
NAND2x1p5_ASAP7_75t_L g524 ( .A(n_463), .B(n_460), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_451), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_421), .B(n_361), .Y(n_526) );
NOR2x1_ASAP7_75t_L g527 ( .A(n_463), .B(n_336), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_421), .B(n_363), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_461), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_427), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_461), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_467), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_393), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_423), .B(n_384), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_460), .B(n_387), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_397), .Y(n_536) );
INVx2_ASAP7_75t_SL g537 ( .A(n_417), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_434), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_465), .Y(n_539) );
AND2x4_ASAP7_75t_SL g540 ( .A(n_455), .B(n_349), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_435), .B(n_350), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_423), .B(n_340), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_435), .B(n_350), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_422), .B(n_389), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_422), .B(n_363), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_464), .B(n_466), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_442), .B(n_350), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_442), .B(n_340), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_438), .B(n_340), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_397), .Y(n_550) );
INVx1_ASAP7_75t_SL g551 ( .A(n_426), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_391), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_398), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_399), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_399), .Y(n_555) );
NAND2x1p5_ASAP7_75t_L g556 ( .A(n_450), .B(n_387), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_401), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_469), .B(n_413), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_487), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_497), .A2(n_412), .B1(n_436), .B2(n_400), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_476), .B(n_413), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_491), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_500), .B(n_438), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_503), .Y(n_564) );
INVx2_ASAP7_75t_SL g565 ( .A(n_540), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_538), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_486), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_530), .B(n_443), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_519), .B(n_413), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_506), .B(n_443), .Y(n_570) );
O2A1O1Ixp33_ASAP7_75t_L g571 ( .A1(n_539), .A2(n_449), .B(n_524), .C(n_496), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_470), .B(n_444), .Y(n_572) );
INVx1_ASAP7_75t_SL g573 ( .A(n_540), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_468), .Y(n_574) );
INVx3_ASAP7_75t_L g575 ( .A(n_485), .Y(n_575) );
AOI221xp5_ASAP7_75t_L g576 ( .A1(n_504), .A2(n_448), .B1(n_446), .B2(n_432), .C(n_444), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_471), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_519), .B(n_394), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_516), .B(n_437), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_473), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_497), .B(n_456), .Y(n_581) );
INVxp67_ASAP7_75t_L g582 ( .A(n_546), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_492), .B(n_394), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_477), .B(n_401), .Y(n_584) );
NOR2x1_ASAP7_75t_L g585 ( .A(n_499), .B(n_437), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_509), .Y(n_586) );
INVxp67_ASAP7_75t_L g587 ( .A(n_522), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_511), .B(n_13), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_474), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_478), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_483), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_506), .B(n_458), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_498), .B(n_394), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_509), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_552), .B(n_426), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_507), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_488), .B(n_402), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_508), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_512), .Y(n_599) );
INVxp67_ASAP7_75t_L g600 ( .A(n_537), .Y(n_600) );
OAI22xp33_ASAP7_75t_L g601 ( .A1(n_556), .A2(n_445), .B1(n_377), .B2(n_459), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_482), .B(n_458), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_472), .B(n_429), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_472), .B(n_484), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_490), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_541), .B(n_429), .Y(n_606) );
AND2x4_ASAP7_75t_L g607 ( .A(n_505), .B(n_448), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_553), .B(n_386), .Y(n_608) );
INVxp67_ASAP7_75t_L g609 ( .A(n_475), .Y(n_609) );
INVxp67_ASAP7_75t_L g610 ( .A(n_475), .Y(n_610) );
OR2x2_ASAP7_75t_L g611 ( .A(n_543), .B(n_386), .Y(n_611) );
OAI21xp33_ASAP7_75t_L g612 ( .A1(n_504), .A2(n_448), .B(n_377), .Y(n_612) );
NAND4xp25_ASAP7_75t_SL g613 ( .A(n_527), .B(n_371), .C(n_439), .D(n_352), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_489), .B(n_402), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_495), .B(n_402), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_520), .B(n_386), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_515), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_515), .Y(n_618) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_517), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_524), .A2(n_386), .B1(n_346), .B2(n_363), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_501), .B(n_386), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_520), .B(n_363), .Y(n_622) );
AOI32xp33_ASAP7_75t_L g623 ( .A1(n_505), .A2(n_346), .A3(n_371), .B1(n_352), .B2(n_351), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_533), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_517), .Y(n_625) );
OAI321xp33_ASAP7_75t_L g626 ( .A1(n_556), .A2(n_459), .A3(n_352), .B1(n_351), .B2(n_148), .C(n_346), .Y(n_626) );
OR2x2_ASAP7_75t_L g627 ( .A(n_523), .B(n_351), .Y(n_627) );
OAI31xp33_ASAP7_75t_L g628 ( .A1(n_485), .A2(n_14), .A3(n_15), .B(n_16), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_518), .B(n_14), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_523), .B(n_16), .Y(n_630) );
OAI32xp33_ASAP7_75t_SL g631 ( .A1(n_609), .A2(n_17), .A3(n_18), .B1(n_19), .B2(n_20), .Y(n_631) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_619), .Y(n_632) );
OAI21xp33_ASAP7_75t_L g633 ( .A1(n_612), .A2(n_542), .B(n_548), .Y(n_633) );
AO22x1_ASAP7_75t_L g634 ( .A1(n_573), .A2(n_513), .B1(n_535), .B2(n_549), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_610), .B(n_544), .Y(n_635) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_560), .A2(n_535), .B1(n_544), .B2(n_481), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_573), .B(n_521), .Y(n_637) );
OAI211xp5_ASAP7_75t_SL g638 ( .A1(n_612), .A2(n_513), .B(n_526), .C(n_479), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_578), .B(n_565), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_617), .B(n_528), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_580), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_618), .B(n_526), .Y(n_642) );
NAND3xp33_ASAP7_75t_L g643 ( .A(n_571), .B(n_481), .C(n_479), .Y(n_643) );
XOR2x2_ASAP7_75t_L g644 ( .A(n_581), .B(n_514), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_587), .B(n_494), .Y(n_645) );
INVx2_ASAP7_75t_SL g646 ( .A(n_584), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_589), .Y(n_647) );
OAI221xp5_ASAP7_75t_L g648 ( .A1(n_560), .A2(n_502), .B1(n_493), .B2(n_528), .C(n_545), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_590), .Y(n_649) );
OAI22xp33_ASAP7_75t_L g650 ( .A1(n_620), .A2(n_493), .B1(n_502), .B2(n_547), .Y(n_650) );
NAND3xp33_ASAP7_75t_SL g651 ( .A(n_628), .B(n_551), .C(n_532), .Y(n_651) );
OAI32xp33_ASAP7_75t_L g652 ( .A1(n_600), .A2(n_575), .A3(n_604), .B1(n_572), .B2(n_570), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_626), .A2(n_480), .B(n_529), .Y(n_653) );
OAI221xp5_ASAP7_75t_SL g654 ( .A1(n_576), .A2(n_545), .B1(n_510), .B2(n_534), .C(n_531), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_620), .A2(n_525), .B1(n_510), .B2(n_554), .Y(n_655) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_602), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_591), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_596), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_625), .B(n_570), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_598), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_599), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_567), .B(n_555), .Y(n_662) );
NOR2x1_ASAP7_75t_L g663 ( .A(n_585), .B(n_536), .Y(n_663) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_588), .A2(n_557), .B1(n_550), .B2(n_533), .C(n_21), .Y(n_664) );
INVxp67_ASAP7_75t_L g665 ( .A(n_574), .Y(n_665) );
BUFx2_ASAP7_75t_L g666 ( .A(n_575), .Y(n_666) );
O2A1O1Ixp33_ASAP7_75t_L g667 ( .A1(n_628), .A2(n_557), .B(n_550), .C(n_20), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_559), .B(n_17), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_577), .Y(n_669) );
INVxp67_ASAP7_75t_L g670 ( .A(n_562), .Y(n_670) );
OAI211xp5_ASAP7_75t_SL g671 ( .A1(n_623), .A2(n_18), .B(n_21), .C(n_181), .Y(n_671) );
OR2x2_ASAP7_75t_L g672 ( .A(n_563), .B(n_23), .Y(n_672) );
OAI22xp33_ASAP7_75t_L g673 ( .A1(n_626), .A2(n_249), .B1(n_241), .B2(n_32), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_564), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_632), .Y(n_675) );
AOI21xp5_ASAP7_75t_L g676 ( .A1(n_634), .A2(n_601), .B(n_613), .Y(n_676) );
OAI221xp5_ASAP7_75t_L g677 ( .A1(n_633), .A2(n_582), .B1(n_566), .B2(n_630), .C(n_579), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_654), .A2(n_648), .B1(n_666), .B2(n_636), .Y(n_678) );
O2A1O1Ixp33_ASAP7_75t_L g679 ( .A1(n_651), .A2(n_629), .B(n_605), .C(n_568), .Y(n_679) );
AOI21xp5_ASAP7_75t_L g680 ( .A1(n_652), .A2(n_592), .B(n_608), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_671), .A2(n_607), .B1(n_569), .B2(n_603), .Y(n_681) );
O2A1O1Ixp33_ASAP7_75t_L g682 ( .A1(n_667), .A2(n_592), .B(n_563), .C(n_595), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g683 ( .A1(n_638), .A2(n_607), .B(n_616), .Y(n_683) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_644), .A2(n_606), .B(n_611), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_662), .Y(n_685) );
O2A1O1Ixp5_ASAP7_75t_SL g686 ( .A1(n_665), .A2(n_624), .B(n_594), .C(n_586), .Y(n_686) );
OAI21xp33_ASAP7_75t_SL g687 ( .A1(n_663), .A2(n_639), .B(n_646), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_643), .A2(n_627), .B1(n_561), .B2(n_558), .Y(n_688) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_631), .A2(n_597), .B1(n_614), .B2(n_622), .C(n_583), .Y(n_689) );
OAI21xp33_ASAP7_75t_SL g690 ( .A1(n_637), .A2(n_593), .B(n_615), .Y(n_690) );
OAI21xp33_ASAP7_75t_L g691 ( .A1(n_659), .A2(n_621), .B(n_181), .Y(n_691) );
A2O1A1Ixp33_ASAP7_75t_L g692 ( .A1(n_645), .A2(n_249), .B(n_241), .C(n_174), .Y(n_692) );
NOR2xp33_ASAP7_75t_SL g693 ( .A(n_673), .B(n_249), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_662), .Y(n_694) );
OA33x2_ASAP7_75t_L g695 ( .A1(n_650), .A2(n_24), .A3(n_31), .B1(n_33), .B2(n_35), .B3(n_36), .Y(n_695) );
OAI221xp5_ASAP7_75t_L g696 ( .A1(n_664), .A2(n_174), .B1(n_159), .B2(n_233), .C(n_48), .Y(n_696) );
OA22x2_ASAP7_75t_L g697 ( .A1(n_655), .A2(n_656), .B1(n_670), .B2(n_668), .Y(n_697) );
OAI21xp33_ASAP7_75t_SL g698 ( .A1(n_659), .A2(n_38), .B(n_40), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_655), .A2(n_43), .B1(n_50), .B2(n_51), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_635), .B(n_52), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_642), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g702 ( .A1(n_640), .A2(n_53), .B1(n_55), .B2(n_56), .Y(n_702) );
OAI211xp5_ASAP7_75t_L g703 ( .A1(n_653), .A2(n_57), .B(n_59), .C(n_60), .Y(n_703) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_642), .B(n_63), .Y(n_704) );
NAND3xp33_ASAP7_75t_SL g705 ( .A(n_672), .B(n_91), .C(n_65), .Y(n_705) );
AOI221x1_ASAP7_75t_L g706 ( .A1(n_641), .A2(n_64), .B1(n_66), .B2(n_68), .C(n_70), .Y(n_706) );
AOI21xp5_ASAP7_75t_L g707 ( .A1(n_674), .A2(n_72), .B(n_75), .Y(n_707) );
NAND2xp5_ASAP7_75t_SL g708 ( .A(n_647), .B(n_77), .Y(n_708) );
OAI322xp33_ASAP7_75t_L g709 ( .A1(n_649), .A2(n_79), .A3(n_82), .B1(n_84), .B2(n_85), .C1(n_86), .C2(n_87), .Y(n_709) );
NAND4xp25_ASAP7_75t_L g710 ( .A(n_693), .B(n_676), .C(n_679), .D(n_682), .Y(n_710) );
NOR3xp33_ASAP7_75t_L g711 ( .A(n_687), .B(n_703), .C(n_678), .Y(n_711) );
NAND5xp2_ASAP7_75t_L g712 ( .A(n_681), .B(n_699), .C(n_696), .D(n_707), .E(n_677), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_690), .B(n_688), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_675), .B(n_694), .Y(n_714) );
AND4x1_ASAP7_75t_L g715 ( .A(n_689), .B(n_700), .C(n_683), .D(n_684), .Y(n_715) );
INVxp67_ASAP7_75t_L g716 ( .A(n_710), .Y(n_716) );
NAND4xp25_ASAP7_75t_SL g717 ( .A(n_711), .B(n_698), .C(n_686), .D(n_680), .Y(n_717) );
NAND4xp75_ASAP7_75t_L g718 ( .A(n_713), .B(n_706), .C(n_697), .D(n_702), .Y(n_718) );
NOR3x1_ASAP7_75t_L g719 ( .A(n_715), .B(n_705), .C(n_697), .Y(n_719) );
AOI21xp5_ASAP7_75t_L g720 ( .A1(n_716), .A2(n_714), .B(n_712), .Y(n_720) );
AND2x4_ASAP7_75t_L g721 ( .A(n_719), .B(n_685), .Y(n_721) );
AND2x2_ASAP7_75t_L g722 ( .A(n_718), .B(n_701), .Y(n_722) );
BUFx3_ASAP7_75t_L g723 ( .A(n_721), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_721), .Y(n_724) );
INVx3_ASAP7_75t_SL g725 ( .A(n_723), .Y(n_725) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_724), .A2(n_720), .B1(n_722), .B2(n_717), .Y(n_726) );
OAI22x1_ASAP7_75t_L g727 ( .A1(n_725), .A2(n_724), .B1(n_723), .B2(n_704), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_726), .B(n_723), .Y(n_728) );
OAI222xp33_ASAP7_75t_L g729 ( .A1(n_728), .A2(n_708), .B1(n_658), .B2(n_660), .C1(n_661), .C2(n_669), .Y(n_729) );
OR2x6_ASAP7_75t_L g730 ( .A(n_729), .B(n_727), .Y(n_730) );
OA21x2_ASAP7_75t_L g731 ( .A1(n_730), .A2(n_691), .B(n_692), .Y(n_731) );
OAI22xp5_ASAP7_75t_SL g732 ( .A1(n_731), .A2(n_657), .B1(n_695), .B2(n_709), .Y(n_732) );
endmodule