module fake_ariane_187_n_2310 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_226, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_229, n_70, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_227, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_232, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_230, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_223, n_35, n_54, n_25, n_2310);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_226;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_229;
input n_70;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_232;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_230;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_223;
input n_35;
input n_54;
input n_25;

output n_2310;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_373;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_2207;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_2248;
wire n_813;
wire n_419;
wire n_1985;
wire n_2288;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2200;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_2233;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_249;
wire n_1108;
wire n_355;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_2185;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_382;
wire n_489;
wire n_2294;
wire n_2274;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_299;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_2262;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_2168;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_502;
wire n_2194;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_604;
wire n_677;
wire n_439;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_2184;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_321;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_2300;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_2266;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2211;
wire n_2292;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_2306;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_2285;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_2173;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2196;
wire n_1038;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_2303;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2270;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_2251;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_399;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_2212;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_2268;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2252;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2260;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_371;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_2209;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

INVx2_ASAP7_75t_L g233 ( 
.A(n_20),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_23),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_228),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_73),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_22),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_26),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_160),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_93),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_53),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_80),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_8),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_22),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_31),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_43),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_79),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_148),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_87),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_53),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_201),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_178),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_186),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_29),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_88),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_66),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_20),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_17),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_227),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_155),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_195),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_56),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_198),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_119),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_3),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_230),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g267 ( 
.A(n_165),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_79),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_92),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_176),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_12),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_108),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_4),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_196),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_37),
.Y(n_275)
);

BUFx2_ASAP7_75t_SL g276 ( 
.A(n_193),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_5),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_132),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_18),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_105),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_169),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_112),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_91),
.Y(n_283)
);

BUFx10_ASAP7_75t_L g284 ( 
.A(n_4),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_102),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_177),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_71),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_15),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_110),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_141),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_163),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_54),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_106),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_207),
.Y(n_294)
);

BUFx10_ASAP7_75t_L g295 ( 
.A(n_167),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_114),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_145),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_174),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_1),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_48),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_17),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_1),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_157),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_32),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_96),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_194),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_97),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_98),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_147),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_164),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_18),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_45),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_213),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_78),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_190),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_162),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_80),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_152),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_27),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_231),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_187),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_73),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_191),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_192),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_137),
.Y(n_325)
);

BUFx5_ASAP7_75t_L g326 ( 
.A(n_117),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_99),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_34),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_135),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_206),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_120),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_65),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_124),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_46),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_57),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_121),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_61),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_15),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_159),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_27),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_151),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_89),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_125),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_221),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_90),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_65),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_6),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_47),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_150),
.Y(n_349)
);

BUFx10_ASAP7_75t_L g350 ( 
.A(n_77),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_199),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_158),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_128),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_16),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_46),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_181),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_212),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_33),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_57),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_60),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_218),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_211),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_173),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_29),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_182),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_170),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_23),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_154),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_116),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_60),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_111),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_156),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_58),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_19),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_66),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_204),
.Y(n_376)
);

BUFx5_ASAP7_75t_L g377 ( 
.A(n_188),
.Y(n_377)
);

BUFx10_ASAP7_75t_L g378 ( 
.A(n_41),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_63),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_123),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_0),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_133),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_229),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_77),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_203),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_83),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_82),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_101),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_8),
.Y(n_389)
);

INVx4_ASAP7_75t_R g390 ( 
.A(n_34),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_3),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_82),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_54),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_200),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_64),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_202),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_33),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_131),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_26),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_94),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_183),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_126),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_217),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_127),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_24),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_47),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_197),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_219),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_138),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_37),
.Y(n_410)
);

BUFx10_ASAP7_75t_L g411 ( 
.A(n_85),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_13),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_2),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_76),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_84),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_161),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_13),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_19),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_32),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_74),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_75),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_41),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_216),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_214),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_109),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_9),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_142),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_130),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_58),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_136),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_9),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_95),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_56),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_172),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_166),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_209),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_224),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_184),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_223),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g440 ( 
.A(n_30),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_100),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_70),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g443 ( 
.A(n_153),
.Y(n_443)
);

BUFx2_ASAP7_75t_L g444 ( 
.A(n_61),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_139),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_215),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_48),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_78),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_5),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_28),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_185),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_84),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_144),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_72),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_68),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_140),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_226),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_386),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_401),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_253),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_305),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_432),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_315),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_267),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_237),
.Y(n_465)
);

INVxp67_ASAP7_75t_SL g466 ( 
.A(n_386),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_267),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_244),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_245),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_254),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_256),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_265),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_273),
.Y(n_473)
);

INVxp67_ASAP7_75t_SL g474 ( 
.A(n_386),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_279),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_440),
.B(n_0),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_281),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_299),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_267),
.Y(n_479)
);

INVxp67_ASAP7_75t_SL g480 ( 
.A(n_386),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_300),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_304),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_316),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_444),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_319),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_351),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_366),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_368),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_386),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_284),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_233),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_233),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_295),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_409),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_334),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_338),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_340),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_295),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_424),
.Y(n_499)
);

NOR2xp67_ASAP7_75t_L g500 ( 
.A(n_241),
.B(n_2),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_240),
.B(n_6),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_370),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_295),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_373),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_234),
.Y(n_505)
);

INVxp67_ASAP7_75t_SL g506 ( 
.A(n_241),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_428),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_257),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_271),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_411),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_379),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_248),
.B(n_7),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_384),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_392),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_411),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_411),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_235),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_R g518 ( 
.A(n_457),
.B(n_86),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_235),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_355),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_284),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_413),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_417),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_421),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_239),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_431),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_442),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_239),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_310),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_249),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_449),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_249),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_251),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_234),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_247),
.Y(n_535)
);

INVxp33_ASAP7_75t_L g536 ( 
.A(n_247),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_312),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_367),
.Y(n_538)
);

NOR2xp67_ASAP7_75t_L g539 ( 
.A(n_312),
.B(n_7),
.Y(n_539)
);

INVx1_ASAP7_75t_SL g540 ( 
.A(n_420),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_251),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_429),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_429),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_236),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_259),
.B(n_10),
.Y(n_545)
);

INVxp33_ASAP7_75t_L g546 ( 
.A(n_447),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_447),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_310),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_455),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_383),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_252),
.Y(n_551)
);

CKINVDCx16_ASAP7_75t_R g552 ( 
.A(n_284),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_252),
.Y(n_553)
);

INVxp33_ASAP7_75t_L g554 ( 
.A(n_455),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_296),
.Y(n_555)
);

INVxp67_ASAP7_75t_SL g556 ( 
.A(n_383),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_350),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_350),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_296),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_236),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_344),
.Y(n_561)
);

NOR2xp67_ASAP7_75t_L g562 ( 
.A(n_238),
.B(n_10),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_255),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_238),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_350),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_378),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_378),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_378),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_255),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_260),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_260),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_242),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_242),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_261),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_269),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_243),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_261),
.Y(n_577)
);

INVxp67_ASAP7_75t_SL g578 ( 
.A(n_344),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_264),
.Y(n_579)
);

INVxp67_ASAP7_75t_L g580 ( 
.A(n_243),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_264),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_458),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_477),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_460),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_458),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_461),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_489),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_463),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_489),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_555),
.Y(n_590)
);

CKINVDCx8_ASAP7_75t_R g591 ( 
.A(n_552),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_555),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_477),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_477),
.Y(n_594)
);

HB1xp67_ASAP7_75t_L g595 ( 
.A(n_573),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_576),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_477),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_477),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_483),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_559),
.Y(n_600)
);

OR2x6_ASAP7_75t_L g601 ( 
.A(n_500),
.B(n_276),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_486),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_536),
.B(n_246),
.Y(n_603)
);

INVx4_ASAP7_75t_L g604 ( 
.A(n_529),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_559),
.Y(n_605)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_540),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_487),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_556),
.B(n_274),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_488),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_561),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_464),
.B(n_266),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_561),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_529),
.B(n_283),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_491),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_464),
.B(n_266),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_491),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_R g617 ( 
.A(n_517),
.B(n_280),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_467),
.B(n_272),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_546),
.B(n_246),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_466),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_578),
.B(n_286),
.Y(n_621)
);

AND2x4_ASAP7_75t_L g622 ( 
.A(n_575),
.B(n_380),
.Y(n_622)
);

BUFx8_ASAP7_75t_L g623 ( 
.A(n_566),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_492),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_492),
.Y(n_625)
);

NAND2xp33_ASAP7_75t_SL g626 ( 
.A(n_462),
.B(n_250),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_494),
.Y(n_627)
);

BUFx10_ASAP7_75t_L g628 ( 
.A(n_459),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_535),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_L g630 ( 
.A(n_517),
.B(n_287),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_508),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_499),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_535),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_474),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_537),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_507),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_512),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_480),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_467),
.B(n_289),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_462),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_519),
.Y(n_641)
);

CKINVDCx20_ASAP7_75t_R g642 ( 
.A(n_509),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_542),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_479),
.B(n_294),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_519),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_543),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_547),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_479),
.B(n_303),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_549),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_493),
.B(n_306),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_465),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_468),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_554),
.B(n_250),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_469),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_470),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_471),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_493),
.B(n_327),
.Y(n_657)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_505),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_525),
.B(n_357),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_472),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_525),
.B(n_330),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_473),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_475),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_478),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_498),
.B(n_333),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_481),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_482),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_498),
.B(n_339),
.Y(n_668)
);

BUFx2_ASAP7_75t_L g669 ( 
.A(n_459),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_528),
.Y(n_670)
);

OA21x2_ASAP7_75t_L g671 ( 
.A1(n_501),
.A2(n_356),
.B(n_341),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_503),
.B(n_361),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_503),
.B(n_272),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_485),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_506),
.B(n_258),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_528),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_510),
.B(n_278),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_530),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_620),
.B(n_530),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_620),
.B(n_532),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_634),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_612),
.Y(n_682)
);

INVx4_ASAP7_75t_L g683 ( 
.A(n_637),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_634),
.B(n_510),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_638),
.B(n_515),
.Y(n_685)
);

BUFx2_ASAP7_75t_L g686 ( 
.A(n_606),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_637),
.B(n_532),
.Y(n_687)
);

INVx1_ASAP7_75t_SL g688 ( 
.A(n_631),
.Y(n_688)
);

AND2x4_ASAP7_75t_L g689 ( 
.A(n_601),
.B(n_567),
.Y(n_689)
);

NAND3xp33_ASAP7_75t_L g690 ( 
.A(n_661),
.B(n_541),
.C(n_533),
.Y(n_690)
);

NAND2xp33_ASAP7_75t_SL g691 ( 
.A(n_641),
.B(n_645),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_638),
.B(n_515),
.Y(n_692)
);

OR2x2_ASAP7_75t_L g693 ( 
.A(n_603),
.B(n_484),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_671),
.A2(n_545),
.B1(n_476),
.B2(n_539),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_659),
.A2(n_541),
.B1(n_551),
.B2(n_533),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_666),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_585),
.Y(n_697)
);

OAI22xp33_ASAP7_75t_L g698 ( 
.A1(n_601),
.A2(n_676),
.B1(n_678),
.B2(n_670),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_666),
.Y(n_699)
);

BUFx4f_ASAP7_75t_L g700 ( 
.A(n_637),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_612),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_656),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_671),
.A2(n_496),
.B1(n_497),
.B2(n_495),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_637),
.B(n_551),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_604),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_651),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_671),
.A2(n_504),
.B1(n_511),
.B2(n_502),
.Y(n_707)
);

NAND2x1p5_ASAP7_75t_L g708 ( 
.A(n_656),
.B(n_513),
.Y(n_708)
);

NAND2xp33_ASAP7_75t_L g709 ( 
.A(n_637),
.B(n_326),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_651),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_603),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_612),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_601),
.A2(n_563),
.B1(n_569),
.B2(n_553),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_637),
.B(n_553),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_585),
.Y(n_715)
);

AND2x6_ASAP7_75t_L g716 ( 
.A(n_622),
.B(n_380),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_584),
.Y(n_717)
);

INVx6_ASAP7_75t_L g718 ( 
.A(n_604),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_604),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_617),
.B(n_563),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_587),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_639),
.B(n_569),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_587),
.Y(n_723)
);

AND2x4_ASAP7_75t_L g724 ( 
.A(n_601),
.B(n_514),
.Y(n_724)
);

AND2x4_ASAP7_75t_L g725 ( 
.A(n_601),
.B(n_522),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_612),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_652),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_604),
.Y(n_728)
);

AND2x6_ASAP7_75t_L g729 ( 
.A(n_622),
.B(n_427),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_612),
.Y(n_730)
);

AND2x6_ASAP7_75t_L g731 ( 
.A(n_622),
.B(n_660),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_644),
.B(n_570),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_656),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_648),
.B(n_570),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_660),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_652),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_650),
.B(n_571),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_654),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_657),
.B(n_571),
.Y(n_739)
);

AND2x6_ASAP7_75t_L g740 ( 
.A(n_622),
.B(n_427),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_586),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_655),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_665),
.B(n_574),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_660),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_612),
.Y(n_745)
);

AND2x2_ASAP7_75t_SL g746 ( 
.A(n_671),
.B(n_363),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_660),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_582),
.Y(n_748)
);

INVx4_ASAP7_75t_SL g749 ( 
.A(n_654),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_662),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_668),
.B(n_516),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_654),
.Y(n_752)
);

AND2x2_ASAP7_75t_SL g753 ( 
.A(n_630),
.B(n_365),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_664),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_672),
.B(n_516),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_614),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_608),
.B(n_574),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_619),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_590),
.A2(n_600),
.B1(n_605),
.B2(n_592),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_621),
.B(n_577),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_611),
.B(n_577),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_654),
.B(n_579),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_614),
.Y(n_763)
);

INVx5_ASAP7_75t_L g764 ( 
.A(n_583),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_582),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_667),
.B(n_523),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_619),
.B(n_490),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_589),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_654),
.B(n_579),
.Y(n_769)
);

INVx4_ASAP7_75t_L g770 ( 
.A(n_654),
.Y(n_770)
);

INVx4_ASAP7_75t_L g771 ( 
.A(n_663),
.Y(n_771)
);

INVxp33_ASAP7_75t_SL g772 ( 
.A(n_640),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_663),
.B(n_581),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_663),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_614),
.Y(n_775)
);

NOR2x1p5_ASAP7_75t_L g776 ( 
.A(n_653),
.B(n_581),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_653),
.B(n_521),
.Y(n_777)
);

OR2x6_ASAP7_75t_L g778 ( 
.A(n_669),
.B(n_534),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_663),
.B(n_369),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_663),
.B(n_372),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_589),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_614),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_675),
.B(n_572),
.Y(n_783)
);

INVxp67_ASAP7_75t_SL g784 ( 
.A(n_613),
.Y(n_784)
);

OAI21xp33_ASAP7_75t_SL g785 ( 
.A1(n_675),
.A2(n_562),
.B(n_526),
.Y(n_785)
);

CKINVDCx20_ASAP7_75t_R g786 ( 
.A(n_642),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_614),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_614),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_658),
.B(n_544),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_663),
.B(n_580),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_674),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_615),
.A2(n_335),
.B1(n_359),
.B2(n_332),
.Y(n_792)
);

INVx3_ASAP7_75t_L g793 ( 
.A(n_674),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_674),
.Y(n_794)
);

INVx4_ASAP7_75t_L g795 ( 
.A(n_674),
.Y(n_795)
);

INVx5_ASAP7_75t_L g796 ( 
.A(n_583),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_618),
.B(n_560),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_674),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_628),
.Y(n_799)
);

OR2x2_ASAP7_75t_L g800 ( 
.A(n_669),
.B(n_564),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_674),
.B(n_548),
.Y(n_801)
);

OR2x2_ASAP7_75t_L g802 ( 
.A(n_595),
.B(n_524),
.Y(n_802)
);

AND2x6_ASAP7_75t_L g803 ( 
.A(n_590),
.B(n_281),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_643),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_616),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_616),
.Y(n_806)
);

BUFx3_ASAP7_75t_L g807 ( 
.A(n_646),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_592),
.B(n_550),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_628),
.B(n_396),
.Y(n_809)
);

INVx4_ASAP7_75t_L g810 ( 
.A(n_646),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_673),
.B(n_677),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_643),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_583),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_628),
.B(n_407),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_646),
.B(n_527),
.Y(n_815)
);

AOI22xp5_ASAP7_75t_L g816 ( 
.A1(n_626),
.A2(n_415),
.B1(n_337),
.B2(n_374),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_628),
.B(n_568),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_600),
.B(n_531),
.Y(n_818)
);

OR2x2_ASAP7_75t_L g819 ( 
.A(n_596),
.B(n_258),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_647),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_SL g821 ( 
.A(n_591),
.B(n_623),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_616),
.Y(n_822)
);

BUFx4f_ASAP7_75t_L g823 ( 
.A(n_647),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_588),
.Y(n_824)
);

HB1xp67_ASAP7_75t_L g825 ( 
.A(n_599),
.Y(n_825)
);

BUFx3_ASAP7_75t_L g826 ( 
.A(n_646),
.Y(n_826)
);

INVx5_ASAP7_75t_L g827 ( 
.A(n_583),
.Y(n_827)
);

OAI22xp5_ASAP7_75t_L g828 ( 
.A1(n_591),
.A2(n_262),
.B1(n_268),
.B2(n_454),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_605),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_610),
.B(n_263),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_616),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_629),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_629),
.B(n_416),
.Y(n_833)
);

INVx5_ASAP7_75t_L g834 ( 
.A(n_583),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_629),
.Y(n_835)
);

O2A1O1Ixp5_ASAP7_75t_L g836 ( 
.A1(n_762),
.A2(n_629),
.B(n_443),
.C(n_453),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_753),
.A2(n_623),
.B1(n_423),
.B2(n_345),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_805),
.Y(n_838)
);

NAND3xp33_ASAP7_75t_L g839 ( 
.A(n_760),
.B(n_623),
.C(n_268),
.Y(n_839)
);

AOI221xp5_ASAP7_75t_L g840 ( 
.A1(n_828),
.A2(n_418),
.B1(n_277),
.B2(n_275),
.C(n_262),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_805),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_806),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_748),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_748),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_686),
.B(n_602),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_753),
.B(n_623),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_760),
.B(n_635),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_806),
.Y(n_848)
);

AOI22xp5_ASAP7_75t_L g849 ( 
.A1(n_722),
.A2(n_345),
.B1(n_423),
.B2(n_430),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_757),
.B(n_722),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_700),
.B(n_278),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_789),
.B(n_607),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_784),
.B(n_624),
.Y(n_853)
);

NAND3xp33_ASAP7_75t_SL g854 ( 
.A(n_695),
.B(n_277),
.C(n_275),
.Y(n_854)
);

BUFx12f_ASAP7_75t_L g855 ( 
.A(n_717),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_734),
.B(n_624),
.Y(n_856)
);

AOI22xp5_ASAP7_75t_L g857 ( 
.A1(n_734),
.A2(n_430),
.B1(n_434),
.B2(n_435),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_737),
.B(n_625),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_737),
.B(n_635),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_743),
.A2(n_434),
.B1(n_435),
.B2(n_436),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_743),
.B(n_649),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_679),
.B(n_625),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_679),
.B(n_633),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_680),
.B(n_633),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_700),
.B(n_436),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_810),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_681),
.B(n_270),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_681),
.B(n_376),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_815),
.B(n_425),
.Y(n_869)
);

INVxp67_ASAP7_75t_L g870 ( 
.A(n_800),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_778),
.Y(n_871)
);

NOR3xp33_ASAP7_75t_L g872 ( 
.A(n_691),
.B(n_636),
.C(n_627),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_751),
.B(n_288),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_724),
.B(n_609),
.Y(n_874)
);

AND2x6_ASAP7_75t_SL g875 ( 
.A(n_778),
.B(n_520),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_755),
.B(n_292),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_732),
.B(n_301),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_682),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_765),
.Y(n_879)
);

INVx4_ASAP7_75t_L g880 ( 
.A(n_731),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_822),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_746),
.A2(n_422),
.B1(n_433),
.B2(n_448),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_831),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_732),
.B(n_302),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_831),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_811),
.B(n_437),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_768),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_815),
.B(n_437),
.Y(n_888)
);

OR2x2_ASAP7_75t_SL g889 ( 
.A(n_825),
.B(n_538),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_811),
.B(n_438),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_815),
.B(n_438),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_832),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_731),
.Y(n_893)
);

NAND2x1_ASAP7_75t_L g894 ( 
.A(n_731),
.B(n_583),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_810),
.B(n_439),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_832),
.Y(n_896)
);

BUFx2_ASAP7_75t_L g897 ( 
.A(n_786),
.Y(n_897)
);

BUFx6f_ASAP7_75t_SL g898 ( 
.A(n_778),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_783),
.B(n_439),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_739),
.B(n_311),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_768),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_724),
.B(n_632),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_724),
.B(n_445),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_767),
.B(n_777),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_725),
.B(n_445),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_746),
.A2(n_414),
.B1(n_433),
.B2(n_426),
.Y(n_906)
);

AOI22xp33_ASAP7_75t_L g907 ( 
.A1(n_694),
.A2(n_729),
.B1(n_740),
.B2(n_716),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_725),
.B(n_446),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_823),
.B(n_446),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_706),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_781),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_710),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_725),
.B(n_451),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_823),
.B(n_451),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_766),
.B(n_456),
.Y(n_915)
);

INVxp67_ASAP7_75t_SL g916 ( 
.A(n_702),
.Y(n_916)
);

INVx2_ASAP7_75t_SL g917 ( 
.A(n_802),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_766),
.B(n_456),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_727),
.Y(n_919)
);

AND2x6_ASAP7_75t_L g920 ( 
.A(n_689),
.B(n_281),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_739),
.B(n_314),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_766),
.B(n_317),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_736),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_697),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_801),
.B(n_322),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_731),
.B(n_328),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_762),
.A2(n_441),
.B(n_593),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_693),
.B(n_557),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_731),
.B(n_346),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_741),
.Y(n_930)
);

A2O1A1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_785),
.A2(n_414),
.B(n_418),
.C(n_419),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_711),
.B(n_347),
.Y(n_932)
);

A2O1A1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_694),
.A2(n_419),
.B(n_422),
.C(n_426),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_682),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_758),
.B(n_348),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_742),
.B(n_354),
.Y(n_936)
);

BUFx2_ASAP7_75t_L g937 ( 
.A(n_786),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_817),
.B(n_558),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_697),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_687),
.B(n_358),
.Y(n_940)
);

AOI22xp5_ASAP7_75t_L g941 ( 
.A1(n_761),
.A2(n_282),
.B1(n_290),
.B2(n_291),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_715),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_683),
.B(n_326),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_718),
.Y(n_944)
);

INVx5_ASAP7_75t_L g945 ( 
.A(n_803),
.Y(n_945)
);

INVxp67_ASAP7_75t_SL g946 ( 
.A(n_702),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_750),
.B(n_360),
.Y(n_947)
);

INVx2_ASAP7_75t_SL g948 ( 
.A(n_776),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_754),
.B(n_364),
.Y(n_949)
);

OAI221xp5_ASAP7_75t_L g950 ( 
.A1(n_792),
.A2(n_448),
.B1(n_450),
.B2(n_452),
.C(n_454),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_715),
.Y(n_951)
);

INVxp67_ASAP7_75t_SL g952 ( 
.A(n_733),
.Y(n_952)
);

AOI22xp33_ASAP7_75t_L g953 ( 
.A1(n_716),
.A2(n_450),
.B1(n_452),
.B2(n_565),
.Y(n_953)
);

NOR2xp67_ASAP7_75t_SL g954 ( 
.A(n_799),
.B(n_375),
.Y(n_954)
);

OR2x4_ASAP7_75t_L g955 ( 
.A(n_761),
.B(n_390),
.Y(n_955)
);

O2A1O1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_687),
.A2(n_405),
.B(n_381),
.C(n_387),
.Y(n_956)
);

BUFx6f_ASAP7_75t_SL g957 ( 
.A(n_824),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_704),
.B(n_389),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_829),
.Y(n_959)
);

OR2x2_ASAP7_75t_L g960 ( 
.A(n_688),
.B(n_391),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_818),
.B(n_393),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_818),
.B(n_830),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_733),
.B(n_395),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_683),
.B(n_326),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_721),
.Y(n_965)
);

INVxp33_ASAP7_75t_L g966 ( 
.A(n_819),
.Y(n_966)
);

AOI22xp5_ASAP7_75t_L g967 ( 
.A1(n_704),
.A2(n_353),
.B1(n_293),
.B2(n_297),
.Y(n_967)
);

NOR2xp67_ASAP7_75t_SL g968 ( 
.A(n_690),
.B(n_397),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_684),
.B(n_399),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_685),
.B(n_692),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_714),
.B(n_406),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_808),
.B(n_410),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_714),
.B(n_797),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_790),
.B(n_412),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_721),
.Y(n_975)
);

NOR2xp67_ASAP7_75t_L g976 ( 
.A(n_713),
.B(n_298),
.Y(n_976)
);

BUFx3_ASAP7_75t_L g977 ( 
.A(n_718),
.Y(n_977)
);

AND2x4_ASAP7_75t_SL g978 ( 
.A(n_689),
.B(n_281),
.Y(n_978)
);

AND2x6_ASAP7_75t_SL g979 ( 
.A(n_797),
.B(n_11),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_804),
.B(n_307),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_809),
.B(n_11),
.Y(n_981)
);

OAI22xp5_ASAP7_75t_L g982 ( 
.A1(n_769),
.A2(n_313),
.B1(n_309),
.B2(n_308),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_835),
.Y(n_983)
);

AOI221xp5_ASAP7_75t_L g984 ( 
.A1(n_698),
.A2(n_518),
.B1(n_318),
.B2(n_362),
.C(n_320),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_812),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_769),
.A2(n_773),
.B(n_719),
.Y(n_986)
);

NOR2x1p5_ASAP7_75t_L g987 ( 
.A(n_689),
.B(n_321),
.Y(n_987)
);

OR2x6_ASAP7_75t_L g988 ( 
.A(n_708),
.B(n_281),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_820),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_718),
.Y(n_990)
);

INVx8_ASAP7_75t_L g991 ( 
.A(n_716),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_696),
.Y(n_992)
);

NAND2xp33_ASAP7_75t_L g993 ( 
.A(n_705),
.B(n_326),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_SL g994 ( 
.A(n_821),
.B(n_323),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_735),
.B(n_324),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_809),
.B(n_12),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_683),
.B(n_326),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_699),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_735),
.B(n_325),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_744),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_850),
.B(n_847),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_841),
.Y(n_1002)
);

INVx1_ASAP7_75t_SL g1003 ( 
.A(n_845),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_910),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_986),
.A2(n_709),
.B(n_773),
.Y(n_1005)
);

O2A1O1Ixp33_ASAP7_75t_SL g1006 ( 
.A1(n_850),
.A2(n_814),
.B(n_720),
.C(n_833),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_893),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_973),
.A2(n_744),
.B(n_747),
.C(n_691),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_893),
.B(n_747),
.Y(n_1009)
);

AOI21x1_ASAP7_75t_L g1010 ( 
.A1(n_943),
.A2(n_791),
.B(n_774),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_970),
.A2(n_720),
.B(n_814),
.C(n_833),
.Y(n_1011)
);

AOI22x1_ASAP7_75t_L g1012 ( 
.A1(n_866),
.A2(n_795),
.B1(n_726),
.B2(n_745),
.Y(n_1012)
);

A2O1A1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_973),
.A2(n_759),
.B(n_707),
.C(n_703),
.Y(n_1013)
);

CKINVDCx10_ASAP7_75t_R g1014 ( 
.A(n_957),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_917),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_993),
.A2(n_719),
.B(n_705),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_856),
.A2(n_728),
.B(n_709),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_858),
.A2(n_728),
.B(n_807),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_912),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_847),
.B(n_708),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_930),
.Y(n_1021)
);

AOI22xp33_ASAP7_75t_L g1022 ( 
.A1(n_882),
.A2(n_906),
.B1(n_907),
.B2(n_981),
.Y(n_1022)
);

O2A1O1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_933),
.A2(n_826),
.B(n_807),
.C(n_772),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_924),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_943),
.A2(n_794),
.B(n_798),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_962),
.A2(n_826),
.B(n_795),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_897),
.Y(n_1027)
);

AOI21x1_ASAP7_75t_L g1028 ( 
.A1(n_964),
.A2(n_726),
.B(n_745),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_975),
.Y(n_1029)
);

AOI21x1_ASAP7_75t_L g1030 ( 
.A1(n_964),
.A2(n_997),
.B(n_927),
.Y(n_1030)
);

O2A1O1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_933),
.A2(n_772),
.B(n_793),
.C(n_738),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_895),
.A2(n_795),
.B(n_738),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_904),
.B(n_816),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_991),
.Y(n_1034)
);

A2O1A1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_981),
.A2(n_759),
.B(n_703),
.C(n_707),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_895),
.A2(n_752),
.B(n_793),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_886),
.B(n_770),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_859),
.B(n_716),
.Y(n_1038)
);

OR2x6_ASAP7_75t_SL g1039 ( 
.A(n_839),
.B(n_329),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_996),
.A2(n_788),
.B(n_787),
.C(n_782),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_862),
.A2(n_752),
.B(n_770),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_880),
.B(n_682),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_975),
.Y(n_1043)
);

AOI22x1_ASAP7_75t_L g1044 ( 
.A1(n_866),
.A2(n_983),
.B1(n_885),
.B2(n_892),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_863),
.A2(n_864),
.B(n_861),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_991),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_852),
.B(n_729),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_997),
.A2(n_771),
.B(n_782),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_838),
.A2(n_771),
.B(n_787),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_843),
.Y(n_1050)
);

INVx2_ASAP7_75t_SL g1051 ( 
.A(n_874),
.Y(n_1051)
);

O2A1O1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_931),
.A2(n_779),
.B(n_780),
.C(n_788),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_987),
.B(n_729),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_939),
.A2(n_723),
.B(n_779),
.Y(n_1054)
);

A2O1A1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_996),
.A2(n_723),
.B(n_780),
.C(n_712),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_842),
.A2(n_730),
.B(n_712),
.Y(n_1056)
);

BUFx2_ASAP7_75t_L g1057 ( 
.A(n_937),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_844),
.Y(n_1058)
);

NOR2x1p5_ASAP7_75t_SL g1059 ( 
.A(n_848),
.B(n_326),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_881),
.A2(n_730),
.B(n_712),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_855),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_931),
.A2(n_854),
.B(n_890),
.C(n_886),
.Y(n_1062)
);

NOR2x1_ASAP7_75t_R g1063 ( 
.A(n_874),
.B(n_331),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_890),
.B(n_682),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_851),
.A2(n_865),
.B(n_995),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_919),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_873),
.B(n_876),
.Y(n_1067)
);

CKINVDCx8_ASAP7_75t_R g1068 ( 
.A(n_875),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_851),
.A2(n_775),
.B(n_712),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_865),
.A2(n_775),
.B(n_756),
.Y(n_1070)
);

O2A1O1Ixp5_ASAP7_75t_L g1071 ( 
.A1(n_836),
.A2(n_749),
.B(n_701),
.C(n_730),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_879),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_880),
.B(n_701),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_873),
.B(n_701),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_942),
.A2(n_965),
.B(n_951),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_999),
.A2(n_775),
.B(n_756),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_974),
.A2(n_775),
.B(n_756),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_977),
.B(n_701),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_870),
.B(n_740),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_876),
.B(n_740),
.Y(n_1080)
);

NOR3xp33_ASAP7_75t_L g1081 ( 
.A(n_877),
.B(n_900),
.C(n_884),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_923),
.Y(n_1082)
);

AO21x1_ASAP7_75t_L g1083 ( 
.A1(n_940),
.A2(n_749),
.B(n_740),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_853),
.A2(n_896),
.B(n_883),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_961),
.B(n_730),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_882),
.A2(n_763),
.B1(n_756),
.B2(n_813),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_977),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_887),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_925),
.B(n_763),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_940),
.A2(n_763),
.B(n_813),
.C(n_827),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_909),
.A2(n_763),
.B(n_813),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_925),
.B(n_749),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_909),
.A2(n_813),
.B(n_827),
.Y(n_1093)
);

AOI21x1_ASAP7_75t_L g1094 ( 
.A1(n_894),
.A2(n_834),
.B(n_827),
.Y(n_1094)
);

AND2x4_ASAP7_75t_L g1095 ( 
.A(n_902),
.B(n_764),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_901),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_991),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_907),
.B(n_764),
.Y(n_1098)
);

AOI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_906),
.A2(n_398),
.B1(n_394),
.B2(n_342),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_SL g1100 ( 
.A1(n_956),
.A2(n_14),
.B(n_16),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_966),
.B(n_14),
.Y(n_1101)
);

AO32x1_ASAP7_75t_L g1102 ( 
.A1(n_911),
.A2(n_803),
.A3(n_377),
.B1(n_326),
.B2(n_594),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_914),
.A2(n_834),
.B(n_764),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_914),
.A2(n_834),
.B(n_764),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_966),
.B(n_21),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_963),
.A2(n_834),
.B(n_796),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_992),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_980),
.A2(n_796),
.B(n_388),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_916),
.A2(n_796),
.B(n_343),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_946),
.A2(n_796),
.B(n_349),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_952),
.A2(n_352),
.B(n_382),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_877),
.A2(n_402),
.B1(n_371),
.B2(n_385),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_867),
.B(n_803),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_928),
.B(n_21),
.Y(n_1114)
);

BUFx2_ASAP7_75t_L g1115 ( 
.A(n_871),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_878),
.B(n_326),
.Y(n_1116)
);

NOR2x1p5_ASAP7_75t_SL g1117 ( 
.A(n_959),
.B(n_377),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_969),
.B(n_24),
.Y(n_1118)
);

AND2x4_ASAP7_75t_L g1119 ( 
.A(n_948),
.B(n_803),
.Y(n_1119)
);

CKINVDCx10_ASAP7_75t_R g1120 ( 
.A(n_957),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_868),
.B(n_803),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_958),
.B(n_403),
.Y(n_1122)
);

HB1xp67_ASAP7_75t_L g1123 ( 
.A(n_988),
.Y(n_1123)
);

AOI21xp33_ASAP7_75t_L g1124 ( 
.A1(n_884),
.A2(n_404),
.B(n_408),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_846),
.B(n_25),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_846),
.B(n_25),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_958),
.B(n_28),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1000),
.A2(n_598),
.B(n_597),
.Y(n_1128)
);

O2A1O1Ixp5_ASAP7_75t_L g1129 ( 
.A1(n_971),
.A2(n_377),
.B(n_597),
.C(n_594),
.Y(n_1129)
);

OAI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_998),
.A2(n_377),
.B(n_597),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_971),
.B(n_30),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_900),
.B(n_31),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_921),
.B(n_35),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_899),
.B(n_35),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_921),
.B(n_36),
.Y(n_1135)
);

NOR2xp67_ASAP7_75t_L g1136 ( 
.A(n_960),
.B(n_837),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_926),
.A2(n_598),
.B(n_597),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_985),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_929),
.A2(n_598),
.B(n_597),
.Y(n_1139)
);

OAI21xp33_ASAP7_75t_L g1140 ( 
.A1(n_849),
.A2(n_285),
.B(n_336),
.Y(n_1140)
);

OR2x2_ASAP7_75t_L g1141 ( 
.A(n_938),
.B(n_36),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_857),
.B(n_38),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_989),
.B(n_38),
.Y(n_1143)
);

AOI22x1_ASAP7_75t_L g1144 ( 
.A1(n_944),
.A2(n_598),
.B1(n_597),
.B2(n_594),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_978),
.Y(n_1145)
);

AOI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_860),
.A2(n_377),
.B1(n_400),
.B2(n_336),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_978),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_944),
.A2(n_598),
.B(n_594),
.Y(n_1148)
);

A2O1A1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_950),
.A2(n_984),
.B(n_932),
.C(n_953),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_990),
.Y(n_1150)
);

OAI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_888),
.A2(n_400),
.B1(n_336),
.B2(n_285),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_990),
.A2(n_598),
.B(n_594),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_936),
.A2(n_377),
.B(n_593),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_891),
.A2(n_594),
.B(n_593),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_889),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_878),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_878),
.B(n_377),
.Y(n_1157)
);

AOI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_953),
.A2(n_377),
.B1(n_400),
.B2(n_336),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_915),
.A2(n_593),
.B(n_400),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_918),
.A2(n_593),
.B(n_400),
.Y(n_1160)
);

A2O1A1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_840),
.A2(n_285),
.B(n_40),
.C(n_42),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_878),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_947),
.A2(n_285),
.B(n_103),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_934),
.Y(n_1164)
);

AOI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_869),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_1165)
);

INVx3_ASAP7_75t_L g1166 ( 
.A(n_934),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_SL g1167 ( 
.A(n_898),
.B(n_994),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_934),
.Y(n_1168)
);

AOI21x1_ASAP7_75t_L g1169 ( 
.A1(n_968),
.A2(n_104),
.B(n_225),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_934),
.B(n_39),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_949),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_922),
.A2(n_232),
.B(n_222),
.Y(n_1172)
);

OAI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_935),
.A2(n_220),
.B(n_210),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_972),
.B(n_43),
.Y(n_1174)
);

INVx3_ASAP7_75t_L g1175 ( 
.A(n_920),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_988),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_903),
.A2(n_208),
.B(n_205),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_920),
.Y(n_1178)
);

NAND2x1_ASAP7_75t_L g1179 ( 
.A(n_920),
.B(n_189),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_920),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_905),
.B(n_44),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_908),
.B(n_44),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_988),
.Y(n_1183)
);

A2O1A1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_976),
.A2(n_45),
.B(n_49),
.C(n_50),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1067),
.A2(n_913),
.B(n_941),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1001),
.A2(n_982),
.B(n_955),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1095),
.B(n_872),
.Y(n_1187)
);

INVx4_ASAP7_75t_L g1188 ( 
.A(n_1021),
.Y(n_1188)
);

INVx4_ASAP7_75t_L g1189 ( 
.A(n_1007),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1045),
.A2(n_955),
.B(n_967),
.Y(n_1190)
);

AOI21xp33_ASAP7_75t_L g1191 ( 
.A1(n_1067),
.A2(n_954),
.B(n_945),
.Y(n_1191)
);

NAND2x1p5_ASAP7_75t_L g1192 ( 
.A(n_1007),
.B(n_945),
.Y(n_1192)
);

NOR2xp67_ASAP7_75t_SL g1193 ( 
.A(n_1061),
.B(n_945),
.Y(n_1193)
);

INVx4_ASAP7_75t_L g1194 ( 
.A(n_1007),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1004),
.Y(n_1195)
);

NAND2xp33_ASAP7_75t_SL g1196 ( 
.A(n_1132),
.B(n_898),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_1034),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1028),
.A2(n_920),
.B(n_945),
.Y(n_1198)
);

NAND2x1p5_ASAP7_75t_L g1199 ( 
.A(n_1007),
.B(n_979),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1033),
.B(n_49),
.Y(n_1200)
);

BUFx2_ASAP7_75t_L g1201 ( 
.A(n_1027),
.Y(n_1201)
);

INVx3_ASAP7_75t_L g1202 ( 
.A(n_1034),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_1057),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1016),
.A2(n_50),
.B(n_51),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1003),
.B(n_1033),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1074),
.A2(n_51),
.B(n_52),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1019),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1017),
.A2(n_52),
.B(n_55),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1066),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1010),
.A2(n_180),
.B(n_179),
.Y(n_1210)
);

OR2x2_ASAP7_75t_L g1211 ( 
.A(n_1015),
.B(n_55),
.Y(n_1211)
);

HB1xp67_ASAP7_75t_L g1212 ( 
.A(n_1015),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_SL g1213 ( 
.A1(n_1133),
.A2(n_59),
.B(n_62),
.Y(n_1213)
);

AOI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1081),
.A2(n_59),
.B1(n_62),
.B2(n_63),
.Y(n_1214)
);

AOI21xp33_ASAP7_75t_L g1215 ( 
.A1(n_1135),
.A2(n_64),
.B(n_67),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1074),
.A2(n_67),
.B(n_68),
.Y(n_1216)
);

AOI21xp33_ASAP7_75t_L g1217 ( 
.A1(n_1022),
.A2(n_69),
.B(n_70),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_1014),
.Y(n_1218)
);

AOI21xp33_ASAP7_75t_L g1219 ( 
.A1(n_1022),
.A2(n_69),
.B(n_71),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1137),
.A2(n_118),
.B(n_171),
.Y(n_1220)
);

OR2x2_ASAP7_75t_L g1221 ( 
.A(n_1051),
.B(n_72),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1082),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1085),
.A2(n_74),
.B(n_75),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1081),
.B(n_76),
.Y(n_1224)
);

NOR2xp67_ASAP7_75t_L g1225 ( 
.A(n_1171),
.B(n_129),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_SL g1226 ( 
.A1(n_1127),
.A2(n_81),
.B(n_83),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1020),
.A2(n_81),
.B(n_107),
.Y(n_1227)
);

INVx1_ASAP7_75t_SL g1228 ( 
.A(n_1115),
.Y(n_1228)
);

AOI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1142),
.A2(n_113),
.B1(n_115),
.B2(n_122),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1114),
.B(n_134),
.Y(n_1230)
);

INVx2_ASAP7_75t_SL g1231 ( 
.A(n_1120),
.Y(n_1231)
);

AOI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1065),
.A2(n_143),
.B(n_146),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1138),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1149),
.B(n_149),
.Y(n_1234)
);

AOI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1089),
.A2(n_1077),
.B(n_1076),
.Y(n_1235)
);

A2O1A1Ixp33_ASAP7_75t_L g1236 ( 
.A1(n_1142),
.A2(n_168),
.B(n_175),
.C(n_1149),
.Y(n_1236)
);

AOI21xp33_ASAP7_75t_L g1237 ( 
.A1(n_1131),
.A2(n_1062),
.B(n_1122),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1136),
.B(n_1047),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1080),
.A2(n_1018),
.B(n_1038),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1139),
.A2(n_1012),
.B(n_1030),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1026),
.A2(n_1005),
.B(n_1011),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1107),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1050),
.Y(n_1243)
);

AO21x1_ASAP7_75t_L g1244 ( 
.A1(n_1173),
.A2(n_1118),
.B(n_1064),
.Y(n_1244)
);

OAI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1040),
.A2(n_1008),
.B(n_1084),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1155),
.B(n_1101),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1095),
.B(n_1053),
.Y(n_1247)
);

INVx4_ASAP7_75t_L g1248 ( 
.A(n_1034),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1013),
.A2(n_1134),
.B1(n_1035),
.B2(n_1118),
.Y(n_1249)
);

CKINVDCx11_ASAP7_75t_R g1250 ( 
.A(n_1068),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1101),
.B(n_1105),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1134),
.A2(n_1174),
.B1(n_1009),
.B2(n_1181),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1041),
.A2(n_1064),
.B(n_1052),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1075),
.A2(n_1054),
.B(n_1091),
.Y(n_1254)
);

AOI21x1_ASAP7_75t_SL g1255 ( 
.A1(n_1182),
.A2(n_1143),
.B(n_1092),
.Y(n_1255)
);

BUFx8_ASAP7_75t_L g1256 ( 
.A(n_1141),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_SL g1257 ( 
.A1(n_1090),
.A2(n_1098),
.B(n_1034),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1044),
.A2(n_1069),
.B(n_1070),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1006),
.A2(n_1049),
.B(n_1154),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1009),
.A2(n_1158),
.B1(n_1161),
.B2(n_1099),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1079),
.B(n_1150),
.Y(n_1261)
);

NAND2x1p5_ASAP7_75t_L g1262 ( 
.A(n_1046),
.B(n_1097),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_1053),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1056),
.A2(n_1060),
.B(n_1094),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1105),
.B(n_1125),
.Y(n_1265)
);

AOI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1125),
.A2(n_1126),
.B1(n_1112),
.B2(n_1124),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1024),
.Y(n_1267)
);

A2O1A1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1126),
.A2(n_1037),
.B(n_1161),
.C(n_1023),
.Y(n_1268)
);

A2O1A1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1037),
.A2(n_1031),
.B(n_1140),
.C(n_1184),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1048),
.A2(n_1036),
.B(n_1153),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1029),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_1087),
.B(n_1063),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1128),
.A2(n_1025),
.B(n_1129),
.Y(n_1273)
);

OAI22x1_ASAP7_75t_L g1274 ( 
.A1(n_1165),
.A2(n_1123),
.B1(n_1170),
.B2(n_1183),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1058),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1129),
.A2(n_1071),
.B(n_1144),
.Y(n_1276)
);

INVxp67_ASAP7_75t_L g1277 ( 
.A(n_1167),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_1046),
.Y(n_1278)
);

INVx3_ASAP7_75t_L g1279 ( 
.A(n_1046),
.Y(n_1279)
);

OAI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1032),
.A2(n_1071),
.B(n_1055),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_SL g1281 ( 
.A(n_1168),
.B(n_1166),
.Y(n_1281)
);

OA22x2_ASAP7_75t_L g1282 ( 
.A1(n_1146),
.A2(n_1100),
.B1(n_1147),
.B2(n_1145),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1087),
.B(n_1176),
.Y(n_1283)
);

A2O1A1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1184),
.A2(n_1055),
.B(n_1172),
.C(n_1177),
.Y(n_1284)
);

AO31x2_ASAP7_75t_L g1285 ( 
.A1(n_1083),
.A2(n_1151),
.A3(n_1160),
.B(n_1159),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1163),
.A2(n_1098),
.B(n_1086),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_SL g1287 ( 
.A1(n_1046),
.A2(n_1097),
.B(n_1042),
.Y(n_1287)
);

INVx2_ASAP7_75t_SL g1288 ( 
.A(n_1119),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1043),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1106),
.A2(n_1116),
.B(n_1157),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1116),
.A2(n_1157),
.B(n_1108),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1093),
.A2(n_1130),
.B(n_1042),
.Y(n_1292)
);

OAI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1073),
.A2(n_1156),
.B(n_1164),
.Y(n_1293)
);

INVx4_ASAP7_75t_L g1294 ( 
.A(n_1097),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_1097),
.B(n_1119),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1072),
.B(n_1096),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1073),
.A2(n_1104),
.B(n_1103),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1148),
.A2(n_1152),
.B(n_1169),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1088),
.B(n_1166),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_L g1300 ( 
.A(n_1162),
.B(n_1039),
.Y(n_1300)
);

BUFx2_ASAP7_75t_L g1301 ( 
.A(n_1162),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1078),
.A2(n_1178),
.B(n_1180),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1175),
.B(n_1168),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1078),
.A2(n_1121),
.B(n_1113),
.Y(n_1304)
);

OAI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1109),
.A2(n_1110),
.B(n_1111),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1170),
.A2(n_1168),
.B(n_1102),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1175),
.B(n_1168),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1102),
.A2(n_1179),
.B(n_1059),
.Y(n_1308)
);

AOI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1117),
.A2(n_1028),
.B(n_1065),
.Y(n_1309)
);

AOI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1102),
.A2(n_1028),
.B(n_1065),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1001),
.A2(n_1045),
.B(n_1067),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1067),
.B(n_1001),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_SL g1313 ( 
.A(n_1081),
.B(n_1067),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1002),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1028),
.A2(n_1010),
.B(n_1137),
.Y(n_1315)
);

OAI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1067),
.A2(n_1001),
.B(n_850),
.Y(n_1316)
);

NAND2x1p5_ASAP7_75t_L g1317 ( 
.A(n_1007),
.B(n_893),
.Y(n_1317)
);

OR2x6_ASAP7_75t_L g1318 ( 
.A(n_1051),
.B(n_991),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1067),
.A2(n_1001),
.B(n_850),
.Y(n_1319)
);

OAI222xp33_ASAP7_75t_L g1320 ( 
.A1(n_1022),
.A2(n_906),
.B1(n_882),
.B2(n_1158),
.C1(n_837),
.C2(n_1067),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1001),
.A2(n_1045),
.B(n_1067),
.Y(n_1321)
);

AOI221xp5_ASAP7_75t_L g1322 ( 
.A1(n_1067),
.A2(n_1001),
.B1(n_1081),
.B2(n_1142),
.C(n_1022),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1028),
.A2(n_1010),
.B(n_1137),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1028),
.A2(n_1010),
.B(n_1137),
.Y(n_1324)
);

O2A1O1Ixp5_ASAP7_75t_L g1325 ( 
.A1(n_1067),
.A2(n_1127),
.B(n_1131),
.C(n_1132),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1028),
.A2(n_1010),
.B(n_1137),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1028),
.A2(n_1010),
.B(n_1137),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1001),
.B(n_850),
.Y(n_1328)
);

AOI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1028),
.A2(n_1065),
.B(n_1089),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1004),
.Y(n_1330)
);

BUFx5_ASAP7_75t_L g1331 ( 
.A(n_1009),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1001),
.B(n_850),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1003),
.B(n_870),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1028),
.A2(n_1010),
.B(n_1137),
.Y(n_1334)
);

INVx1_ASAP7_75t_SL g1335 ( 
.A(n_1027),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1001),
.A2(n_1045),
.B(n_1067),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_SL g1337 ( 
.A1(n_1132),
.A2(n_1135),
.B(n_1133),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1001),
.A2(n_1045),
.B(n_1067),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1001),
.B(n_850),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1001),
.A2(n_1045),
.B(n_1067),
.Y(n_1340)
);

INVx2_ASAP7_75t_SL g1341 ( 
.A(n_1021),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1028),
.A2(n_1010),
.B(n_1137),
.Y(n_1342)
);

INVxp67_ASAP7_75t_L g1343 ( 
.A(n_1333),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1195),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1312),
.A2(n_1322),
.B1(n_1316),
.B2(n_1319),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1207),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1311),
.A2(n_1336),
.B(n_1321),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1312),
.B(n_1328),
.Y(n_1348)
);

INVx1_ASAP7_75t_SL g1349 ( 
.A(n_1335),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_SL g1350 ( 
.A(n_1322),
.B(n_1266),
.Y(n_1350)
);

BUFx6f_ASAP7_75t_L g1351 ( 
.A(n_1247),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1240),
.A2(n_1298),
.B(n_1254),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1338),
.A2(n_1340),
.B(n_1313),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1338),
.A2(n_1340),
.B(n_1313),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1332),
.B(n_1339),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1251),
.A2(n_1265),
.B1(n_1205),
.B2(n_1249),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1212),
.B(n_1246),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1242),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1200),
.A2(n_1224),
.B1(n_1185),
.B2(n_1236),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1331),
.B(n_1238),
.Y(n_1360)
);

INVx5_ASAP7_75t_L g1361 ( 
.A(n_1318),
.Y(n_1361)
);

INVx4_ASAP7_75t_SL g1362 ( 
.A(n_1318),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1212),
.B(n_1201),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1203),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1244),
.A2(n_1237),
.B(n_1286),
.Y(n_1365)
);

A2O1A1Ixp33_ASAP7_75t_SL g1366 ( 
.A1(n_1208),
.A2(n_1241),
.B(n_1305),
.C(n_1191),
.Y(n_1366)
);

BUFx2_ASAP7_75t_SL g1367 ( 
.A(n_1188),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1228),
.Y(n_1368)
);

AND2x6_ASAP7_75t_L g1369 ( 
.A(n_1303),
.B(n_1307),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1247),
.B(n_1318),
.Y(n_1370)
);

BUFx12f_ASAP7_75t_L g1371 ( 
.A(n_1250),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1209),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1222),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1211),
.B(n_1341),
.Y(n_1374)
);

BUFx6f_ASAP7_75t_SL g1375 ( 
.A(n_1218),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1233),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1330),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1315),
.A2(n_1342),
.B(n_1323),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1243),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1256),
.A2(n_1217),
.B1(n_1219),
.B2(n_1275),
.Y(n_1380)
);

NAND2xp33_ASAP7_75t_L g1381 ( 
.A(n_1236),
.B(n_1331),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1248),
.Y(n_1382)
);

INVx4_ASAP7_75t_L g1383 ( 
.A(n_1188),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1199),
.B(n_1187),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1263),
.B(n_1295),
.Y(n_1385)
);

O2A1O1Ixp5_ASAP7_75t_SL g1386 ( 
.A1(n_1215),
.A2(n_1252),
.B(n_1281),
.C(n_1280),
.Y(n_1386)
);

INVx8_ASAP7_75t_L g1387 ( 
.A(n_1295),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1331),
.B(n_1268),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1286),
.A2(n_1239),
.B(n_1297),
.Y(n_1389)
);

INVxp67_ASAP7_75t_SL g1390 ( 
.A(n_1331),
.Y(n_1390)
);

INVx4_ASAP7_75t_L g1391 ( 
.A(n_1248),
.Y(n_1391)
);

INVx3_ASAP7_75t_L g1392 ( 
.A(n_1294),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1324),
.A2(n_1334),
.B(n_1327),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1239),
.A2(n_1297),
.B(n_1284),
.Y(n_1394)
);

BUFx2_ASAP7_75t_L g1395 ( 
.A(n_1256),
.Y(n_1395)
);

INVx1_ASAP7_75t_SL g1396 ( 
.A(n_1301),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1331),
.B(n_1186),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1296),
.Y(n_1398)
);

AOI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1196),
.A2(n_1187),
.B1(n_1272),
.B2(n_1277),
.Y(n_1399)
);

NAND3xp33_ASAP7_75t_L g1400 ( 
.A(n_1214),
.B(n_1206),
.C(n_1216),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1284),
.A2(n_1253),
.B(n_1325),
.Y(n_1401)
);

AOI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1325),
.A2(n_1270),
.B(n_1245),
.Y(n_1402)
);

INVx1_ASAP7_75t_SL g1403 ( 
.A(n_1283),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1270),
.A2(n_1259),
.B(n_1337),
.Y(n_1404)
);

AND2x4_ASAP7_75t_L g1405 ( 
.A(n_1277),
.B(n_1288),
.Y(n_1405)
);

INVx3_ASAP7_75t_L g1406 ( 
.A(n_1294),
.Y(n_1406)
);

O2A1O1Ixp5_ASAP7_75t_L g1407 ( 
.A1(n_1320),
.A2(n_1234),
.B(n_1190),
.C(n_1290),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1331),
.B(n_1186),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1326),
.A2(n_1258),
.B(n_1264),
.Y(n_1409)
);

HB1xp67_ASAP7_75t_L g1410 ( 
.A(n_1221),
.Y(n_1410)
);

NAND2x1p5_ASAP7_75t_L g1411 ( 
.A(n_1189),
.B(n_1194),
.Y(n_1411)
);

CKINVDCx20_ASAP7_75t_R g1412 ( 
.A(n_1231),
.Y(n_1412)
);

NAND3xp33_ASAP7_75t_L g1413 ( 
.A(n_1206),
.B(n_1216),
.C(n_1229),
.Y(n_1413)
);

AOI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1272),
.A2(n_1260),
.B1(n_1300),
.B2(n_1230),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1300),
.B(n_1261),
.Y(n_1415)
);

OAI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1320),
.A2(n_1190),
.B(n_1269),
.Y(n_1416)
);

NOR2x1_ASAP7_75t_L g1417 ( 
.A(n_1278),
.B(n_1189),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1267),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1274),
.A2(n_1271),
.B1(n_1314),
.B2(n_1289),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1261),
.A2(n_1225),
.B1(n_1299),
.B2(n_1282),
.Y(n_1420)
);

A2O1A1Ixp33_ASAP7_75t_L g1421 ( 
.A1(n_1227),
.A2(n_1204),
.B(n_1223),
.C(n_1306),
.Y(n_1421)
);

AND2x4_ASAP7_75t_L g1422 ( 
.A(n_1303),
.B(n_1307),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1299),
.B(n_1317),
.Y(n_1423)
);

BUFx2_ASAP7_75t_SL g1424 ( 
.A(n_1194),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1235),
.A2(n_1329),
.B(n_1309),
.Y(n_1425)
);

INVx5_ASAP7_75t_L g1426 ( 
.A(n_1197),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1317),
.B(n_1257),
.Y(n_1427)
);

INVx3_ASAP7_75t_L g1428 ( 
.A(n_1262),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1223),
.Y(n_1429)
);

INVx1_ASAP7_75t_SL g1430 ( 
.A(n_1281),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1197),
.B(n_1279),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1291),
.A2(n_1276),
.B(n_1292),
.Y(n_1432)
);

NOR2x1_ASAP7_75t_SL g1433 ( 
.A(n_1232),
.B(n_1310),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1202),
.B(n_1293),
.Y(n_1434)
);

NAND2x1_ASAP7_75t_SL g1435 ( 
.A(n_1202),
.B(n_1193),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1287),
.B(n_1262),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1192),
.B(n_1204),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_R g1438 ( 
.A(n_1192),
.B(n_1255),
.Y(n_1438)
);

NOR2xp67_ASAP7_75t_L g1439 ( 
.A(n_1227),
.B(n_1306),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1282),
.Y(n_1440)
);

O2A1O1Ixp5_ASAP7_75t_L g1441 ( 
.A1(n_1308),
.A2(n_1255),
.B(n_1285),
.C(n_1273),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1304),
.B(n_1302),
.Y(n_1442)
);

OAI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1308),
.A2(n_1220),
.B(n_1210),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1198),
.A2(n_1213),
.B(n_1226),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1285),
.B(n_1312),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_L g1446 ( 
.A(n_1312),
.B(n_772),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1195),
.Y(n_1447)
);

INVx1_ASAP7_75t_SL g1448 ( 
.A(n_1335),
.Y(n_1448)
);

INVxp67_ASAP7_75t_L g1449 ( 
.A(n_1333),
.Y(n_1449)
);

BUFx12f_ASAP7_75t_L g1450 ( 
.A(n_1250),
.Y(n_1450)
);

NAND2x1_ASAP7_75t_L g1451 ( 
.A(n_1287),
.B(n_1162),
.Y(n_1451)
);

O2A1O1Ixp5_ASAP7_75t_L g1452 ( 
.A1(n_1244),
.A2(n_1067),
.B(n_1313),
.C(n_1249),
.Y(n_1452)
);

BUFx6f_ASAP7_75t_L g1453 ( 
.A(n_1247),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1205),
.B(n_1333),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1240),
.A2(n_1298),
.B(n_1254),
.Y(n_1455)
);

AOI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1311),
.A2(n_1340),
.B(n_1336),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1205),
.B(n_1333),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1195),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1242),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_SL g1460 ( 
.A1(n_1312),
.A2(n_786),
.B1(n_1142),
.B2(n_889),
.Y(n_1460)
);

BUFx2_ASAP7_75t_L g1461 ( 
.A(n_1201),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1312),
.B(n_1316),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1195),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1312),
.B(n_1316),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1195),
.Y(n_1465)
);

A2O1A1Ixp33_ASAP7_75t_L g1466 ( 
.A1(n_1322),
.A2(n_1067),
.B(n_1081),
.C(n_850),
.Y(n_1466)
);

AOI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1312),
.A2(n_1067),
.B1(n_1081),
.B2(n_1322),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1201),
.Y(n_1468)
);

AND2x4_ASAP7_75t_L g1469 ( 
.A(n_1247),
.B(n_1318),
.Y(n_1469)
);

OAI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1265),
.A2(n_1067),
.B1(n_1266),
.B2(n_1200),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1247),
.B(n_1318),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_SL g1472 ( 
.A(n_1322),
.B(n_1081),
.Y(n_1472)
);

BUFx6f_ASAP7_75t_L g1473 ( 
.A(n_1247),
.Y(n_1473)
);

INVx2_ASAP7_75t_SL g1474 ( 
.A(n_1201),
.Y(n_1474)
);

OAI221xp5_ASAP7_75t_L g1475 ( 
.A1(n_1322),
.A2(n_1312),
.B1(n_1067),
.B2(n_1319),
.C(n_1316),
.Y(n_1475)
);

INVx2_ASAP7_75t_SL g1476 ( 
.A(n_1201),
.Y(n_1476)
);

AO21x1_ASAP7_75t_L g1477 ( 
.A1(n_1249),
.A2(n_1067),
.B(n_1081),
.Y(n_1477)
);

A2O1A1Ixp33_ASAP7_75t_L g1478 ( 
.A1(n_1322),
.A2(n_1067),
.B(n_1081),
.C(n_850),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1205),
.B(n_1333),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1195),
.Y(n_1480)
);

BUFx2_ASAP7_75t_L g1481 ( 
.A(n_1201),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1195),
.Y(n_1482)
);

INVx3_ASAP7_75t_L g1483 ( 
.A(n_1248),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1205),
.B(n_1333),
.Y(n_1484)
);

A2O1A1Ixp33_ASAP7_75t_L g1485 ( 
.A1(n_1322),
.A2(n_1067),
.B(n_1081),
.C(n_850),
.Y(n_1485)
);

INVx2_ASAP7_75t_SL g1486 ( 
.A(n_1201),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_1250),
.Y(n_1487)
);

BUFx3_ASAP7_75t_L g1488 ( 
.A(n_1201),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1242),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1195),
.Y(n_1490)
);

A2O1A1Ixp33_ASAP7_75t_L g1491 ( 
.A1(n_1322),
.A2(n_1067),
.B(n_1081),
.C(n_850),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1312),
.A2(n_1001),
.B1(n_1322),
.B2(n_1319),
.Y(n_1492)
);

INVx1_ASAP7_75t_SL g1493 ( 
.A(n_1335),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1322),
.A2(n_1067),
.B1(n_1081),
.B2(n_1022),
.Y(n_1494)
);

AOI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1311),
.A2(n_1340),
.B(n_1336),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1242),
.Y(n_1496)
);

OAI21x1_ASAP7_75t_L g1497 ( 
.A1(n_1240),
.A2(n_1298),
.B(n_1254),
.Y(n_1497)
);

NAND2x1_ASAP7_75t_L g1498 ( 
.A(n_1287),
.B(n_1162),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1195),
.Y(n_1499)
);

BUFx6f_ASAP7_75t_L g1500 ( 
.A(n_1247),
.Y(n_1500)
);

BUFx3_ASAP7_75t_L g1501 ( 
.A(n_1201),
.Y(n_1501)
);

AND2x4_ASAP7_75t_L g1502 ( 
.A(n_1247),
.B(n_1318),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1205),
.B(n_1335),
.Y(n_1503)
);

BUFx8_ASAP7_75t_L g1504 ( 
.A(n_1218),
.Y(n_1504)
);

INVx3_ASAP7_75t_L g1505 ( 
.A(n_1248),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1248),
.Y(n_1506)
);

INVx3_ASAP7_75t_L g1507 ( 
.A(n_1248),
.Y(n_1507)
);

BUFx10_ASAP7_75t_L g1508 ( 
.A(n_1218),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1357),
.B(n_1454),
.Y(n_1509)
);

INVx3_ASAP7_75t_L g1510 ( 
.A(n_1437),
.Y(n_1510)
);

AOI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1359),
.A2(n_1350),
.B(n_1365),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1429),
.Y(n_1512)
);

BUFx12f_ASAP7_75t_L g1513 ( 
.A(n_1487),
.Y(n_1513)
);

BUFx2_ASAP7_75t_SL g1514 ( 
.A(n_1375),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1344),
.Y(n_1515)
);

INVx1_ASAP7_75t_SL g1516 ( 
.A(n_1349),
.Y(n_1516)
);

BUFx2_ASAP7_75t_L g1517 ( 
.A(n_1468),
.Y(n_1517)
);

BUFx2_ASAP7_75t_R g1518 ( 
.A(n_1395),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1445),
.B(n_1472),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1346),
.Y(n_1520)
);

INVx3_ASAP7_75t_L g1521 ( 
.A(n_1426),
.Y(n_1521)
);

OA21x2_ASAP7_75t_L g1522 ( 
.A1(n_1389),
.A2(n_1394),
.B(n_1347),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1475),
.A2(n_1460),
.B1(n_1467),
.B2(n_1494),
.Y(n_1523)
);

OAI21x1_ASAP7_75t_L g1524 ( 
.A1(n_1352),
.A2(n_1497),
.B(n_1455),
.Y(n_1524)
);

CKINVDCx20_ASAP7_75t_R g1525 ( 
.A(n_1412),
.Y(n_1525)
);

AND2x4_ASAP7_75t_L g1526 ( 
.A(n_1362),
.B(n_1361),
.Y(n_1526)
);

BUFx8_ASAP7_75t_L g1527 ( 
.A(n_1375),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1363),
.Y(n_1528)
);

BUFx12f_ASAP7_75t_L g1529 ( 
.A(n_1371),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1372),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1373),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1376),
.Y(n_1532)
);

HB1xp67_ASAP7_75t_L g1533 ( 
.A(n_1368),
.Y(n_1533)
);

INVx8_ASAP7_75t_L g1534 ( 
.A(n_1387),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1397),
.Y(n_1535)
);

INVxp67_ASAP7_75t_SL g1536 ( 
.A(n_1423),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1377),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_L g1538 ( 
.A(n_1475),
.B(n_1446),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1348),
.B(n_1355),
.Y(n_1539)
);

BUFx12f_ASAP7_75t_L g1540 ( 
.A(n_1450),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1447),
.Y(n_1541)
);

AOI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1492),
.A2(n_1470),
.B1(n_1345),
.B2(n_1359),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1458),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1463),
.Y(n_1544)
);

AOI21xp5_ASAP7_75t_L g1545 ( 
.A1(n_1466),
.A2(n_1485),
.B(n_1478),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1465),
.Y(n_1546)
);

OAI21x1_ASAP7_75t_L g1547 ( 
.A1(n_1409),
.A2(n_1425),
.B(n_1432),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1348),
.B(n_1355),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1480),
.Y(n_1549)
);

AOI222xp33_ASAP7_75t_L g1550 ( 
.A1(n_1492),
.A2(n_1345),
.B1(n_1416),
.B2(n_1356),
.C1(n_1491),
.C2(n_1464),
.Y(n_1550)
);

BUFx2_ASAP7_75t_L g1551 ( 
.A(n_1488),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1482),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1396),
.Y(n_1553)
);

CKINVDCx20_ASAP7_75t_R g1554 ( 
.A(n_1504),
.Y(n_1554)
);

INVx5_ASAP7_75t_L g1555 ( 
.A(n_1369),
.Y(n_1555)
);

BUFx2_ASAP7_75t_L g1556 ( 
.A(n_1501),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1416),
.A2(n_1477),
.B1(n_1457),
.B2(n_1484),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1490),
.Y(n_1558)
);

OAI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1414),
.A2(n_1464),
.B1(n_1462),
.B2(n_1399),
.Y(n_1559)
);

AO21x1_ASAP7_75t_SL g1560 ( 
.A1(n_1388),
.A2(n_1442),
.B(n_1420),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1499),
.Y(n_1561)
);

INVxp33_ASAP7_75t_L g1562 ( 
.A(n_1479),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_SL g1563 ( 
.A1(n_1440),
.A2(n_1400),
.B1(n_1413),
.B2(n_1381),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1379),
.Y(n_1564)
);

BUFx6f_ASAP7_75t_L g1565 ( 
.A(n_1387),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1358),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1459),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1462),
.B(n_1349),
.Y(n_1568)
);

AOI21x1_ASAP7_75t_L g1569 ( 
.A1(n_1444),
.A2(n_1404),
.B(n_1354),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1489),
.Y(n_1570)
);

INVxp67_ASAP7_75t_SL g1571 ( 
.A(n_1423),
.Y(n_1571)
);

AO21x2_ASAP7_75t_L g1572 ( 
.A1(n_1443),
.A2(n_1421),
.B(n_1439),
.Y(n_1572)
);

CKINVDCx6p67_ASAP7_75t_R g1573 ( 
.A(n_1508),
.Y(n_1573)
);

OA21x2_ASAP7_75t_L g1574 ( 
.A1(n_1347),
.A2(n_1456),
.B(n_1495),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_1504),
.Y(n_1575)
);

AOI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1415),
.A2(n_1380),
.B1(n_1374),
.B2(n_1448),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1496),
.Y(n_1577)
);

CKINVDCx6p67_ASAP7_75t_R g1578 ( 
.A(n_1508),
.Y(n_1578)
);

NAND2x1p5_ASAP7_75t_L g1579 ( 
.A(n_1426),
.B(n_1370),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1418),
.Y(n_1580)
);

INVx4_ASAP7_75t_L g1581 ( 
.A(n_1384),
.Y(n_1581)
);

INVx4_ASAP7_75t_L g1582 ( 
.A(n_1370),
.Y(n_1582)
);

INVx3_ASAP7_75t_L g1583 ( 
.A(n_1411),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1343),
.A2(n_1449),
.B1(n_1503),
.B2(n_1410),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1396),
.Y(n_1585)
);

INVx1_ASAP7_75t_SL g1586 ( 
.A(n_1448),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1398),
.Y(n_1587)
);

BUFx2_ASAP7_75t_R g1588 ( 
.A(n_1367),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1403),
.Y(n_1589)
);

OAI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1493),
.A2(n_1360),
.B1(n_1388),
.B2(n_1476),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1403),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1434),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1431),
.Y(n_1593)
);

OAI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1360),
.A2(n_1474),
.B1(n_1486),
.B2(n_1500),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1364),
.B(n_1461),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_SL g1596 ( 
.A1(n_1405),
.A2(n_1401),
.B1(n_1502),
.B2(n_1471),
.Y(n_1596)
);

NOR2x1_ASAP7_75t_R g1597 ( 
.A(n_1383),
.B(n_1481),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_1383),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1419),
.A2(n_1469),
.B1(n_1502),
.B2(n_1385),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1430),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1431),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1422),
.B(n_1351),
.Y(n_1602)
);

CKINVDCx11_ASAP7_75t_R g1603 ( 
.A(n_1351),
.Y(n_1603)
);

BUFx12f_ASAP7_75t_L g1604 ( 
.A(n_1453),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1430),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1452),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1441),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1436),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1436),
.Y(n_1609)
);

INVx5_ASAP7_75t_L g1610 ( 
.A(n_1369),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1453),
.B(n_1473),
.Y(n_1611)
);

INVx8_ASAP7_75t_L g1612 ( 
.A(n_1369),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1422),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1433),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1427),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1427),
.Y(n_1616)
);

OAI21x1_ASAP7_75t_L g1617 ( 
.A1(n_1456),
.A2(n_1393),
.B(n_1378),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1407),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1390),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1428),
.Y(n_1620)
);

INVx1_ASAP7_75t_SL g1621 ( 
.A(n_1453),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1428),
.Y(n_1622)
);

AO21x1_ASAP7_75t_SL g1623 ( 
.A1(n_1443),
.A2(n_1386),
.B(n_1366),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1353),
.Y(n_1624)
);

NAND2x1p5_ASAP7_75t_L g1625 ( 
.A(n_1451),
.B(n_1498),
.Y(n_1625)
);

CKINVDCx16_ASAP7_75t_R g1626 ( 
.A(n_1473),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1353),
.B(n_1402),
.Y(n_1627)
);

OAI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1382),
.A2(n_1507),
.B1(n_1392),
.B2(n_1406),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1424),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1382),
.Y(n_1630)
);

INVx6_ASAP7_75t_L g1631 ( 
.A(n_1500),
.Y(n_1631)
);

OAI21x1_ASAP7_75t_L g1632 ( 
.A1(n_1411),
.A2(n_1435),
.B(n_1392),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1406),
.Y(n_1633)
);

BUFx6f_ASAP7_75t_SL g1634 ( 
.A(n_1391),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1483),
.Y(n_1635)
);

INVx3_ASAP7_75t_L g1636 ( 
.A(n_1483),
.Y(n_1636)
);

OAI21x1_ASAP7_75t_SL g1637 ( 
.A1(n_1391),
.A2(n_1417),
.B(n_1438),
.Y(n_1637)
);

BUFx3_ASAP7_75t_L g1638 ( 
.A(n_1507),
.Y(n_1638)
);

INVx2_ASAP7_75t_SL g1639 ( 
.A(n_1505),
.Y(n_1639)
);

AO22x1_ASAP7_75t_L g1640 ( 
.A1(n_1505),
.A2(n_1081),
.B1(n_1067),
.B2(n_1142),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1506),
.A2(n_1350),
.B1(n_1322),
.B2(n_1081),
.Y(n_1641)
);

BUFx3_ASAP7_75t_L g1642 ( 
.A(n_1506),
.Y(n_1642)
);

AO21x2_ASAP7_75t_L g1643 ( 
.A1(n_1443),
.A2(n_1416),
.B(n_1421),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1344),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_SL g1645 ( 
.A1(n_1460),
.A2(n_1067),
.B1(n_461),
.B2(n_463),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1344),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1344),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1348),
.B(n_1312),
.Y(n_1648)
);

OAI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1467),
.A2(n_1067),
.B1(n_1312),
.B2(n_1475),
.Y(n_1649)
);

OAI21x1_ASAP7_75t_L g1650 ( 
.A1(n_1352),
.A2(n_1497),
.B(n_1455),
.Y(n_1650)
);

OAI22xp5_ASAP7_75t_SL g1651 ( 
.A1(n_1460),
.A2(n_1446),
.B1(n_1467),
.B2(n_1475),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1357),
.B(n_1454),
.Y(n_1652)
);

BUFx6f_ASAP7_75t_L g1653 ( 
.A(n_1387),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1344),
.Y(n_1654)
);

AOI22xp33_ASAP7_75t_L g1655 ( 
.A1(n_1350),
.A2(n_1322),
.B1(n_1081),
.B2(n_1022),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1445),
.B(n_1472),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1344),
.Y(n_1657)
);

AND2x4_ASAP7_75t_L g1658 ( 
.A(n_1362),
.B(n_1361),
.Y(n_1658)
);

CKINVDCx20_ASAP7_75t_R g1659 ( 
.A(n_1412),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1344),
.Y(n_1660)
);

CKINVDCx11_ASAP7_75t_R g1661 ( 
.A(n_1371),
.Y(n_1661)
);

BUFx3_ASAP7_75t_L g1662 ( 
.A(n_1468),
.Y(n_1662)
);

OAI21x1_ASAP7_75t_L g1663 ( 
.A1(n_1352),
.A2(n_1497),
.B(n_1455),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1344),
.Y(n_1664)
);

OAI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1467),
.A2(n_1067),
.B1(n_1312),
.B2(n_1475),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1363),
.Y(n_1666)
);

AO21x1_ASAP7_75t_SL g1667 ( 
.A1(n_1494),
.A2(n_1416),
.B(n_1408),
.Y(n_1667)
);

BUFx2_ASAP7_75t_R g1668 ( 
.A(n_1487),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1344),
.Y(n_1669)
);

BUFx12f_ASAP7_75t_L g1670 ( 
.A(n_1487),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_SL g1671 ( 
.A1(n_1460),
.A2(n_1067),
.B1(n_461),
.B2(n_463),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1344),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1344),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1350),
.A2(n_1322),
.B1(n_1081),
.B2(n_1022),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1344),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1350),
.A2(n_1322),
.B1(n_1081),
.B2(n_1022),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1648),
.B(n_1525),
.Y(n_1677)
);

BUFx6f_ASAP7_75t_L g1678 ( 
.A(n_1555),
.Y(n_1678)
);

OR2x6_ASAP7_75t_L g1679 ( 
.A(n_1612),
.B(n_1526),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1519),
.B(n_1656),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_1553),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1525),
.B(n_1659),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1512),
.Y(n_1683)
);

OR2x6_ASAP7_75t_L g1684 ( 
.A(n_1612),
.B(n_1526),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1519),
.B(n_1656),
.Y(n_1685)
);

AO21x2_ASAP7_75t_L g1686 ( 
.A1(n_1511),
.A2(n_1618),
.B(n_1542),
.Y(n_1686)
);

INVx4_ASAP7_75t_L g1687 ( 
.A(n_1521),
.Y(n_1687)
);

BUFx3_ASAP7_75t_L g1688 ( 
.A(n_1662),
.Y(n_1688)
);

HB1xp67_ASAP7_75t_L g1689 ( 
.A(n_1585),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1568),
.B(n_1539),
.Y(n_1690)
);

BUFx3_ASAP7_75t_L g1691 ( 
.A(n_1662),
.Y(n_1691)
);

INVx3_ASAP7_75t_L g1692 ( 
.A(n_1614),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1515),
.Y(n_1693)
);

AO21x2_ASAP7_75t_L g1694 ( 
.A1(n_1618),
.A2(n_1606),
.B(n_1624),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1510),
.B(n_1667),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1520),
.Y(n_1696)
);

BUFx3_ASAP7_75t_L g1697 ( 
.A(n_1517),
.Y(n_1697)
);

OR2x6_ASAP7_75t_L g1698 ( 
.A(n_1612),
.B(n_1526),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1548),
.B(n_1509),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1652),
.B(n_1538),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1510),
.B(n_1627),
.Y(n_1701)
);

BUFx2_ASAP7_75t_L g1702 ( 
.A(n_1614),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1538),
.B(n_1649),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1592),
.Y(n_1704)
);

BUFx3_ASAP7_75t_L g1705 ( 
.A(n_1551),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1615),
.Y(n_1706)
);

OAI21x1_ASAP7_75t_L g1707 ( 
.A1(n_1569),
.A2(n_1617),
.B(n_1547),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_SL g1708 ( 
.A1(n_1651),
.A2(n_1665),
.B1(n_1545),
.B2(n_1612),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1616),
.Y(n_1709)
);

HB1xp67_ASAP7_75t_L g1710 ( 
.A(n_1533),
.Y(n_1710)
);

AND2x4_ASAP7_75t_L g1711 ( 
.A(n_1510),
.B(n_1555),
.Y(n_1711)
);

INVx3_ASAP7_75t_L g1712 ( 
.A(n_1535),
.Y(n_1712)
);

BUFx3_ASAP7_75t_L g1713 ( 
.A(n_1556),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1608),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1609),
.Y(n_1715)
);

INVx1_ASAP7_75t_SL g1716 ( 
.A(n_1518),
.Y(n_1716)
);

INVx3_ASAP7_75t_L g1717 ( 
.A(n_1572),
.Y(n_1717)
);

INVx3_ASAP7_75t_L g1718 ( 
.A(n_1572),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1559),
.B(n_1528),
.Y(n_1719)
);

CKINVDCx20_ASAP7_75t_R g1720 ( 
.A(n_1659),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1530),
.Y(n_1721)
);

HB1xp67_ASAP7_75t_L g1722 ( 
.A(n_1666),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1531),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1532),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1600),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_L g1726 ( 
.A(n_1575),
.B(n_1554),
.Y(n_1726)
);

AND2x4_ASAP7_75t_L g1727 ( 
.A(n_1555),
.B(n_1610),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1575),
.B(n_1554),
.Y(n_1728)
);

OAI21x1_ASAP7_75t_L g1729 ( 
.A1(n_1524),
.A2(n_1663),
.B(n_1650),
.Y(n_1729)
);

INVx4_ASAP7_75t_L g1730 ( 
.A(n_1521),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1537),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1541),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_SL g1733 ( 
.A(n_1590),
.B(n_1594),
.Y(n_1733)
);

CKINVDCx5p33_ASAP7_75t_R g1734 ( 
.A(n_1661),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1627),
.B(n_1643),
.Y(n_1735)
);

HB1xp67_ASAP7_75t_SL g1736 ( 
.A(n_1527),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1593),
.Y(n_1737)
);

AOI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1523),
.A2(n_1676),
.B1(n_1674),
.B2(n_1655),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1516),
.B(n_1586),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1543),
.B(n_1544),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1601),
.Y(n_1741)
);

INVx3_ASAP7_75t_L g1742 ( 
.A(n_1521),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1546),
.B(n_1549),
.Y(n_1743)
);

NAND2x1_ASAP7_75t_L g1744 ( 
.A(n_1637),
.B(n_1607),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1536),
.B(n_1571),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1605),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1605),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1552),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_SL g1749 ( 
.A(n_1668),
.B(n_1588),
.Y(n_1749)
);

HB1xp67_ASAP7_75t_L g1750 ( 
.A(n_1595),
.Y(n_1750)
);

BUFx2_ASAP7_75t_L g1751 ( 
.A(n_1619),
.Y(n_1751)
);

OAI21x1_ASAP7_75t_L g1752 ( 
.A1(n_1625),
.A2(n_1522),
.B(n_1574),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1558),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1564),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1561),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1644),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1550),
.B(n_1641),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1646),
.Y(n_1758)
);

INVxp67_ASAP7_75t_L g1759 ( 
.A(n_1597),
.Y(n_1759)
);

OAI21x1_ASAP7_75t_L g1760 ( 
.A1(n_1625),
.A2(n_1522),
.B(n_1574),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1647),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1654),
.B(n_1657),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1660),
.Y(n_1763)
);

INVx2_ASAP7_75t_SL g1764 ( 
.A(n_1638),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1664),
.Y(n_1765)
);

AO21x1_ASAP7_75t_L g1766 ( 
.A1(n_1669),
.A2(n_1675),
.B(n_1673),
.Y(n_1766)
);

INVx2_ASAP7_75t_SL g1767 ( 
.A(n_1638),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1672),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1580),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1589),
.Y(n_1770)
);

BUFx3_ASAP7_75t_L g1771 ( 
.A(n_1598),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1587),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1591),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1522),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1630),
.Y(n_1775)
);

INVxp67_ASAP7_75t_L g1776 ( 
.A(n_1613),
.Y(n_1776)
);

HB1xp67_ASAP7_75t_L g1777 ( 
.A(n_1633),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1566),
.Y(n_1778)
);

AOI21x1_ASAP7_75t_L g1779 ( 
.A1(n_1640),
.A2(n_1574),
.B(n_1628),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1567),
.Y(n_1780)
);

AO21x2_ASAP7_75t_L g1781 ( 
.A1(n_1570),
.A2(n_1577),
.B(n_1620),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1622),
.Y(n_1782)
);

INVx3_ASAP7_75t_L g1783 ( 
.A(n_1632),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1563),
.Y(n_1784)
);

HB1xp67_ASAP7_75t_L g1785 ( 
.A(n_1635),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1636),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1560),
.B(n_1557),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_L g1788 ( 
.A(n_1598),
.B(n_1578),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1557),
.B(n_1562),
.Y(n_1789)
);

INVx3_ASAP7_75t_L g1790 ( 
.A(n_1636),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1636),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1642),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1581),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1581),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1639),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1562),
.B(n_1641),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1523),
.B(n_1676),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1581),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_SL g1799 ( 
.A(n_1596),
.B(n_1674),
.Y(n_1799)
);

AND2x4_ASAP7_75t_L g1800 ( 
.A(n_1610),
.B(n_1658),
.Y(n_1800)
);

AO21x2_ASAP7_75t_L g1801 ( 
.A1(n_1576),
.A2(n_1611),
.B(n_1623),
.Y(n_1801)
);

AND2x4_ASAP7_75t_L g1802 ( 
.A(n_1610),
.B(n_1582),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1639),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1642),
.Y(n_1804)
);

CKINVDCx6p67_ASAP7_75t_R g1805 ( 
.A(n_1661),
.Y(n_1805)
);

INVxp67_ASAP7_75t_L g1806 ( 
.A(n_1602),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1584),
.B(n_1655),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1582),
.B(n_1584),
.Y(n_1808)
);

BUFx2_ASAP7_75t_L g1809 ( 
.A(n_1583),
.Y(n_1809)
);

HB1xp67_ASAP7_75t_L g1810 ( 
.A(n_1694),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1735),
.B(n_1582),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1735),
.B(n_1629),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1766),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1701),
.B(n_1610),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1680),
.B(n_1514),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1766),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1701),
.B(n_1583),
.Y(n_1817)
);

BUFx2_ASAP7_75t_L g1818 ( 
.A(n_1702),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1706),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1706),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1709),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1703),
.B(n_1599),
.Y(n_1822)
);

OR2x2_ASAP7_75t_L g1823 ( 
.A(n_1680),
.B(n_1626),
.Y(n_1823)
);

OR2x2_ASAP7_75t_L g1824 ( 
.A(n_1685),
.B(n_1579),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1694),
.B(n_1573),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1709),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1737),
.B(n_1573),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1683),
.Y(n_1828)
);

OR2x2_ASAP7_75t_L g1829 ( 
.A(n_1685),
.B(n_1578),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1745),
.B(n_1621),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1683),
.Y(n_1831)
);

INVx4_ASAP7_75t_L g1832 ( 
.A(n_1678),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_1751),
.Y(n_1833)
);

INVx2_ASAP7_75t_SL g1834 ( 
.A(n_1783),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1774),
.B(n_1631),
.Y(n_1835)
);

HB1xp67_ASAP7_75t_L g1836 ( 
.A(n_1751),
.Y(n_1836)
);

INVxp67_ASAP7_75t_L g1837 ( 
.A(n_1801),
.Y(n_1837)
);

HB1xp67_ASAP7_75t_L g1838 ( 
.A(n_1761),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1686),
.B(n_1631),
.Y(n_1839)
);

OR2x6_ASAP7_75t_L g1840 ( 
.A(n_1727),
.B(n_1534),
.Y(n_1840)
);

INVxp67_ASAP7_75t_L g1841 ( 
.A(n_1801),
.Y(n_1841)
);

OR2x2_ASAP7_75t_L g1842 ( 
.A(n_1745),
.B(n_1565),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1737),
.B(n_1671),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1741),
.B(n_1645),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1686),
.B(n_1631),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1722),
.B(n_1653),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1686),
.B(n_1603),
.Y(n_1847)
);

HB1xp67_ASAP7_75t_L g1848 ( 
.A(n_1681),
.Y(n_1848)
);

HB1xp67_ASAP7_75t_L g1849 ( 
.A(n_1689),
.Y(n_1849)
);

NOR2x1_ASAP7_75t_L g1850 ( 
.A(n_1801),
.B(n_1653),
.Y(n_1850)
);

NOR2xp33_ASAP7_75t_L g1851 ( 
.A(n_1677),
.B(n_1513),
.Y(n_1851)
);

INVx2_ASAP7_75t_SL g1852 ( 
.A(n_1783),
.Y(n_1852)
);

HB1xp67_ASAP7_75t_L g1853 ( 
.A(n_1710),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1712),
.B(n_1603),
.Y(n_1854)
);

BUFx2_ASAP7_75t_L g1855 ( 
.A(n_1702),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1748),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1773),
.B(n_1534),
.Y(n_1857)
);

INVxp67_ASAP7_75t_SL g1858 ( 
.A(n_1717),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1717),
.B(n_1540),
.Y(n_1859)
);

OR2x2_ASAP7_75t_L g1860 ( 
.A(n_1773),
.B(n_1534),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1748),
.Y(n_1861)
);

NOR2xp33_ASAP7_75t_L g1862 ( 
.A(n_1771),
.B(n_1513),
.Y(n_1862)
);

HB1xp67_ASAP7_75t_L g1863 ( 
.A(n_1750),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1717),
.B(n_1540),
.Y(n_1864)
);

BUFx2_ASAP7_75t_L g1865 ( 
.A(n_1695),
.Y(n_1865)
);

HB1xp67_ASAP7_75t_L g1866 ( 
.A(n_1775),
.Y(n_1866)
);

HB1xp67_ASAP7_75t_L g1867 ( 
.A(n_1777),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1718),
.B(n_1529),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1718),
.B(n_1529),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1741),
.B(n_1690),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1718),
.B(n_1670),
.Y(n_1871)
);

AND2x4_ASAP7_75t_L g1872 ( 
.A(n_1711),
.B(n_1783),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1740),
.B(n_1527),
.Y(n_1873)
);

BUFx2_ASAP7_75t_L g1874 ( 
.A(n_1695),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1752),
.B(n_1670),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1752),
.B(n_1604),
.Y(n_1876)
);

BUFx2_ASAP7_75t_L g1877 ( 
.A(n_1692),
.Y(n_1877)
);

BUFx3_ASAP7_75t_L g1878 ( 
.A(n_1688),
.Y(n_1878)
);

NOR2xp33_ASAP7_75t_L g1879 ( 
.A(n_1771),
.B(n_1527),
.Y(n_1879)
);

AOI21xp33_ASAP7_75t_L g1880 ( 
.A1(n_1757),
.A2(n_1604),
.B(n_1534),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1865),
.B(n_1697),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1863),
.B(n_1700),
.Y(n_1882)
);

OAI21xp5_ASAP7_75t_SL g1883 ( 
.A1(n_1875),
.A2(n_1708),
.B(n_1738),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1838),
.B(n_1740),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1838),
.Y(n_1885)
);

NAND4xp25_ASAP7_75t_L g1886 ( 
.A(n_1827),
.B(n_1719),
.C(n_1697),
.D(n_1713),
.Y(n_1886)
);

AOI221xp5_ASAP7_75t_L g1887 ( 
.A1(n_1813),
.A2(n_1784),
.B1(n_1797),
.B2(n_1789),
.C(n_1799),
.Y(n_1887)
);

NAND3xp33_ASAP7_75t_L g1888 ( 
.A(n_1813),
.B(n_1733),
.C(n_1784),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1812),
.B(n_1787),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1848),
.B(n_1743),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1848),
.B(n_1743),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_SL g1892 ( 
.A(n_1825),
.B(n_1764),
.Y(n_1892)
);

AOI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1816),
.A2(n_1744),
.B(n_1787),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1849),
.B(n_1762),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1812),
.B(n_1692),
.Y(n_1895)
);

OAI221xp5_ASAP7_75t_SL g1896 ( 
.A1(n_1816),
.A2(n_1807),
.B1(n_1796),
.B2(n_1789),
.C(n_1808),
.Y(n_1896)
);

AOI221xp5_ASAP7_75t_L g1897 ( 
.A1(n_1843),
.A2(n_1807),
.B1(n_1770),
.B2(n_1763),
.C(n_1721),
.Y(n_1897)
);

OAI221xp5_ASAP7_75t_SL g1898 ( 
.A1(n_1837),
.A2(n_1796),
.B1(n_1808),
.B2(n_1776),
.C(n_1759),
.Y(n_1898)
);

OAI21xp5_ASAP7_75t_SL g1899 ( 
.A1(n_1875),
.A2(n_1788),
.B(n_1716),
.Y(n_1899)
);

OAI221xp5_ASAP7_75t_L g1900 ( 
.A1(n_1822),
.A2(n_1844),
.B1(n_1843),
.B2(n_1837),
.C(n_1841),
.Y(n_1900)
);

AOI21xp5_ASAP7_75t_L g1901 ( 
.A1(n_1850),
.A2(n_1744),
.B(n_1760),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1849),
.B(n_1762),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1853),
.B(n_1699),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1853),
.B(n_1705),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1866),
.B(n_1867),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_SL g1906 ( 
.A(n_1825),
.B(n_1764),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_SL g1907 ( 
.A(n_1825),
.B(n_1767),
.Y(n_1907)
);

NOR3xp33_ASAP7_75t_L g1908 ( 
.A(n_1841),
.B(n_1804),
.C(n_1779),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1812),
.B(n_1705),
.Y(n_1909)
);

NOR2xp33_ASAP7_75t_L g1910 ( 
.A(n_1827),
.B(n_1713),
.Y(n_1910)
);

OAI22xp5_ASAP7_75t_L g1911 ( 
.A1(n_1822),
.A2(n_1815),
.B1(n_1829),
.B2(n_1873),
.Y(n_1911)
);

OAI21xp5_ASAP7_75t_SL g1912 ( 
.A1(n_1875),
.A2(n_1779),
.B(n_1682),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1870),
.B(n_1739),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1856),
.Y(n_1914)
);

NOR3xp33_ASAP7_75t_L g1915 ( 
.A(n_1859),
.B(n_1804),
.C(n_1792),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1856),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1870),
.B(n_1693),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1833),
.B(n_1696),
.Y(n_1918)
);

OA211x2_ASAP7_75t_L g1919 ( 
.A1(n_1879),
.A2(n_1749),
.B(n_1726),
.C(n_1728),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1865),
.B(n_1688),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1833),
.B(n_1723),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1836),
.B(n_1724),
.Y(n_1922)
);

AOI22xp5_ASAP7_75t_L g1923 ( 
.A1(n_1847),
.A2(n_1684),
.B1(n_1698),
.B2(n_1679),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1836),
.B(n_1819),
.Y(n_1924)
);

AOI221xp5_ASAP7_75t_L g1925 ( 
.A1(n_1844),
.A2(n_1753),
.B1(n_1732),
.B2(n_1755),
.C(n_1756),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1819),
.B(n_1731),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1820),
.B(n_1758),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1874),
.B(n_1692),
.Y(n_1928)
);

NAND3xp33_ASAP7_75t_L g1929 ( 
.A(n_1850),
.B(n_1785),
.C(n_1795),
.Y(n_1929)
);

AOI22xp33_ASAP7_75t_L g1930 ( 
.A1(n_1847),
.A2(n_1805),
.B1(n_1772),
.B2(n_1780),
.Y(n_1930)
);

OAI21xp33_ASAP7_75t_L g1931 ( 
.A1(n_1835),
.A2(n_1795),
.B(n_1803),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1874),
.B(n_1765),
.Y(n_1932)
);

NAND4xp25_ASAP7_75t_L g1933 ( 
.A(n_1829),
.B(n_1803),
.C(n_1786),
.D(n_1791),
.Y(n_1933)
);

OAI22xp5_ASAP7_75t_L g1934 ( 
.A1(n_1815),
.A2(n_1720),
.B1(n_1805),
.B2(n_1691),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1820),
.B(n_1768),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1811),
.B(n_1691),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1811),
.B(n_1767),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1821),
.B(n_1754),
.Y(n_1938)
);

OAI221xp5_ASAP7_75t_L g1939 ( 
.A1(n_1847),
.A2(n_1754),
.B1(n_1772),
.B2(n_1782),
.C(n_1806),
.Y(n_1939)
);

OAI21xp33_ASAP7_75t_L g1940 ( 
.A1(n_1835),
.A2(n_1786),
.B(n_1791),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1821),
.B(n_1782),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1826),
.B(n_1714),
.Y(n_1942)
);

NOR2xp33_ASAP7_75t_L g1943 ( 
.A(n_1873),
.B(n_1809),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1826),
.B(n_1714),
.Y(n_1944)
);

OAI21xp5_ASAP7_75t_SL g1945 ( 
.A1(n_1871),
.A2(n_1802),
.B(n_1736),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_SL g1946 ( 
.A(n_1818),
.B(n_1793),
.Y(n_1946)
);

OAI22xp5_ASAP7_75t_L g1947 ( 
.A1(n_1823),
.A2(n_1720),
.B1(n_1794),
.B2(n_1793),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1817),
.B(n_1794),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1830),
.B(n_1715),
.Y(n_1949)
);

NOR2xp33_ASAP7_75t_L g1950 ( 
.A(n_1871),
.B(n_1798),
.Y(n_1950)
);

AOI22xp33_ASAP7_75t_L g1951 ( 
.A1(n_1839),
.A2(n_1778),
.B1(n_1780),
.B2(n_1781),
.Y(n_1951)
);

AOI211xp5_ASAP7_75t_L g1952 ( 
.A1(n_1871),
.A2(n_1734),
.B(n_1798),
.C(n_1778),
.Y(n_1952)
);

OA21x2_ASAP7_75t_L g1953 ( 
.A1(n_1858),
.A2(n_1729),
.B(n_1707),
.Y(n_1953)
);

OAI22xp5_ASAP7_75t_L g1954 ( 
.A1(n_1823),
.A2(n_1734),
.B1(n_1790),
.B2(n_1634),
.Y(n_1954)
);

AND2x2_ASAP7_75t_SL g1955 ( 
.A(n_1818),
.B(n_1800),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1830),
.B(n_1715),
.Y(n_1956)
);

NOR2xp33_ASAP7_75t_SL g1957 ( 
.A(n_1851),
.B(n_1802),
.Y(n_1957)
);

AOI221x1_ASAP7_75t_SL g1958 ( 
.A1(n_1861),
.A2(n_1769),
.B1(n_1746),
.B2(n_1747),
.C(n_1704),
.Y(n_1958)
);

NAND3xp33_ASAP7_75t_L g1959 ( 
.A(n_1842),
.B(n_1747),
.C(n_1746),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1861),
.B(n_1790),
.Y(n_1960)
);

NOR3xp33_ASAP7_75t_L g1961 ( 
.A(n_1859),
.B(n_1742),
.C(n_1730),
.Y(n_1961)
);

NAND3xp33_ASAP7_75t_L g1962 ( 
.A(n_1842),
.B(n_1769),
.C(n_1725),
.Y(n_1962)
);

OA211x2_ASAP7_75t_L g1963 ( 
.A1(n_1862),
.A2(n_1634),
.B(n_1730),
.C(n_1687),
.Y(n_1963)
);

OAI221xp5_ASAP7_75t_L g1964 ( 
.A1(n_1839),
.A2(n_1845),
.B1(n_1880),
.B2(n_1860),
.C(n_1857),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1855),
.B(n_1878),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1889),
.B(n_1872),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1889),
.B(n_1872),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1914),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1958),
.B(n_1855),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1881),
.B(n_1920),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1955),
.B(n_1872),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1916),
.Y(n_1972)
);

AND2x4_ASAP7_75t_L g1973 ( 
.A(n_1961),
.B(n_1872),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1953),
.Y(n_1974)
);

AND2x4_ASAP7_75t_SL g1975 ( 
.A(n_1923),
.B(n_1840),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1885),
.B(n_1828),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1953),
.Y(n_1977)
);

HB1xp67_ASAP7_75t_L g1978 ( 
.A(n_1924),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1941),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1955),
.B(n_1878),
.Y(n_1980)
);

INVxp67_ASAP7_75t_L g1981 ( 
.A(n_1905),
.Y(n_1981)
);

AND2x4_ASAP7_75t_L g1982 ( 
.A(n_1928),
.B(n_1892),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1953),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1936),
.B(n_1878),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1938),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1913),
.B(n_1859),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1936),
.B(n_1864),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1918),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1921),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1882),
.B(n_1864),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1895),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1932),
.B(n_1864),
.Y(n_1992)
);

HB1xp67_ASAP7_75t_L g1993 ( 
.A(n_1932),
.Y(n_1993)
);

AND2x4_ASAP7_75t_L g1994 ( 
.A(n_1892),
.B(n_1834),
.Y(n_1994)
);

AND2x4_ASAP7_75t_L g1995 ( 
.A(n_1906),
.B(n_1834),
.Y(n_1995)
);

OR2x2_ASAP7_75t_L g1996 ( 
.A(n_1890),
.B(n_1846),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1922),
.Y(n_1997)
);

AND2x4_ASAP7_75t_L g1998 ( 
.A(n_1906),
.B(n_1852),
.Y(n_1998)
);

OR2x2_ASAP7_75t_L g1999 ( 
.A(n_1891),
.B(n_1846),
.Y(n_1999)
);

NOR2xp33_ASAP7_75t_L g2000 ( 
.A(n_1899),
.B(n_1934),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1942),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1944),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1960),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1937),
.B(n_1868),
.Y(n_2004)
);

AND2x4_ASAP7_75t_SL g2005 ( 
.A(n_1915),
.B(n_1840),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1948),
.B(n_1869),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1926),
.Y(n_2007)
);

INVx2_ASAP7_75t_L g2008 ( 
.A(n_1927),
.Y(n_2008)
);

NOR2xp33_ASAP7_75t_L g2009 ( 
.A(n_1910),
.B(n_1854),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1935),
.Y(n_2010)
);

OR2x2_ASAP7_75t_SL g2011 ( 
.A(n_1888),
.B(n_1824),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1943),
.B(n_1814),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1903),
.B(n_1877),
.Y(n_2013)
);

BUFx2_ASAP7_75t_L g2014 ( 
.A(n_1965),
.Y(n_2014)
);

NOR2xp33_ASAP7_75t_L g2015 ( 
.A(n_1910),
.B(n_1854),
.Y(n_2015)
);

NOR2xp33_ASAP7_75t_SL g2016 ( 
.A(n_1883),
.B(n_1832),
.Y(n_2016)
);

AND2x4_ASAP7_75t_L g2017 ( 
.A(n_1907),
.B(n_1929),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1917),
.B(n_1884),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1894),
.B(n_1877),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1959),
.Y(n_2020)
);

OR2x2_ASAP7_75t_L g2021 ( 
.A(n_1902),
.B(n_1824),
.Y(n_2021)
);

OR2x2_ASAP7_75t_L g2022 ( 
.A(n_1949),
.B(n_1828),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1943),
.B(n_1814),
.Y(n_2023)
);

HB1xp67_ASAP7_75t_L g2024 ( 
.A(n_1904),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1909),
.B(n_1814),
.Y(n_2025)
);

INVxp67_ASAP7_75t_L g2026 ( 
.A(n_1911),
.Y(n_2026)
);

OR2x2_ASAP7_75t_L g2027 ( 
.A(n_1956),
.B(n_1831),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1925),
.B(n_1835),
.Y(n_2028)
);

AND2x4_ASAP7_75t_L g2029 ( 
.A(n_1907),
.B(n_1852),
.Y(n_2029)
);

INVx6_ASAP7_75t_L g2030 ( 
.A(n_1963),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1962),
.Y(n_2031)
);

INVx1_ASAP7_75t_SL g2032 ( 
.A(n_1946),
.Y(n_2032)
);

INVxp67_ASAP7_75t_L g2033 ( 
.A(n_1886),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1939),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1968),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1974),
.Y(n_2036)
);

BUFx12f_ASAP7_75t_L g2037 ( 
.A(n_2030),
.Y(n_2037)
);

NOR2x1_ASAP7_75t_L g2038 ( 
.A(n_2000),
.B(n_2017),
.Y(n_2038)
);

HB1xp67_ASAP7_75t_L g2039 ( 
.A(n_2031),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1968),
.Y(n_2040)
);

INVx3_ASAP7_75t_R g2041 ( 
.A(n_2017),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_2020),
.B(n_1893),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1971),
.B(n_1912),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1974),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_2020),
.B(n_1897),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_1971),
.B(n_1950),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1972),
.Y(n_2047)
);

INVxp67_ASAP7_75t_L g2048 ( 
.A(n_1969),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_1966),
.B(n_1950),
.Y(n_2049)
);

INVxp67_ASAP7_75t_SL g2050 ( 
.A(n_2020),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1972),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1976),
.Y(n_2052)
);

OR2x2_ASAP7_75t_L g2053 ( 
.A(n_2031),
.B(n_1900),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_1974),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_1966),
.B(n_1952),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1976),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1988),
.B(n_1989),
.Y(n_2057)
);

AOI21xp5_ASAP7_75t_L g2058 ( 
.A1(n_2016),
.A2(n_1896),
.B(n_1898),
.Y(n_2058)
);

INVxp67_ASAP7_75t_SL g2059 ( 
.A(n_2033),
.Y(n_2059)
);

OR2x2_ASAP7_75t_L g2060 ( 
.A(n_1978),
.B(n_1988),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2007),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_1967),
.B(n_1930),
.Y(n_2062)
);

NAND2x1_ASAP7_75t_L g2063 ( 
.A(n_2017),
.B(n_1852),
.Y(n_2063)
);

AND2x4_ASAP7_75t_L g2064 ( 
.A(n_2005),
.B(n_1973),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1989),
.B(n_1931),
.Y(n_2065)
);

INVx3_ASAP7_75t_L g2066 ( 
.A(n_1994),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1979),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1979),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1985),
.Y(n_2069)
);

INVxp67_ASAP7_75t_L g2070 ( 
.A(n_2016),
.Y(n_2070)
);

OR2x2_ASAP7_75t_L g2071 ( 
.A(n_1997),
.B(n_1933),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_1997),
.B(n_1940),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1977),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_1977),
.Y(n_2074)
);

OR2x2_ASAP7_75t_L g2075 ( 
.A(n_2008),
.B(n_1946),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1985),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2008),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_2008),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_1977),
.Y(n_2079)
);

INVxp67_ASAP7_75t_SL g2080 ( 
.A(n_2017),
.Y(n_2080)
);

OR2x2_ASAP7_75t_L g2081 ( 
.A(n_2022),
.B(n_1964),
.Y(n_2081)
);

AND2x4_ASAP7_75t_L g2082 ( 
.A(n_2005),
.B(n_1908),
.Y(n_2082)
);

INVx2_ASAP7_75t_L g2083 ( 
.A(n_1983),
.Y(n_2083)
);

NOR2x1_ASAP7_75t_L g2084 ( 
.A(n_2007),
.B(n_2010),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_2010),
.B(n_1930),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_2026),
.B(n_1947),
.Y(n_2086)
);

OR2x2_ASAP7_75t_L g2087 ( 
.A(n_2022),
.B(n_1951),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1983),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_1983),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2027),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_2036),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2035),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_2038),
.B(n_1967),
.Y(n_2093)
);

NAND2x1p5_ASAP7_75t_L g2094 ( 
.A(n_2063),
.B(n_1980),
.Y(n_2094)
);

HB1xp67_ASAP7_75t_L g2095 ( 
.A(n_2071),
.Y(n_2095)
);

INVx2_ASAP7_75t_SL g2096 ( 
.A(n_2064),
.Y(n_2096)
);

OR2x2_ASAP7_75t_L g2097 ( 
.A(n_2060),
.B(n_2018),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_2043),
.B(n_2014),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_2043),
.B(n_2014),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2035),
.Y(n_2100)
);

INVx1_ASAP7_75t_SL g2101 ( 
.A(n_2042),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2050),
.B(n_1981),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_2039),
.B(n_2028),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2047),
.Y(n_2104)
);

NOR3xp33_ASAP7_75t_L g2105 ( 
.A(n_2048),
.B(n_2032),
.C(n_2034),
.Y(n_2105)
);

OR2x2_ASAP7_75t_L g2106 ( 
.A(n_2060),
.B(n_2027),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_2059),
.B(n_2032),
.Y(n_2107)
);

OR2x2_ASAP7_75t_L g2108 ( 
.A(n_2090),
.B(n_2057),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_2036),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2047),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_2045),
.B(n_2003),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2080),
.B(n_2012),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2051),
.Y(n_2113)
);

INVx4_ASAP7_75t_L g2114 ( 
.A(n_2037),
.Y(n_2114)
);

OR2x2_ASAP7_75t_L g2115 ( 
.A(n_2090),
.B(n_2003),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2051),
.Y(n_2116)
);

INVx2_ASAP7_75t_SL g2117 ( 
.A(n_2064),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_2065),
.B(n_2003),
.Y(n_2118)
);

INVxp67_ASAP7_75t_L g2119 ( 
.A(n_2053),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_2055),
.B(n_2012),
.Y(n_2120)
);

OR2x2_ASAP7_75t_L g2121 ( 
.A(n_2071),
.B(n_2081),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_2044),
.Y(n_2122)
);

OR2x2_ASAP7_75t_L g2123 ( 
.A(n_2081),
.B(n_1996),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_2044),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_2055),
.B(n_2023),
.Y(n_2125)
);

OR2x2_ASAP7_75t_L g2126 ( 
.A(n_2072),
.B(n_1996),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_2054),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_2062),
.B(n_2023),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_2086),
.B(n_1993),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2040),
.Y(n_2130)
);

HB1xp67_ASAP7_75t_L g2131 ( 
.A(n_2084),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_2054),
.Y(n_2132)
);

OAI21xp33_ASAP7_75t_L g2133 ( 
.A1(n_2053),
.A2(n_2013),
.B(n_2024),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_2073),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2067),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_2062),
.B(n_1980),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2067),
.Y(n_2137)
);

AOI22xp5_ASAP7_75t_L g2138 ( 
.A1(n_2058),
.A2(n_1887),
.B1(n_2034),
.B2(n_1975),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2064),
.B(n_1982),
.Y(n_2139)
);

NAND2x1_ASAP7_75t_L g2140 ( 
.A(n_2066),
.B(n_1982),
.Y(n_2140)
);

NOR2xp33_ASAP7_75t_L g2141 ( 
.A(n_2041),
.B(n_2009),
.Y(n_2141)
);

OAI21xp5_ASAP7_75t_SL g2142 ( 
.A1(n_2066),
.A2(n_2070),
.B(n_1945),
.Y(n_2142)
);

NOR2xp67_ASAP7_75t_L g2143 ( 
.A(n_2066),
.B(n_1982),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2068),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_2073),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_2061),
.B(n_2085),
.Y(n_2146)
);

OR2x2_ASAP7_75t_L g2147 ( 
.A(n_2106),
.B(n_2052),
.Y(n_2147)
);

NOR2x1_ASAP7_75t_R g2148 ( 
.A(n_2114),
.B(n_2037),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_2128),
.B(n_2049),
.Y(n_2149)
);

CKINVDCx16_ASAP7_75t_R g2150 ( 
.A(n_2114),
.Y(n_2150)
);

NAND2x1_ASAP7_75t_L g2151 ( 
.A(n_2139),
.B(n_2082),
.Y(n_2151)
);

AND2x4_ASAP7_75t_SL g2152 ( 
.A(n_2114),
.B(n_2082),
.Y(n_2152)
);

AOI22xp33_ASAP7_75t_L g2153 ( 
.A1(n_2105),
.A2(n_2121),
.B1(n_2119),
.B2(n_2034),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_2112),
.Y(n_2154)
);

HB1xp67_ASAP7_75t_L g2155 ( 
.A(n_2095),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2130),
.Y(n_2156)
);

INVx3_ASAP7_75t_SL g2157 ( 
.A(n_2096),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_2128),
.B(n_2049),
.Y(n_2158)
);

CKINVDCx16_ASAP7_75t_R g2159 ( 
.A(n_2121),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_2120),
.B(n_2063),
.Y(n_2160)
);

AOI21xp5_ASAP7_75t_L g2161 ( 
.A1(n_2103),
.A2(n_2087),
.B(n_2082),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2130),
.Y(n_2162)
);

OR2x2_ASAP7_75t_L g2163 ( 
.A(n_2106),
.B(n_2052),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2104),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_2112),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2104),
.Y(n_2166)
);

AND2x4_ASAP7_75t_L g2167 ( 
.A(n_2096),
.B(n_2056),
.Y(n_2167)
);

OR2x2_ASAP7_75t_L g2168 ( 
.A(n_2097),
.B(n_2056),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_2091),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_2101),
.B(n_2068),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_2120),
.B(n_2046),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2110),
.Y(n_2172)
);

AOI21xp5_ASAP7_75t_SL g2173 ( 
.A1(n_2107),
.A2(n_2041),
.B(n_1634),
.Y(n_2173)
);

OR2x2_ASAP7_75t_L g2174 ( 
.A(n_2097),
.B(n_2069),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2110),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2113),
.Y(n_2176)
);

INVx1_ASAP7_75t_SL g2177 ( 
.A(n_2117),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2113),
.Y(n_2178)
);

OR2x2_ASAP7_75t_L g2179 ( 
.A(n_2126),
.B(n_2069),
.Y(n_2179)
);

INVx1_ASAP7_75t_SL g2180 ( 
.A(n_2117),
.Y(n_2180)
);

OR2x2_ASAP7_75t_L g2181 ( 
.A(n_2126),
.B(n_2076),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2116),
.Y(n_2182)
);

CKINVDCx16_ASAP7_75t_R g2183 ( 
.A(n_2098),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_2146),
.B(n_2076),
.Y(n_2184)
);

AND2x4_ASAP7_75t_L g2185 ( 
.A(n_2093),
.B(n_2005),
.Y(n_2185)
);

INVxp67_ASAP7_75t_SL g2186 ( 
.A(n_2131),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2125),
.B(n_2046),
.Y(n_2187)
);

INVx2_ASAP7_75t_SL g2188 ( 
.A(n_2139),
.Y(n_2188)
);

OAI321xp33_ASAP7_75t_L g2189 ( 
.A1(n_2153),
.A2(n_2138),
.A3(n_2111),
.B1(n_2133),
.B2(n_2141),
.C(n_2102),
.Y(n_2189)
);

NOR2xp67_ASAP7_75t_SL g2190 ( 
.A(n_2150),
.B(n_2030),
.Y(n_2190)
);

AND2x2_ASAP7_75t_L g2191 ( 
.A(n_2183),
.B(n_2125),
.Y(n_2191)
);

OR2x2_ASAP7_75t_L g2192 ( 
.A(n_2159),
.B(n_2154),
.Y(n_2192)
);

OAI332xp33_ASAP7_75t_L g2193 ( 
.A1(n_2186),
.A2(n_2123),
.A3(n_2087),
.B1(n_2129),
.B2(n_2118),
.B3(n_2108),
.C1(n_2122),
.C2(n_2132),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_SL g2194 ( 
.A(n_2185),
.B(n_2143),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_2155),
.B(n_2154),
.Y(n_2195)
);

OAI22xp33_ASAP7_75t_L g2196 ( 
.A1(n_2161),
.A2(n_2123),
.B1(n_2142),
.B2(n_2098),
.Y(n_2196)
);

NAND3xp33_ASAP7_75t_L g2197 ( 
.A(n_2170),
.B(n_2137),
.C(n_2135),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2164),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2166),
.Y(n_2199)
);

NOR3xp33_ASAP7_75t_L g2200 ( 
.A(n_2177),
.B(n_2099),
.C(n_2135),
.Y(n_2200)
);

OAI222xp33_ASAP7_75t_L g2201 ( 
.A1(n_2184),
.A2(n_2099),
.B1(n_2136),
.B2(n_2091),
.C1(n_2134),
.C2(n_2109),
.Y(n_2201)
);

AO21x1_ASAP7_75t_L g2202 ( 
.A1(n_2152),
.A2(n_2140),
.B(n_2137),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_2165),
.B(n_2136),
.Y(n_2203)
);

INVxp67_ASAP7_75t_L g2204 ( 
.A(n_2148),
.Y(n_2204)
);

NAND3xp33_ASAP7_75t_L g2205 ( 
.A(n_2167),
.B(n_2144),
.C(n_2108),
.Y(n_2205)
);

NAND2x1_ASAP7_75t_L g2206 ( 
.A(n_2160),
.B(n_2185),
.Y(n_2206)
);

A2O1A1Ixp33_ASAP7_75t_L g2207 ( 
.A1(n_2152),
.A2(n_2093),
.B(n_2140),
.C(n_2089),
.Y(n_2207)
);

OR2x2_ASAP7_75t_L g2208 ( 
.A(n_2165),
.B(n_2092),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_2149),
.B(n_2100),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_2149),
.B(n_2158),
.Y(n_2210)
);

OAI21xp5_ASAP7_75t_L g2211 ( 
.A1(n_2180),
.A2(n_2167),
.B(n_2188),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_2158),
.Y(n_2212)
);

AOI22xp5_ASAP7_75t_SL g2213 ( 
.A1(n_2185),
.A2(n_2094),
.B1(n_1919),
.B2(n_2144),
.Y(n_2213)
);

NOR2x1_ASAP7_75t_L g2214 ( 
.A(n_2151),
.B(n_2116),
.Y(n_2214)
);

OR2x2_ASAP7_75t_L g2215 ( 
.A(n_2179),
.B(n_2181),
.Y(n_2215)
);

AOI22xp33_ASAP7_75t_L g2216 ( 
.A1(n_2169),
.A2(n_2145),
.B1(n_2134),
.B2(n_2132),
.Y(n_2216)
);

OAI21xp33_ASAP7_75t_SL g2217 ( 
.A1(n_2160),
.A2(n_1970),
.B(n_2015),
.Y(n_2217)
);

AOI311xp33_ASAP7_75t_L g2218 ( 
.A1(n_2156),
.A2(n_2019),
.A3(n_1954),
.B(n_2094),
.C(n_1992),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2172),
.Y(n_2219)
);

AOI22xp5_ASAP7_75t_L g2220 ( 
.A1(n_2196),
.A2(n_2188),
.B1(n_2169),
.B2(n_2157),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2215),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_2191),
.B(n_2171),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_2210),
.B(n_2171),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2208),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2203),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2209),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_2212),
.B(n_2187),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2195),
.Y(n_2228)
);

AOI22xp33_ASAP7_75t_L g2229 ( 
.A1(n_2196),
.A2(n_2122),
.B1(n_2109),
.B2(n_2124),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2198),
.Y(n_2230)
);

INVxp67_ASAP7_75t_L g2231 ( 
.A(n_2192),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2193),
.B(n_2187),
.Y(n_2232)
);

AND2x2_ASAP7_75t_L g2233 ( 
.A(n_2211),
.B(n_2157),
.Y(n_2233)
);

NOR2xp33_ASAP7_75t_L g2234 ( 
.A(n_2204),
.B(n_2179),
.Y(n_2234)
);

NOR2xp33_ASAP7_75t_L g2235 ( 
.A(n_2204),
.B(n_2181),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2199),
.Y(n_2236)
);

AND2x4_ASAP7_75t_SL g2237 ( 
.A(n_2200),
.B(n_2167),
.Y(n_2237)
);

INVx2_ASAP7_75t_L g2238 ( 
.A(n_2214),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2219),
.Y(n_2239)
);

INVx1_ASAP7_75t_SL g2240 ( 
.A(n_2206),
.Y(n_2240)
);

NOR2xp33_ASAP7_75t_L g2241 ( 
.A(n_2201),
.B(n_2174),
.Y(n_2241)
);

AOI22xp33_ASAP7_75t_SL g2242 ( 
.A1(n_2213),
.A2(n_2162),
.B1(n_2178),
.B2(n_2176),
.Y(n_2242)
);

HB1xp67_ASAP7_75t_L g2243 ( 
.A(n_2200),
.Y(n_2243)
);

A2O1A1Ixp33_ASAP7_75t_L g2244 ( 
.A1(n_2241),
.A2(n_2189),
.B(n_2205),
.C(n_2197),
.Y(n_2244)
);

HB1xp67_ASAP7_75t_L g2245 ( 
.A(n_2222),
.Y(n_2245)
);

AOI221xp5_ASAP7_75t_L g2246 ( 
.A1(n_2241),
.A2(n_2201),
.B1(n_2216),
.B2(n_2202),
.C(n_2207),
.Y(n_2246)
);

OAI21xp33_ASAP7_75t_L g2247 ( 
.A1(n_2232),
.A2(n_2194),
.B(n_2217),
.Y(n_2247)
);

AOI322xp5_ASAP7_75t_L g2248 ( 
.A1(n_2243),
.A2(n_2218),
.A3(n_2124),
.B1(n_2127),
.B2(n_2145),
.C1(n_2074),
.C2(n_2079),
.Y(n_2248)
);

AOI32xp33_ASAP7_75t_L g2249 ( 
.A1(n_2229),
.A2(n_2182),
.A3(n_2175),
.B1(n_2174),
.B2(n_2168),
.Y(n_2249)
);

OAI21xp5_ASAP7_75t_SL g2250 ( 
.A1(n_2220),
.A2(n_2094),
.B(n_2147),
.Y(n_2250)
);

O2A1O1Ixp5_ASAP7_75t_L g2251 ( 
.A1(n_2238),
.A2(n_2190),
.B(n_2147),
.C(n_2163),
.Y(n_2251)
);

O2A1O1Ixp33_ASAP7_75t_L g2252 ( 
.A1(n_2238),
.A2(n_2168),
.B(n_2163),
.C(n_2127),
.Y(n_2252)
);

AOI21xp5_ASAP7_75t_L g2253 ( 
.A1(n_2237),
.A2(n_2173),
.B(n_2079),
.Y(n_2253)
);

OR2x2_ASAP7_75t_L g2254 ( 
.A(n_2223),
.B(n_2227),
.Y(n_2254)
);

AOI21xp33_ASAP7_75t_SL g2255 ( 
.A1(n_2234),
.A2(n_2115),
.B(n_2075),
.Y(n_2255)
);

OAI21xp5_ASAP7_75t_SL g2256 ( 
.A1(n_2242),
.A2(n_1973),
.B(n_1994),
.Y(n_2256)
);

A2O1A1Ixp33_ASAP7_75t_L g2257 ( 
.A1(n_2237),
.A2(n_2089),
.B(n_2088),
.C(n_2083),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_SL g2258 ( 
.A(n_2222),
.B(n_2115),
.Y(n_2258)
);

AOI22xp5_ASAP7_75t_L g2259 ( 
.A1(n_2234),
.A2(n_2074),
.B1(n_2083),
.B2(n_2088),
.Y(n_2259)
);

OAI322xp33_ASAP7_75t_L g2260 ( 
.A1(n_2255),
.A2(n_2235),
.A3(n_2231),
.B1(n_2228),
.B2(n_2221),
.C1(n_2224),
.C2(n_2226),
.Y(n_2260)
);

NAND4xp75_ASAP7_75t_L g2261 ( 
.A(n_2246),
.B(n_2235),
.C(n_2233),
.D(n_2225),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2245),
.Y(n_2262)
);

OAI21x1_ASAP7_75t_SL g2263 ( 
.A1(n_2252),
.A2(n_2236),
.B(n_2230),
.Y(n_2263)
);

AOI21xp33_ASAP7_75t_L g2264 ( 
.A1(n_2244),
.A2(n_2247),
.B(n_2251),
.Y(n_2264)
);

AOI21xp5_ASAP7_75t_L g2265 ( 
.A1(n_2253),
.A2(n_2250),
.B(n_2258),
.Y(n_2265)
);

NOR3x1_ASAP7_75t_L g2266 ( 
.A(n_2254),
.B(n_2239),
.C(n_2240),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_2259),
.Y(n_2267)
);

NAND4xp75_ASAP7_75t_L g2268 ( 
.A(n_2248),
.B(n_2233),
.C(n_2173),
.D(n_2078),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_2249),
.B(n_2075),
.Y(n_2269)
);

NOR2xp33_ASAP7_75t_L g2270 ( 
.A(n_2256),
.B(n_2030),
.Y(n_2270)
);

NOR3xp33_ASAP7_75t_L g2271 ( 
.A(n_2257),
.B(n_2078),
.C(n_2077),
.Y(n_2271)
);

OA22x2_ASAP7_75t_L g2272 ( 
.A1(n_2250),
.A2(n_1973),
.B1(n_1998),
.B2(n_2029),
.Y(n_2272)
);

NAND3xp33_ASAP7_75t_L g2273 ( 
.A(n_2264),
.B(n_2077),
.C(n_1957),
.Y(n_2273)
);

NAND4xp25_ASAP7_75t_SL g2274 ( 
.A(n_2265),
.B(n_1984),
.C(n_1987),
.D(n_2030),
.Y(n_2274)
);

AOI221xp5_ASAP7_75t_L g2275 ( 
.A1(n_2263),
.A2(n_1951),
.B1(n_2001),
.B2(n_2002),
.C(n_2011),
.Y(n_2275)
);

AND2x2_ASAP7_75t_L g2276 ( 
.A(n_2266),
.B(n_1970),
.Y(n_2276)
);

OAI21xp33_ASAP7_75t_L g2277 ( 
.A1(n_2270),
.A2(n_1995),
.B(n_1994),
.Y(n_2277)
);

AOI211xp5_ASAP7_75t_L g2278 ( 
.A1(n_2260),
.A2(n_1880),
.B(n_1994),
.C(n_2029),
.Y(n_2278)
);

AOI221xp5_ASAP7_75t_L g2279 ( 
.A1(n_2269),
.A2(n_2002),
.B1(n_2001),
.B2(n_2011),
.C(n_1986),
.Y(n_2279)
);

NOR2x1_ASAP7_75t_L g2280 ( 
.A(n_2261),
.B(n_1982),
.Y(n_2280)
);

AOI22xp5_ASAP7_75t_L g2281 ( 
.A1(n_2276),
.A2(n_2268),
.B1(n_2267),
.B2(n_2272),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2280),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_SL g2283 ( 
.A(n_2273),
.B(n_2262),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_2274),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2278),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2279),
.Y(n_2286)
);

OAI22xp5_ASAP7_75t_L g2287 ( 
.A1(n_2277),
.A2(n_2266),
.B1(n_2271),
.B2(n_2030),
.Y(n_2287)
);

AOI22xp5_ASAP7_75t_L g2288 ( 
.A1(n_2275),
.A2(n_1975),
.B1(n_2029),
.B2(n_1995),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2282),
.Y(n_2289)
);

OAI21xp33_ASAP7_75t_SL g2290 ( 
.A1(n_2283),
.A2(n_1984),
.B(n_2004),
.Y(n_2290)
);

AOI22xp5_ASAP7_75t_L g2291 ( 
.A1(n_2281),
.A2(n_2029),
.B1(n_1998),
.B2(n_1995),
.Y(n_2291)
);

NAND4xp75_ASAP7_75t_L g2292 ( 
.A(n_2285),
.B(n_1901),
.C(n_1854),
.D(n_1990),
.Y(n_2292)
);

NOR3xp33_ASAP7_75t_L g2293 ( 
.A(n_2286),
.B(n_2002),
.C(n_2001),
.Y(n_2293)
);

AND2x4_ASAP7_75t_L g2294 ( 
.A(n_2284),
.B(n_1973),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2289),
.Y(n_2295)
);

AND2x4_ASAP7_75t_L g2296 ( 
.A(n_2294),
.B(n_2288),
.Y(n_2296)
);

INVxp67_ASAP7_75t_L g2297 ( 
.A(n_2292),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2290),
.Y(n_2298)
);

AOI22xp5_ASAP7_75t_L g2299 ( 
.A1(n_2297),
.A2(n_2287),
.B1(n_2291),
.B2(n_2293),
.Y(n_2299)
);

OAI322xp33_ASAP7_75t_L g2300 ( 
.A1(n_2299),
.A2(n_2298),
.A3(n_2295),
.B1(n_2296),
.B2(n_2021),
.C1(n_1999),
.C2(n_1857),
.Y(n_2300)
);

INVx2_ASAP7_75t_SL g2301 ( 
.A(n_2300),
.Y(n_2301)
);

AO22x1_ASAP7_75t_L g2302 ( 
.A1(n_2300),
.A2(n_2296),
.B1(n_1998),
.B2(n_1995),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_2302),
.Y(n_2303)
);

AND2x4_ASAP7_75t_L g2304 ( 
.A(n_2301),
.B(n_1991),
.Y(n_2304)
);

AOI21xp33_ASAP7_75t_L g2305 ( 
.A1(n_2303),
.A2(n_1810),
.B(n_1781),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2304),
.B(n_1810),
.Y(n_2306)
);

NAND2x1p5_ASAP7_75t_SL g2307 ( 
.A(n_2305),
.B(n_1876),
.Y(n_2307)
);

AOI22xp33_ASAP7_75t_L g2308 ( 
.A1(n_2307),
.A2(n_2306),
.B1(n_1876),
.B2(n_1975),
.Y(n_2308)
);

AOI221xp5_ASAP7_75t_L g2309 ( 
.A1(n_2308),
.A2(n_2025),
.B1(n_1998),
.B2(n_2006),
.C(n_1987),
.Y(n_2309)
);

AOI211xp5_ASAP7_75t_L g2310 ( 
.A1(n_2309),
.A2(n_1999),
.B(n_2021),
.C(n_2025),
.Y(n_2310)
);


endmodule