module real_aes_6358_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_314;
wire n_252;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_359;
wire n_156;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_0), .B(n_112), .C(n_113), .Y(n_111) );
INVx1_ASAP7_75t_L g451 ( .A(n_0), .Y(n_451) );
INVx1_ASAP7_75t_L g544 ( .A(n_1), .Y(n_544) );
INVx1_ASAP7_75t_L g158 ( .A(n_2), .Y(n_158) );
AOI222xp33_ASAP7_75t_L g457 ( .A1(n_3), .A2(n_458), .B1(n_742), .B2(n_743), .C1(n_752), .C2(n_754), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_4), .A2(n_39), .B1(n_183), .B2(n_490), .Y(n_513) );
AOI21xp33_ASAP7_75t_L g190 ( .A1(n_5), .A2(n_174), .B(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_6), .B(n_172), .Y(n_556) );
AND2x6_ASAP7_75t_L g151 ( .A(n_7), .B(n_152), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_8), .A2(n_261), .B(n_262), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_9), .B(n_110), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_9), .B(n_40), .Y(n_452) );
INVx1_ASAP7_75t_L g196 ( .A(n_10), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_11), .B(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g143 ( .A(n_12), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_13), .B(n_164), .Y(n_499) );
INVx1_ASAP7_75t_L g267 ( .A(n_14), .Y(n_267) );
INVx1_ASAP7_75t_L g538 ( .A(n_15), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_16), .B(n_139), .Y(n_527) );
AO32x2_ASAP7_75t_L g511 ( .A1(n_17), .A2(n_138), .A3(n_172), .B1(n_492), .B2(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_18), .B(n_183), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_19), .B(n_179), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_20), .B(n_139), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_21), .A2(n_50), .B1(n_183), .B2(n_490), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_22), .B(n_174), .Y(n_224) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_23), .A2(n_100), .B1(n_749), .B2(n_750), .Y(n_748) );
INVx1_ASAP7_75t_L g750 ( .A(n_23), .Y(n_750) );
AOI22xp33_ASAP7_75t_SL g491 ( .A1(n_24), .A2(n_77), .B1(n_164), .B2(n_183), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_25), .B(n_183), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_26), .B(n_186), .Y(n_185) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_27), .A2(n_265), .B(n_266), .C(n_268), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_28), .B(n_454), .Y(n_453) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_29), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_30), .B(n_169), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_31), .B(n_162), .Y(n_161) );
OAI22xp5_ASAP7_75t_SL g128 ( .A1(n_32), .A2(n_90), .B1(n_129), .B2(n_130), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_32), .Y(n_129) );
INVx1_ASAP7_75t_L g211 ( .A(n_33), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_34), .B(n_169), .Y(n_483) );
INVx2_ASAP7_75t_L g149 ( .A(n_35), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_36), .B(n_183), .Y(n_560) );
OAI22xp5_ASAP7_75t_SL g124 ( .A1(n_37), .A2(n_70), .B1(n_125), .B2(n_126), .Y(n_124) );
CKINVDCx16_ASAP7_75t_R g125 ( .A(n_37), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_37), .B(n_169), .Y(n_504) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_38), .A2(n_151), .B(n_154), .C(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g110 ( .A(n_40), .Y(n_110) );
INVx1_ASAP7_75t_L g209 ( .A(n_41), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_42), .B(n_162), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_43), .B(n_183), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_44), .A2(n_88), .B1(n_231), .B2(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_45), .B(n_183), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_46), .B(n_183), .Y(n_539) );
CKINVDCx16_ASAP7_75t_R g212 ( .A(n_47), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_48), .B(n_543), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_49), .B(n_174), .Y(n_255) );
AOI22xp33_ASAP7_75t_SL g531 ( .A1(n_51), .A2(n_62), .B1(n_164), .B2(n_183), .Y(n_531) );
OAI22xp5_ASAP7_75t_SL g746 ( .A1(n_52), .A2(n_747), .B1(n_748), .B2(n_751), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_52), .Y(n_751) );
AOI22xp5_ASAP7_75t_L g206 ( .A1(n_53), .A2(n_154), .B1(n_164), .B2(n_207), .Y(n_206) );
CKINVDCx20_ASAP7_75t_R g234 ( .A(n_54), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_55), .B(n_183), .Y(n_498) );
CKINVDCx16_ASAP7_75t_R g145 ( .A(n_56), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_57), .B(n_183), .Y(n_564) );
A2O1A1Ixp33_ASAP7_75t_L g193 ( .A1(n_58), .A2(n_182), .B(n_194), .C(n_195), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g244 ( .A(n_59), .Y(n_244) );
INVx1_ASAP7_75t_L g192 ( .A(n_60), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_61), .A2(n_105), .B1(n_116), .B2(n_758), .Y(n_104) );
INVx1_ASAP7_75t_L g152 ( .A(n_63), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_64), .B(n_183), .Y(n_545) );
INVx1_ASAP7_75t_L g142 ( .A(n_65), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_66), .Y(n_121) );
AO32x2_ASAP7_75t_L g487 ( .A1(n_67), .A2(n_172), .A3(n_247), .B1(n_488), .B2(n_492), .Y(n_487) );
INVx1_ASAP7_75t_L g563 ( .A(n_68), .Y(n_563) );
INVx1_ASAP7_75t_L g478 ( .A(n_69), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_70), .Y(n_126) );
A2O1A1Ixp33_ASAP7_75t_SL g178 ( .A1(n_71), .A2(n_179), .B(n_180), .C(n_182), .Y(n_178) );
INVxp67_ASAP7_75t_L g181 ( .A(n_72), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_73), .B(n_164), .Y(n_479) );
INVx1_ASAP7_75t_L g115 ( .A(n_74), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g214 ( .A(n_75), .Y(n_214) );
INVx1_ASAP7_75t_L g237 ( .A(n_76), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_78), .A2(n_151), .B(n_154), .C(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_79), .B(n_490), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_80), .B(n_164), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_81), .A2(n_744), .B1(n_745), .B2(n_746), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_81), .Y(n_744) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_82), .B(n_159), .Y(n_227) );
INVx2_ASAP7_75t_L g140 ( .A(n_83), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_84), .B(n_179), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_85), .B(n_164), .Y(n_552) );
A2O1A1Ixp33_ASAP7_75t_L g153 ( .A1(n_86), .A2(n_151), .B(n_154), .C(n_157), .Y(n_153) );
INVx2_ASAP7_75t_L g112 ( .A(n_87), .Y(n_112) );
OR2x2_ASAP7_75t_L g448 ( .A(n_87), .B(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g461 ( .A(n_87), .B(n_450), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_89), .A2(n_103), .B1(n_164), .B2(n_165), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_90), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_91), .B(n_169), .Y(n_197) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_92), .Y(n_167) );
A2O1A1Ixp33_ASAP7_75t_L g249 ( .A1(n_93), .A2(n_151), .B(n_154), .C(n_250), .Y(n_249) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_94), .Y(n_257) );
INVx1_ASAP7_75t_L g177 ( .A(n_95), .Y(n_177) );
CKINVDCx16_ASAP7_75t_R g263 ( .A(n_96), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_97), .B(n_159), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_98), .B(n_164), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_99), .B(n_172), .Y(n_269) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_100), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_101), .B(n_115), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_102), .A2(n_174), .B(n_175), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx12_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_SL g759 ( .A(n_108), .Y(n_759) );
OR2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
OR2x2_ASAP7_75t_L g465 ( .A(n_112), .B(n_450), .Y(n_465) );
NOR2x2_ASAP7_75t_L g756 ( .A(n_112), .B(n_449), .Y(n_756) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
AO21x1_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_122), .B(n_456), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_SL g757 ( .A(n_120), .Y(n_757) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI21xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_445), .B(n_453), .Y(n_122) );
AOI22xp33_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_127), .B1(n_443), .B2(n_444), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_124), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_127), .Y(n_444) );
XNOR2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_131), .Y(n_127) );
INVx1_ASAP7_75t_L g462 ( .A(n_131), .Y(n_462) );
OAI22xp5_ASAP7_75t_SL g752 ( .A1(n_131), .A2(n_463), .B1(n_467), .B2(n_753), .Y(n_752) );
NAND2x1_ASAP7_75t_L g131 ( .A(n_132), .B(n_359), .Y(n_131) );
NOR5xp2_ASAP7_75t_L g132 ( .A(n_133), .B(n_282), .C(n_314), .D(n_329), .E(n_346), .Y(n_132) );
A2O1A1Ixp33_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_198), .B(n_219), .C(n_270), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_170), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_135), .B(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_135), .B(n_334), .Y(n_397) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_136), .B(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_136), .B(n_216), .Y(n_283) );
AND2x2_ASAP7_75t_L g324 ( .A(n_136), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_136), .B(n_293), .Y(n_328) );
OR2x2_ASAP7_75t_L g365 ( .A(n_136), .B(n_204), .Y(n_365) );
INVx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g203 ( .A(n_137), .B(n_204), .Y(n_203) );
INVx3_ASAP7_75t_L g273 ( .A(n_137), .Y(n_273) );
OR2x2_ASAP7_75t_L g436 ( .A(n_137), .B(n_276), .Y(n_436) );
AO21x2_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_144), .B(n_166), .Y(n_137) );
AO21x2_ASAP7_75t_L g204 ( .A1(n_138), .A2(n_205), .B(n_213), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_138), .B(n_214), .Y(n_213) );
INVx2_ASAP7_75t_L g232 ( .A(n_138), .Y(n_232) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_139), .Y(n_172) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x2_ASAP7_75t_SL g169 ( .A(n_140), .B(n_141), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
OAI21xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_146), .B(n_153), .Y(n_144) );
OAI22xp33_ASAP7_75t_L g205 ( .A1(n_146), .A2(n_184), .B1(n_206), .B2(n_212), .Y(n_205) );
OAI21xp5_ASAP7_75t_L g236 ( .A1(n_146), .A2(n_237), .B(n_238), .Y(n_236) );
NAND2x1p5_ASAP7_75t_L g146 ( .A(n_147), .B(n_151), .Y(n_146) );
AND2x4_ASAP7_75t_L g174 ( .A(n_147), .B(n_151), .Y(n_174) );
AND2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_150), .Y(n_147) );
INVx1_ASAP7_75t_L g543 ( .A(n_148), .Y(n_543) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g155 ( .A(n_149), .Y(n_155) );
INVx1_ASAP7_75t_L g165 ( .A(n_149), .Y(n_165) );
INVx1_ASAP7_75t_L g156 ( .A(n_150), .Y(n_156) );
INVx3_ASAP7_75t_L g160 ( .A(n_150), .Y(n_160) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_150), .Y(n_162) );
INVx1_ASAP7_75t_L g179 ( .A(n_150), .Y(n_179) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_150), .Y(n_208) );
INVx4_ASAP7_75t_SL g184 ( .A(n_151), .Y(n_184) );
OAI21xp5_ASAP7_75t_L g476 ( .A1(n_151), .A2(n_477), .B(n_480), .Y(n_476) );
BUFx3_ASAP7_75t_L g492 ( .A(n_151), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g496 ( .A1(n_151), .A2(n_497), .B(n_501), .Y(n_496) );
OAI21xp5_ASAP7_75t_L g536 ( .A1(n_151), .A2(n_537), .B(n_541), .Y(n_536) );
OAI21xp5_ASAP7_75t_L g549 ( .A1(n_151), .A2(n_550), .B(n_553), .Y(n_549) );
INVx5_ASAP7_75t_L g176 ( .A(n_154), .Y(n_176) );
AND2x6_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_155), .Y(n_183) );
BUFx3_ASAP7_75t_L g231 ( .A(n_155), .Y(n_231) );
INVx1_ASAP7_75t_L g490 ( .A(n_155), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_159), .B(n_161), .C(n_163), .Y(n_157) );
O2A1O1Ixp5_ASAP7_75t_SL g477 ( .A1(n_159), .A2(n_182), .B(n_478), .C(n_479), .Y(n_477) );
INVx2_ASAP7_75t_L g514 ( .A(n_159), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_159), .A2(n_551), .B(n_552), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_159), .A2(n_560), .B(n_561), .Y(n_559) );
INVx5_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_160), .B(n_181), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_160), .B(n_196), .Y(n_195) );
OAI22xp5_ASAP7_75t_SL g488 ( .A1(n_160), .A2(n_162), .B1(n_489), .B2(n_491), .Y(n_488) );
INVx2_ASAP7_75t_L g194 ( .A(n_162), .Y(n_194) );
INVx4_ASAP7_75t_L g253 ( .A(n_162), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_162), .A2(n_513), .B1(n_514), .B2(n_515), .Y(n_512) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_162), .A2(n_514), .B1(n_530), .B2(n_531), .Y(n_529) );
O2A1O1Ixp33_ASAP7_75t_L g537 ( .A1(n_163), .A2(n_538), .B(n_539), .C(n_540), .Y(n_537) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_168), .B(n_244), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_168), .B(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g247 ( .A(n_169), .Y(n_247) );
OA21x2_ASAP7_75t_L g259 ( .A1(n_169), .A2(n_260), .B(n_269), .Y(n_259) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_169), .A2(n_476), .B(n_483), .Y(n_475) );
OA21x2_ASAP7_75t_L g495 ( .A1(n_169), .A2(n_496), .B(n_504), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g338 ( .A1(n_170), .A2(n_339), .B1(n_340), .B2(n_343), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_170), .B(n_273), .Y(n_422) );
AND2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_188), .Y(n_170) );
AND2x2_ASAP7_75t_L g218 ( .A(n_171), .B(n_204), .Y(n_218) );
AND2x2_ASAP7_75t_L g275 ( .A(n_171), .B(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g280 ( .A(n_171), .Y(n_280) );
INVx3_ASAP7_75t_L g293 ( .A(n_171), .Y(n_293) );
OR2x2_ASAP7_75t_L g313 ( .A(n_171), .B(n_276), .Y(n_313) );
AND2x2_ASAP7_75t_L g332 ( .A(n_171), .B(n_189), .Y(n_332) );
BUFx2_ASAP7_75t_L g364 ( .A(n_171), .Y(n_364) );
OA21x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_185), .Y(n_171) );
INVx4_ASAP7_75t_L g187 ( .A(n_172), .Y(n_187) );
OA21x2_ASAP7_75t_L g548 ( .A1(n_172), .A2(n_549), .B(n_556), .Y(n_548) );
BUFx2_ASAP7_75t_L g261 ( .A(n_174), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_178), .C(n_184), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_L g191 ( .A1(n_176), .A2(n_184), .B(n_192), .C(n_193), .Y(n_191) );
O2A1O1Ixp33_ASAP7_75t_L g262 ( .A1(n_176), .A2(n_184), .B(n_263), .C(n_264), .Y(n_262) );
INVx1_ASAP7_75t_L g500 ( .A(n_179), .Y(n_500) );
INVx3_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_183), .Y(n_254) );
OA21x2_ASAP7_75t_L g189 ( .A1(n_186), .A2(n_190), .B(n_197), .Y(n_189) );
INVx3_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NOR2xp33_ASAP7_75t_SL g233 ( .A(n_187), .B(n_234), .Y(n_233) );
NAND3xp33_ASAP7_75t_L g528 ( .A(n_187), .B(n_492), .C(n_529), .Y(n_528) );
AO21x1_ASAP7_75t_L g618 ( .A1(n_187), .A2(n_529), .B(n_619), .Y(n_618) );
AND2x4_ASAP7_75t_L g279 ( .A(n_188), .B(n_280), .Y(n_279) );
INVx1_ASAP7_75t_SL g188 ( .A(n_189), .Y(n_188) );
BUFx2_ASAP7_75t_L g202 ( .A(n_189), .Y(n_202) );
INVx2_ASAP7_75t_L g217 ( .A(n_189), .Y(n_217) );
OR2x2_ASAP7_75t_L g295 ( .A(n_189), .B(n_276), .Y(n_295) );
AND2x2_ASAP7_75t_L g325 ( .A(n_189), .B(n_204), .Y(n_325) );
AND2x2_ASAP7_75t_L g342 ( .A(n_189), .B(n_273), .Y(n_342) );
AND2x2_ASAP7_75t_L g382 ( .A(n_189), .B(n_293), .Y(n_382) );
AND2x2_ASAP7_75t_SL g418 ( .A(n_189), .B(n_218), .Y(n_418) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_194), .A2(n_502), .B(n_503), .Y(n_501) );
O2A1O1Ixp5_ASAP7_75t_L g562 ( .A1(n_194), .A2(n_542), .B(n_563), .C(n_564), .Y(n_562) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NAND2xp33_ASAP7_75t_SL g199 ( .A(n_200), .B(n_215), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_201), .B(n_203), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_201), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g201 ( .A(n_202), .Y(n_201) );
OAI21xp33_ASAP7_75t_L g356 ( .A1(n_202), .A2(n_218), .B(n_357), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_202), .B(n_204), .Y(n_412) );
AND2x2_ASAP7_75t_L g348 ( .A(n_203), .B(n_349), .Y(n_348) );
INVx3_ASAP7_75t_L g276 ( .A(n_204), .Y(n_276) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_204), .Y(n_374) );
OAI22xp5_ASAP7_75t_SL g207 ( .A1(n_208), .A2(n_209), .B1(n_210), .B2(n_211), .Y(n_207) );
INVx2_ASAP7_75t_L g210 ( .A(n_208), .Y(n_210) );
INVx4_ASAP7_75t_L g265 ( .A(n_208), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_215), .B(n_273), .Y(n_441) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_216), .A2(n_384), .B1(n_385), .B2(n_390), .Y(n_383) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
AND2x2_ASAP7_75t_L g274 ( .A(n_217), .B(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g312 ( .A(n_217), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_SL g349 ( .A(n_217), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_218), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g403 ( .A(n_218), .Y(n_403) );
CKINVDCx16_ASAP7_75t_R g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_245), .Y(n_220) );
INVx4_ASAP7_75t_L g289 ( .A(n_221), .Y(n_289) );
AND2x2_ASAP7_75t_L g367 ( .A(n_221), .B(n_334), .Y(n_367) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_235), .Y(n_221) );
INVx3_ASAP7_75t_L g286 ( .A(n_222), .Y(n_286) );
AND2x2_ASAP7_75t_L g300 ( .A(n_222), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g304 ( .A(n_222), .Y(n_304) );
INVx2_ASAP7_75t_L g318 ( .A(n_222), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_222), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g375 ( .A(n_222), .B(n_370), .Y(n_375) );
AND2x2_ASAP7_75t_L g440 ( .A(n_222), .B(n_410), .Y(n_440) );
OR2x6_ASAP7_75t_L g222 ( .A(n_223), .B(n_233), .Y(n_222) );
AOI21xp5_ASAP7_75t_SL g223 ( .A1(n_224), .A2(n_225), .B(n_232), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_229), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_229), .A2(n_240), .B(n_241), .Y(n_239) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g268 ( .A(n_231), .Y(n_268) );
INVx1_ASAP7_75t_L g242 ( .A(n_232), .Y(n_242) );
OA21x2_ASAP7_75t_L g535 ( .A1(n_232), .A2(n_536), .B(n_546), .Y(n_535) );
OA21x2_ASAP7_75t_L g557 ( .A1(n_232), .A2(n_558), .B(n_565), .Y(n_557) );
AND2x2_ASAP7_75t_L g281 ( .A(n_235), .B(n_259), .Y(n_281) );
INVx2_ASAP7_75t_L g301 ( .A(n_235), .Y(n_301) );
AO21x2_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_242), .B(n_243), .Y(n_235) );
INVx1_ASAP7_75t_L g306 ( .A(n_245), .Y(n_306) );
AND2x2_ASAP7_75t_L g352 ( .A(n_245), .B(n_300), .Y(n_352) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_258), .Y(n_245) );
INVx2_ASAP7_75t_L g291 ( .A(n_246), .Y(n_291) );
INVx1_ASAP7_75t_L g299 ( .A(n_246), .Y(n_299) );
AND2x2_ASAP7_75t_L g317 ( .A(n_246), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_246), .B(n_301), .Y(n_355) );
AO21x2_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_248), .B(n_256), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_249), .B(n_255), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_252), .B(n_254), .Y(n_250) );
AND2x2_ASAP7_75t_L g334 ( .A(n_258), .B(n_291), .Y(n_334) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g287 ( .A(n_259), .Y(n_287) );
AND2x2_ASAP7_75t_L g370 ( .A(n_259), .B(n_301), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_265), .B(n_267), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_265), .A2(n_481), .B(n_482), .Y(n_480) );
INVx1_ASAP7_75t_L g540 ( .A(n_265), .Y(n_540) );
OAI21xp5_ASAP7_75t_SL g270 ( .A1(n_271), .A2(n_277), .B(n_281), .Y(n_270) );
INVx1_ASAP7_75t_SL g315 ( .A(n_271), .Y(n_315) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_272), .B(n_279), .Y(n_372) );
INVx1_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g321 ( .A(n_273), .B(n_276), .Y(n_321) );
AND2x2_ASAP7_75t_L g350 ( .A(n_273), .B(n_294), .Y(n_350) );
OR2x2_ASAP7_75t_L g353 ( .A(n_273), .B(n_313), .Y(n_353) );
AOI222xp33_ASAP7_75t_L g417 ( .A1(n_274), .A2(n_366), .B1(n_418), .B2(n_419), .C1(n_421), .C2(n_423), .Y(n_417) );
BUFx2_ASAP7_75t_L g331 ( .A(n_276), .Y(n_331) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g320 ( .A(n_279), .B(n_321), .Y(n_320) );
INVx3_ASAP7_75t_SL g337 ( .A(n_279), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_279), .B(n_331), .Y(n_391) );
AND2x2_ASAP7_75t_L g326 ( .A(n_281), .B(n_286), .Y(n_326) );
INVx1_ASAP7_75t_L g345 ( .A(n_281), .Y(n_345) );
OAI221xp5_ASAP7_75t_SL g282 ( .A1(n_283), .A2(n_284), .B1(n_288), .B2(n_292), .C(n_296), .Y(n_282) );
OR2x2_ASAP7_75t_L g354 ( .A(n_284), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
AND2x2_ASAP7_75t_L g339 ( .A(n_286), .B(n_309), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_286), .B(n_299), .Y(n_379) );
AND2x2_ASAP7_75t_L g384 ( .A(n_286), .B(n_334), .Y(n_384) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_286), .Y(n_394) );
NAND2x1_ASAP7_75t_SL g405 ( .A(n_286), .B(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g290 ( .A(n_287), .B(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g310 ( .A(n_287), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_287), .B(n_305), .Y(n_336) );
INVx1_ASAP7_75t_L g402 ( .A(n_287), .Y(n_402) );
INVx1_ASAP7_75t_L g377 ( .A(n_288), .Y(n_377) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
INVx1_ASAP7_75t_L g389 ( .A(n_289), .Y(n_389) );
NOR2xp67_ASAP7_75t_L g401 ( .A(n_289), .B(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g406 ( .A(n_290), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_290), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g309 ( .A(n_291), .B(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_291), .B(n_301), .Y(n_322) );
INVx1_ASAP7_75t_L g388 ( .A(n_291), .Y(n_388) );
INVx1_ASAP7_75t_L g409 ( .A(n_292), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OAI21xp5_ASAP7_75t_SL g296 ( .A1(n_297), .A2(n_302), .B(n_311), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_300), .Y(n_297) );
AND2x2_ASAP7_75t_L g442 ( .A(n_298), .B(n_375), .Y(n_442) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g410 ( .A(n_299), .B(n_370), .Y(n_410) );
AOI32xp33_ASAP7_75t_L g323 ( .A1(n_300), .A2(n_306), .A3(n_324), .B1(n_326), .B2(n_327), .Y(n_323) );
AOI322xp5_ASAP7_75t_L g425 ( .A1(n_300), .A2(n_332), .A3(n_415), .B1(n_426), .B2(n_427), .C1(n_428), .C2(n_430), .Y(n_425) );
INVx2_ASAP7_75t_L g305 ( .A(n_301), .Y(n_305) );
INVx1_ASAP7_75t_L g415 ( .A(n_301), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_306), .B1(n_307), .B2(n_308), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_303), .B(n_309), .Y(n_358) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_304), .B(n_370), .Y(n_420) );
INVx1_ASAP7_75t_L g307 ( .A(n_305), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_305), .B(n_334), .Y(n_424) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_313), .B(n_408), .Y(n_407) );
OAI221xp5_ASAP7_75t_SL g314 ( .A1(n_315), .A2(n_316), .B1(n_319), .B2(n_322), .C(n_323), .Y(n_314) );
OR2x2_ASAP7_75t_L g335 ( .A(n_316), .B(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g344 ( .A(n_316), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g369 ( .A(n_317), .B(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g373 ( .A(n_327), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OAI221xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_333), .B1(n_335), .B2(n_337), .C(n_338), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_331), .A2(n_362), .B1(n_366), .B2(n_367), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_332), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g437 ( .A(n_332), .Y(n_437) );
INVx1_ASAP7_75t_L g431 ( .A(n_334), .Y(n_431) );
INVx1_ASAP7_75t_SL g366 ( .A(n_335), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_337), .B(n_365), .Y(n_427) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_342), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_SL g408 ( .A(n_342), .Y(n_408) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
OAI221xp5_ASAP7_75t_SL g346 ( .A1(n_347), .A2(n_351), .B1(n_353), .B2(n_354), .C(n_356), .Y(n_346) );
NOR2xp33_ASAP7_75t_SL g347 ( .A(n_348), .B(n_350), .Y(n_347) );
AOI22xp5_ASAP7_75t_L g411 ( .A1(n_348), .A2(n_366), .B1(n_412), .B2(n_413), .Y(n_411) );
CKINVDCx14_ASAP7_75t_R g351 ( .A(n_352), .Y(n_351) );
OAI21xp33_ASAP7_75t_L g430 ( .A1(n_353), .A2(n_431), .B(n_432), .Y(n_430) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NOR3xp33_ASAP7_75t_SL g359 ( .A(n_360), .B(n_392), .C(n_416), .Y(n_359) );
NAND4xp25_ASAP7_75t_L g360 ( .A(n_361), .B(n_368), .C(n_376), .D(n_383), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
INVx1_ASAP7_75t_L g439 ( .A(n_364), .Y(n_439) );
INVx3_ASAP7_75t_SL g433 ( .A(n_365), .Y(n_433) );
OR2x2_ASAP7_75t_L g438 ( .A(n_365), .B(n_439), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_371), .B1(n_373), .B2(n_375), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_370), .B(n_388), .Y(n_429) );
INVxp67_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OAI21xp5_ASAP7_75t_SL g376 ( .A1(n_377), .A2(n_378), .B(n_380), .Y(n_376) );
INVxp67_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_389), .Y(n_386) );
INVxp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OAI211xp5_ASAP7_75t_SL g392 ( .A1(n_393), .A2(n_395), .B(n_398), .C(n_411), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g426 ( .A(n_397), .Y(n_426) );
AOI222xp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_403), .B1(n_404), .B2(n_407), .C1(n_409), .C2(n_410), .Y(n_398) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NAND4xp25_ASAP7_75t_SL g435 ( .A(n_408), .B(n_436), .C(n_437), .D(n_438), .Y(n_435) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NAND3xp33_ASAP7_75t_SL g416 ( .A(n_417), .B(n_425), .C(n_434), .Y(n_416) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_440), .B1(n_441), .B2(n_442), .Y(n_434) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
BUFx2_ASAP7_75t_L g455 ( .A(n_448), .Y(n_455) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
AOI21xp33_ASAP7_75t_L g456 ( .A1(n_453), .A2(n_457), .B(n_757), .Y(n_456) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_462), .B1(n_463), .B2(n_466), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g753 ( .A(n_460), .Y(n_753) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_663), .Y(n_467) );
NAND3xp33_ASAP7_75t_L g468 ( .A(n_469), .B(n_612), .C(n_654), .Y(n_468) );
AOI211xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_521), .B(n_566), .C(n_588), .Y(n_469) );
OAI211xp5_ASAP7_75t_SL g470 ( .A1(n_471), .A2(n_484), .B(n_505), .C(n_516), .Y(n_470) );
INVxp67_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_472), .B(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g675 ( .A(n_472), .B(n_592), .Y(n_675) );
BUFx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g577 ( .A(n_473), .B(n_508), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_473), .B(n_495), .Y(n_694) );
INVx1_ASAP7_75t_L g712 ( .A(n_473), .Y(n_712) );
AND2x2_ASAP7_75t_L g721 ( .A(n_473), .B(n_609), .Y(n_721) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
OR2x2_ASAP7_75t_L g604 ( .A(n_474), .B(n_495), .Y(n_604) );
AND2x2_ASAP7_75t_L g662 ( .A(n_474), .B(n_609), .Y(n_662) );
INVx1_ASAP7_75t_L g706 ( .A(n_474), .Y(n_706) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
OR2x2_ASAP7_75t_L g583 ( .A(n_475), .B(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g591 ( .A(n_475), .Y(n_591) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_475), .Y(n_631) );
INVxp67_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_486), .B(n_493), .Y(n_485) );
AND2x2_ASAP7_75t_L g570 ( .A(n_486), .B(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g603 ( .A(n_486), .Y(n_603) );
OR2x2_ASAP7_75t_L g729 ( .A(n_486), .B(n_730), .Y(n_729) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_486), .B(n_495), .Y(n_733) );
BUFx6f_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g508 ( .A(n_487), .Y(n_508) );
INVx1_ASAP7_75t_L g519 ( .A(n_487), .Y(n_519) );
AND2x2_ASAP7_75t_L g592 ( .A(n_487), .B(n_510), .Y(n_592) );
AND2x2_ASAP7_75t_L g632 ( .A(n_487), .B(n_511), .Y(n_632) );
OAI21xp5_ASAP7_75t_L g558 ( .A1(n_492), .A2(n_559), .B(n_562), .Y(n_558) );
INVxp67_ASAP7_75t_L g674 ( .A(n_493), .Y(n_674) );
AND2x4_ASAP7_75t_L g699 ( .A(n_493), .B(n_592), .Y(n_699) );
BUFx3_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_SL g590 ( .A(n_494), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g509 ( .A(n_495), .B(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g578 ( .A(n_495), .B(n_511), .Y(n_578) );
INVx1_ASAP7_75t_L g584 ( .A(n_495), .Y(n_584) );
INVx2_ASAP7_75t_L g610 ( .A(n_495), .Y(n_610) );
AND2x2_ASAP7_75t_L g626 ( .A(n_495), .B(n_627), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_499), .B(n_500), .Y(n_497) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_506), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_509), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx2_ASAP7_75t_L g581 ( .A(n_508), .Y(n_581) );
AND2x2_ASAP7_75t_L g689 ( .A(n_508), .B(n_510), .Y(n_689) );
AND2x2_ASAP7_75t_L g606 ( .A(n_509), .B(n_591), .Y(n_606) );
AND2x2_ASAP7_75t_L g705 ( .A(n_509), .B(n_706), .Y(n_705) );
NOR2xp67_ASAP7_75t_L g627 ( .A(n_510), .B(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g730 ( .A(n_510), .B(n_591), .Y(n_730) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx2_ASAP7_75t_L g520 ( .A(n_511), .Y(n_520) );
AND2x2_ASAP7_75t_L g609 ( .A(n_511), .B(n_610), .Y(n_609) );
O2A1O1Ixp33_ASAP7_75t_L g541 ( .A1(n_514), .A2(n_542), .B(n_544), .C(n_545), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_514), .A2(n_554), .B(n_555), .Y(n_553) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_520), .Y(n_517) );
AND2x2_ASAP7_75t_L g655 ( .A(n_518), .B(n_590), .Y(n_655) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_519), .B(n_591), .Y(n_640) );
INVx2_ASAP7_75t_L g639 ( .A(n_520), .Y(n_639) );
OAI222xp33_ASAP7_75t_L g643 ( .A1(n_520), .A2(n_583), .B1(n_644), .B2(n_646), .C1(n_647), .C2(n_650), .Y(n_643) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_532), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g568 ( .A(n_525), .Y(n_568) );
OR2x2_ASAP7_75t_L g679 ( .A(n_525), .B(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx3_ASAP7_75t_L g601 ( .A(n_526), .Y(n_601) );
NOR2x1_ASAP7_75t_L g652 ( .A(n_526), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g658 ( .A(n_526), .B(n_572), .Y(n_658) );
AND2x4_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
INVx1_ASAP7_75t_L g619 ( .A(n_527), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_532), .A2(n_622), .B1(n_661), .B2(n_662), .Y(n_660) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_547), .Y(n_532) );
INVx3_ASAP7_75t_L g594 ( .A(n_533), .Y(n_594) );
OR2x2_ASAP7_75t_L g727 ( .A(n_533), .B(n_603), .Y(n_727) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g600 ( .A(n_534), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g616 ( .A(n_534), .B(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g624 ( .A(n_534), .B(n_572), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_534), .B(n_548), .Y(n_680) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g571 ( .A(n_535), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g575 ( .A(n_535), .B(n_548), .Y(n_575) );
AND2x2_ASAP7_75t_L g651 ( .A(n_535), .B(n_598), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_535), .B(n_557), .Y(n_691) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_547), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g607 ( .A(n_547), .B(n_568), .Y(n_607) );
AND2x2_ASAP7_75t_L g611 ( .A(n_547), .B(n_601), .Y(n_611) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_557), .Y(n_547) );
INVx3_ASAP7_75t_L g572 ( .A(n_548), .Y(n_572) );
AND2x2_ASAP7_75t_L g597 ( .A(n_548), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g732 ( .A(n_548), .B(n_715), .Y(n_732) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_557), .Y(n_586) );
INVx2_ASAP7_75t_L g598 ( .A(n_557), .Y(n_598) );
AND2x2_ASAP7_75t_L g642 ( .A(n_557), .B(n_618), .Y(n_642) );
INVx1_ASAP7_75t_L g685 ( .A(n_557), .Y(n_685) );
OR2x2_ASAP7_75t_L g716 ( .A(n_557), .B(n_618), .Y(n_716) );
AND2x2_ASAP7_75t_L g736 ( .A(n_557), .B(n_572), .Y(n_736) );
OAI21xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_569), .B(n_573), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g574 ( .A(n_568), .B(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_568), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g693 ( .A(n_570), .Y(n_693) );
INVx2_ASAP7_75t_SL g587 ( .A(n_571), .Y(n_587) );
AND2x2_ASAP7_75t_L g707 ( .A(n_571), .B(n_601), .Y(n_707) );
INVx2_ASAP7_75t_L g653 ( .A(n_572), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_572), .B(n_685), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_576), .B1(n_579), .B2(n_585), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_575), .B(n_720), .Y(n_719) );
INVx1_ASAP7_75t_SL g741 ( .A(n_575), .Y(n_741) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
INVx1_ASAP7_75t_L g666 ( .A(n_577), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_577), .B(n_609), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_578), .B(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g682 ( .A(n_578), .B(n_631), .Y(n_682) );
INVx2_ASAP7_75t_L g738 ( .A(n_578), .Y(n_738) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
AND2x2_ASAP7_75t_L g608 ( .A(n_581), .B(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_581), .B(n_626), .Y(n_659) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_583), .B(n_603), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
INVx1_ASAP7_75t_L g720 ( .A(n_586), .Y(n_720) );
O2A1O1Ixp33_ASAP7_75t_SL g670 ( .A1(n_587), .A2(n_671), .B(n_673), .C(n_676), .Y(n_670) );
OR2x2_ASAP7_75t_L g697 ( .A(n_587), .B(n_601), .Y(n_697) );
OAI221xp5_ASAP7_75t_SL g588 ( .A1(n_589), .A2(n_593), .B1(n_595), .B2(n_602), .C(n_605), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_590), .B(n_592), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_590), .B(n_639), .Y(n_646) );
AND2x2_ASAP7_75t_L g688 ( .A(n_590), .B(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g724 ( .A(n_590), .Y(n_724) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_591), .Y(n_615) );
INVx1_ASAP7_75t_L g628 ( .A(n_591), .Y(n_628) );
NOR2xp67_ASAP7_75t_L g648 ( .A(n_594), .B(n_649), .Y(n_648) );
INVxp67_ASAP7_75t_L g702 ( .A(n_594), .Y(n_702) );
NAND2xp5_ASAP7_75t_SL g718 ( .A(n_594), .B(n_642), .Y(n_718) );
INVx2_ASAP7_75t_L g704 ( .A(n_595), .Y(n_704) );
OR2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_599), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g645 ( .A(n_597), .B(n_616), .Y(n_645) );
O2A1O1Ixp33_ASAP7_75t_L g654 ( .A1(n_597), .A2(n_613), .B(n_655), .C(n_656), .Y(n_654) );
AND2x2_ASAP7_75t_L g623 ( .A(n_598), .B(n_618), .Y(n_623) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_602), .B(n_701), .Y(n_700) );
OR2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
OR2x2_ASAP7_75t_L g671 ( .A(n_603), .B(n_672), .Y(n_671) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_607), .B1(n_608), .B2(n_611), .Y(n_605) );
INVx1_ASAP7_75t_L g725 ( .A(n_607), .Y(n_725) );
INVx1_ASAP7_75t_L g672 ( .A(n_609), .Y(n_672) );
INVx1_ASAP7_75t_L g723 ( .A(n_611), .Y(n_723) );
AOI211xp5_ASAP7_75t_SL g612 ( .A1(n_613), .A2(n_616), .B(n_620), .C(n_643), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g635 ( .A(n_615), .B(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g686 ( .A(n_616), .Y(n_686) );
AND2x2_ASAP7_75t_L g735 ( .A(n_616), .B(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OAI21xp33_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_625), .B(n_633), .Y(n_620) );
INVx1_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
INVx2_ASAP7_75t_L g649 ( .A(n_623), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_623), .B(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g641 ( .A(n_624), .B(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g717 ( .A(n_624), .Y(n_717) );
OAI32xp33_ASAP7_75t_L g728 ( .A1(n_624), .A2(n_676), .A3(n_683), .B1(n_724), .B2(n_729), .Y(n_728) );
NOR2xp33_ASAP7_75t_SL g625 ( .A(n_626), .B(n_629), .Y(n_625) );
INVx1_ASAP7_75t_SL g696 ( .A(n_626), .Y(n_696) );
AND2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_SL g636 ( .A(n_632), .Y(n_636) );
OAI21xp33_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_637), .B(n_641), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OAI22xp33_ASAP7_75t_L g708 ( .A1(n_635), .A2(n_683), .B1(n_709), .B2(n_711), .Y(n_708) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_639), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g676 ( .A(n_642), .Y(n_676) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND2x1p5_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
INVx1_ASAP7_75t_L g669 ( .A(n_653), .Y(n_669) );
OAI21xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_659), .B(n_660), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_662), .A2(n_704), .B1(n_705), .B2(n_707), .C(n_708), .Y(n_703) );
NAND5xp2_ASAP7_75t_L g663 ( .A(n_664), .B(n_687), .C(n_703), .D(n_713), .E(n_731), .Y(n_663) );
AOI211xp5_ASAP7_75t_SL g664 ( .A1(n_665), .A2(n_667), .B(n_670), .C(n_677), .Y(n_664) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g734 ( .A(n_671), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
OAI22xp33_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_679), .B1(n_681), .B2(n_683), .Y(n_677) );
INVx1_ASAP7_75t_SL g710 ( .A(n_680), .Y(n_710) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
OAI322xp33_ASAP7_75t_L g692 ( .A1(n_683), .A2(n_693), .A3(n_694), .B1(n_695), .B2(n_696), .C1(n_697), .C2(n_698), .Y(n_692) );
OR2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_686), .Y(n_683) );
INVx1_ASAP7_75t_L g695 ( .A(n_685), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_685), .B(n_710), .Y(n_709) );
AOI211xp5_ASAP7_75t_SL g687 ( .A1(n_688), .A2(n_690), .B(n_692), .C(n_700), .Y(n_687) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
OAI22xp33_ASAP7_75t_L g722 ( .A1(n_696), .A2(n_723), .B1(n_724), .B2(n_725), .Y(n_722) );
INVx1_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g739 ( .A(n_706), .Y(n_739) );
AOI221xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_721), .B1(n_722), .B2(n_726), .C(n_728), .Y(n_713) );
OAI211xp5_ASAP7_75t_SL g714 ( .A1(n_715), .A2(n_717), .B(n_718), .C(n_719), .Y(n_714) );
INVx1_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
OR2x2_ASAP7_75t_L g740 ( .A(n_716), .B(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
AOI221xp5_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_733), .B1(n_734), .B2(n_735), .C(n_737), .Y(n_731) );
AOI21xp33_ASAP7_75t_SL g737 ( .A1(n_738), .A2(n_739), .B(n_740), .Y(n_737) );
CKINVDCx16_ASAP7_75t_R g742 ( .A(n_743), .Y(n_742) );
CKINVDCx16_ASAP7_75t_R g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
INVx3_ASAP7_75t_SL g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
endmodule