module fake_jpeg_30456_n_24 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_24);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_24;

wire n_13;
wire n_21;
wire n_23;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_16;
wire n_11;
wire n_17;
wire n_12;
wire n_15;

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_4),
.B(n_6),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_12),
.A2(n_10),
.B1(n_9),
.B2(n_8),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_15),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_0),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_16),
.B(n_17),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_0),
.C(n_1),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_19),
.B(n_17),
.C(n_14),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_20),
.A2(n_21),
.B(n_2),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_18),
.B(n_1),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_22),
.B(n_2),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_23),
.B(n_3),
.C(n_4),
.Y(n_24)
);


endmodule