module fake_aes_8721_n_747 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_747);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_747;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_466;
wire n_302;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_146;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g82 ( .A(n_34), .Y(n_82) );
BUFx6f_ASAP7_75t_L g83 ( .A(n_65), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_77), .Y(n_84) );
INVxp33_ASAP7_75t_SL g85 ( .A(n_15), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_16), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_23), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_42), .Y(n_88) );
BUFx3_ASAP7_75t_L g89 ( .A(n_35), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_78), .Y(n_90) );
CKINVDCx20_ASAP7_75t_R g91 ( .A(n_73), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_11), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_47), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_43), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_60), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_54), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_2), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_6), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_14), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_0), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_59), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_44), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_10), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_21), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_1), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_39), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_37), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_49), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_14), .Y(n_109) );
INVxp33_ASAP7_75t_L g110 ( .A(n_1), .Y(n_110) );
CKINVDCx14_ASAP7_75t_R g111 ( .A(n_41), .Y(n_111) );
BUFx3_ASAP7_75t_L g112 ( .A(n_50), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_61), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_81), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_45), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_66), .Y(n_116) );
INVxp67_ASAP7_75t_L g117 ( .A(n_9), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_6), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_25), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_74), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_38), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_63), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_21), .Y(n_123) );
INVxp67_ASAP7_75t_SL g124 ( .A(n_2), .Y(n_124) );
INVxp67_ASAP7_75t_SL g125 ( .A(n_15), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_12), .Y(n_126) );
INVxp33_ASAP7_75t_SL g127 ( .A(n_12), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_9), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_24), .Y(n_129) );
INVxp67_ASAP7_75t_SL g130 ( .A(n_27), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_26), .Y(n_131) );
INVx6_ASAP7_75t_L g132 ( .A(n_83), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_82), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_82), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_84), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_84), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_83), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_87), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_94), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_118), .Y(n_140) );
AND2x6_ASAP7_75t_L g141 ( .A(n_89), .B(n_40), .Y(n_141) );
NAND2x1_ASAP7_75t_L g142 ( .A(n_86), .B(n_0), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_110), .B(n_3), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g144 ( .A(n_85), .B(n_3), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_87), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_118), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_95), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_95), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_117), .B(n_4), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_94), .B(n_4), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_102), .B(n_5), .Y(n_151) );
OAI21x1_ASAP7_75t_L g152 ( .A1(n_102), .A2(n_48), .B(n_79), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_107), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_127), .B(n_5), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_107), .B(n_7), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_108), .B(n_7), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_96), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_83), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_113), .B(n_8), .Y(n_159) );
OAI22xp5_ASAP7_75t_SL g160 ( .A1(n_109), .A2(n_8), .B1(n_10), .B2(n_11), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_83), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_96), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_101), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_131), .B(n_13), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_101), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_86), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_106), .B(n_13), .Y(n_167) );
BUFx3_ASAP7_75t_L g168 ( .A(n_89), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_106), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_115), .Y(n_170) );
AND2x6_ASAP7_75t_L g171 ( .A(n_112), .B(n_53), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_115), .Y(n_172) );
AND2x4_ASAP7_75t_L g173 ( .A(n_92), .B(n_16), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_83), .B(n_17), .Y(n_174) );
AND2x4_ASAP7_75t_L g175 ( .A(n_92), .B(n_17), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_112), .Y(n_176) );
BUFx3_ASAP7_75t_L g177 ( .A(n_168), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_176), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_173), .Y(n_179) );
INVxp67_ASAP7_75t_L g180 ( .A(n_143), .Y(n_180) );
INVxp67_ASAP7_75t_L g181 ( .A(n_143), .Y(n_181) );
CKINVDCx5p33_ASAP7_75t_R g182 ( .A(n_141), .Y(n_182) );
AND2x4_ASAP7_75t_L g183 ( .A(n_173), .B(n_98), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_133), .B(n_114), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_139), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_166), .B(n_133), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_139), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_173), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_175), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_168), .B(n_111), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_137), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_176), .Y(n_192) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_134), .Y(n_193) );
INVx3_ASAP7_75t_L g194 ( .A(n_175), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_134), .B(n_99), .Y(n_195) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_137), .Y(n_196) );
AND2x6_ASAP7_75t_L g197 ( .A(n_175), .B(n_116), .Y(n_197) );
AND2x4_ASAP7_75t_SL g198 ( .A(n_144), .B(n_91), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_176), .Y(n_199) );
INVx4_ASAP7_75t_L g200 ( .A(n_141), .Y(n_200) );
NAND3xp33_ASAP7_75t_L g201 ( .A(n_149), .B(n_103), .C(n_104), .Y(n_201) );
INVx3_ASAP7_75t_L g202 ( .A(n_153), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_153), .Y(n_203) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_137), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_135), .B(n_99), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_135), .B(n_98), .Y(n_206) );
AND2x4_ASAP7_75t_L g207 ( .A(n_136), .B(n_100), .Y(n_207) );
INVx4_ASAP7_75t_L g208 ( .A(n_141), .Y(n_208) );
BUFx3_ASAP7_75t_L g209 ( .A(n_176), .Y(n_209) );
OR2x2_ASAP7_75t_L g210 ( .A(n_136), .B(n_97), .Y(n_210) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_137), .Y(n_211) );
AND2x6_ASAP7_75t_L g212 ( .A(n_138), .B(n_119), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_162), .Y(n_213) );
BUFx3_ASAP7_75t_L g214 ( .A(n_176), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_162), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_138), .B(n_119), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_145), .B(n_88), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_145), .B(n_103), .Y(n_218) );
AND2x4_ASAP7_75t_L g219 ( .A(n_147), .B(n_100), .Y(n_219) );
AND2x4_ASAP7_75t_L g220 ( .A(n_147), .B(n_148), .Y(n_220) );
OA22x2_ASAP7_75t_L g221 ( .A1(n_142), .A2(n_123), .B1(n_104), .B2(n_128), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_141), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_148), .B(n_123), .Y(n_223) );
AND2x4_ASAP7_75t_L g224 ( .A(n_157), .B(n_105), .Y(n_224) );
BUFx3_ASAP7_75t_L g225 ( .A(n_141), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_137), .Y(n_226) );
INVx3_ASAP7_75t_L g227 ( .A(n_170), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_170), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_157), .B(n_105), .Y(n_229) );
INVxp67_ASAP7_75t_L g230 ( .A(n_154), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_163), .B(n_90), .Y(n_231) );
AND2x4_ASAP7_75t_L g232 ( .A(n_163), .B(n_97), .Y(n_232) );
AND2x2_ASAP7_75t_L g233 ( .A(n_165), .B(n_128), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_165), .B(n_122), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_141), .Y(n_235) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_169), .A2(n_125), .B1(n_124), .B2(n_116), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_169), .B(n_93), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_172), .B(n_129), .Y(n_238) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_158), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_132), .Y(n_240) );
AND2x2_ASAP7_75t_L g241 ( .A(n_172), .B(n_129), .Y(n_241) );
NAND3xp33_ASAP7_75t_L g242 ( .A(n_159), .B(n_164), .C(n_156), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_140), .B(n_122), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_152), .Y(n_244) );
INVx4_ASAP7_75t_L g245 ( .A(n_141), .Y(n_245) );
BUFx10_ASAP7_75t_L g246 ( .A(n_171), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_220), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_193), .B(n_146), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_198), .Y(n_249) );
BUFx2_ASAP7_75t_L g250 ( .A(n_212), .Y(n_250) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_246), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_178), .Y(n_252) );
OR2x2_ASAP7_75t_SL g253 ( .A(n_242), .B(n_160), .Y(n_253) );
INVx5_ASAP7_75t_L g254 ( .A(n_197), .Y(n_254) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_246), .Y(n_255) );
BUFx3_ASAP7_75t_L g256 ( .A(n_225), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_178), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_220), .B(n_167), .Y(n_258) );
NOR2x1_ASAP7_75t_R g259 ( .A(n_183), .B(n_130), .Y(n_259) );
AND2x4_ASAP7_75t_L g260 ( .A(n_183), .B(n_142), .Y(n_260) );
INVx1_ASAP7_75t_SL g261 ( .A(n_210), .Y(n_261) );
BUFx4f_ASAP7_75t_L g262 ( .A(n_197), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_220), .Y(n_263) );
AND2x4_ASAP7_75t_L g264 ( .A(n_183), .B(n_140), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_197), .A2(n_171), .B1(n_150), .B2(n_151), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_215), .Y(n_266) );
INVxp67_ASAP7_75t_SL g267 ( .A(n_225), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_186), .B(n_155), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_215), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_228), .Y(n_270) );
BUFx4f_ASAP7_75t_L g271 ( .A(n_197), .Y(n_271) );
AND2x4_ASAP7_75t_L g272 ( .A(n_180), .B(n_140), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_228), .Y(n_273) );
INVx5_ASAP7_75t_L g274 ( .A(n_197), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_186), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_206), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_230), .B(n_146), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g278 ( .A1(n_197), .A2(n_171), .B1(n_174), .B2(n_146), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_192), .Y(n_279) );
AOI22xp5_ASAP7_75t_L g280 ( .A1(n_181), .A2(n_171), .B1(n_126), .B2(n_120), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_206), .Y(n_281) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_246), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_198), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_192), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_206), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_207), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_231), .B(n_171), .Y(n_287) );
AND2x4_ASAP7_75t_L g288 ( .A(n_201), .B(n_152), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_207), .Y(n_289) );
INVx6_ASAP7_75t_L g290 ( .A(n_177), .Y(n_290) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_207), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_219), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_199), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_219), .Y(n_294) );
BUFx3_ASAP7_75t_L g295 ( .A(n_200), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_219), .B(n_171), .Y(n_296) );
INVx1_ASAP7_75t_SL g297 ( .A(n_210), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_223), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_212), .Y(n_299) );
BUFx2_ASAP7_75t_L g300 ( .A(n_212), .Y(n_300) );
AND2x6_ASAP7_75t_L g301 ( .A(n_194), .B(n_121), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_199), .Y(n_302) );
NOR2xp33_ASAP7_75t_R g303 ( .A(n_182), .B(n_171), .Y(n_303) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_200), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_223), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_223), .Y(n_306) );
INVx4_ASAP7_75t_L g307 ( .A(n_200), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_224), .B(n_121), .Y(n_308) );
BUFx3_ASAP7_75t_L g309 ( .A(n_208), .Y(n_309) );
BUFx3_ASAP7_75t_L g310 ( .A(n_208), .Y(n_310) );
BUFx3_ASAP7_75t_L g311 ( .A(n_208), .Y(n_311) );
BUFx2_ASAP7_75t_L g312 ( .A(n_212), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_212), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_224), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_224), .Y(n_315) );
INVxp67_ASAP7_75t_SL g316 ( .A(n_194), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_229), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_184), .B(n_120), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_229), .B(n_132), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_229), .B(n_132), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_232), .B(n_132), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_261), .B(n_195), .Y(n_322) );
BUFx2_ASAP7_75t_SL g323 ( .A(n_254), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_266), .Y(n_324) );
AOI21xp5_ASAP7_75t_L g325 ( .A1(n_287), .A2(n_245), .B(n_244), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_269), .Y(n_326) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_297), .Y(n_327) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_291), .Y(n_328) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_298), .Y(n_329) );
O2A1O1Ixp33_ASAP7_75t_L g330 ( .A1(n_268), .A2(n_188), .B(n_179), .C(n_189), .Y(n_330) );
BUFx12f_ASAP7_75t_L g331 ( .A(n_249), .Y(n_331) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_304), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_258), .B(n_260), .Y(n_333) );
INVx4_ASAP7_75t_L g334 ( .A(n_262), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_270), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_273), .Y(n_336) );
INVx2_ASAP7_75t_SL g337 ( .A(n_254), .Y(n_337) );
CKINVDCx8_ASAP7_75t_R g338 ( .A(n_249), .Y(n_338) );
NAND2xp33_ASAP7_75t_L g339 ( .A(n_303), .B(n_182), .Y(n_339) );
AOI22xp33_ASAP7_75t_SL g340 ( .A1(n_283), .A2(n_221), .B1(n_212), .B2(n_232), .Y(n_340) );
A2O1A1Ixp33_ASAP7_75t_L g341 ( .A1(n_276), .A2(n_194), .B(n_234), .C(n_216), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_275), .B(n_195), .Y(n_342) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_304), .Y(n_343) );
INVx2_ASAP7_75t_SL g344 ( .A(n_254), .Y(n_344) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_304), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_259), .B(n_217), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_252), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_247), .Y(n_348) );
NOR2x1_ASAP7_75t_L g349 ( .A(n_263), .B(n_177), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_248), .B(n_233), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_248), .B(n_233), .Y(n_351) );
INVx3_ASAP7_75t_L g352 ( .A(n_307), .Y(n_352) );
AO21x2_ASAP7_75t_L g353 ( .A1(n_288), .A2(n_244), .B(n_238), .Y(n_353) );
OR2x6_ASAP7_75t_L g354 ( .A(n_300), .B(n_250), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_252), .Y(n_355) );
INVx3_ASAP7_75t_L g356 ( .A(n_307), .Y(n_356) );
AOI22xp5_ASAP7_75t_L g357 ( .A1(n_281), .A2(n_221), .B1(n_232), .B2(n_241), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_285), .Y(n_358) );
AND2x4_ASAP7_75t_L g359 ( .A(n_260), .B(n_241), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_286), .Y(n_360) );
AOI21xp33_ASAP7_75t_L g361 ( .A1(n_280), .A2(n_222), .B(n_235), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_257), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_260), .B(n_205), .Y(n_363) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_301), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_289), .B(n_238), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_292), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_257), .Y(n_367) );
OR2x6_ASAP7_75t_SL g368 ( .A(n_283), .B(n_235), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_294), .B(n_218), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_305), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_279), .Y(n_371) );
NAND2xp5_ASAP7_75t_SL g372 ( .A(n_254), .B(n_245), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_306), .B(n_218), .Y(n_373) );
BUFx2_ASAP7_75t_L g374 ( .A(n_301), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_314), .B(n_315), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_262), .A2(n_222), .B1(n_245), .B2(n_236), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_317), .Y(n_377) );
NOR2xp67_ASAP7_75t_L g378 ( .A(n_254), .B(n_202), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_253), .B(n_205), .Y(n_379) );
OAI221xp5_ASAP7_75t_L g380 ( .A1(n_379), .A2(n_277), .B1(n_318), .B2(n_308), .C(n_265), .Y(n_380) );
O2A1O1Ixp33_ASAP7_75t_L g381 ( .A1(n_341), .A2(n_277), .B(n_318), .C(n_272), .Y(n_381) );
OAI21xp5_ASAP7_75t_L g382 ( .A1(n_325), .A2(n_288), .B(n_296), .Y(n_382) );
CKINVDCx11_ASAP7_75t_R g383 ( .A(n_338), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_324), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_327), .A2(n_301), .B1(n_272), .B2(n_264), .Y(n_385) );
A2O1A1Ixp33_ASAP7_75t_L g386 ( .A1(n_330), .A2(n_288), .B(n_271), .C(n_262), .Y(n_386) );
INVx6_ASAP7_75t_L g387 ( .A(n_332), .Y(n_387) );
AND2x4_ASAP7_75t_L g388 ( .A(n_359), .B(n_274), .Y(n_388) );
AOI22xp33_ASAP7_75t_SL g389 ( .A1(n_322), .A2(n_301), .B1(n_271), .B2(n_221), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_347), .Y(n_390) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_322), .Y(n_391) );
OAI21x1_ASAP7_75t_L g392 ( .A1(n_324), .A2(n_278), .B(n_284), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_359), .A2(n_301), .B1(n_272), .B2(n_264), .Y(n_393) );
BUFx3_ASAP7_75t_L g394 ( .A(n_332), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_363), .B(n_264), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_359), .A2(n_301), .B1(n_316), .B2(n_271), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_324), .Y(n_397) );
CKINVDCx20_ASAP7_75t_R g398 ( .A(n_338), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_335), .Y(n_399) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_359), .Y(n_400) );
AOI222xp33_ASAP7_75t_L g401 ( .A1(n_350), .A2(n_253), .B1(n_243), .B2(n_213), .C1(n_237), .C2(n_185), .Y(n_401) );
CKINVDCx5p33_ASAP7_75t_R g402 ( .A(n_331), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_335), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_335), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_336), .Y(n_405) );
AOI21xp5_ASAP7_75t_L g406 ( .A1(n_353), .A2(n_267), .B(n_307), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_328), .Y(n_407) );
INVx3_ASAP7_75t_L g408 ( .A(n_334), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_347), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_379), .A2(n_243), .B1(n_227), .B2(n_185), .Y(n_410) );
BUFx4_ASAP7_75t_SL g411 ( .A(n_374), .Y(n_411) );
CKINVDCx11_ASAP7_75t_R g412 ( .A(n_331), .Y(n_412) );
BUFx12f_ASAP7_75t_L g413 ( .A(n_331), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_363), .B(n_227), .Y(n_414) );
AOI21xp5_ASAP7_75t_L g415 ( .A1(n_353), .A2(n_309), .B(n_295), .Y(n_415) );
OAI22xp33_ASAP7_75t_L g416 ( .A1(n_391), .A2(n_368), .B1(n_374), .B2(n_357), .Y(n_416) );
NAND2xp5_ASAP7_75t_SL g417 ( .A(n_384), .B(n_336), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_401), .A2(n_340), .B1(n_351), .B2(n_350), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_410), .B(n_351), .Y(n_419) );
A2O1A1Ixp33_ASAP7_75t_L g420 ( .A1(n_381), .A2(n_357), .B(n_326), .C(n_336), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_384), .B(n_353), .Y(n_421) );
BUFx3_ASAP7_75t_L g422 ( .A(n_413), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_380), .A2(n_342), .B1(n_369), .B2(n_326), .Y(n_423) );
AOI21xp5_ASAP7_75t_L g424 ( .A1(n_386), .A2(n_382), .B(n_390), .Y(n_424) );
OAI22xp33_ASAP7_75t_L g425 ( .A1(n_410), .A2(n_368), .B1(n_333), .B2(n_354), .Y(n_425) );
AND2x4_ASAP7_75t_L g426 ( .A(n_397), .B(n_348), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_397), .B(n_342), .Y(n_427) );
BUFx4f_ASAP7_75t_SL g428 ( .A(n_413), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_399), .B(n_369), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_399), .A2(n_375), .B1(n_377), .B2(n_360), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_390), .Y(n_431) );
AO31x2_ASAP7_75t_L g432 ( .A1(n_403), .A2(n_370), .A3(n_377), .B(n_358), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_389), .A2(n_329), .B1(n_346), .B2(n_360), .Y(n_433) );
OR2x6_ASAP7_75t_L g434 ( .A(n_403), .B(n_354), .Y(n_434) );
OAI22xp33_ASAP7_75t_L g435 ( .A1(n_398), .A2(n_354), .B1(n_365), .B2(n_364), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_400), .A2(n_370), .B1(n_366), .B2(n_358), .Y(n_436) );
INVx1_ASAP7_75t_SL g437 ( .A(n_390), .Y(n_437) );
INVx2_ASAP7_75t_SL g438 ( .A(n_411), .Y(n_438) );
OAI221xp5_ASAP7_75t_L g439 ( .A1(n_385), .A2(n_373), .B1(n_366), .B2(n_348), .C(n_361), .Y(n_439) );
AOI221xp5_ASAP7_75t_SL g440 ( .A1(n_404), .A2(n_375), .B1(n_187), .B2(n_203), .C(n_320), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_407), .A2(n_349), .B1(n_353), .B2(n_356), .Y(n_441) );
AOI222xp33_ASAP7_75t_L g442 ( .A1(n_395), .A2(n_187), .B1(n_203), .B2(n_376), .C1(n_227), .C2(n_202), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_409), .Y(n_443) );
AOI221xp5_ASAP7_75t_SL g444 ( .A1(n_404), .A2(n_319), .B1(n_321), .B2(n_190), .C(n_202), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_393), .A2(n_349), .B1(n_352), .B2(n_356), .Y(n_445) );
AOI221xp5_ASAP7_75t_L g446 ( .A1(n_423), .A2(n_414), .B1(n_405), .B2(n_402), .C(n_396), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_427), .B(n_405), .Y(n_447) );
AOI33xp33_ASAP7_75t_L g448 ( .A1(n_418), .A2(n_240), .A3(n_388), .B1(n_20), .B2(n_18), .B3(n_19), .Y(n_448) );
BUFx3_ASAP7_75t_L g449 ( .A(n_434), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_431), .Y(n_450) );
INVx3_ASAP7_75t_L g451 ( .A(n_426), .Y(n_451) );
BUFx3_ASAP7_75t_L g452 ( .A(n_434), .Y(n_452) );
OAI211xp5_ASAP7_75t_L g453 ( .A1(n_433), .A2(n_383), .B(n_412), .C(n_402), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_431), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_425), .A2(n_409), .B1(n_388), .B2(n_408), .Y(n_455) );
AOI211xp5_ASAP7_75t_L g456 ( .A1(n_416), .A2(n_388), .B(n_409), .C(n_415), .Y(n_456) );
OAI221xp5_ASAP7_75t_L g457 ( .A1(n_419), .A2(n_430), .B1(n_436), .B2(n_440), .C(n_420), .Y(n_457) );
AOI22xp33_ASAP7_75t_SL g458 ( .A1(n_438), .A2(n_408), .B1(n_388), .B2(n_394), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_443), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_435), .A2(n_408), .B1(n_406), .B2(n_352), .Y(n_460) );
OAI31xp33_ASAP7_75t_L g461 ( .A1(n_427), .A2(n_408), .A3(n_352), .B(n_356), .Y(n_461) );
OAI221xp5_ASAP7_75t_L g462 ( .A1(n_430), .A2(n_354), .B1(n_367), .B2(n_362), .C(n_347), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_434), .A2(n_354), .B1(n_387), .B2(n_394), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_443), .Y(n_464) );
AOI211xp5_ASAP7_75t_L g465 ( .A1(n_438), .A2(n_378), .B(n_355), .C(n_362), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_437), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_442), .A2(n_352), .B1(n_356), .B2(n_394), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_437), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_422), .B(n_387), .Y(n_469) );
AOI33xp33_ASAP7_75t_L g470 ( .A1(n_441), .A2(n_240), .A3(n_18), .B1(n_19), .B2(n_20), .B3(n_355), .Y(n_470) );
AOI221xp5_ASAP7_75t_L g471 ( .A1(n_429), .A2(n_371), .B1(n_367), .B2(n_362), .C(n_355), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_421), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_422), .B(n_387), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_429), .B(n_367), .Y(n_474) );
OAI22xp33_ASAP7_75t_L g475 ( .A1(n_434), .A2(n_334), .B1(n_313), .B2(n_299), .Y(n_475) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_444), .A2(n_392), .B(n_371), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_442), .A2(n_334), .B1(n_387), .B2(n_290), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_421), .Y(n_478) );
OAI31xp33_ASAP7_75t_L g479 ( .A1(n_439), .A2(n_300), .A3(n_312), .B(n_371), .Y(n_479) );
AOI221xp5_ASAP7_75t_L g480 ( .A1(n_440), .A2(n_158), .B1(n_161), .B2(n_214), .C(n_209), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_432), .Y(n_481) );
OAI222xp33_ASAP7_75t_L g482 ( .A1(n_434), .A2(n_334), .B1(n_299), .B2(n_313), .C1(n_337), .C2(n_344), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_426), .B(n_392), .Y(n_483) );
INVx2_ASAP7_75t_SL g484 ( .A(n_451), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_481), .Y(n_485) );
BUFx3_ASAP7_75t_L g486 ( .A(n_451), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_474), .B(n_426), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_481), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_481), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_450), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_472), .B(n_432), .Y(n_491) );
INVx1_ASAP7_75t_SL g492 ( .A(n_466), .Y(n_492) );
AOI221xp5_ASAP7_75t_L g493 ( .A1(n_457), .A2(n_444), .B1(n_426), .B2(n_424), .C(n_445), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_472), .B(n_432), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_450), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_478), .Y(n_496) );
INVx2_ASAP7_75t_SL g497 ( .A(n_451), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_450), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_478), .B(n_432), .Y(n_499) );
INVxp67_ASAP7_75t_L g500 ( .A(n_474), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_454), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_454), .Y(n_502) );
NAND4xp25_ASAP7_75t_L g503 ( .A(n_448), .B(n_209), .C(n_214), .D(n_417), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_454), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_459), .Y(n_505) );
AOI33xp33_ASAP7_75t_L g506 ( .A1(n_458), .A2(n_428), .A3(n_293), .B1(n_302), .B2(n_279), .B3(n_284), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_447), .B(n_432), .Y(n_507) );
NOR2x1_ASAP7_75t_L g508 ( .A(n_462), .B(n_378), .Y(n_508) );
OAI211xp5_ASAP7_75t_SL g509 ( .A1(n_453), .A2(n_302), .B(n_293), .C(n_372), .Y(n_509) );
INVx3_ASAP7_75t_L g510 ( .A(n_459), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_459), .B(n_158), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_464), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_446), .A2(n_345), .B1(n_343), .B2(n_332), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_447), .B(n_345), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_464), .B(n_158), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_464), .B(n_451), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_465), .B(n_345), .Y(n_517) );
INVx4_ASAP7_75t_L g518 ( .A(n_449), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_483), .Y(n_519) );
OAI31xp33_ASAP7_75t_L g520 ( .A1(n_462), .A2(n_344), .A3(n_337), .B(n_310), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_466), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_466), .Y(n_522) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_476), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_483), .B(n_161), .Y(n_524) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_468), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_468), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_468), .B(n_345), .Y(n_527) );
OAI221xp5_ASAP7_75t_SL g528 ( .A1(n_470), .A2(n_22), .B1(n_28), .B2(n_29), .C(n_30), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_476), .Y(n_529) );
NAND3xp33_ASAP7_75t_L g530 ( .A(n_465), .B(n_161), .C(n_158), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_449), .B(n_161), .Y(n_531) );
AOI33xp33_ASAP7_75t_L g532 ( .A1(n_458), .A2(n_161), .A3(n_32), .B1(n_33), .B2(n_36), .B3(n_46), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_455), .A2(n_345), .B1(n_343), .B2(n_332), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_476), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_453), .B(n_290), .Y(n_535) );
INVxp67_ASAP7_75t_SL g536 ( .A(n_463), .Y(n_536) );
OAI322xp33_ASAP7_75t_L g537 ( .A1(n_500), .A2(n_457), .A3(n_455), .B1(n_469), .B2(n_473), .C1(n_463), .C2(n_475), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_530), .A2(n_480), .B(n_461), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_510), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_496), .Y(n_540) );
NOR2x1_ASAP7_75t_L g541 ( .A(n_530), .B(n_452), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_496), .Y(n_542) );
OAI322xp33_ASAP7_75t_L g543 ( .A1(n_494), .A2(n_446), .A3(n_461), .B1(n_456), .B2(n_204), .C1(n_196), .C2(n_211), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_487), .B(n_449), .Y(n_544) );
INVx3_ASAP7_75t_L g545 ( .A(n_518), .Y(n_545) );
NAND4xp25_ASAP7_75t_L g546 ( .A(n_493), .B(n_456), .C(n_479), .D(n_460), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_491), .B(n_452), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_519), .B(n_452), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_519), .B(n_471), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_491), .B(n_476), .Y(n_550) );
INVxp67_ASAP7_75t_L g551 ( .A(n_507), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_494), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_507), .B(n_476), .Y(n_553) );
INVx2_ASAP7_75t_SL g554 ( .A(n_518), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_535), .B(n_482), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_499), .B(n_479), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_499), .B(n_480), .Y(n_557) );
NAND4xp25_ASAP7_75t_L g558 ( .A(n_503), .B(n_467), .C(n_477), .D(n_471), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_501), .B(n_31), .Y(n_559) );
BUFx2_ASAP7_75t_L g560 ( .A(n_518), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_510), .Y(n_561) );
AND2x4_ASAP7_75t_L g562 ( .A(n_518), .B(n_51), .Y(n_562) );
OAI211xp5_ASAP7_75t_SL g563 ( .A1(n_506), .A2(n_339), .B(n_482), .C(n_56), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_501), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_510), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_509), .B(n_52), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_536), .B(n_345), .Y(n_567) );
NAND2x1p5_ASAP7_75t_L g568 ( .A(n_508), .B(n_343), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_489), .B(n_502), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_502), .Y(n_570) );
OAI31xp33_ASAP7_75t_SL g571 ( .A1(n_508), .A2(n_55), .A3(n_57), .B(n_58), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_504), .Y(n_572) );
NAND3xp33_ASAP7_75t_L g573 ( .A(n_532), .B(n_239), .C(n_226), .Y(n_573) );
NOR2xp67_ASAP7_75t_L g574 ( .A(n_503), .B(n_62), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_489), .B(n_343), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_516), .B(n_64), .Y(n_576) );
AND2x2_ASAP7_75t_SL g577 ( .A(n_513), .B(n_343), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_504), .Y(n_578) );
NAND4xp25_ASAP7_75t_SL g579 ( .A(n_520), .B(n_67), .C(n_68), .D(n_69), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_510), .Y(n_580) );
INVx1_ASAP7_75t_SL g581 ( .A(n_492), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_516), .B(n_70), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_505), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_512), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_486), .B(n_71), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_524), .B(n_72), .Y(n_586) );
NAND4xp25_ASAP7_75t_L g587 ( .A(n_528), .B(n_295), .C(n_309), .D(n_310), .Y(n_587) );
NAND2x1p5_ASAP7_75t_L g588 ( .A(n_517), .B(n_343), .Y(n_588) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_520), .A2(n_332), .B(n_274), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_490), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_512), .Y(n_591) );
AND2x4_ASAP7_75t_L g592 ( .A(n_486), .B(n_75), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_490), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_490), .B(n_76), .Y(n_594) );
NAND2xp33_ASAP7_75t_L g595 ( .A(n_484), .B(n_332), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_485), .B(n_290), .Y(n_596) );
NAND2x1p5_ASAP7_75t_L g597 ( .A(n_486), .B(n_274), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_495), .B(n_80), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_590), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_551), .B(n_495), .Y(n_600) );
AOI211xp5_ASAP7_75t_L g601 ( .A1(n_571), .A2(n_533), .B(n_531), .C(n_524), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_548), .B(n_488), .Y(n_602) );
NAND2x1p5_ASAP7_75t_L g603 ( .A(n_562), .B(n_484), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_540), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_552), .B(n_488), .Y(n_605) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_560), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_549), .B(n_542), .Y(n_607) );
OAI21xp5_ASAP7_75t_SL g608 ( .A1(n_571), .A2(n_533), .B(n_531), .Y(n_608) );
AOI211x1_ASAP7_75t_SL g609 ( .A1(n_563), .A2(n_485), .B(n_488), .C(n_514), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_555), .B(n_497), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_564), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_547), .B(n_521), .Y(n_612) );
INVx1_ASAP7_75t_SL g613 ( .A(n_545), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_570), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_550), .B(n_521), .Y(n_615) );
INVx1_ASAP7_75t_SL g616 ( .A(n_545), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_550), .B(n_525), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_539), .B(n_521), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_556), .B(n_526), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_537), .B(n_558), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_572), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_556), .B(n_526), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_561), .B(n_522), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_565), .B(n_522), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_578), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_546), .B(n_497), .Y(n_626) );
NOR2x1_ASAP7_75t_L g627 ( .A(n_574), .B(n_498), .Y(n_627) );
NAND3xp33_ASAP7_75t_L g628 ( .A(n_566), .B(n_523), .C(n_529), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_568), .A2(n_498), .B1(n_495), .B2(n_492), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_580), .B(n_522), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_569), .B(n_498), .Y(n_631) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_554), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_593), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_553), .B(n_526), .Y(n_634) );
OR2x2_ASAP7_75t_L g635 ( .A(n_569), .B(n_527), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_583), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_541), .B(n_523), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_584), .Y(n_638) );
AOI31xp33_ASAP7_75t_SL g639 ( .A1(n_538), .A2(n_534), .A3(n_527), .B(n_523), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_591), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_544), .B(n_529), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_553), .B(n_534), .Y(n_642) );
INVxp67_ASAP7_75t_SL g643 ( .A(n_581), .Y(n_643) );
OR2x2_ASAP7_75t_L g644 ( .A(n_581), .B(n_575), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_557), .B(n_534), .Y(n_645) );
INVxp67_ASAP7_75t_SL g646 ( .A(n_595), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_575), .Y(n_647) );
OR2x2_ASAP7_75t_L g648 ( .A(n_567), .B(n_523), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_557), .B(n_515), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_567), .Y(n_650) );
INVx2_ASAP7_75t_SL g651 ( .A(n_562), .Y(n_651) );
AND4x1_ASAP7_75t_L g652 ( .A(n_585), .B(n_515), .C(n_511), .D(n_323), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_604), .Y(n_653) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_606), .Y(n_654) );
INVx1_ASAP7_75t_SL g655 ( .A(n_632), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_607), .B(n_568), .Y(n_656) );
AND2x4_ASAP7_75t_L g657 ( .A(n_613), .B(n_592), .Y(n_657) );
OAI221xp5_ASAP7_75t_L g658 ( .A1(n_620), .A2(n_626), .B1(n_608), .B2(n_610), .C(n_639), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_619), .B(n_577), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g660 ( .A1(n_637), .A2(n_543), .B(n_579), .Y(n_660) );
NAND2xp33_ASAP7_75t_L g661 ( .A(n_603), .B(n_588), .Y(n_661) );
AOI322xp5_ASAP7_75t_L g662 ( .A1(n_620), .A2(n_582), .A3(n_576), .B1(n_592), .B2(n_586), .C1(n_511), .C2(n_596), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_626), .A2(n_587), .B1(n_573), .B2(n_588), .Y(n_663) );
OAI211xp5_ASAP7_75t_L g664 ( .A1(n_601), .A2(n_589), .B(n_559), .C(n_598), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_610), .B(n_596), .Y(n_665) );
AND3x1_ASAP7_75t_L g666 ( .A(n_651), .B(n_597), .C(n_594), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_611), .Y(n_667) );
NAND3xp33_ASAP7_75t_L g668 ( .A(n_628), .B(n_523), .C(n_196), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_622), .B(n_523), .Y(n_669) );
INVx1_ASAP7_75t_SL g670 ( .A(n_616), .Y(n_670) );
XNOR2xp5_ASAP7_75t_L g671 ( .A(n_652), .B(n_597), .Y(n_671) );
XOR2x2_ASAP7_75t_L g672 ( .A(n_603), .B(n_323), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_612), .B(n_191), .Y(n_673) );
NAND2xp5_ASAP7_75t_SL g674 ( .A(n_627), .B(n_274), .Y(n_674) );
AOI222xp33_ASAP7_75t_L g675 ( .A1(n_650), .A2(n_191), .B1(n_196), .B2(n_204), .C1(n_211), .C2(n_226), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_612), .B(n_191), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_642), .B(n_196), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_645), .B(n_196), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_614), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_642), .B(n_204), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_602), .B(n_204), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_621), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_602), .B(n_204), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_615), .B(n_211), .Y(n_684) );
INVxp67_ASAP7_75t_L g685 ( .A(n_643), .Y(n_685) );
OR2x2_ASAP7_75t_L g686 ( .A(n_617), .B(n_211), .Y(n_686) );
NAND2xp5_ASAP7_75t_SL g687 ( .A(n_646), .B(n_274), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_625), .Y(n_688) );
AOI22x1_ASAP7_75t_L g689 ( .A1(n_609), .A2(n_226), .B1(n_239), .B2(n_304), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_634), .B(n_226), .Y(n_690) );
INVxp67_ASAP7_75t_SL g691 ( .A(n_637), .Y(n_691) );
OAI22xp33_ASAP7_75t_L g692 ( .A1(n_649), .A2(n_290), .B1(n_226), .B2(n_239), .Y(n_692) );
OAI221xp5_ASAP7_75t_L g693 ( .A1(n_644), .A2(n_239), .B1(n_311), .B2(n_256), .C(n_255), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_634), .B(n_641), .Y(n_694) );
AOI22xp33_ASAP7_75t_SL g695 ( .A1(n_629), .A2(n_251), .B1(n_255), .B2(n_282), .Y(n_695) );
OAI21xp5_ASAP7_75t_SL g696 ( .A1(n_617), .A2(n_251), .B(n_255), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_636), .Y(n_697) );
AOI211xp5_ASAP7_75t_L g698 ( .A1(n_635), .A2(n_251), .B(n_282), .C(n_640), .Y(n_698) );
XNOR2x1_ASAP7_75t_L g699 ( .A(n_631), .B(n_251), .Y(n_699) );
OAI22xp33_ASAP7_75t_L g700 ( .A1(n_600), .A2(n_282), .B1(n_647), .B2(n_638), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_633), .Y(n_701) );
OA21x2_ASAP7_75t_L g702 ( .A1(n_648), .A2(n_282), .B(n_647), .Y(n_702) );
OAI221xp5_ASAP7_75t_SL g703 ( .A1(n_648), .A2(n_605), .B1(n_633), .B2(n_599), .C(n_623), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_605), .B(n_618), .Y(n_704) );
AND2x2_ASAP7_75t_L g705 ( .A(n_618), .B(n_623), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_630), .B(n_624), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_624), .B(n_630), .Y(n_707) );
AOI221xp5_ASAP7_75t_L g708 ( .A1(n_599), .A2(n_620), .B1(n_626), .B2(n_607), .C(n_610), .Y(n_708) );
OAI21xp33_ASAP7_75t_L g709 ( .A1(n_620), .A2(n_626), .B(n_571), .Y(n_709) );
NAND3x1_ASAP7_75t_L g710 ( .A(n_620), .B(n_571), .C(n_652), .Y(n_710) );
INVx1_ASAP7_75t_SL g711 ( .A(n_655), .Y(n_711) );
A2O1A1Ixp33_ASAP7_75t_L g712 ( .A1(n_709), .A2(n_658), .B(n_660), .C(n_708), .Y(n_712) );
AOI211xp5_ASAP7_75t_L g713 ( .A1(n_664), .A2(n_696), .B(n_703), .C(n_660), .Y(n_713) );
OAI21xp5_ASAP7_75t_SL g714 ( .A1(n_671), .A2(n_664), .B(n_662), .Y(n_714) );
AND2x4_ASAP7_75t_L g715 ( .A(n_691), .B(n_666), .Y(n_715) );
AOI21xp33_ASAP7_75t_L g716 ( .A1(n_710), .A2(n_686), .B(n_691), .Y(n_716) );
INVx2_ASAP7_75t_L g717 ( .A(n_702), .Y(n_717) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_665), .A2(n_670), .B1(n_663), .B2(n_656), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_654), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_654), .Y(n_720) );
OAI211xp5_ASAP7_75t_L g721 ( .A1(n_698), .A2(n_685), .B(n_689), .C(n_659), .Y(n_721) );
AND2x2_ASAP7_75t_L g722 ( .A(n_694), .B(n_705), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_685), .B(n_697), .Y(n_723) );
NOR2x1_ASAP7_75t_L g724 ( .A(n_661), .B(n_668), .Y(n_724) );
AOI21xp33_ASAP7_75t_SL g725 ( .A1(n_699), .A2(n_700), .B(n_657), .Y(n_725) );
OAI221xp5_ASAP7_75t_L g726 ( .A1(n_712), .A2(n_653), .B1(n_688), .B2(n_667), .C(n_682), .Y(n_726) );
AOI221xp5_ASAP7_75t_L g727 ( .A1(n_716), .A2(n_679), .B1(n_700), .B2(n_669), .C(n_701), .Y(n_727) );
OA22x2_ASAP7_75t_L g728 ( .A1(n_714), .A2(n_704), .B1(n_706), .B2(n_707), .Y(n_728) );
OAI211xp5_ASAP7_75t_L g729 ( .A1(n_716), .A2(n_695), .B(n_675), .C(n_674), .Y(n_729) );
OAI211xp5_ASAP7_75t_SL g730 ( .A1(n_713), .A2(n_687), .B(n_673), .C(n_676), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_711), .Y(n_731) );
AOI211xp5_ASAP7_75t_L g732 ( .A1(n_725), .A2(n_692), .B(n_693), .C(n_683), .Y(n_732) );
OAI211xp5_ASAP7_75t_SL g733 ( .A1(n_718), .A2(n_695), .B(n_680), .C(n_677), .Y(n_733) );
AOI221xp5_ASAP7_75t_L g734 ( .A1(n_726), .A2(n_727), .B1(n_731), .B2(n_730), .C(n_715), .Y(n_734) );
AOI211xp5_ASAP7_75t_L g735 ( .A1(n_729), .A2(n_721), .B(n_720), .C(n_719), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_728), .A2(n_724), .B1(n_723), .B2(n_717), .Y(n_736) );
NOR3xp33_ASAP7_75t_L g737 ( .A(n_733), .B(n_690), .C(n_684), .Y(n_737) );
NOR2xp67_ASAP7_75t_L g738 ( .A(n_736), .B(n_722), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_735), .B(n_732), .Y(n_739) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_734), .A2(n_672), .B1(n_681), .B2(n_678), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_739), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_740), .Y(n_742) );
BUFx2_ASAP7_75t_L g743 ( .A(n_741), .Y(n_743) );
INVxp67_ASAP7_75t_SL g744 ( .A(n_742), .Y(n_744) );
INVxp67_ASAP7_75t_SL g745 ( .A(n_743), .Y(n_745) );
BUFx2_ASAP7_75t_SL g746 ( .A(n_745), .Y(n_746) );
AOI221xp5_ASAP7_75t_L g747 ( .A1(n_746), .A2(n_744), .B1(n_743), .B2(n_737), .C(n_738), .Y(n_747) );
endmodule