module fake_jpeg_1440_n_144 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_144);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_26),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_21),
.B(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_45),
.B(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_53),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_1),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_52),
.B(n_57),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_44),
.B(n_1),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_3),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_2),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_54),
.A2(n_47),
.B1(n_55),
.B2(n_52),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_64),
.B1(n_65),
.B2(n_41),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_62),
.B(n_67),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_55),
.B1(n_47),
.B2(n_40),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_57),
.A2(n_39),
.B1(n_49),
.B2(n_37),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_50),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_40),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_42),
.Y(n_74)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_SL g70 ( 
.A1(n_64),
.A2(n_51),
.B(n_42),
.C(n_49),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_81),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_68),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_72),
.B(n_79),
.Y(n_84)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_74),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_53),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_4),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_78),
.B1(n_61),
.B2(n_43),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_50),
.B1(n_46),
.B2(n_38),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_63),
.B(n_46),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_63),
.B(n_38),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_5),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_70),
.A2(n_62),
.B1(n_61),
.B2(n_66),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_83),
.A2(n_88),
.B1(n_94),
.B2(n_85),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_69),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_77),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_74),
.A2(n_3),
.B(n_4),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_90),
.A2(n_7),
.B(n_8),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_91),
.B(n_92),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_5),
.B(n_6),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_75),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_99),
.B(n_101),
.Y(n_124)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_71),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_81),
.C(n_19),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_103),
.C(n_110),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_88),
.C(n_93),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_96),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_105),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_6),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_25),
.B1(n_32),
.B2(n_31),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_109),
.Y(n_119)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_108),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_95),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_20),
.C(n_33),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_8),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_118),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_SL g117 ( 
.A(n_112),
.B(n_10),
.C(n_12),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_14),
.C(n_16),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_110),
.A2(n_97),
.B1(n_109),
.B2(n_102),
.Y(n_120)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_23),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_121),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_98),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_123),
.A2(n_16),
.B(n_27),
.C(n_28),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_127),
.C(n_131),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_18),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_130),
.A2(n_113),
.B1(n_128),
.B2(n_132),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_30),
.C(n_34),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_122),
.C(n_115),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_134),
.B(n_135),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_119),
.C(n_125),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_117),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_124),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_137),
.C(n_133),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_140),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_141),
.A2(n_125),
.B(n_138),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_130),
.B(n_121),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_116),
.Y(n_144)
);


endmodule