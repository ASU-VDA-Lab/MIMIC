module fake_netlist_6_2446_n_1630 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1630);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1630;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_163;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_148;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_147;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_149;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_L g147 ( 
.A(n_27),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_84),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_124),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_13),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_76),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_83),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_144),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_129),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_69),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_92),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_137),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_74),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_62),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_79),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_66),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_36),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_135),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_37),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_34),
.Y(n_165)
);

BUFx10_ASAP7_75t_L g166 ( 
.A(n_12),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_60),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_0),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_20),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_63),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_95),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_115),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_119),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_96),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_38),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_68),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_18),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_24),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_89),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_71),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_130),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_136),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_20),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_143),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_6),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_6),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_31),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_34),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_41),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_21),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_87),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_107),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_104),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_58),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_27),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_99),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_3),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_112),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_9),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_26),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_105),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_80),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_59),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_94),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_75),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_8),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_106),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_78),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_23),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_142),
.Y(n_211)
);

BUFx10_ASAP7_75t_L g212 ( 
.A(n_86),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_82),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_40),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_91),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_90),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_10),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_38),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_118),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_37),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_127),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_110),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_49),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_49),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_7),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_51),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_88),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_55),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_139),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_48),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_77),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_17),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_31),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_24),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_100),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_50),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_3),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_11),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_32),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_28),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_53),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_35),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_102),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_46),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_93),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_33),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_12),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_36),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_145),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_56),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_126),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_81),
.Y(n_252)
);

BUFx10_ASAP7_75t_L g253 ( 
.A(n_109),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_113),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_98),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_61),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_128),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_19),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_9),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_120),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_141),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_15),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_13),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_42),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_101),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_19),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_15),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_64),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_32),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_138),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_28),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_65),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_21),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_39),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_39),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_122),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_7),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_121),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_11),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_97),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_70),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_33),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_52),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_5),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_42),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_8),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_17),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_26),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_146),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_67),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_2),
.Y(n_291)
);

INVxp67_ASAP7_75t_SL g292 ( 
.A(n_123),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_29),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_114),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_269),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_190),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_190),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_178),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_239),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_239),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_190),
.Y(n_301)
);

INVxp33_ASAP7_75t_SL g302 ( 
.A(n_150),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_205),
.Y(n_303)
);

INVx4_ASAP7_75t_R g304 ( 
.A(n_153),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_190),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_166),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_190),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_209),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_147),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_166),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_147),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_169),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_184),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_188),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_169),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_210),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_210),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_220),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_220),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_170),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_176),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_186),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_191),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_152),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_189),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_198),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_166),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_214),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_150),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_234),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_237),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_196),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_201),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_259),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_264),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_226),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_267),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_241),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_243),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_207),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_273),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_277),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_282),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_284),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_215),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_286),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_291),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_293),
.Y(n_348)
);

INVxp33_ASAP7_75t_SL g349 ( 
.A(n_162),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_159),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_218),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_165),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_167),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_171),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_251),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_268),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_180),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_172),
.Y(n_358)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_212),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_173),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_223),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_224),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_225),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_177),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_194),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_197),
.Y(n_366)
);

INVxp33_ASAP7_75t_SL g367 ( 
.A(n_162),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_164),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_298),
.B(n_313),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_296),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_296),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_295),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_307),
.Y(n_373)
);

NAND3xp33_ASAP7_75t_L g374 ( 
.A(n_299),
.B(n_300),
.C(n_325),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_307),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_352),
.A2(n_271),
.B1(n_247),
.B2(n_232),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_357),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_297),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_298),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_297),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_301),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_313),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_329),
.Y(n_383)
);

AND2x4_ASAP7_75t_L g384 ( 
.A(n_324),
.B(n_153),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_350),
.B(n_229),
.Y(n_385)
);

INVx4_ASAP7_75t_L g386 ( 
.A(n_345),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_314),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_305),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_345),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_355),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_355),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_320),
.Y(n_392)
);

BUFx8_ASAP7_75t_L g393 ( 
.A(n_359),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_345),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_303),
.A2(n_275),
.B1(n_187),
.B2(n_200),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_353),
.B(n_229),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_345),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_345),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_309),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_309),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_308),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_320),
.Y(n_402)
);

NAND2x1p5_ASAP7_75t_L g403 ( 
.A(n_354),
.B(n_156),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_302),
.A2(n_217),
.B1(n_285),
.B2(n_287),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_314),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_311),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_323),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_321),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_358),
.B(n_251),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_360),
.B(n_148),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_364),
.B(n_256),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_311),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_323),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_332),
.B(n_181),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_321),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_312),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_365),
.B(n_256),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_312),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_322),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_315),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g421 ( 
.A(n_332),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_322),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_366),
.B(n_199),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_315),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_336),
.A2(n_258),
.B1(n_164),
.B2(n_274),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_316),
.B(n_208),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_334),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_333),
.B(n_257),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_316),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_334),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_317),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_333),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_340),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_340),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_351),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_317),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_378),
.Y(n_437)
);

BUFx4f_ASAP7_75t_L g438 ( 
.A(n_394),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_378),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_370),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_380),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_414),
.B(n_306),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_384),
.B(n_318),
.Y(n_443)
);

INVx2_ASAP7_75t_SL g444 ( 
.A(n_384),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_370),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_384),
.B(n_351),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_398),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g448 ( 
.A(n_401),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_380),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_384),
.B(n_361),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_418),
.Y(n_451)
);

BUFx10_ASAP7_75t_L g452 ( 
.A(n_369),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_394),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_418),
.Y(n_454)
);

INVx1_ASAP7_75t_SL g455 ( 
.A(n_405),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_371),
.Y(n_456)
);

INVxp33_ASAP7_75t_L g457 ( 
.A(n_372),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_371),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_373),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_428),
.B(n_361),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_373),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_398),
.B(n_362),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_L g463 ( 
.A1(n_426),
.A2(n_302),
.B1(n_367),
.B2(n_349),
.Y(n_463)
);

INVx2_ASAP7_75t_SL g464 ( 
.A(n_403),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_375),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_418),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_403),
.B(n_327),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_394),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_383),
.Y(n_469)
);

INVxp33_ASAP7_75t_L g470 ( 
.A(n_395),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_394),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_418),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_418),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_403),
.B(n_362),
.Y(n_474)
);

AND2x6_ASAP7_75t_L g475 ( 
.A(n_426),
.B(n_215),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_L g476 ( 
.A1(n_426),
.A2(n_349),
.B1(n_367),
.B2(n_343),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_426),
.B(n_390),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_418),
.Y(n_478)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_394),
.Y(n_479)
);

INVx2_ASAP7_75t_SL g480 ( 
.A(n_410),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_398),
.B(n_363),
.Y(n_481)
);

BUFx6f_ASAP7_75t_SL g482 ( 
.A(n_393),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_394),
.Y(n_483)
);

AOI22xp33_ASAP7_75t_L g484 ( 
.A1(n_423),
.A2(n_337),
.B1(n_348),
.B2(n_347),
.Y(n_484)
);

INVxp33_ASAP7_75t_L g485 ( 
.A(n_395),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_381),
.Y(n_486)
);

INVx2_ASAP7_75t_SL g487 ( 
.A(n_410),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_386),
.Y(n_488)
);

INVx1_ASAP7_75t_SL g489 ( 
.A(n_405),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_398),
.B(n_363),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_420),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_420),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_393),
.B(n_368),
.Y(n_493)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_386),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_393),
.B(n_339),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_393),
.B(n_356),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_382),
.B(n_310),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_420),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_420),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_420),
.Y(n_500)
);

INVx2_ASAP7_75t_SL g501 ( 
.A(n_379),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_420),
.Y(n_502)
);

AND3x2_ASAP7_75t_L g503 ( 
.A(n_421),
.B(n_179),
.C(n_292),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_386),
.Y(n_504)
);

INVx5_ASAP7_75t_L g505 ( 
.A(n_386),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_388),
.B(n_270),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_389),
.B(n_182),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_389),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_392),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_389),
.B(n_183),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_397),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_392),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_402),
.B(n_222),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_413),
.B(n_212),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_397),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_397),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_390),
.B(n_318),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_402),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_399),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_408),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_408),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_415),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_399),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_415),
.Y(n_524)
);

INVx2_ASAP7_75t_SL g525 ( 
.A(n_407),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_419),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_391),
.B(n_185),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_419),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_432),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_422),
.Y(n_530)
);

CKINVDCx6p67_ASAP7_75t_R g531 ( 
.A(n_421),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_391),
.B(n_192),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_399),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_422),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_400),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_400),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_R g537 ( 
.A(n_377),
.B(n_338),
.Y(n_537)
);

BUFx2_ASAP7_75t_L g538 ( 
.A(n_434),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_435),
.B(n_212),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_400),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_433),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_406),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_406),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_406),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_427),
.Y(n_545)
);

BUFx6f_ASAP7_75t_SL g546 ( 
.A(n_427),
.Y(n_546)
);

NAND3xp33_ASAP7_75t_L g547 ( 
.A(n_404),
.B(n_346),
.C(n_344),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_412),
.Y(n_548)
);

INVx4_ASAP7_75t_L g549 ( 
.A(n_412),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_412),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_430),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_416),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_416),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_387),
.B(n_385),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_404),
.B(n_253),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_416),
.Y(n_556)
);

OR2x6_ASAP7_75t_L g557 ( 
.A(n_374),
.B(n_396),
.Y(n_557)
);

BUFx10_ASAP7_75t_L g558 ( 
.A(n_430),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_424),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_424),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_424),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_425),
.B(n_253),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_429),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_429),
.Y(n_564)
);

INVx1_ASAP7_75t_SL g565 ( 
.A(n_376),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_425),
.A2(n_376),
.B1(n_149),
.B2(n_151),
.Y(n_566)
);

INVx4_ASAP7_75t_L g567 ( 
.A(n_429),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_431),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_431),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_396),
.B(n_253),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_431),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_436),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_436),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_436),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_409),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_411),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_417),
.Y(n_577)
);

OR2x6_ASAP7_75t_L g578 ( 
.A(n_403),
.B(n_231),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_384),
.B(n_193),
.Y(n_579)
);

INVx5_ASAP7_75t_L g580 ( 
.A(n_394),
.Y(n_580)
);

NOR3xp33_ASAP7_75t_L g581 ( 
.A(n_376),
.B(n_244),
.C(n_246),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_480),
.B(n_149),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_444),
.B(n_480),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_L g584 ( 
.A1(n_487),
.A2(n_255),
.B1(n_294),
.B2(n_272),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_537),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_437),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_487),
.B(n_276),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_437),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_509),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_455),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_464),
.B(n_215),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_575),
.B(n_278),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_575),
.B(n_281),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_576),
.B(n_289),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_576),
.B(n_195),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_460),
.B(n_151),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_464),
.B(n_558),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_558),
.B(n_154),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_446),
.B(n_450),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_501),
.B(n_342),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_SL g601 ( 
.A(n_482),
.B(n_154),
.Y(n_601)
);

INVxp67_ASAP7_75t_L g602 ( 
.A(n_469),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_501),
.B(n_341),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_577),
.B(n_202),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_521),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_554),
.A2(n_477),
.B1(n_443),
.B2(n_578),
.Y(n_606)
);

AND2x4_ASAP7_75t_SL g607 ( 
.A(n_531),
.B(n_558),
.Y(n_607)
);

OR2x2_ASAP7_75t_L g608 ( 
.A(n_489),
.B(n_326),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_577),
.B(n_203),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_521),
.B(n_204),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_521),
.B(n_206),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_442),
.B(n_155),
.Y(n_612)
);

OR2x2_ASAP7_75t_L g613 ( 
.A(n_565),
.B(n_328),
.Y(n_613)
);

INVx6_ASAP7_75t_L g614 ( 
.A(n_558),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_530),
.B(n_155),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_439),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_530),
.B(n_211),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_525),
.B(n_330),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_530),
.B(n_213),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_439),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_579),
.B(n_157),
.Y(n_621)
);

O2A1O1Ixp33_ASAP7_75t_L g622 ( 
.A1(n_557),
.A2(n_335),
.B(n_331),
.C(n_319),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_462),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_512),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_477),
.B(n_216),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_481),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_439),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_443),
.A2(n_252),
.B1(n_215),
.B2(n_287),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_557),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_578),
.A2(n_219),
.B1(n_227),
.B2(n_228),
.Y(n_630)
);

O2A1O1Ixp5_ASAP7_75t_L g631 ( 
.A1(n_518),
.A2(n_319),
.B(n_304),
.C(n_215),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_441),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_520),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_490),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_522),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_525),
.Y(n_636)
);

NAND3xp33_ASAP7_75t_L g637 ( 
.A(n_476),
.B(n_230),
.C(n_233),
.Y(n_637)
);

OR2x2_ASAP7_75t_L g638 ( 
.A(n_529),
.B(n_258),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_524),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_463),
.B(n_157),
.Y(n_640)
);

NOR2x1p5_ASAP7_75t_L g641 ( 
.A(n_531),
.B(n_262),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_555),
.B(n_158),
.Y(n_642)
);

AO221x1_ASAP7_75t_L g643 ( 
.A1(n_524),
.A2(n_252),
.B1(n_262),
.B2(n_263),
.C(n_266),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_526),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_526),
.B(n_235),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_L g646 ( 
.A1(n_578),
.A2(n_249),
.B1(n_245),
.B2(n_250),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_529),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_528),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_578),
.A2(n_254),
.B1(n_158),
.B2(n_283),
.Y(n_649)
);

OAI22x1_ASAP7_75t_R g650 ( 
.A1(n_448),
.A2(n_274),
.B1(n_288),
.B2(n_263),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_441),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_452),
.B(n_160),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_538),
.B(n_236),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_474),
.B(n_290),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_528),
.B(n_534),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_557),
.A2(n_551),
.B1(n_545),
.B2(n_534),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_457),
.B(n_288),
.Y(n_657)
);

BUFx8_ASAP7_75t_L g658 ( 
.A(n_482),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_452),
.B(n_290),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_452),
.B(n_160),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_452),
.B(n_283),
.Y(n_661)
);

NAND2xp33_ASAP7_75t_L g662 ( 
.A(n_475),
.B(n_252),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_441),
.Y(n_663)
);

BUFx6f_ASAP7_75t_SL g664 ( 
.A(n_578),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_557),
.B(n_280),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_545),
.B(n_252),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_449),
.Y(n_667)
);

NOR2x1p5_ASAP7_75t_L g668 ( 
.A(n_547),
.B(n_279),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_557),
.A2(n_252),
.B1(n_279),
.B2(n_266),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_551),
.B(n_280),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_513),
.B(n_72),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_549),
.B(n_265),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_513),
.A2(n_238),
.B1(n_240),
.B2(n_242),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_549),
.B(n_175),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_506),
.B(n_175),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_517),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_447),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_517),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_440),
.B(n_261),
.Y(n_679)
);

INVx4_ASAP7_75t_L g680 ( 
.A(n_494),
.Y(n_680)
);

INVxp67_ASAP7_75t_L g681 ( 
.A(n_497),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_527),
.B(n_261),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_532),
.B(n_467),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_449),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_447),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_449),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_573),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_514),
.B(n_260),
.Y(n_688)
);

O2A1O1Ixp33_ASAP7_75t_L g689 ( 
.A1(n_445),
.A2(n_260),
.B(n_221),
.C(n_174),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_573),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_541),
.B(n_221),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_445),
.B(n_456),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_539),
.B(n_174),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_486),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_456),
.B(n_168),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_458),
.B(n_168),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_458),
.B(n_163),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_573),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_519),
.Y(n_699)
);

NOR2xp67_ASAP7_75t_L g700 ( 
.A(n_566),
.B(n_161),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_570),
.B(n_163),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_503),
.Y(n_702)
);

INVxp67_ASAP7_75t_SL g703 ( 
.A(n_488),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_459),
.B(n_248),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_459),
.B(n_0),
.Y(n_705)
);

BUFx4_ASAP7_75t_L g706 ( 
.A(n_482),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_519),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_513),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_461),
.B(n_140),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_447),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_581),
.B(n_1),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_519),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_535),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_465),
.B(n_4),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_535),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_549),
.B(n_567),
.Y(n_716)
);

NOR2xp67_ASAP7_75t_L g717 ( 
.A(n_493),
.B(n_133),
.Y(n_717)
);

INVx1_ASAP7_75t_SL g718 ( 
.A(n_562),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_535),
.Y(n_719)
);

OAI221xp5_ASAP7_75t_L g720 ( 
.A1(n_484),
.A2(n_10),
.B1(n_14),
.B2(n_16),
.C(n_18),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_540),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_507),
.B(n_14),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_560),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_560),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_546),
.B(n_16),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_561),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_510),
.B(n_22),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_549),
.B(n_54),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_SL g729 ( 
.A(n_482),
.B(n_22),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_572),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_567),
.B(n_57),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_572),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_567),
.B(n_132),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_488),
.B(n_23),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_687),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_606),
.B(n_488),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_590),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_656),
.B(n_488),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_639),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_585),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_608),
.B(n_470),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_599),
.B(n_485),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_687),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_599),
.B(n_567),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_639),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_583),
.B(n_546),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_656),
.B(n_504),
.Y(n_747)
);

NOR3xp33_ASAP7_75t_SL g748 ( 
.A(n_720),
.B(n_496),
.C(n_495),
.Y(n_748)
);

OAI22xp5_ASAP7_75t_L g749 ( 
.A1(n_669),
.A2(n_546),
.B1(n_494),
.B2(n_515),
.Y(n_749)
);

AND2x6_ASAP7_75t_L g750 ( 
.A(n_671),
.B(n_451),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_596),
.B(n_494),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_589),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_R g753 ( 
.A(n_658),
.B(n_546),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_690),
.Y(n_754)
);

INVx5_ASAP7_75t_L g755 ( 
.A(n_680),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_703),
.B(n_623),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_690),
.Y(n_757)
);

OR2x2_ASAP7_75t_L g758 ( 
.A(n_613),
.B(n_508),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_624),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_669),
.A2(n_475),
.B1(n_574),
.B2(n_571),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_626),
.B(n_634),
.Y(n_761)
);

O2A1O1Ixp5_ASAP7_75t_L g762 ( 
.A1(n_592),
.A2(n_515),
.B(n_508),
.C(n_516),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_708),
.A2(n_475),
.B1(n_574),
.B2(n_571),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_633),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_SL g765 ( 
.A1(n_729),
.A2(n_475),
.B1(n_29),
.B2(n_30),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_658),
.Y(n_766)
);

INVx5_ASAP7_75t_L g767 ( 
.A(n_680),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_682),
.B(n_494),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_635),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_600),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_682),
.B(n_523),
.Y(n_771)
);

AND2x6_ASAP7_75t_L g772 ( 
.A(n_671),
.B(n_451),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_644),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_698),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_629),
.A2(n_475),
.B1(n_454),
.B2(n_500),
.Y(n_775)
);

A2O1A1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_708),
.A2(n_665),
.B(n_714),
.C(n_705),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_582),
.B(n_523),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_665),
.A2(n_475),
.B1(n_454),
.B2(n_500),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_582),
.B(n_523),
.Y(n_779)
);

BUFx3_ASAP7_75t_L g780 ( 
.A(n_607),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_681),
.B(n_523),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_677),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_603),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_648),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_586),
.Y(n_785)
);

INVx4_ASAP7_75t_L g786 ( 
.A(n_614),
.Y(n_786)
);

NAND3xp33_ASAP7_75t_SL g787 ( 
.A(n_654),
.B(n_550),
.C(n_540),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_605),
.Y(n_788)
);

O2A1O1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_734),
.A2(n_553),
.B(n_571),
.C(n_569),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_586),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_588),
.Y(n_791)
);

INVx3_ASAP7_75t_L g792 ( 
.A(n_677),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_723),
.Y(n_793)
);

AO21x1_ASAP7_75t_L g794 ( 
.A1(n_731),
.A2(n_473),
.B(n_472),
.Y(n_794)
);

INVx3_ASAP7_75t_L g795 ( 
.A(n_677),
.Y(n_795)
);

BUFx12f_ASAP7_75t_L g796 ( 
.A(n_636),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_676),
.B(n_451),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_678),
.B(n_492),
.Y(n_798)
);

BUFx8_ASAP7_75t_L g799 ( 
.A(n_664),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_677),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_694),
.B(n_492),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_628),
.A2(n_475),
.B1(n_569),
.B2(n_568),
.Y(n_802)
);

HB1xp67_ASAP7_75t_L g803 ( 
.A(n_647),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_718),
.B(n_536),
.Y(n_804)
);

A2O1A1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_705),
.A2(n_552),
.B(n_569),
.C(n_568),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_616),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_618),
.B(n_553),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_685),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_607),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_602),
.B(n_638),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_621),
.B(n_533),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_621),
.B(n_655),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_616),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_724),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_726),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_657),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_664),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_692),
.B(n_595),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_620),
.Y(n_819)
);

BUFx3_ASAP7_75t_L g820 ( 
.A(n_685),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_604),
.B(n_453),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_620),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_609),
.B(n_453),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_695),
.B(n_453),
.Y(n_824)
);

NOR3xp33_ASAP7_75t_SL g825 ( 
.A(n_640),
.B(n_25),
.C(n_30),
.Y(n_825)
);

BUFx6f_ASAP7_75t_L g826 ( 
.A(n_685),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_627),
.Y(n_827)
);

INVx3_ASAP7_75t_L g828 ( 
.A(n_685),
.Y(n_828)
);

INVx1_ASAP7_75t_SL g829 ( 
.A(n_653),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_652),
.Y(n_830)
);

INVx4_ASAP7_75t_L g831 ( 
.A(n_614),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_668),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_625),
.B(n_542),
.Y(n_833)
);

BUFx2_ASAP7_75t_L g834 ( 
.A(n_711),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_696),
.B(n_615),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_627),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_683),
.A2(n_654),
.B1(n_642),
.B2(n_612),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_612),
.B(n_542),
.Y(n_838)
);

NOR3xp33_ASAP7_75t_SL g839 ( 
.A(n_637),
.B(n_25),
.C(n_35),
.Y(n_839)
);

BUFx3_ASAP7_75t_L g840 ( 
.A(n_710),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_730),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_732),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_696),
.B(n_615),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_632),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_642),
.B(n_542),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_614),
.A2(n_508),
.B1(n_511),
.B2(n_515),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_587),
.B(n_659),
.Y(n_847)
);

INVx2_ASAP7_75t_SL g848 ( 
.A(n_702),
.Y(n_848)
);

AND2x6_ASAP7_75t_L g849 ( 
.A(n_725),
.B(n_473),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_593),
.B(n_483),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_594),
.B(n_483),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_660),
.B(n_559),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_710),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_651),
.Y(n_854)
);

INVxp67_ASAP7_75t_L g855 ( 
.A(n_714),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_663),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_661),
.B(n_559),
.Y(n_857)
);

OAI22xp33_ASAP7_75t_L g858 ( 
.A1(n_717),
.A2(n_543),
.B1(n_568),
.B2(n_564),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_663),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_667),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_628),
.B(n_468),
.Y(n_861)
);

HB1xp67_ASAP7_75t_L g862 ( 
.A(n_710),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_SL g863 ( 
.A1(n_688),
.A2(n_475),
.B1(n_41),
.B2(n_43),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_704),
.B(n_483),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_SL g865 ( 
.A1(n_693),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_865)
);

AND3x1_ASAP7_75t_L g866 ( 
.A(n_693),
.B(n_511),
.C(n_516),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_667),
.Y(n_867)
);

OR2x2_ASAP7_75t_L g868 ( 
.A(n_691),
.B(n_516),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_709),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_716),
.A2(n_438),
.B(n_505),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_597),
.A2(n_511),
.B1(n_491),
.B2(n_502),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_643),
.A2(n_552),
.B1(n_564),
.B2(n_563),
.Y(n_872)
);

AND2x4_ASAP7_75t_SL g873 ( 
.A(n_630),
.B(n_472),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_684),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_641),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_684),
.Y(n_876)
);

INVx5_ASAP7_75t_L g877 ( 
.A(n_686),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_649),
.Y(n_878)
);

INVx5_ASAP7_75t_L g879 ( 
.A(n_686),
.Y(n_879)
);

INVxp67_ASAP7_75t_SL g880 ( 
.A(n_699),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_699),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_728),
.Y(n_882)
);

AND2x6_ASAP7_75t_SL g883 ( 
.A(n_725),
.B(n_44),
.Y(n_883)
);

BUFx3_ASAP7_75t_L g884 ( 
.A(n_707),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_645),
.B(n_471),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_733),
.B(n_622),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_707),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_712),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_679),
.B(n_471),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_731),
.A2(n_673),
.B1(n_727),
.B2(n_722),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_697),
.B(n_468),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_610),
.B(n_540),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_670),
.Y(n_893)
);

OAI22xp5_ASAP7_75t_L g894 ( 
.A1(n_835),
.A2(n_673),
.B1(n_646),
.B2(n_619),
.Y(n_894)
);

INVx5_ASAP7_75t_L g895 ( 
.A(n_796),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_L g896 ( 
.A1(n_843),
.A2(n_700),
.B1(n_670),
.B2(n_584),
.Y(n_896)
);

A2O1A1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_837),
.A2(n_776),
.B(n_742),
.C(n_847),
.Y(n_897)
);

A2O1A1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_776),
.A2(n_689),
.B(n_598),
.C(n_631),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_742),
.A2(n_890),
.B1(n_893),
.B2(n_849),
.Y(n_899)
);

O2A1O1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_855),
.A2(n_675),
.B(n_701),
.C(n_591),
.Y(n_900)
);

XOR2x2_ASAP7_75t_SL g901 ( 
.A(n_765),
.B(n_650),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_741),
.B(n_611),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_R g903 ( 
.A(n_740),
.B(n_817),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_744),
.A2(n_438),
.B(n_591),
.Y(n_904)
);

O2A1O1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_855),
.A2(n_672),
.B(n_674),
.C(n_617),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_752),
.Y(n_906)
);

A2O1A1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_847),
.A2(n_674),
.B(n_672),
.C(n_601),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_737),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_812),
.B(n_721),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_818),
.B(n_721),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_829),
.B(n_719),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_770),
.B(n_719),
.Y(n_912)
);

INVx1_ASAP7_75t_SL g913 ( 
.A(n_737),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_782),
.Y(n_914)
);

AO32x2_ASAP7_75t_L g915 ( 
.A1(n_749),
.A2(n_479),
.A3(n_666),
.B1(n_712),
.B2(n_713),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_750),
.A2(n_662),
.B1(n_715),
.B2(n_713),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_768),
.A2(n_438),
.B(n_505),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_759),
.Y(n_918)
);

OR2x6_ASAP7_75t_SL g919 ( 
.A(n_878),
.B(n_706),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_782),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_807),
.B(n_543),
.Y(n_921)
);

INVx4_ASAP7_75t_L g922 ( 
.A(n_786),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_764),
.Y(n_923)
);

O2A1O1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_748),
.A2(n_543),
.B(n_564),
.C(n_563),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_769),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_783),
.B(n_542),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_763),
.A2(n_559),
.B1(n_472),
.B2(n_466),
.Y(n_927)
);

CKINVDCx20_ASAP7_75t_R g928 ( 
.A(n_753),
.Y(n_928)
);

INVx4_ASAP7_75t_L g929 ( 
.A(n_786),
.Y(n_929)
);

OR2x2_ASAP7_75t_SL g930 ( 
.A(n_803),
.B(n_466),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_782),
.Y(n_931)
);

OA22x2_ASAP7_75t_L g932 ( 
.A1(n_832),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_799),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_763),
.A2(n_559),
.B1(n_473),
.B2(n_466),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_803),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_766),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_761),
.B(n_491),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_756),
.B(n_550),
.Y(n_938)
);

OR2x2_ASAP7_75t_L g939 ( 
.A(n_758),
.B(n_552),
.Y(n_939)
);

AOI21xp33_ASAP7_75t_L g940 ( 
.A1(n_890),
.A2(n_478),
.B(n_491),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_781),
.B(n_553),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_773),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_784),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_781),
.B(n_739),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_810),
.B(n_478),
.Y(n_945)
);

A2O1A1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_748),
.A2(n_502),
.B(n_498),
.C(n_499),
.Y(n_946)
);

BUFx4f_ASAP7_75t_L g947 ( 
.A(n_849),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_745),
.B(n_548),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_751),
.A2(n_580),
.B(n_478),
.Y(n_949)
);

HB1xp67_ASAP7_75t_SL g950 ( 
.A(n_799),
.Y(n_950)
);

AOI22xp5_ASAP7_75t_L g951 ( 
.A1(n_750),
.A2(n_544),
.B1(n_563),
.B2(n_556),
.Y(n_951)
);

NAND3xp33_ASAP7_75t_SL g952 ( 
.A(n_830),
.B(n_498),
.C(n_499),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_793),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_780),
.B(n_499),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_884),
.Y(n_955)
);

O2A1O1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_816),
.A2(n_825),
.B(n_839),
.C(n_746),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_750),
.A2(n_556),
.B1(n_548),
.B2(n_544),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_782),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_808),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_814),
.Y(n_960)
);

INVxp67_ASAP7_75t_L g961 ( 
.A(n_834),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_SL g962 ( 
.A(n_831),
.B(n_498),
.Y(n_962)
);

INVx3_ASAP7_75t_L g963 ( 
.A(n_808),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_815),
.Y(n_964)
);

NOR3xp33_ASAP7_75t_L g965 ( 
.A(n_848),
.B(n_556),
.C(n_544),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_808),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_808),
.Y(n_967)
);

OR2x6_ASAP7_75t_L g968 ( 
.A(n_780),
.B(n_103),
.Y(n_968)
);

O2A1O1Ixp5_ASAP7_75t_SL g969 ( 
.A1(n_886),
.A2(n_45),
.B(n_47),
.C(n_48),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_884),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_738),
.A2(n_580),
.B(n_73),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_809),
.B(n_116),
.Y(n_972)
);

AND2x6_ASAP7_75t_L g973 ( 
.A(n_869),
.B(n_85),
.Y(n_973)
);

BUFx3_ASAP7_75t_L g974 ( 
.A(n_809),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_841),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_826),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_842),
.Y(n_977)
);

BUFx2_ASAP7_75t_L g978 ( 
.A(n_788),
.Y(n_978)
);

BUFx2_ASAP7_75t_L g979 ( 
.A(n_788),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_844),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_833),
.A2(n_108),
.B(n_111),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_738),
.A2(n_117),
.B(n_125),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_804),
.B(n_50),
.Y(n_983)
);

AOI221xp5_ASAP7_75t_L g984 ( 
.A1(n_863),
.A2(n_131),
.B1(n_765),
.B2(n_825),
.C(n_839),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_747),
.A2(n_767),
.B(n_755),
.Y(n_985)
);

OR2x6_ASAP7_75t_L g986 ( 
.A(n_831),
.B(n_826),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_736),
.A2(n_804),
.B(n_805),
.C(n_747),
.Y(n_987)
);

BUFx2_ASAP7_75t_L g988 ( 
.A(n_753),
.Y(n_988)
);

CKINVDCx8_ASAP7_75t_R g989 ( 
.A(n_875),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_859),
.Y(n_990)
);

OR2x2_ASAP7_75t_L g991 ( 
.A(n_868),
.B(n_797),
.Y(n_991)
);

NOR3xp33_ASAP7_75t_SL g992 ( 
.A(n_883),
.B(n_865),
.C(n_852),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_838),
.A2(n_845),
.B1(n_760),
.B2(n_771),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_L g994 ( 
.A1(n_750),
.A2(n_772),
.B1(n_863),
.B2(n_849),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_838),
.B(n_845),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_820),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_887),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_826),
.Y(n_998)
);

INVx3_ASAP7_75t_SL g999 ( 
.A(n_849),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_821),
.A2(n_823),
.B(n_892),
.Y(n_1000)
);

A2O1A1Ixp33_ASAP7_75t_SL g1001 ( 
.A1(n_852),
.A2(n_857),
.B(n_872),
.C(n_811),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_820),
.Y(n_1002)
);

BUFx2_ASAP7_75t_SL g1003 ( 
.A(n_840),
.Y(n_1003)
);

NAND2x1p5_ASAP7_75t_L g1004 ( 
.A(n_840),
.B(n_792),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_792),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_862),
.B(n_869),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_860),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_862),
.B(n_798),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_857),
.A2(n_864),
.B(n_889),
.C(n_891),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_885),
.A2(n_870),
.B(n_880),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_772),
.B(n_880),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_887),
.Y(n_1012)
);

OAI21x1_ASAP7_75t_L g1013 ( 
.A1(n_762),
.A2(n_789),
.B(n_871),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_R g1014 ( 
.A(n_795),
.B(n_800),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_R g1015 ( 
.A(n_795),
.B(n_800),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_850),
.A2(n_851),
.B(n_802),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_760),
.A2(n_802),
.B1(n_861),
.B2(n_824),
.Y(n_1017)
);

INVx5_ASAP7_75t_L g1018 ( 
.A(n_986),
.Y(n_1018)
);

AOI21xp33_ASAP7_75t_SL g1019 ( 
.A1(n_932),
.A2(n_872),
.B(n_853),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_1005),
.Y(n_1020)
);

AOI22xp33_ASAP7_75t_SL g1021 ( 
.A1(n_894),
.A2(n_873),
.B1(n_882),
.B2(n_777),
.Y(n_1021)
);

AOI221xp5_ASAP7_75t_L g1022 ( 
.A1(n_984),
.A2(n_866),
.B1(n_787),
.B2(n_858),
.C(n_779),
.Y(n_1022)
);

AOI221x1_ASAP7_75t_L g1023 ( 
.A1(n_907),
.A2(n_882),
.B1(n_846),
.B2(n_876),
.C(n_867),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_896),
.A2(n_778),
.B(n_775),
.C(n_801),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_908),
.Y(n_1025)
);

BUFx3_ASAP7_75t_L g1026 ( 
.A(n_974),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_902),
.B(n_961),
.Y(n_1027)
);

OAI21xp33_ASAP7_75t_L g1028 ( 
.A1(n_983),
.A2(n_992),
.B(n_899),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_1005),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_903),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_900),
.A2(n_882),
.B(n_743),
.C(n_754),
.Y(n_1031)
);

NOR2x1_ASAP7_75t_SL g1032 ( 
.A(n_986),
.B(n_879),
.Y(n_1032)
);

OAI21xp33_ASAP7_75t_SL g1033 ( 
.A1(n_994),
.A2(n_971),
.B(n_995),
.Y(n_1033)
);

AO21x2_ASAP7_75t_L g1034 ( 
.A1(n_1001),
.A2(n_881),
.B(n_757),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_1000),
.A2(n_882),
.B(n_879),
.Y(n_1035)
);

OAI21x1_ASAP7_75t_L g1036 ( 
.A1(n_949),
.A2(n_827),
.B(n_874),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_909),
.B(n_735),
.Y(n_1037)
);

INVx1_ASAP7_75t_SL g1038 ( 
.A(n_913),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_931),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_918),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_931),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_911),
.B(n_774),
.Y(n_1042)
);

AO31x2_ASAP7_75t_L g1043 ( 
.A1(n_993),
.A2(n_898),
.A3(n_1009),
.B(n_946),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_945),
.B(n_785),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_910),
.B(n_790),
.Y(n_1045)
);

OAI21x1_ASAP7_75t_SL g1046 ( 
.A1(n_994),
.A2(n_791),
.B(n_806),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_1008),
.B(n_879),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_935),
.Y(n_1048)
);

INVx1_ASAP7_75t_SL g1049 ( 
.A(n_978),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_923),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_979),
.B(n_853),
.Y(n_1051)
);

INVxp67_ASAP7_75t_SL g1052 ( 
.A(n_1006),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_925),
.Y(n_1053)
);

AOI21x1_ASAP7_75t_L g1054 ( 
.A1(n_904),
.A2(n_813),
.B(n_819),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_895),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_905),
.A2(n_822),
.B(n_856),
.C(n_836),
.Y(n_1056)
);

BUFx10_ASAP7_75t_L g1057 ( 
.A(n_936),
.Y(n_1057)
);

AOI221xp5_ASAP7_75t_SL g1058 ( 
.A1(n_956),
.A2(n_854),
.B1(n_888),
.B2(n_828),
.C(n_877),
.Y(n_1058)
);

AOI21x1_ASAP7_75t_L g1059 ( 
.A1(n_1016),
.A2(n_877),
.B(n_828),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_1008),
.B(n_888),
.Y(n_1060)
);

CKINVDCx14_ASAP7_75t_R g1061 ( 
.A(n_919),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_944),
.B(n_937),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_991),
.B(n_912),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_942),
.B(n_943),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_917),
.A2(n_924),
.B(n_987),
.Y(n_1065)
);

AO31x2_ASAP7_75t_L g1066 ( 
.A1(n_1017),
.A2(n_934),
.A3(n_927),
.B(n_941),
.Y(n_1066)
);

INVx2_ASAP7_75t_SL g1067 ( 
.A(n_895),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_955),
.B(n_970),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_953),
.Y(n_1069)
);

OAI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_940),
.A2(n_969),
.B(n_982),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_960),
.B(n_964),
.Y(n_1071)
);

OAI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_981),
.A2(n_951),
.B(n_957),
.Y(n_1072)
);

AO31x2_ASAP7_75t_L g1073 ( 
.A1(n_1011),
.A2(n_915),
.A3(n_938),
.B(n_990),
.Y(n_1073)
);

OAI21x1_ASAP7_75t_L g1074 ( 
.A1(n_948),
.A2(n_921),
.B(n_916),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_901),
.B(n_947),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_975),
.B(n_977),
.Y(n_1076)
);

NOR4xp25_ASAP7_75t_L g1077 ( 
.A(n_952),
.B(n_1007),
.C(n_980),
.D(n_926),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_962),
.A2(n_986),
.B(n_939),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_895),
.Y(n_1079)
);

OA22x2_ASAP7_75t_L g1080 ( 
.A1(n_968),
.A2(n_972),
.B1(n_988),
.B2(n_999),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_931),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_916),
.A2(n_914),
.B(n_963),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_997),
.B(n_1012),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_922),
.A2(n_929),
.B(n_954),
.Y(n_1084)
);

NAND3xp33_ASAP7_75t_L g1085 ( 
.A(n_965),
.B(n_968),
.C(n_954),
.Y(n_1085)
);

AO31x2_ASAP7_75t_L g1086 ( 
.A1(n_915),
.A2(n_922),
.A3(n_929),
.B(n_930),
.Y(n_1086)
);

OR2x2_ASAP7_75t_L g1087 ( 
.A(n_996),
.B(n_1002),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_1004),
.A2(n_958),
.B(n_920),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_958),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_959),
.A2(n_998),
.B(n_967),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_SL g1091 ( 
.A1(n_973),
.A2(n_968),
.B(n_1015),
.Y(n_1091)
);

BUFx2_ASAP7_75t_L g1092 ( 
.A(n_1014),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_1005),
.B(n_989),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_959),
.A2(n_967),
.B(n_963),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_915),
.A2(n_973),
.B(n_1003),
.Y(n_1095)
);

OA22x2_ASAP7_75t_L g1096 ( 
.A1(n_950),
.A2(n_973),
.B1(n_933),
.B2(n_928),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_973),
.B(n_966),
.Y(n_1097)
);

AO31x2_ASAP7_75t_L g1098 ( 
.A1(n_966),
.A2(n_993),
.A3(n_776),
.B(n_805),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_976),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_897),
.B(n_742),
.Y(n_1100)
);

INVx2_ASAP7_75t_SL g1101 ( 
.A(n_908),
.Y(n_1101)
);

BUFx2_ASAP7_75t_L g1102 ( 
.A(n_908),
.Y(n_1102)
);

OA22x2_ASAP7_75t_L g1103 ( 
.A1(n_901),
.A2(n_566),
.B1(n_395),
.B2(n_376),
.Y(n_1103)
);

OAI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_897),
.A2(n_995),
.B(n_776),
.Y(n_1104)
);

AO31x2_ASAP7_75t_L g1105 ( 
.A1(n_993),
.A2(n_776),
.A3(n_805),
.B(n_794),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_897),
.B(n_742),
.Y(n_1106)
);

AO31x2_ASAP7_75t_L g1107 ( 
.A1(n_993),
.A2(n_776),
.A3(n_805),
.B(n_794),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_903),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_902),
.B(n_742),
.Y(n_1109)
);

INVx5_ASAP7_75t_L g1110 ( 
.A(n_986),
.Y(n_1110)
);

NAND2x1_ASAP7_75t_L g1111 ( 
.A(n_986),
.B(n_750),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_902),
.B(n_742),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_897),
.B(n_742),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_897),
.B(n_742),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_1010),
.A2(n_985),
.B(n_1013),
.Y(n_1115)
);

AOI221x1_ASAP7_75t_L g1116 ( 
.A1(n_897),
.A2(n_776),
.B1(n_907),
.B2(n_894),
.C(n_843),
.Y(n_1116)
);

INVx6_ASAP7_75t_SL g1117 ( 
.A(n_968),
.Y(n_1117)
);

OAI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_897),
.A2(n_995),
.B(n_776),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_908),
.B(n_829),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_897),
.B(n_742),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_1010),
.A2(n_985),
.B(n_1013),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_906),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_908),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_902),
.B(n_742),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_897),
.B(n_742),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_906),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_1010),
.A2(n_985),
.B(n_1013),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_906),
.Y(n_1128)
);

OR2x2_ASAP7_75t_L g1129 ( 
.A(n_913),
.B(n_741),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_906),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_897),
.B(n_742),
.Y(n_1131)
);

NAND2x1p5_ASAP7_75t_L g1132 ( 
.A(n_947),
.B(n_786),
.Y(n_1132)
);

INVxp67_ASAP7_75t_SL g1133 ( 
.A(n_935),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1010),
.A2(n_985),
.B(n_1013),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_931),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_1010),
.A2(n_985),
.B(n_1013),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_SL g1137 ( 
.A1(n_994),
.A2(n_982),
.B(n_985),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_995),
.A2(n_1000),
.B(n_744),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_906),
.Y(n_1139)
);

A2O1A1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_897),
.A2(n_837),
.B(n_776),
.C(n_835),
.Y(n_1140)
);

NOR2xp67_ASAP7_75t_L g1141 ( 
.A(n_961),
.B(n_602),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_906),
.Y(n_1142)
);

O2A1O1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_1028),
.A2(n_1112),
.B(n_1140),
.C(n_1120),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_SL g1144 ( 
.A1(n_1091),
.A2(n_1032),
.B(n_1046),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_1100),
.B(n_1106),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1071),
.Y(n_1146)
);

AND2x4_ASAP7_75t_L g1147 ( 
.A(n_1060),
.B(n_1018),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1071),
.Y(n_1148)
);

NAND2x1p5_ASAP7_75t_L g1149 ( 
.A(n_1018),
.B(n_1110),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1109),
.B(n_1124),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1134),
.A2(n_1136),
.B(n_1054),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1059),
.A2(n_1036),
.B(n_1035),
.Y(n_1152)
);

OA21x2_ASAP7_75t_L g1153 ( 
.A1(n_1023),
.A2(n_1065),
.B(n_1116),
.Y(n_1153)
);

OA21x2_ASAP7_75t_L g1154 ( 
.A1(n_1070),
.A2(n_1095),
.B(n_1138),
.Y(n_1154)
);

AO21x2_ASAP7_75t_L g1155 ( 
.A1(n_1070),
.A2(n_1137),
.B(n_1118),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_1018),
.B(n_1110),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1050),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1076),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_1018),
.Y(n_1159)
);

BUFx4f_ASAP7_75t_SL g1160 ( 
.A(n_1117),
.Y(n_1160)
);

OAI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_1103),
.A2(n_1106),
.B1(n_1113),
.B2(n_1131),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1063),
.B(n_1051),
.Y(n_1162)
);

HB1xp67_ASAP7_75t_L g1163 ( 
.A(n_1098),
.Y(n_1163)
);

OR2x2_ASAP7_75t_L g1164 ( 
.A(n_1129),
.B(n_1063),
.Y(n_1164)
);

NAND2x1p5_ASAP7_75t_L g1165 ( 
.A(n_1110),
.B(n_1111),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_1102),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_1100),
.B(n_1113),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1114),
.A2(n_1131),
.B(n_1125),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1052),
.B(n_1027),
.Y(n_1169)
);

NAND2x1p5_ASAP7_75t_L g1170 ( 
.A(n_1110),
.B(n_1047),
.Y(n_1170)
);

AO21x2_ASAP7_75t_L g1171 ( 
.A1(n_1104),
.A2(n_1118),
.B(n_1077),
.Y(n_1171)
);

AO21x2_ASAP7_75t_L g1172 ( 
.A1(n_1104),
.A2(n_1077),
.B(n_1072),
.Y(n_1172)
);

NAND3xp33_ASAP7_75t_L g1173 ( 
.A(n_1114),
.B(n_1120),
.C(n_1085),
.Y(n_1173)
);

OR2x2_ASAP7_75t_L g1174 ( 
.A(n_1049),
.B(n_1068),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_SL g1175 ( 
.A1(n_1103),
.A2(n_1061),
.B1(n_1080),
.B2(n_1096),
.Y(n_1175)
);

AOI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_1033),
.A2(n_1080),
.B1(n_1022),
.B2(n_1075),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_1082),
.A2(n_1074),
.B(n_1072),
.Y(n_1177)
);

CKINVDCx11_ASAP7_75t_R g1178 ( 
.A(n_1057),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1126),
.Y(n_1179)
);

AOI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1096),
.A2(n_1085),
.B1(n_1141),
.B2(n_1119),
.Y(n_1180)
);

AO21x2_ASAP7_75t_L g1181 ( 
.A1(n_1031),
.A2(n_1056),
.B(n_1024),
.Y(n_1181)
);

OAI222xp33_ASAP7_75t_L g1182 ( 
.A1(n_1049),
.A2(n_1038),
.B1(n_1062),
.B2(n_1042),
.C1(n_1021),
.C2(n_1133),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1076),
.Y(n_1183)
);

OAI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1062),
.A2(n_1078),
.B(n_1044),
.Y(n_1184)
);

INVx1_ASAP7_75t_SL g1185 ( 
.A(n_1038),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_SL g1186 ( 
.A1(n_1019),
.A2(n_1097),
.B(n_1088),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1064),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1040),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_1048),
.B(n_1025),
.Y(n_1189)
);

INVx1_ASAP7_75t_SL g1190 ( 
.A(n_1087),
.Y(n_1190)
);

OA21x2_ASAP7_75t_L g1191 ( 
.A1(n_1058),
.A2(n_1037),
.B(n_1045),
.Y(n_1191)
);

BUFx4f_ASAP7_75t_L g1192 ( 
.A(n_1132),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_1123),
.Y(n_1193)
);

BUFx12f_ASAP7_75t_L g1194 ( 
.A(n_1057),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1117),
.A2(n_1142),
.B1(n_1139),
.B2(n_1053),
.Y(n_1195)
);

O2A1O1Ixp33_ASAP7_75t_SL g1196 ( 
.A1(n_1097),
.A2(n_1037),
.B(n_1045),
.C(n_1089),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1069),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1122),
.Y(n_1198)
);

OR2x6_ASAP7_75t_L g1199 ( 
.A(n_1132),
.B(n_1084),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1128),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1090),
.A2(n_1094),
.B(n_1083),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_1020),
.B(n_1029),
.Y(n_1202)
);

AND2x4_ASAP7_75t_L g1203 ( 
.A(n_1020),
.B(n_1029),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1130),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1034),
.A2(n_1066),
.B(n_1043),
.Y(n_1205)
);

OR2x6_ASAP7_75t_L g1206 ( 
.A(n_1093),
.B(n_1067),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1099),
.A2(n_1098),
.B(n_1034),
.Y(n_1207)
);

AO21x2_ASAP7_75t_L g1208 ( 
.A1(n_1043),
.A2(n_1066),
.B(n_1107),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1101),
.A2(n_1092),
.B1(n_1030),
.B2(n_1108),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1055),
.A2(n_1079),
.B(n_1066),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_1086),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1105),
.A2(n_1107),
.B(n_1073),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1105),
.A2(n_1073),
.B(n_1086),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1039),
.B(n_1041),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1081),
.Y(n_1215)
);

AO21x2_ASAP7_75t_L g1216 ( 
.A1(n_1081),
.A2(n_1070),
.B(n_1059),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1135),
.B(n_1112),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1135),
.A2(n_1121),
.B(n_1115),
.Y(n_1218)
);

AOI21xp33_ASAP7_75t_L g1219 ( 
.A1(n_1112),
.A2(n_843),
.B(n_835),
.Y(n_1219)
);

INVxp67_ASAP7_75t_SL g1220 ( 
.A(n_1058),
.Y(n_1220)
);

INVx2_ASAP7_75t_SL g1221 ( 
.A(n_1087),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1112),
.A2(n_1028),
.B1(n_1103),
.B2(n_1100),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1112),
.A2(n_1028),
.B1(n_1103),
.B2(n_1100),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1054),
.A2(n_1121),
.B(n_1115),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1054),
.A2(n_1121),
.B(n_1115),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1060),
.B(n_1018),
.Y(n_1226)
);

INVx2_ASAP7_75t_SL g1227 ( 
.A(n_1087),
.Y(n_1227)
);

INVx5_ASAP7_75t_L g1228 ( 
.A(n_1018),
.Y(n_1228)
);

AND2x4_ASAP7_75t_L g1229 ( 
.A(n_1060),
.B(n_1018),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1071),
.Y(n_1230)
);

NAND3xp33_ASAP7_75t_SL g1231 ( 
.A(n_1112),
.B(n_837),
.C(n_460),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_SL g1232 ( 
.A1(n_1061),
.A2(n_1112),
.B1(n_395),
.B2(n_830),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_SL g1233 ( 
.A1(n_1091),
.A2(n_1032),
.B(n_1046),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1050),
.Y(n_1234)
);

AOI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1112),
.A2(n_308),
.B1(n_336),
.B2(n_303),
.Y(n_1235)
);

HB1xp67_ASAP7_75t_L g1236 ( 
.A(n_1098),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1115),
.A2(n_1127),
.B(n_1121),
.Y(n_1237)
);

OAI222xp33_ASAP7_75t_L g1238 ( 
.A1(n_1103),
.A2(n_865),
.B1(n_669),
.B2(n_765),
.C1(n_863),
.C2(n_837),
.Y(n_1238)
);

O2A1O1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1028),
.A2(n_897),
.B(n_776),
.C(n_843),
.Y(n_1239)
);

A2O1A1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_1140),
.A2(n_776),
.B(n_897),
.C(n_742),
.Y(n_1240)
);

OR2x6_ASAP7_75t_L g1241 ( 
.A(n_1091),
.B(n_1080),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1071),
.Y(n_1242)
);

BUFx4f_ASAP7_75t_SL g1243 ( 
.A(n_1117),
.Y(n_1243)
);

OA21x2_ASAP7_75t_L g1244 ( 
.A1(n_1023),
.A2(n_1065),
.B(n_1116),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1112),
.B(n_1109),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1054),
.A2(n_1121),
.B(n_1115),
.Y(n_1246)
);

AOI21xp33_ASAP7_75t_L g1247 ( 
.A1(n_1112),
.A2(n_843),
.B(n_835),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1026),
.Y(n_1248)
);

AOI21xp33_ASAP7_75t_SL g1249 ( 
.A1(n_1103),
.A2(n_377),
.B(n_585),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1050),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1109),
.B(n_1124),
.Y(n_1251)
);

A2O1A1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_1140),
.A2(n_776),
.B(n_897),
.C(n_742),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1054),
.A2(n_1121),
.B(n_1115),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1112),
.B(n_1109),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1054),
.A2(n_1121),
.B(n_1115),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1109),
.B(n_1124),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1050),
.Y(n_1257)
);

AO21x1_ASAP7_75t_L g1258 ( 
.A1(n_1100),
.A2(n_843),
.B(n_835),
.Y(n_1258)
);

OR2x2_ASAP7_75t_L g1259 ( 
.A(n_1164),
.B(n_1174),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_SL g1260 ( 
.A1(n_1240),
.A2(n_1252),
.B(n_1156),
.Y(n_1260)
);

AND2x4_ASAP7_75t_L g1261 ( 
.A(n_1147),
.B(n_1226),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1222),
.A2(n_1223),
.B1(n_1175),
.B2(n_1176),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_1178),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_1178),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_1248),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1167),
.B(n_1168),
.Y(n_1266)
);

O2A1O1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1238),
.A2(n_1219),
.B(n_1247),
.C(n_1231),
.Y(n_1267)
);

CKINVDCx20_ASAP7_75t_R g1268 ( 
.A(n_1160),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_SL g1269 ( 
.A1(n_1232),
.A2(n_1223),
.B1(n_1222),
.B2(n_1176),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_SL g1270 ( 
.A1(n_1240),
.A2(n_1252),
.B(n_1156),
.Y(n_1270)
);

OR2x2_ASAP7_75t_L g1271 ( 
.A(n_1162),
.B(n_1190),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1167),
.B(n_1146),
.Y(n_1272)
);

O2A1O1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1143),
.A2(n_1239),
.B(n_1161),
.C(n_1182),
.Y(n_1273)
);

OR2x2_ASAP7_75t_L g1274 ( 
.A(n_1150),
.B(n_1169),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1220),
.A2(n_1184),
.B(n_1181),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1220),
.A2(n_1181),
.B(n_1145),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_1194),
.Y(n_1277)
);

AOI221x1_ASAP7_75t_SL g1278 ( 
.A1(n_1161),
.A2(n_1245),
.B1(n_1254),
.B2(n_1173),
.C(n_1187),
.Y(n_1278)
);

AOI221x1_ASAP7_75t_SL g1279 ( 
.A1(n_1217),
.A2(n_1189),
.B1(n_1183),
.B2(n_1158),
.C(n_1148),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1251),
.B(n_1256),
.Y(n_1280)
);

BUFx4f_ASAP7_75t_L g1281 ( 
.A(n_1194),
.Y(n_1281)
);

HB1xp67_ASAP7_75t_L g1282 ( 
.A(n_1189),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_1166),
.Y(n_1283)
);

A2O1A1Ixp33_ASAP7_75t_SL g1284 ( 
.A1(n_1210),
.A2(n_1195),
.B(n_1205),
.C(n_1180),
.Y(n_1284)
);

OA22x2_ASAP7_75t_L g1285 ( 
.A1(n_1206),
.A2(n_1186),
.B1(n_1241),
.B2(n_1242),
.Y(n_1285)
);

OAI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1195),
.A2(n_1235),
.B1(n_1206),
.B2(n_1185),
.Y(n_1286)
);

INVxp67_ASAP7_75t_L g1287 ( 
.A(n_1221),
.Y(n_1287)
);

INVxp67_ASAP7_75t_L g1288 ( 
.A(n_1227),
.Y(n_1288)
);

OA21x2_ASAP7_75t_L g1289 ( 
.A1(n_1177),
.A2(n_1151),
.B(n_1255),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1230),
.Y(n_1290)
);

OA21x2_ASAP7_75t_L g1291 ( 
.A1(n_1177),
.A2(n_1151),
.B(n_1253),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1145),
.B(n_1171),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1171),
.B(n_1258),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1193),
.Y(n_1294)
);

A2O1A1Ixp33_ASAP7_75t_L g1295 ( 
.A1(n_1249),
.A2(n_1192),
.B(n_1198),
.C(n_1197),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1188),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1191),
.B(n_1172),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1191),
.B(n_1172),
.Y(n_1298)
);

AOI221x1_ASAP7_75t_SL g1299 ( 
.A1(n_1209),
.A2(n_1204),
.B1(n_1200),
.B2(n_1257),
.C(n_1250),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_1248),
.Y(n_1300)
);

AOI221x1_ASAP7_75t_SL g1301 ( 
.A1(n_1157),
.A2(n_1257),
.B1(n_1179),
.B2(n_1234),
.C(n_1250),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_1160),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1191),
.B(n_1155),
.Y(n_1303)
);

NOR2x1_ASAP7_75t_SL g1304 ( 
.A(n_1241),
.B(n_1199),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1206),
.A2(n_1241),
.B1(n_1243),
.B2(n_1170),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1229),
.B(n_1202),
.Y(n_1306)
);

BUFx3_ASAP7_75t_L g1307 ( 
.A(n_1243),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_SL g1308 ( 
.A1(n_1149),
.A2(n_1159),
.B(n_1199),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1229),
.B(n_1202),
.Y(n_1309)
);

INVx1_ASAP7_75t_SL g1310 ( 
.A(n_1214),
.Y(n_1310)
);

OR2x2_ASAP7_75t_L g1311 ( 
.A(n_1155),
.B(n_1236),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1163),
.B(n_1236),
.Y(n_1312)
);

O2A1O1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1196),
.A2(n_1144),
.B(n_1233),
.C(n_1170),
.Y(n_1313)
);

AOI21x1_ASAP7_75t_SL g1314 ( 
.A1(n_1211),
.A2(n_1203),
.B(n_1163),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_SL g1315 ( 
.A1(n_1149),
.A2(n_1159),
.B(n_1199),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1208),
.B(n_1211),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1207),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1215),
.A2(n_1228),
.B1(n_1165),
.B2(n_1159),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1208),
.B(n_1212),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1215),
.B(n_1159),
.Y(n_1320)
);

CKINVDCx20_ASAP7_75t_R g1321 ( 
.A(n_1228),
.Y(n_1321)
);

OA21x2_ASAP7_75t_L g1322 ( 
.A1(n_1224),
.A2(n_1225),
.B(n_1246),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1212),
.B(n_1244),
.Y(n_1323)
);

NAND2x1_ASAP7_75t_L g1324 ( 
.A(n_1154),
.B(n_1244),
.Y(n_1324)
);

INVx1_ASAP7_75t_SL g1325 ( 
.A(n_1216),
.Y(n_1325)
);

OR2x2_ASAP7_75t_L g1326 ( 
.A(n_1213),
.B(n_1153),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1201),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1153),
.A2(n_1154),
.B1(n_1152),
.B2(n_1218),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1154),
.Y(n_1329)
);

OA21x2_ASAP7_75t_L g1330 ( 
.A1(n_1237),
.A2(n_1205),
.B(n_1023),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1237),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1162),
.B(n_1251),
.Y(n_1332)
);

O2A1O1Ixp33_ASAP7_75t_L g1333 ( 
.A1(n_1238),
.A2(n_1247),
.B(n_1219),
.C(n_1231),
.Y(n_1333)
);

INVx5_ASAP7_75t_L g1334 ( 
.A(n_1228),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1162),
.B(n_1251),
.Y(n_1335)
);

INVx1_ASAP7_75t_SL g1336 ( 
.A(n_1190),
.Y(n_1336)
);

INVxp33_ASAP7_75t_L g1337 ( 
.A(n_1282),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1292),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1292),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1266),
.B(n_1272),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1326),
.B(n_1329),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1327),
.Y(n_1342)
);

OR2x2_ASAP7_75t_L g1343 ( 
.A(n_1297),
.B(n_1298),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1297),
.B(n_1298),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1323),
.B(n_1303),
.Y(n_1345)
);

OR2x6_ASAP7_75t_L g1346 ( 
.A(n_1275),
.B(n_1308),
.Y(n_1346)
);

OAI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1267),
.A2(n_1333),
.B(n_1273),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1323),
.B(n_1303),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1319),
.B(n_1266),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1311),
.B(n_1324),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1272),
.B(n_1290),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1267),
.B(n_1333),
.Y(n_1352)
);

AND2x4_ASAP7_75t_L g1353 ( 
.A(n_1304),
.B(n_1317),
.Y(n_1353)
);

HB1xp67_ASAP7_75t_L g1354 ( 
.A(n_1316),
.Y(n_1354)
);

OR2x2_ASAP7_75t_L g1355 ( 
.A(n_1293),
.B(n_1316),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1269),
.B(n_1286),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_SL g1357 ( 
.A1(n_1273),
.A2(n_1295),
.B(n_1262),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1325),
.Y(n_1358)
);

OR2x2_ASAP7_75t_L g1359 ( 
.A(n_1312),
.B(n_1328),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1331),
.Y(n_1360)
);

AO21x2_ASAP7_75t_L g1361 ( 
.A1(n_1276),
.A2(n_1284),
.B(n_1312),
.Y(n_1361)
);

OR2x2_ASAP7_75t_L g1362 ( 
.A(n_1276),
.B(n_1330),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1259),
.B(n_1289),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1301),
.Y(n_1364)
);

OR2x2_ASAP7_75t_L g1365 ( 
.A(n_1291),
.B(n_1296),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1285),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1285),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1322),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1260),
.B(n_1270),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1322),
.Y(n_1370)
);

BUFx6f_ASAP7_75t_L g1371 ( 
.A(n_1334),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1313),
.Y(n_1372)
);

OR2x6_ASAP7_75t_L g1373 ( 
.A(n_1315),
.B(n_1313),
.Y(n_1373)
);

AO21x2_ASAP7_75t_L g1374 ( 
.A1(n_1305),
.A2(n_1314),
.B(n_1318),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1332),
.B(n_1335),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1279),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1360),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1363),
.B(n_1271),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1349),
.B(n_1280),
.Y(n_1379)
);

BUFx3_ASAP7_75t_L g1380 ( 
.A(n_1353),
.Y(n_1380)
);

INVx5_ASAP7_75t_L g1381 ( 
.A(n_1346),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1358),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1353),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1365),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1363),
.B(n_1274),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1363),
.B(n_1283),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1343),
.B(n_1336),
.Y(n_1387)
);

OAI221xp5_ASAP7_75t_L g1388 ( 
.A1(n_1356),
.A2(n_1278),
.B1(n_1299),
.B2(n_1287),
.C(n_1288),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1360),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1343),
.B(n_1310),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1343),
.B(n_1294),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1365),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1353),
.Y(n_1393)
);

NOR2xp67_ASAP7_75t_L g1394 ( 
.A(n_1365),
.B(n_1344),
.Y(n_1394)
);

AND2x4_ASAP7_75t_L g1395 ( 
.A(n_1353),
.B(n_1261),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1342),
.Y(n_1396)
);

INVxp67_ASAP7_75t_SL g1397 ( 
.A(n_1358),
.Y(n_1397)
);

INVxp67_ASAP7_75t_L g1398 ( 
.A(n_1351),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1349),
.B(n_1265),
.Y(n_1399)
);

AND2x2_ASAP7_75t_SL g1400 ( 
.A(n_1369),
.B(n_1281),
.Y(n_1400)
);

NOR2x1_ASAP7_75t_L g1401 ( 
.A(n_1373),
.B(n_1321),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1338),
.B(n_1320),
.Y(n_1402)
);

INVxp67_ASAP7_75t_L g1403 ( 
.A(n_1351),
.Y(n_1403)
);

INVx4_ASAP7_75t_L g1404 ( 
.A(n_1371),
.Y(n_1404)
);

AOI221xp5_ASAP7_75t_L g1405 ( 
.A1(n_1352),
.A2(n_1300),
.B1(n_1309),
.B2(n_1306),
.C(n_1264),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1368),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1386),
.B(n_1344),
.Y(n_1407)
);

AOI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1388),
.A2(n_1356),
.B1(n_1352),
.B2(n_1347),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1406),
.Y(n_1409)
);

NOR2x1p5_ASAP7_75t_L g1410 ( 
.A(n_1404),
.B(n_1376),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1386),
.B(n_1344),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1377),
.Y(n_1412)
);

AND2x4_ASAP7_75t_L g1413 ( 
.A(n_1380),
.B(n_1353),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1382),
.Y(n_1414)
);

INVx3_ASAP7_75t_L g1415 ( 
.A(n_1380),
.Y(n_1415)
);

INVxp67_ASAP7_75t_SL g1416 ( 
.A(n_1394),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1383),
.B(n_1345),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1383),
.B(n_1345),
.Y(n_1418)
);

OAI33xp33_ASAP7_75t_L g1419 ( 
.A1(n_1398),
.A2(n_1376),
.A3(n_1355),
.B1(n_1340),
.B2(n_1372),
.B3(n_1339),
.Y(n_1419)
);

AOI221xp5_ASAP7_75t_L g1420 ( 
.A1(n_1403),
.A2(n_1357),
.B1(n_1347),
.B2(n_1337),
.C(n_1364),
.Y(n_1420)
);

OAI221xp5_ASAP7_75t_SL g1421 ( 
.A1(n_1405),
.A2(n_1346),
.B1(n_1373),
.B2(n_1340),
.C(n_1367),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1377),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1384),
.B(n_1348),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1384),
.B(n_1348),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1390),
.B(n_1337),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1400),
.A2(n_1366),
.B1(n_1346),
.B2(n_1374),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1392),
.B(n_1348),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1397),
.Y(n_1428)
);

OAI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1400),
.A2(n_1364),
.B1(n_1373),
.B2(n_1346),
.Y(n_1429)
);

NAND2xp33_ASAP7_75t_R g1430 ( 
.A(n_1390),
.B(n_1263),
.Y(n_1430)
);

AOI221xp5_ASAP7_75t_L g1431 ( 
.A1(n_1402),
.A2(n_1372),
.B1(n_1375),
.B2(n_1354),
.C(n_1361),
.Y(n_1431)
);

AND2x4_ASAP7_75t_L g1432 ( 
.A(n_1380),
.B(n_1341),
.Y(n_1432)
);

INVx1_ASAP7_75t_SL g1433 ( 
.A(n_1378),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1385),
.B(n_1359),
.Y(n_1434)
);

INVx1_ASAP7_75t_SL g1435 ( 
.A(n_1378),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1393),
.B(n_1350),
.Y(n_1436)
);

INVx2_ASAP7_75t_SL g1437 ( 
.A(n_1393),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1401),
.A2(n_1346),
.B1(n_1374),
.B2(n_1373),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1436),
.B(n_1379),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1412),
.Y(n_1440)
);

OR2x6_ASAP7_75t_L g1441 ( 
.A(n_1429),
.B(n_1346),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1425),
.B(n_1379),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1413),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1414),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1436),
.B(n_1395),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1412),
.Y(n_1446)
);

OAI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1408),
.A2(n_1420),
.B(n_1431),
.Y(n_1447)
);

BUFx2_ASAP7_75t_L g1448 ( 
.A(n_1410),
.Y(n_1448)
);

INVx1_ASAP7_75t_SL g1449 ( 
.A(n_1428),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1422),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1409),
.Y(n_1451)
);

AOI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1409),
.A2(n_1370),
.B(n_1396),
.Y(n_1452)
);

INVx1_ASAP7_75t_SL g1453 ( 
.A(n_1433),
.Y(n_1453)
);

BUFx8_ASAP7_75t_L g1454 ( 
.A(n_1437),
.Y(n_1454)
);

INVx1_ASAP7_75t_SL g1455 ( 
.A(n_1435),
.Y(n_1455)
);

INVxp67_ASAP7_75t_SL g1456 ( 
.A(n_1410),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1413),
.B(n_1381),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_1408),
.B(n_1277),
.Y(n_1458)
);

OA21x2_ASAP7_75t_L g1459 ( 
.A1(n_1438),
.A2(n_1362),
.B(n_1389),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1434),
.B(n_1385),
.Y(n_1460)
);

INVx4_ASAP7_75t_SL g1461 ( 
.A(n_1437),
.Y(n_1461)
);

NOR2x1p5_ASAP7_75t_L g1462 ( 
.A(n_1416),
.B(n_1404),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1435),
.B(n_1391),
.Y(n_1463)
);

INVx3_ASAP7_75t_L g1464 ( 
.A(n_1415),
.Y(n_1464)
);

NAND4xp25_ASAP7_75t_L g1465 ( 
.A(n_1447),
.B(n_1426),
.C(n_1421),
.D(n_1430),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1460),
.B(n_1434),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1460),
.B(n_1407),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1448),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1449),
.B(n_1423),
.Y(n_1469)
);

INVx4_ASAP7_75t_L g1470 ( 
.A(n_1448),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_L g1471 ( 
.A(n_1458),
.B(n_1307),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1449),
.B(n_1423),
.Y(n_1472)
);

INVxp67_ASAP7_75t_L g1473 ( 
.A(n_1444),
.Y(n_1473)
);

NOR2xp33_ASAP7_75t_L g1474 ( 
.A(n_1442),
.B(n_1447),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1462),
.B(n_1415),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1462),
.B(n_1432),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1456),
.B(n_1445),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1452),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1440),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1453),
.B(n_1407),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1453),
.B(n_1424),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1455),
.Y(n_1482)
);

INVx3_ASAP7_75t_L g1483 ( 
.A(n_1452),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1461),
.B(n_1381),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1440),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1446),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1441),
.A2(n_1429),
.B1(n_1401),
.B2(n_1381),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1455),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1457),
.B(n_1417),
.Y(n_1489)
);

NOR2xp67_ASAP7_75t_L g1490 ( 
.A(n_1443),
.B(n_1381),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1451),
.Y(n_1491)
);

INVx2_ASAP7_75t_SL g1492 ( 
.A(n_1454),
.Y(n_1492)
);

INVx2_ASAP7_75t_SL g1493 ( 
.A(n_1454),
.Y(n_1493)
);

INVx1_ASAP7_75t_SL g1494 ( 
.A(n_1461),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1446),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1463),
.B(n_1411),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1450),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1457),
.B(n_1461),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1457),
.B(n_1417),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1465),
.B(n_1419),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1482),
.B(n_1391),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1468),
.Y(n_1502)
);

NAND2x1p5_ASAP7_75t_L g1503 ( 
.A(n_1470),
.B(n_1381),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1465),
.B(n_1268),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1474),
.A2(n_1459),
.B1(n_1361),
.B2(n_1441),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1488),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1473),
.B(n_1439),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1473),
.B(n_1439),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1468),
.Y(n_1509)
);

AND2x4_ASAP7_75t_SL g1510 ( 
.A(n_1488),
.B(n_1457),
.Y(n_1510)
);

AND2x4_ASAP7_75t_L g1511 ( 
.A(n_1498),
.B(n_1461),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1479),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1477),
.B(n_1375),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1477),
.B(n_1375),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1498),
.B(n_1461),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1479),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1469),
.B(n_1427),
.Y(n_1517)
);

INVxp67_ASAP7_75t_L g1518 ( 
.A(n_1492),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1485),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1485),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1469),
.B(n_1472),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1472),
.B(n_1427),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1480),
.B(n_1387),
.Y(n_1523)
);

NAND3xp33_ASAP7_75t_L g1524 ( 
.A(n_1470),
.B(n_1459),
.C(n_1441),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1470),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1492),
.B(n_1443),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1480),
.B(n_1399),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1496),
.B(n_1399),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1496),
.B(n_1402),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1470),
.B(n_1418),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1481),
.B(n_1418),
.Y(n_1531)
);

AND2x2_ASAP7_75t_SL g1532 ( 
.A(n_1487),
.B(n_1281),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1486),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1486),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1515),
.B(n_1476),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1515),
.B(n_1476),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1500),
.B(n_1489),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1512),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1502),
.Y(n_1539)
);

CKINVDCx16_ASAP7_75t_R g1540 ( 
.A(n_1504),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1516),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1511),
.B(n_1475),
.Y(n_1542)
);

AOI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1500),
.A2(n_1493),
.B1(n_1492),
.B2(n_1441),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1506),
.B(n_1467),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1511),
.B(n_1475),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1502),
.B(n_1467),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1509),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1509),
.B(n_1466),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1519),
.Y(n_1549)
);

AO21x2_ASAP7_75t_L g1550 ( 
.A1(n_1524),
.A2(n_1490),
.B(n_1478),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1511),
.B(n_1494),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1520),
.Y(n_1552)
);

AOI22xp5_ASAP7_75t_SL g1553 ( 
.A1(n_1504),
.A2(n_1493),
.B1(n_1471),
.B2(n_1494),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1510),
.B(n_1526),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1518),
.B(n_1489),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1518),
.B(n_1499),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1533),
.Y(n_1557)
);

INVxp67_ASAP7_75t_L g1558 ( 
.A(n_1525),
.Y(n_1558)
);

OR2x6_ASAP7_75t_L g1559 ( 
.A(n_1525),
.B(n_1493),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1546),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1546),
.Y(n_1561)
);

OAI221xp5_ASAP7_75t_L g1562 ( 
.A1(n_1543),
.A2(n_1505),
.B1(n_1521),
.B2(n_1503),
.C(n_1507),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1548),
.B(n_1537),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1548),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1539),
.Y(n_1565)
);

CKINVDCx20_ASAP7_75t_R g1566 ( 
.A(n_1540),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1539),
.Y(n_1567)
);

AND2x4_ASAP7_75t_SL g1568 ( 
.A(n_1554),
.B(n_1484),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1542),
.B(n_1510),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1547),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1542),
.B(n_1508),
.Y(n_1571)
);

INVx2_ASAP7_75t_SL g1572 ( 
.A(n_1554),
.Y(n_1572)
);

NOR2x1_ASAP7_75t_L g1573 ( 
.A(n_1559),
.B(n_1534),
.Y(n_1573)
);

INVxp33_ASAP7_75t_L g1574 ( 
.A(n_1553),
.Y(n_1574)
);

INVx1_ASAP7_75t_SL g1575 ( 
.A(n_1551),
.Y(n_1575)
);

O2A1O1Ixp33_ASAP7_75t_L g1576 ( 
.A1(n_1547),
.A2(n_1505),
.B(n_1503),
.C(n_1530),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1544),
.B(n_1513),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1544),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1575),
.B(n_1558),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1560),
.Y(n_1580)
);

XNOR2x1_ASAP7_75t_L g1581 ( 
.A(n_1563),
.B(n_1302),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1561),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1566),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1571),
.B(n_1551),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1564),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1578),
.Y(n_1586)
);

AOI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1574),
.A2(n_1535),
.B1(n_1536),
.B2(n_1532),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1571),
.B(n_1555),
.Y(n_1588)
);

O2A1O1Ixp33_ASAP7_75t_L g1589 ( 
.A1(n_1579),
.A2(n_1562),
.B(n_1576),
.C(n_1573),
.Y(n_1589)
);

NAND3xp33_ASAP7_75t_L g1590 ( 
.A(n_1587),
.B(n_1573),
.C(n_1572),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1579),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_SL g1592 ( 
.A(n_1583),
.B(n_1569),
.Y(n_1592)
);

OAI221xp5_ASAP7_75t_SL g1593 ( 
.A1(n_1584),
.A2(n_1577),
.B1(n_1559),
.B2(n_1545),
.C(n_1556),
.Y(n_1593)
);

NOR3xp33_ASAP7_75t_SL g1594 ( 
.A(n_1588),
.B(n_1567),
.C(n_1565),
.Y(n_1594)
);

NOR2x1_ASAP7_75t_L g1595 ( 
.A(n_1581),
.B(n_1559),
.Y(n_1595)
);

AOI211xp5_ASAP7_75t_L g1596 ( 
.A1(n_1580),
.A2(n_1569),
.B(n_1570),
.C(n_1545),
.Y(n_1596)
);

NOR3x1_ASAP7_75t_L g1597 ( 
.A(n_1582),
.B(n_1549),
.C(n_1538),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1591),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1596),
.B(n_1586),
.Y(n_1599)
);

NAND3xp33_ASAP7_75t_L g1600 ( 
.A(n_1594),
.B(n_1585),
.C(n_1559),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1592),
.B(n_1568),
.Y(n_1601)
);

OAI21xp33_ASAP7_75t_L g1602 ( 
.A1(n_1595),
.A2(n_1536),
.B(n_1535),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1598),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1602),
.B(n_1590),
.Y(n_1604)
);

INVxp33_ASAP7_75t_SL g1605 ( 
.A(n_1601),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1599),
.Y(n_1606)
);

NOR3xp33_ASAP7_75t_L g1607 ( 
.A(n_1600),
.B(n_1593),
.C(n_1589),
.Y(n_1607)
);

NAND3xp33_ASAP7_75t_L g1608 ( 
.A(n_1600),
.B(n_1557),
.C(n_1552),
.Y(n_1608)
);

AOI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1607),
.A2(n_1541),
.B1(n_1557),
.B2(n_1552),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_R g1610 ( 
.A(n_1606),
.B(n_1597),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1608),
.Y(n_1611)
);

NOR2xp67_ASAP7_75t_SL g1612 ( 
.A(n_1603),
.B(n_1541),
.Y(n_1612)
);

A2O1A1Ixp33_ASAP7_75t_L g1613 ( 
.A1(n_1604),
.A2(n_1490),
.B(n_1483),
.C(n_1532),
.Y(n_1613)
);

NOR3xp33_ASAP7_75t_SL g1614 ( 
.A(n_1611),
.B(n_1605),
.C(n_1550),
.Y(n_1614)
);

OAI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1609),
.A2(n_1613),
.B1(n_1501),
.B2(n_1523),
.Y(n_1615)
);

AOI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1610),
.A2(n_1550),
.B(n_1514),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1615),
.B(n_1550),
.Y(n_1617)
);

AOI322xp5_ASAP7_75t_L g1618 ( 
.A1(n_1617),
.A2(n_1614),
.A3(n_1612),
.B1(n_1616),
.B2(n_1483),
.C1(n_1478),
.C2(n_1484),
.Y(n_1618)
);

INVx1_ASAP7_75t_SL g1619 ( 
.A(n_1618),
.Y(n_1619)
);

OR5x1_ASAP7_75t_L g1620 ( 
.A(n_1618),
.B(n_1483),
.C(n_1491),
.D(n_1478),
.E(n_1464),
.Y(n_1620)
);

AO22x2_ASAP7_75t_L g1621 ( 
.A1(n_1619),
.A2(n_1491),
.B1(n_1483),
.B2(n_1495),
.Y(n_1621)
);

HB1xp67_ASAP7_75t_L g1622 ( 
.A(n_1620),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1621),
.Y(n_1623)
);

CKINVDCx20_ASAP7_75t_R g1624 ( 
.A(n_1622),
.Y(n_1624)
);

OAI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1624),
.A2(n_1491),
.B1(n_1517),
.B2(n_1522),
.Y(n_1625)
);

AOI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1625),
.A2(n_1623),
.B(n_1531),
.Y(n_1626)
);

NOR2xp33_ASAP7_75t_L g1627 ( 
.A(n_1626),
.B(n_1527),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1627),
.A2(n_1484),
.B1(n_1495),
.B2(n_1497),
.Y(n_1628)
);

AOI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1628),
.A2(n_1484),
.B1(n_1497),
.B2(n_1499),
.Y(n_1629)
);

AOI211xp5_ASAP7_75t_L g1630 ( 
.A1(n_1629),
.A2(n_1481),
.B(n_1529),
.C(n_1528),
.Y(n_1630)
);


endmodule