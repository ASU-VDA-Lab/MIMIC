module fake_ariane_2182_n_938 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_938);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_938;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_516;
wire n_307;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_678;
wire n_651;
wire n_936;
wire n_347;
wire n_423;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_285;
wire n_473;
wire n_801;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_557;
wire n_405;
wire n_858;
wire n_242;
wire n_645;
wire n_320;
wire n_331;
wire n_559;
wire n_309;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_600;
wire n_721;
wire n_481;
wire n_840;
wire n_398;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_839;
wire n_821;
wire n_928;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_914;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_301;
wire n_248;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_365;
wire n_238;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_889;
wire n_935;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_543;
wire n_362;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_747;
wire n_741;
wire n_772;
wire n_847;
wire n_371;
wire n_845;
wire n_888;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_922;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_896;
wire n_409;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_915;
wire n_252;
wire n_215;
wire n_664;
wire n_629;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_213;
wire n_895;
wire n_304;
wire n_862;
wire n_659;
wire n_583;
wire n_509;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_751;
wire n_615;
wire n_521;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_580;
wire n_358;
wire n_892;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_882;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_749;
wire n_289;
wire n_542;
wire n_548;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_129),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_91),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_165),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_209),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_85),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_10),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_83),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_81),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_25),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_88),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_166),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_38),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_153),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_175),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_194),
.Y(n_227)
);

CKINVDCx11_ASAP7_75t_R g228 ( 
.A(n_45),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_109),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_108),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_159),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_103),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_189),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_140),
.B(n_124),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_162),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_183),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_96),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_199),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_19),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_146),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_147),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_196),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_134),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_127),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_47),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_200),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_137),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_133),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_128),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_24),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_23),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_130),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_173),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_75),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_160),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_6),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_117),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_107),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_41),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_54),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_142),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_211),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_131),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_138),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_17),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_212),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_139),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_118),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_52),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_5),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_80),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_56),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_148),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_66),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_105),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_74),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_113),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_110),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_161),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_41),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_14),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_73),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_6),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_178),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_57),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_145),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_207),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_51),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_51),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_198),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_193),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_101),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_40),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_115),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_19),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_120),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_77),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_99),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_125),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_180),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_121),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_3),
.Y(n_303)
);

BUFx10_ASAP7_75t_L g304 ( 
.A(n_84),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_182),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_43),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_111),
.Y(n_307)
);

BUFx5_ASAP7_75t_L g308 ( 
.A(n_42),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_82),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_136),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_36),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_27),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_116),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_197),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_46),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_53),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_201),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_58),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_44),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_11),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_144),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_55),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_36),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_152),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_190),
.Y(n_325)
);

BUFx10_ASAP7_75t_L g326 ( 
.A(n_155),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_149),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_86),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_163),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_168),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_94),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_35),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_186),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_21),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_89),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_192),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_177),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_104),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_122),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_64),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_169),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_126),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_97),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_202),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_98),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_179),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_16),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_187),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_38),
.Y(n_349)
);

CKINVDCx14_ASAP7_75t_R g350 ( 
.A(n_14),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_154),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_68),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_119),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_10),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_93),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_48),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_50),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_176),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_45),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_114),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_20),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_112),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_20),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_156),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_1),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_79),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_12),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_70),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_228),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_260),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_260),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_350),
.B(n_0),
.Y(n_372)
);

BUFx6f_ASAP7_75t_SL g373 ( 
.A(n_304),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_350),
.Y(n_374)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_296),
.B(n_0),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_252),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_334),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_308),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_308),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_320),
.Y(n_380)
);

INVxp67_ASAP7_75t_SL g381 ( 
.A(n_281),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_216),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_220),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_261),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_276),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_308),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_308),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_267),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_308),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_308),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_333),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_263),
.B(n_2),
.Y(n_392)
);

INVxp67_ASAP7_75t_SL g393 ( 
.A(n_281),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_251),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_221),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_311),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_224),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_218),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_227),
.B(n_231),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_354),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_332),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_349),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_236),
.B(n_4),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_240),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_246),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_353),
.B(n_4),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_361),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_363),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_257),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_267),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_304),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_266),
.Y(n_412)
);

NOR2xp67_ASAP7_75t_L g413 ( 
.A(n_271),
.B(n_282),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_284),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_289),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_326),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_326),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_326),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_275),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_237),
.B(n_7),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_329),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_290),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_294),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_253),
.Y(n_424)
);

NOR2xp67_ASAP7_75t_L g425 ( 
.A(n_303),
.B(n_7),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_256),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_264),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g428 ( 
.A(n_306),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_274),
.B(n_8),
.Y(n_429)
);

INVxp67_ASAP7_75t_SL g430 ( 
.A(n_275),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_277),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_278),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_319),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_295),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_312),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_285),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_315),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_323),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_293),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_298),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_299),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_300),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_347),
.Y(n_443)
);

INVxp33_ASAP7_75t_SL g444 ( 
.A(n_356),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_301),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_302),
.B(n_8),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_305),
.Y(n_447)
);

NOR2xp67_ASAP7_75t_L g448 ( 
.A(n_357),
.B(n_9),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_359),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_310),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_316),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_327),
.Y(n_452)
);

INVxp67_ASAP7_75t_SL g453 ( 
.A(n_295),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_313),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_328),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_330),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_335),
.B(n_337),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_339),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_365),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_341),
.B(n_9),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_367),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_213),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_343),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_214),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_346),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_215),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_217),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_222),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_223),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_348),
.Y(n_470)
);

INVxp67_ASAP7_75t_SL g471 ( 
.A(n_314),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_225),
.Y(n_472)
);

INVxp67_ASAP7_75t_SL g473 ( 
.A(n_314),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_352),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_226),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_229),
.Y(n_476)
);

CKINVDCx16_ASAP7_75t_R g477 ( 
.A(n_232),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_230),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_232),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_233),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_479),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_477),
.B(n_355),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_479),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_479),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_479),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_378),
.Y(n_486)
);

OA21x2_ASAP7_75t_L g487 ( 
.A1(n_379),
.A2(n_364),
.B(n_368),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_416),
.B(n_219),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_386),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_387),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_412),
.A2(n_239),
.B1(n_283),
.B2(n_248),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_389),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_412),
.A2(n_317),
.B1(n_331),
.B2(n_318),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_390),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_434),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_434),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_394),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_388),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_372),
.B(n_336),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_433),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_388),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_419),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_396),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_424),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_426),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_427),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_401),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_419),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_428),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_410),
.B(n_344),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_372),
.B(n_344),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_402),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_376),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_407),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_408),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_381),
.B(n_360),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_431),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_432),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_380),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_430),
.B(n_238),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_393),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_436),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_371),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_370),
.B(n_232),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_377),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_439),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_440),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_441),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_442),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_445),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_447),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_450),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_451),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_453),
.B(n_232),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_452),
.Y(n_535)
);

OA21x2_ASAP7_75t_L g536 ( 
.A1(n_403),
.A2(n_234),
.B(n_242),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_398),
.A2(n_244),
.B1(n_245),
.B2(n_243),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_417),
.B(n_418),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_455),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_462),
.B(n_247),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_456),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_458),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_375),
.A2(n_250),
.B1(n_254),
.B2(n_249),
.Y(n_543)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_438),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_465),
.Y(n_545)
);

INVx4_ASAP7_75t_L g546 ( 
.A(n_464),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_471),
.B(n_235),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_470),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_454),
.B(n_255),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_473),
.B(n_463),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_400),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_474),
.B(n_235),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_400),
.Y(n_553)
);

INVx1_ASAP7_75t_SL g554 ( 
.A(n_461),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_399),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_411),
.B(n_258),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_466),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_469),
.B(n_259),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_406),
.Y(n_559)
);

OA21x2_ASAP7_75t_L g560 ( 
.A1(n_420),
.A2(n_268),
.B(n_262),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_406),
.B(n_366),
.Y(n_561)
);

OA21x2_ASAP7_75t_L g562 ( 
.A1(n_457),
.A2(n_270),
.B(n_269),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_489),
.Y(n_563)
);

NAND3xp33_ASAP7_75t_L g564 ( 
.A(n_555),
.B(n_475),
.C(n_472),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_500),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_509),
.B(n_395),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_495),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_498),
.Y(n_568)
);

INVx4_ASAP7_75t_SL g569 ( 
.A(n_557),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_544),
.B(n_550),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_498),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_523),
.Y(n_572)
);

BUFx4f_ASAP7_75t_L g573 ( 
.A(n_498),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_496),
.Y(n_574)
);

OR2x2_ASAP7_75t_L g575 ( 
.A(n_554),
.B(n_382),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_540),
.B(n_444),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_557),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_494),
.Y(n_578)
);

AO21x2_ASAP7_75t_L g579 ( 
.A1(n_499),
.A2(n_448),
.B(n_425),
.Y(n_579)
);

BUFx4f_ASAP7_75t_L g580 ( 
.A(n_501),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_496),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_525),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_558),
.B(n_476),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_534),
.B(n_478),
.Y(n_584)
);

OAI22xp33_ASAP7_75t_L g585 ( 
.A1(n_491),
.A2(n_405),
.B1(n_414),
.B2(n_409),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_508),
.B(n_413),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_497),
.Y(n_587)
);

INVx4_ASAP7_75t_SL g588 ( 
.A(n_537),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_503),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_501),
.Y(n_590)
);

AND2x6_ASAP7_75t_L g591 ( 
.A(n_524),
.B(n_235),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_520),
.B(n_423),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_552),
.B(n_467),
.Y(n_593)
);

OR2x2_ASAP7_75t_SL g594 ( 
.A(n_513),
.B(n_397),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_501),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g596 ( 
.A(n_501),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_546),
.B(n_435),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_502),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_502),
.Y(n_599)
);

INVx5_ASAP7_75t_L g600 ( 
.A(n_502),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_502),
.Y(n_601)
);

BUFx4f_ASAP7_75t_L g602 ( 
.A(n_562),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_492),
.Y(n_603)
);

OR2x6_ASAP7_75t_L g604 ( 
.A(n_513),
.B(n_404),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_549),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_486),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_559),
.B(n_482),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_490),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_499),
.A2(n_392),
.B1(n_446),
.B2(n_429),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_492),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_534),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_L g612 ( 
.A(n_561),
.B(n_449),
.Y(n_612)
);

INVx1_ASAP7_75t_SL g613 ( 
.A(n_519),
.Y(n_613)
);

AND2x6_ASAP7_75t_L g614 ( 
.A(n_524),
.B(n_235),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_538),
.B(n_459),
.Y(n_615)
);

INVxp67_ASAP7_75t_SL g616 ( 
.A(n_547),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_553),
.Y(n_617)
);

INVx4_ASAP7_75t_L g618 ( 
.A(n_547),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_511),
.A2(n_392),
.B1(n_446),
.B2(n_429),
.Y(n_619)
);

OR2x2_ASAP7_75t_L g620 ( 
.A(n_519),
.B(n_383),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_507),
.Y(n_621)
);

AND2x4_ASAP7_75t_L g622 ( 
.A(n_552),
.B(n_468),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_512),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_516),
.B(n_415),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_551),
.Y(n_625)
);

NOR2xp67_ASAP7_75t_L g626 ( 
.A(n_565),
.B(n_384),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_607),
.B(n_516),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_563),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_625),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_611),
.Y(n_630)
);

OAI221xp5_ASAP7_75t_L g631 ( 
.A1(n_609),
.A2(n_511),
.B1(n_460),
.B2(n_493),
.C(n_488),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_567),
.Y(n_632)
);

AO22x2_ASAP7_75t_L g633 ( 
.A1(n_588),
.A2(n_622),
.B1(n_593),
.B2(n_575),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_577),
.Y(n_634)
);

NAND2x1p5_ASAP7_75t_L g635 ( 
.A(n_618),
.B(n_514),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_616),
.Y(n_636)
);

AO22x2_ASAP7_75t_L g637 ( 
.A1(n_588),
.A2(n_622),
.B1(n_593),
.B2(n_620),
.Y(n_637)
);

NAND2x1p5_ASAP7_75t_L g638 ( 
.A(n_618),
.B(n_515),
.Y(n_638)
);

OAI221xp5_ASAP7_75t_L g639 ( 
.A1(n_619),
.A2(n_543),
.B1(n_527),
.B2(n_529),
.C(n_528),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_615),
.B(n_385),
.Y(n_640)
);

OAI221xp5_ASAP7_75t_L g641 ( 
.A1(n_624),
.A2(n_530),
.B1(n_532),
.B2(n_531),
.C(n_526),
.Y(n_641)
);

AO22x2_ASAP7_75t_L g642 ( 
.A1(n_613),
.A2(n_391),
.B1(n_561),
.B2(n_374),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_569),
.B(n_521),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_570),
.B(n_437),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_604),
.B(n_510),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_606),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_608),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_569),
.B(n_522),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_563),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_566),
.B(n_443),
.Y(n_650)
);

AO22x2_ASAP7_75t_L g651 ( 
.A1(n_605),
.A2(n_535),
.B1(n_545),
.B2(n_533),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_604),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_574),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_581),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_578),
.Y(n_655)
);

AO22x2_ASAP7_75t_L g656 ( 
.A1(n_587),
.A2(n_505),
.B1(n_506),
.B2(n_504),
.Y(n_656)
);

OAI221xp5_ASAP7_75t_L g657 ( 
.A1(n_584),
.A2(n_539),
.B1(n_517),
.B2(n_518),
.C(n_504),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_L g658 ( 
.A1(n_576),
.A2(n_556),
.B1(n_480),
.B2(n_422),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_572),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_583),
.B(n_421),
.Y(n_660)
);

A2O1A1Ixp33_ASAP7_75t_L g661 ( 
.A1(n_592),
.A2(n_517),
.B(n_541),
.C(n_518),
.Y(n_661)
);

INVxp67_ASAP7_75t_L g662 ( 
.A(n_586),
.Y(n_662)
);

OAI221xp5_ASAP7_75t_L g663 ( 
.A1(n_589),
.A2(n_542),
.B1(n_548),
.B2(n_536),
.C(n_562),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_582),
.Y(n_664)
);

AOI22x1_ASAP7_75t_L g665 ( 
.A1(n_617),
.A2(n_484),
.B1(n_483),
.B2(n_485),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_621),
.Y(n_666)
);

OAI221xp5_ASAP7_75t_L g667 ( 
.A1(n_623),
.A2(n_536),
.B1(n_562),
.B2(n_560),
.C(n_487),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_SL g668 ( 
.A1(n_594),
.A2(n_369),
.B1(n_536),
.B2(n_560),
.Y(n_668)
);

AO22x2_ASAP7_75t_L g669 ( 
.A1(n_564),
.A2(n_373),
.B1(n_560),
.B2(n_487),
.Y(n_669)
);

CKINVDCx20_ASAP7_75t_R g670 ( 
.A(n_597),
.Y(n_670)
);

NAND2x1_ASAP7_75t_L g671 ( 
.A(n_610),
.B(n_487),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_579),
.B(n_272),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_579),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_603),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_568),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_571),
.Y(n_676)
);

AOI22xp5_ASAP7_75t_L g677 ( 
.A1(n_612),
.A2(n_279),
.B1(n_280),
.B2(n_273),
.Y(n_677)
);

INVxp67_ASAP7_75t_L g678 ( 
.A(n_585),
.Y(n_678)
);

AO22x2_ASAP7_75t_L g679 ( 
.A1(n_602),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_571),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_610),
.Y(n_681)
);

NAND2xp33_ASAP7_75t_SL g682 ( 
.A(n_627),
.B(n_590),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_640),
.B(n_573),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_636),
.B(n_591),
.Y(n_684)
);

NAND2xp33_ASAP7_75t_SL g685 ( 
.A(n_650),
.B(n_590),
.Y(n_685)
);

AND2x4_ASAP7_75t_L g686 ( 
.A(n_643),
.B(n_595),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_644),
.B(n_598),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_634),
.B(n_573),
.Y(n_688)
);

NAND2xp33_ASAP7_75t_SL g689 ( 
.A(n_658),
.B(n_590),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_648),
.B(n_580),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_648),
.B(n_580),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_SL g692 ( 
.A(n_626),
.B(n_602),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_646),
.B(n_591),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_660),
.B(n_599),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_647),
.B(n_614),
.Y(n_695)
);

NAND2xp33_ASAP7_75t_SL g696 ( 
.A(n_670),
.B(n_601),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_678),
.B(n_601),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_662),
.B(n_600),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_635),
.B(n_600),
.Y(n_699)
);

NAND2xp33_ASAP7_75t_SL g700 ( 
.A(n_659),
.B(n_287),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_638),
.B(n_596),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_668),
.B(n_291),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_652),
.B(n_292),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_630),
.B(n_297),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_664),
.B(n_485),
.Y(n_705)
);

AND2x4_ASAP7_75t_L g706 ( 
.A(n_666),
.B(n_485),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_677),
.B(n_307),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_645),
.B(n_309),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_641),
.B(n_13),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_681),
.B(n_628),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_672),
.B(n_321),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_631),
.B(n_322),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_655),
.B(n_324),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_649),
.B(n_325),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_651),
.B(n_338),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_661),
.B(n_340),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_675),
.B(n_342),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_676),
.B(n_345),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_633),
.B(n_15),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_680),
.B(n_351),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_673),
.B(n_358),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_629),
.B(n_362),
.Y(n_722)
);

OAI21x1_ASAP7_75t_L g723 ( 
.A1(n_716),
.A2(n_671),
.B(n_665),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_683),
.A2(n_657),
.B(n_639),
.Y(n_724)
);

OA21x2_ASAP7_75t_L g725 ( 
.A1(n_697),
.A2(n_663),
.B(n_667),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_687),
.B(n_651),
.Y(n_726)
);

OAI21x1_ASAP7_75t_L g727 ( 
.A1(n_710),
.A2(n_665),
.B(n_674),
.Y(n_727)
);

OAI21x1_ASAP7_75t_L g728 ( 
.A1(n_693),
.A2(n_695),
.B(n_705),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_709),
.B(n_637),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_709),
.B(n_656),
.Y(n_730)
);

INVx5_ASAP7_75t_L g731 ( 
.A(n_686),
.Y(n_731)
);

OAI21x1_ASAP7_75t_L g732 ( 
.A1(n_684),
.A2(n_699),
.B(n_721),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_719),
.B(n_642),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_706),
.Y(n_734)
);

OAI21x1_ASAP7_75t_L g735 ( 
.A1(n_701),
.A2(n_653),
.B(n_632),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_706),
.Y(n_736)
);

OAI21x1_ASAP7_75t_L g737 ( 
.A1(n_711),
.A2(n_654),
.B(n_484),
.Y(n_737)
);

OAI21x1_ASAP7_75t_L g738 ( 
.A1(n_694),
.A2(n_669),
.B(n_679),
.Y(n_738)
);

AOI21xp5_ASAP7_75t_L g739 ( 
.A1(n_712),
.A2(n_265),
.B(n_241),
.Y(n_739)
);

OAI21x1_ASAP7_75t_L g740 ( 
.A1(n_690),
.A2(n_691),
.B(n_702),
.Y(n_740)
);

AOI21xp5_ASAP7_75t_L g741 ( 
.A1(n_682),
.A2(n_265),
.B(n_241),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_689),
.B(n_481),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_714),
.A2(n_265),
.B(n_241),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_L g744 ( 
.A1(n_707),
.A2(n_288),
.B1(n_286),
.B2(n_241),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_698),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_688),
.Y(n_746)
);

INVx1_ASAP7_75t_SL g747 ( 
.A(n_696),
.Y(n_747)
);

OAI21x1_ASAP7_75t_L g748 ( 
.A1(n_717),
.A2(n_60),
.B(n_59),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_703),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_685),
.B(n_715),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_708),
.B(n_18),
.Y(n_751)
);

OA21x2_ASAP7_75t_L g752 ( 
.A1(n_713),
.A2(n_62),
.B(n_61),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_700),
.B(n_22),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_704),
.B(n_26),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_718),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_720),
.Y(n_756)
);

NAND2x1_ASAP7_75t_L g757 ( 
.A(n_692),
.B(n_63),
.Y(n_757)
);

OAI21x1_ASAP7_75t_L g758 ( 
.A1(n_723),
.A2(n_722),
.B(n_65),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_729),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_759)
);

OAI21x1_ASAP7_75t_L g760 ( 
.A1(n_728),
.A2(n_69),
.B(n_67),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_730),
.B(n_724),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_731),
.Y(n_762)
);

OAI21x1_ASAP7_75t_L g763 ( 
.A1(n_737),
.A2(n_72),
.B(n_71),
.Y(n_763)
);

HB1xp67_ASAP7_75t_L g764 ( 
.A(n_734),
.Y(n_764)
);

BUFx3_ASAP7_75t_L g765 ( 
.A(n_731),
.Y(n_765)
);

OAI21x1_ASAP7_75t_L g766 ( 
.A1(n_727),
.A2(n_78),
.B(n_76),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_747),
.B(n_30),
.Y(n_767)
);

BUFx2_ASAP7_75t_L g768 ( 
.A(n_731),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_735),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_SL g770 ( 
.A1(n_733),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_746),
.Y(n_771)
);

INVx4_ASAP7_75t_SL g772 ( 
.A(n_754),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_747),
.B(n_31),
.Y(n_773)
);

HB1xp67_ASAP7_75t_L g774 ( 
.A(n_736),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_726),
.B(n_32),
.Y(n_775)
);

CKINVDCx20_ASAP7_75t_R g776 ( 
.A(n_749),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_745),
.Y(n_777)
);

A2O1A1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_751),
.A2(n_34),
.B(n_37),
.C(n_39),
.Y(n_778)
);

OA21x2_ASAP7_75t_L g779 ( 
.A1(n_739),
.A2(n_738),
.B(n_732),
.Y(n_779)
);

OR2x6_ASAP7_75t_L g780 ( 
.A(n_740),
.B(n_37),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_755),
.B(n_87),
.Y(n_781)
);

OA21x2_ASAP7_75t_L g782 ( 
.A1(n_750),
.A2(n_143),
.B(n_210),
.Y(n_782)
);

AND2x6_ASAP7_75t_L g783 ( 
.A(n_756),
.B(n_90),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_753),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_757),
.Y(n_785)
);

OAI21x1_ASAP7_75t_L g786 ( 
.A1(n_741),
.A2(n_150),
.B(n_208),
.Y(n_786)
);

AO21x2_ASAP7_75t_L g787 ( 
.A1(n_742),
.A2(n_151),
.B(n_206),
.Y(n_787)
);

OAI21x1_ASAP7_75t_L g788 ( 
.A1(n_748),
.A2(n_141),
.B(n_205),
.Y(n_788)
);

AOI21xp33_ASAP7_75t_L g789 ( 
.A1(n_744),
.A2(n_48),
.B(n_49),
.Y(n_789)
);

INVx1_ASAP7_75t_SL g790 ( 
.A(n_725),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_752),
.Y(n_791)
);

NAND2x1p5_ASAP7_75t_L g792 ( 
.A(n_752),
.B(n_92),
.Y(n_792)
);

OAI21x1_ASAP7_75t_L g793 ( 
.A1(n_743),
.A2(n_158),
.B(n_204),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_779),
.Y(n_794)
);

BUFx2_ASAP7_75t_L g795 ( 
.A(n_780),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_774),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_761),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_779),
.Y(n_798)
);

OAI21x1_ASAP7_75t_L g799 ( 
.A1(n_758),
.A2(n_157),
.B(n_203),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_761),
.Y(n_800)
);

CKINVDCx20_ASAP7_75t_R g801 ( 
.A(n_776),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_771),
.B(n_777),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_775),
.B(n_95),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_790),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_769),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_780),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_791),
.Y(n_807)
);

HB1xp67_ASAP7_75t_L g808 ( 
.A(n_764),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_784),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_767),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_765),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_782),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_773),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_772),
.Y(n_814)
);

OR2x6_ASAP7_75t_L g815 ( 
.A(n_781),
.B(n_100),
.Y(n_815)
);

OAI21x1_ASAP7_75t_L g816 ( 
.A1(n_760),
.A2(n_102),
.B(n_106),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_772),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_787),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_792),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_763),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_766),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_788),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_783),
.Y(n_823)
);

CKINVDCx20_ASAP7_75t_R g824 ( 
.A(n_801),
.Y(n_824)
);

HB1xp67_ASAP7_75t_L g825 ( 
.A(n_796),
.Y(n_825)
);

BUFx4f_ASAP7_75t_L g826 ( 
.A(n_815),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_802),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_810),
.B(n_770),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_813),
.B(n_809),
.Y(n_829)
);

AND2x4_ASAP7_75t_L g830 ( 
.A(n_796),
.B(n_768),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_795),
.B(n_762),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_R g832 ( 
.A(n_811),
.B(n_785),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_808),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_797),
.B(n_759),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_800),
.B(n_778),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_817),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_795),
.B(n_786),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_806),
.B(n_793),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_806),
.B(n_814),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_803),
.B(n_789),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_807),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_807),
.Y(n_842)
);

AND2x4_ASAP7_75t_L g843 ( 
.A(n_823),
.B(n_123),
.Y(n_843)
);

NAND2xp33_ASAP7_75t_R g844 ( 
.A(n_804),
.B(n_132),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_833),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_829),
.B(n_805),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_826),
.Y(n_847)
);

INVxp67_ASAP7_75t_SL g848 ( 
.A(n_825),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_827),
.B(n_794),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_840),
.B(n_798),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_830),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_839),
.B(n_819),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_838),
.B(n_818),
.Y(n_853)
);

INVx3_ASAP7_75t_L g854 ( 
.A(n_838),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_837),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_837),
.B(n_812),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_841),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_830),
.B(n_812),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_835),
.B(n_822),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_842),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_834),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_831),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_831),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_828),
.B(n_821),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_836),
.B(n_820),
.Y(n_865)
);

INVx2_ASAP7_75t_SL g866 ( 
.A(n_832),
.Y(n_866)
);

AND2x4_ASAP7_75t_L g867 ( 
.A(n_843),
.B(n_820),
.Y(n_867)
);

AND2x4_ASAP7_75t_SL g868 ( 
.A(n_847),
.B(n_824),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_848),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_850),
.B(n_816),
.Y(n_870)
);

INVx3_ASAP7_75t_SL g871 ( 
.A(n_866),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_854),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_857),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_854),
.B(n_799),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_849),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_857),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_854),
.B(n_844),
.Y(n_877)
);

BUFx2_ASAP7_75t_L g878 ( 
.A(n_855),
.Y(n_878)
);

BUFx2_ASAP7_75t_L g879 ( 
.A(n_855),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_878),
.B(n_855),
.Y(n_880)
);

AND3x2_ASAP7_75t_L g881 ( 
.A(n_877),
.B(n_861),
.C(n_863),
.Y(n_881)
);

INVxp67_ASAP7_75t_SL g882 ( 
.A(n_869),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_878),
.B(n_845),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_872),
.B(n_853),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_879),
.B(n_845),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_873),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_879),
.B(n_851),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_872),
.B(n_851),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_872),
.B(n_870),
.Y(n_889)
);

AND2x4_ASAP7_75t_L g890 ( 
.A(n_874),
.B(n_853),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_873),
.Y(n_891)
);

OR2x2_ASAP7_75t_L g892 ( 
.A(n_875),
.B(n_864),
.Y(n_892)
);

OR2x2_ASAP7_75t_L g893 ( 
.A(n_875),
.B(n_859),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_882),
.B(n_871),
.Y(n_894)
);

NAND2xp33_ASAP7_75t_SL g895 ( 
.A(n_883),
.B(n_877),
.Y(n_895)
);

INVx2_ASAP7_75t_SL g896 ( 
.A(n_885),
.Y(n_896)
);

INVxp67_ASAP7_75t_L g897 ( 
.A(n_887),
.Y(n_897)
);

INVxp67_ASAP7_75t_L g898 ( 
.A(n_887),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_SL g899 ( 
.A(n_881),
.B(n_868),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_884),
.Y(n_900)
);

NAND2xp33_ASAP7_75t_SL g901 ( 
.A(n_880),
.B(n_865),
.Y(n_901)
);

INVxp67_ASAP7_75t_L g902 ( 
.A(n_894),
.Y(n_902)
);

OR2x2_ASAP7_75t_L g903 ( 
.A(n_897),
.B(n_893),
.Y(n_903)
);

BUFx2_ASAP7_75t_L g904 ( 
.A(n_895),
.Y(n_904)
);

AND3x1_ASAP7_75t_L g905 ( 
.A(n_899),
.B(n_880),
.C(n_888),
.Y(n_905)
);

OR2x2_ASAP7_75t_L g906 ( 
.A(n_898),
.B(n_892),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_896),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_901),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_903),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_902),
.B(n_900),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_905),
.B(n_908),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_906),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_909),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_912),
.B(n_902),
.Y(n_914)
);

NOR2x1_ASAP7_75t_L g915 ( 
.A(n_911),
.B(n_904),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_910),
.B(n_907),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_914),
.Y(n_917)
);

INVx1_ASAP7_75t_SL g918 ( 
.A(n_915),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_913),
.Y(n_919)
);

INVx2_ASAP7_75t_SL g920 ( 
.A(n_916),
.Y(n_920)
);

NOR3xp33_ASAP7_75t_L g921 ( 
.A(n_918),
.B(n_917),
.C(n_920),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_919),
.B(n_889),
.Y(n_922)
);

OAI21xp5_ASAP7_75t_SL g923 ( 
.A1(n_921),
.A2(n_890),
.B(n_874),
.Y(n_923)
);

NOR3xp33_ASAP7_75t_SL g924 ( 
.A(n_922),
.B(n_862),
.C(n_846),
.Y(n_924)
);

NOR2x1_ASAP7_75t_L g925 ( 
.A(n_923),
.B(n_847),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_924),
.B(n_891),
.Y(n_926)
);

OAI21x1_ASAP7_75t_L g927 ( 
.A1(n_925),
.A2(n_886),
.B(n_858),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_R g928 ( 
.A(n_926),
.B(n_135),
.Y(n_928)
);

OAI22x1_ASAP7_75t_L g929 ( 
.A1(n_928),
.A2(n_867),
.B1(n_852),
.B2(n_858),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_927),
.B(n_856),
.Y(n_930)
);

NOR4xp25_ASAP7_75t_L g931 ( 
.A(n_930),
.B(n_929),
.C(n_876),
.D(n_860),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_931),
.B(n_164),
.Y(n_932)
);

AOI31xp33_ASAP7_75t_L g933 ( 
.A1(n_932),
.A2(n_167),
.A3(n_170),
.B(n_171),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_933),
.B(n_172),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_934),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_935),
.Y(n_936)
);

AOI22xp5_ASAP7_75t_L g937 ( 
.A1(n_936),
.A2(n_174),
.B1(n_184),
.B2(n_185),
.Y(n_937)
);

AOI211xp5_ASAP7_75t_L g938 ( 
.A1(n_937),
.A2(n_188),
.B(n_191),
.C(n_195),
.Y(n_938)
);


endmodule