module real_jpeg_12159_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_176;
wire n_221;
wire n_166;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_213;
wire n_167;
wire n_179;
wire n_216;
wire n_133;
wire n_202;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_89;

BUFx10_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_3),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_3),
.A2(n_46),
.B1(n_60),
.B2(n_64),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_3),
.A2(n_29),
.B1(n_35),
.B2(n_46),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_5),
.A2(n_66),
.B1(n_67),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_5),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_5),
.A2(n_60),
.B1(n_64),
.B2(n_70),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_5),
.A2(n_43),
.B1(n_44),
.B2(n_70),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_5),
.A2(n_29),
.B1(n_35),
.B2(n_70),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_6),
.A2(n_66),
.B1(n_67),
.B2(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_6),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_6),
.A2(n_60),
.B1(n_64),
.B2(n_139),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_6),
.A2(n_43),
.B1(n_44),
.B2(n_139),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_6),
.A2(n_29),
.B1(n_35),
.B2(n_139),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_7),
.A2(n_29),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_7),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_9),
.A2(n_29),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_9),
.A2(n_36),
.B1(n_43),
.B2(n_44),
.Y(n_87)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_11),
.A2(n_60),
.B1(n_64),
.B2(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_11),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_11),
.A2(n_43),
.B1(n_44),
.B2(n_81),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_11),
.A2(n_66),
.B1(n_67),
.B2(n_81),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_11),
.A2(n_29),
.B1(n_35),
.B2(n_81),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_12),
.A2(n_66),
.B1(n_67),
.B2(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_12),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_12),
.A2(n_60),
.B1(n_64),
.B2(n_104),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_12),
.A2(n_43),
.B1(n_44),
.B2(n_104),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_12),
.A2(n_29),
.B1(n_35),
.B2(n_104),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_13),
.A2(n_66),
.B1(n_67),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_13),
.A2(n_60),
.B1(n_64),
.B2(n_72),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_13),
.A2(n_43),
.B1(n_44),
.B2(n_72),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_13),
.A2(n_29),
.B1(n_35),
.B2(n_72),
.Y(n_194)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

AOI21xp33_ASAP7_75t_L g134 ( 
.A1(n_15),
.A2(n_66),
.B(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_15),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_15),
.B(n_161),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_L g205 ( 
.A1(n_15),
.A2(n_43),
.B1(n_44),
.B2(n_137),
.Y(n_205)
);

O2A1O1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_15),
.A2(n_43),
.B(n_49),
.C(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_15),
.B(n_111),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_15),
.B(n_32),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_15),
.B(n_54),
.Y(n_232)
);

A2O1A1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_15),
.A2(n_64),
.B(n_75),
.C(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_16),
.A2(n_43),
.B1(n_44),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_16),
.A2(n_29),
.B1(n_35),
.B2(n_53),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_16),
.A2(n_53),
.B1(n_60),
.B2(n_64),
.Y(n_110)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_127),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_126),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_105),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_22),
.B(n_105),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_83),
.C(n_89),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_23),
.B(n_83),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_55),
.B2(n_56),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_24),
.B(n_57),
.C(n_73),
.Y(n_125)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_39),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_26),
.A2(n_27),
.B1(n_39),
.B2(n_40),
.Y(n_260)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_28),
.A2(n_32),
.B(n_37),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_28),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_28),
.A2(n_32),
.B1(n_95),
.B2(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_28),
.A2(n_32),
.B1(n_151),
.B2(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_28),
.A2(n_32),
.B1(n_163),
.B2(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_28),
.A2(n_32),
.B1(n_194),
.B2(n_215),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_28),
.A2(n_32),
.B1(n_137),
.B2(n_227),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_28),
.A2(n_32),
.B1(n_220),
.B2(n_227),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_29),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_29),
.A2(n_35),
.B1(n_49),
.B2(n_50),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_29),
.B(n_229),
.Y(n_228)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_31),
.A2(n_34),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_31),
.A2(n_93),
.B1(n_219),
.B2(n_221),
.Y(n_218)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI21xp33_ASAP7_75t_L g208 ( 
.A1(n_35),
.A2(n_50),
.B(n_137),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_47),
.B1(n_52),
.B2(n_54),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_42),
.A2(n_51),
.B1(n_97),
.B2(n_99),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_44),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_43),
.A2(n_44),
.B1(n_77),
.B2(n_78),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_43),
.B(n_78),
.Y(n_192)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI32xp33_ASAP7_75t_L g190 ( 
.A1(n_44),
.A2(n_64),
.A3(n_77),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_47),
.A2(n_52),
.B1(n_54),
.B2(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_47),
.A2(n_54),
.B1(n_87),
.B2(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_47),
.A2(n_54),
.B1(n_98),
.B2(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_47),
.A2(n_54),
.B1(n_145),
.B2(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_47),
.A2(n_54),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_47),
.A2(n_54),
.B1(n_206),
.B2(n_213),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_51),
.A2(n_99),
.B1(n_186),
.B2(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_73),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_69),
.B2(n_71),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_58),
.A2(n_59),
.B1(n_69),
.B2(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_58),
.A2(n_59),
.B1(n_71),
.B2(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_58),
.A2(n_59),
.B1(n_134),
.B2(n_138),
.Y(n_133)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_58),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_65),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_59),
.Y(n_161)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_60),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_60),
.A2(n_64),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

OAI32xp33_ASAP7_75t_L g153 ( 
.A1(n_60),
.A2(n_63),
.A3(n_66),
.B1(n_136),
.B2(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_60),
.B(n_137),
.Y(n_191)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_62),
.A2(n_63),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_62),
.B(n_64),
.Y(n_154)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_67),
.B(n_137),
.Y(n_136)
);

BUFx16f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_79),
.B1(n_80),
.B2(n_82),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_74),
.A2(n_79),
.B1(n_80),
.B2(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_74),
.A2(n_79),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_75),
.A2(n_111),
.B1(n_157),
.B2(n_159),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_75),
.A2(n_111),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_79),
.A2(n_158),
.B(n_241),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_86),
.B2(n_88),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_88),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_84),
.A2(n_85),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_89),
.B(n_271),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_100),
.C(n_102),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_90),
.A2(n_91),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_96),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_92),
.B(n_96),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_100),
.B(n_102),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_101),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_103),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_125),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_115),
.B1(n_116),
.B2(n_124),
.Y(n_106)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_112),
.B(n_114),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_112),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_123),
.Y(n_116)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_268),
.B(n_272),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_178),
.B(n_256),
.C(n_267),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_164),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_130),
.B(n_164),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_148),
.C(n_155),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_131),
.A2(n_132),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_140),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_141),
.C(n_147),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_140)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_141),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_142),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_144),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_148),
.B(n_155),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_152),
.B2(n_153),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_149),
.B(n_153),
.Y(n_177)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_160),
.C(n_162),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_156),
.B(n_183),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_162),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_161),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_166),
.B(n_167),
.C(n_168),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_177),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_170),
.B(n_173),
.C(n_177),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_255),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_198),
.B(n_254),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_195),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_181),
.B(n_195),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.C(n_187),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_182),
.B(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_184),
.A2(n_187),
.B1(n_188),
.B2(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_184),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_193),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_189),
.A2(n_190),
.B1(n_193),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_191),
.Y(n_242)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_193),
.Y(n_246)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_196),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_248),
.B(n_253),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_236),
.B(n_247),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_216),
.B(n_235),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_209),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_202),
.B(n_209),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_207),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_203),
.A2(n_204),
.B1(n_207),
.B2(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_214),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_212),
.C(n_214),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_213),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_215),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_224),
.B(n_234),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_218),
.B(n_222),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_230),
.B(n_233),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_231),
.B(n_232),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_237),
.B(n_238),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_245),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_243),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_243),
.C(n_245),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_249),
.B(n_250),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_258),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_266),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_264),
.B2(n_265),
.Y(n_259)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_260),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_265),
.C(n_266),
.Y(n_269)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_261),
.Y(n_265)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_270),
.Y(n_272)
);


endmodule