module fake_ibex_1551_n_15 (n_4, n_2, n_0, n_3, n_1, n_15);

input n_4;
input n_2;
input n_0;
input n_3;
input n_1;

output n_15;

wire n_13;
wire n_7;
wire n_5;
wire n_11;
wire n_8;
wire n_6;
wire n_14;
wire n_10;
wire n_9;
wire n_12;

INVx2_ASAP7_75t_L g5 ( 
.A(n_1),
.Y(n_5)
);

INVx1_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

INVx4_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_1),
.B(n_0),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_5),
.B(n_0),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_9),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

OAI21xp33_ASAP7_75t_L g12 ( 
.A1(n_11),
.A2(n_8),
.B(n_6),
.Y(n_12)
);

AND3x4_ASAP7_75t_L g13 ( 
.A(n_12),
.B(n_7),
.C(n_4),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_14),
.Y(n_15)
);


endmodule