module real_aes_1483_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_449;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g519 ( .A(n_0), .B(n_216), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_1), .B(n_109), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_2), .Y(n_123) );
INVx1_ASAP7_75t_L g150 ( .A(n_3), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_4), .B(n_522), .Y(n_541) );
NAND2xp33_ASAP7_75t_SL g512 ( .A(n_5), .B(n_171), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_6), .B(n_184), .Y(n_207) );
INVx1_ASAP7_75t_L g504 ( .A(n_7), .Y(n_504) );
INVx1_ASAP7_75t_L g241 ( .A(n_8), .Y(n_241) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_9), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_10), .Y(n_258) );
AND2x2_ASAP7_75t_L g539 ( .A(n_11), .B(n_140), .Y(n_539) );
INVx2_ASAP7_75t_L g141 ( .A(n_12), .Y(n_141) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_13), .Y(n_110) );
INVx1_ASAP7_75t_L g217 ( .A(n_14), .Y(n_217) );
AOI221x1_ASAP7_75t_L g507 ( .A1(n_15), .A2(n_173), .B1(n_508), .B2(n_510), .C(n_511), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g100 ( .A1(n_16), .A2(n_101), .B1(n_111), .B2(n_807), .Y(n_100) );
NAND2xp5_ASAP7_75t_SL g575 ( .A(n_17), .B(n_522), .Y(n_575) );
INVx1_ASAP7_75t_L g106 ( .A(n_18), .Y(n_106) );
INVx1_ASAP7_75t_L g214 ( .A(n_19), .Y(n_214) );
INVx1_ASAP7_75t_SL g162 ( .A(n_20), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_21), .B(n_165), .Y(n_187) );
AOI33xp33_ASAP7_75t_L g232 ( .A1(n_22), .A2(n_50), .A3(n_147), .B1(n_158), .B2(n_233), .B3(n_234), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_23), .A2(n_510), .B(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_24), .B(n_216), .Y(n_544) );
AOI221xp5_ASAP7_75t_SL g584 ( .A1(n_25), .A2(n_40), .B1(n_510), .B2(n_522), .C(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g251 ( .A(n_26), .Y(n_251) );
OR2x2_ASAP7_75t_L g142 ( .A(n_27), .B(n_88), .Y(n_142) );
OA21x2_ASAP7_75t_L g175 ( .A1(n_27), .A2(n_88), .B(n_141), .Y(n_175) );
INVxp67_ASAP7_75t_L g506 ( .A(n_28), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_29), .B(n_219), .Y(n_579) );
AND2x2_ASAP7_75t_L g533 ( .A(n_30), .B(n_139), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_31), .B(n_145), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_32), .A2(n_510), .B(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_33), .B(n_219), .Y(n_586) );
AND2x2_ASAP7_75t_L g152 ( .A(n_34), .B(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g157 ( .A(n_34), .Y(n_157) );
AND2x2_ASAP7_75t_L g171 ( .A(n_34), .B(n_150), .Y(n_171) );
NOR3xp33_ASAP7_75t_L g107 ( .A(n_35), .B(n_108), .C(n_110), .Y(n_107) );
OR2x6_ASAP7_75t_L g121 ( .A(n_35), .B(n_122), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g253 ( .A(n_36), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_37), .B(n_145), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_38), .A2(n_174), .B1(n_180), .B2(n_184), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_39), .B(n_189), .Y(n_188) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_41), .A2(n_80), .B1(n_155), .B2(n_510), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_42), .B(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_43), .B(n_216), .Y(n_531) );
AOI22xp33_ASAP7_75t_SL g787 ( .A1(n_44), .A2(n_786), .B1(n_788), .B2(n_790), .Y(n_787) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_45), .B(n_191), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_46), .B(n_165), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_47), .Y(n_183) );
AND2x2_ASAP7_75t_L g523 ( .A(n_48), .B(n_139), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_49), .B(n_139), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_51), .B(n_165), .Y(n_282) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_52), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g804 ( .A1(n_52), .A2(n_62), .B1(n_430), .B2(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g148 ( .A(n_53), .Y(n_148) );
INVx1_ASAP7_75t_L g167 ( .A(n_53), .Y(n_167) );
AND2x2_ASAP7_75t_L g283 ( .A(n_54), .B(n_139), .Y(n_283) );
AOI221xp5_ASAP7_75t_L g239 ( .A1(n_55), .A2(n_73), .B1(n_145), .B2(n_155), .C(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_56), .B(n_145), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_57), .B(n_522), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_58), .B(n_174), .Y(n_260) );
AOI21xp5_ASAP7_75t_SL g196 ( .A1(n_59), .A2(n_155), .B(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g560 ( .A(n_60), .B(n_139), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_61), .B(n_219), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_62), .Y(n_805) );
INVx1_ASAP7_75t_L g210 ( .A(n_63), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_64), .B(n_216), .Y(n_558) );
AND2x2_ASAP7_75t_SL g580 ( .A(n_65), .B(n_140), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_66), .A2(n_510), .B(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g281 ( .A(n_67), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_68), .B(n_219), .Y(n_545) );
AND2x2_ASAP7_75t_SL g552 ( .A(n_69), .B(n_191), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_70), .A2(n_155), .B(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g153 ( .A(n_71), .Y(n_153) );
INVx1_ASAP7_75t_L g169 ( .A(n_71), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_72), .B(n_145), .Y(n_235) );
AND2x2_ASAP7_75t_L g172 ( .A(n_74), .B(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g211 ( .A(n_75), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_76), .A2(n_155), .B(n_161), .Y(n_154) );
A2O1A1Ixp33_ASAP7_75t_L g185 ( .A1(n_77), .A2(n_155), .B(n_186), .C(n_190), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g550 ( .A1(n_78), .A2(n_83), .B1(n_145), .B2(n_522), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_79), .B(n_522), .Y(n_559) );
INVx1_ASAP7_75t_L g105 ( .A(n_81), .Y(n_105) );
AND2x2_ASAP7_75t_SL g194 ( .A(n_82), .B(n_173), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g229 ( .A1(n_84), .A2(n_155), .B1(n_230), .B2(n_231), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_85), .B(n_216), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_86), .B(n_216), .Y(n_587) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_87), .A2(n_510), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g198 ( .A(n_89), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_90), .B(n_219), .Y(n_557) );
AND2x2_ASAP7_75t_L g236 ( .A(n_91), .B(n_173), .Y(n_236) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_92), .A2(n_249), .B(n_250), .C(n_252), .Y(n_248) );
INVxp67_ASAP7_75t_L g509 ( .A(n_93), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_94), .B(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_95), .B(n_219), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_96), .A2(n_510), .B(n_577), .Y(n_576) );
BUFx2_ASAP7_75t_L g115 ( .A(n_97), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_98), .B(n_165), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_99), .Y(n_786) );
INVx1_ASAP7_75t_SL g807 ( .A(n_101), .Y(n_807) );
INVx2_ASAP7_75t_R g101 ( .A(n_102), .Y(n_101) );
INVx3_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
AND2x2_ASAP7_75t_SL g103 ( .A(n_104), .B(n_107), .Y(n_103) );
NOR2xp33_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_105), .B(n_106), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_110), .B(n_120), .Y(n_119) );
AND2x6_ASAP7_75t_SL g494 ( .A(n_110), .B(n_121), .Y(n_494) );
OR2x6_ASAP7_75t_SL g785 ( .A(n_110), .B(n_120), .Y(n_785) );
OR2x2_ASAP7_75t_L g793 ( .A(n_110), .B(n_121), .Y(n_793) );
OA21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_124), .B(n_794), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_116), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_114), .B(n_795), .Y(n_794) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_115), .Y(n_114) );
INVxp67_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g795 ( .A1(n_117), .A2(n_796), .B(n_806), .Y(n_795) );
NOR2xp33_ASAP7_75t_SL g117 ( .A(n_118), .B(n_123), .Y(n_117) );
BUFx2_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g806 ( .A(n_119), .Y(n_806) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_121), .Y(n_120) );
OAI21xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_786), .B(n_787), .Y(n_124) );
INVxp67_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OAI22x1_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_493), .B1(n_495), .B2(n_783), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
OAI22xp5_ASAP7_75t_L g788 ( .A1(n_128), .A2(n_493), .B1(n_496), .B2(n_789), .Y(n_788) );
AND3x1_ASAP7_75t_L g128 ( .A(n_129), .B(n_487), .C(n_490), .Y(n_128) );
NAND5xp2_ASAP7_75t_L g129 ( .A(n_130), .B(n_387), .C(n_417), .D(n_431), .E(n_457), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OAI21xp33_ASAP7_75t_L g487 ( .A1(n_131), .A2(n_430), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g801 ( .A(n_131), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_336), .Y(n_131) );
NOR3xp33_ASAP7_75t_SL g132 ( .A(n_133), .B(n_284), .C(n_318), .Y(n_132) );
A2O1A1Ixp33_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_201), .B(n_223), .C(n_262), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_176), .Y(n_134) );
BUFx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_136), .B(n_274), .Y(n_339) );
AND2x2_ASAP7_75t_L g426 ( .A(n_136), .B(n_204), .Y(n_426) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
OR2x2_ASAP7_75t_L g222 ( .A(n_137), .B(n_193), .Y(n_222) );
INVx1_ASAP7_75t_L g264 ( .A(n_137), .Y(n_264) );
INVx2_ASAP7_75t_L g269 ( .A(n_137), .Y(n_269) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_137), .Y(n_297) );
INVx1_ASAP7_75t_L g311 ( .A(n_137), .Y(n_311) );
AND2x2_ASAP7_75t_L g315 ( .A(n_137), .B(n_206), .Y(n_315) );
AND2x2_ASAP7_75t_L g396 ( .A(n_137), .B(n_205), .Y(n_396) );
AO21x2_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_143), .B(n_172), .Y(n_137) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_138), .A2(n_527), .B(n_533), .Y(n_526) );
AO21x2_ASAP7_75t_L g553 ( .A1(n_138), .A2(n_554), .B(n_560), .Y(n_553) );
AO21x2_ASAP7_75t_L g591 ( .A1(n_138), .A2(n_527), .B(n_533), .Y(n_591) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_139), .Y(n_138) );
OA21x2_ASAP7_75t_L g583 ( .A1(n_139), .A2(n_584), .B(n_588), .Y(n_583) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_SL g140 ( .A(n_141), .B(n_142), .Y(n_140) );
AND2x4_ASAP7_75t_L g184 ( .A(n_141), .B(n_142), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_154), .Y(n_143) );
INVx1_ASAP7_75t_L g261 ( .A(n_145), .Y(n_261) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_145), .A2(n_155), .B1(n_503), .B2(n_505), .Y(n_502) );
AND2x4_ASAP7_75t_L g145 ( .A(n_146), .B(n_151), .Y(n_145) );
INVx1_ASAP7_75t_L g181 ( .A(n_146), .Y(n_181) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_149), .Y(n_146) );
OR2x6_ASAP7_75t_L g163 ( .A(n_147), .B(n_159), .Y(n_163) );
INVxp33_ASAP7_75t_L g233 ( .A(n_147), .Y(n_233) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x2_ASAP7_75t_L g160 ( .A(n_148), .B(n_150), .Y(n_160) );
AND2x4_ASAP7_75t_L g219 ( .A(n_148), .B(n_168), .Y(n_219) );
HB1xp67_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g182 ( .A(n_151), .Y(n_182) );
BUFx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AND2x6_ASAP7_75t_L g510 ( .A(n_152), .B(n_160), .Y(n_510) );
INVx2_ASAP7_75t_L g159 ( .A(n_153), .Y(n_159) );
AND2x6_ASAP7_75t_L g216 ( .A(n_153), .B(n_166), .Y(n_216) );
INVxp67_ASAP7_75t_L g259 ( .A(n_155), .Y(n_259) );
AND2x4_ASAP7_75t_L g155 ( .A(n_156), .B(n_160), .Y(n_155) );
NOR2x1p5_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
INVx1_ASAP7_75t_L g234 ( .A(n_158), .Y(n_234) );
INVx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
O2A1O1Ixp33_ASAP7_75t_SL g161 ( .A1(n_162), .A2(n_163), .B(n_164), .C(n_170), .Y(n_161) );
INVx2_ASAP7_75t_L g189 ( .A(n_163), .Y(n_189) );
O2A1O1Ixp33_ASAP7_75t_L g197 ( .A1(n_163), .A2(n_170), .B(n_198), .C(n_199), .Y(n_197) );
OAI22xp5_ASAP7_75t_L g209 ( .A1(n_163), .A2(n_210), .B1(n_211), .B2(n_212), .Y(n_209) );
O2A1O1Ixp33_ASAP7_75t_SL g240 ( .A1(n_163), .A2(n_170), .B(n_241), .C(n_242), .Y(n_240) );
INVxp67_ASAP7_75t_L g249 ( .A(n_163), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_L g280 ( .A1(n_163), .A2(n_170), .B(n_281), .C(n_282), .Y(n_280) );
INVx1_ASAP7_75t_L g212 ( .A(n_165), .Y(n_212) );
AND2x4_ASAP7_75t_L g522 ( .A(n_165), .B(n_171), .Y(n_522) );
AND2x4_ASAP7_75t_L g165 ( .A(n_166), .B(n_168), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_170), .A2(n_187), .B(n_188), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_170), .B(n_184), .Y(n_220) );
INVx1_ASAP7_75t_L g230 ( .A(n_170), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_170), .A2(n_519), .B(n_520), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_170), .A2(n_530), .B(n_531), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_170), .A2(n_544), .B(n_545), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_170), .A2(n_557), .B(n_558), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_170), .A2(n_578), .B(n_579), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_170), .A2(n_586), .B(n_587), .Y(n_585) );
INVx5_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_171), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g247 ( .A1(n_173), .A2(n_248), .B1(n_253), .B2(n_254), .Y(n_247) );
INVx3_ASAP7_75t_L g254 ( .A(n_173), .Y(n_254) );
INVx4_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_174), .B(n_257), .Y(n_256) );
AOI21x1_ASAP7_75t_L g515 ( .A1(n_174), .A2(n_516), .B(n_523), .Y(n_515) );
INVx3_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
BUFx4f_ASAP7_75t_L g191 ( .A(n_175), .Y(n_191) );
AND2x4_ASAP7_75t_SL g176 ( .A(n_177), .B(n_192), .Y(n_176) );
HB1xp67_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g221 ( .A(n_178), .Y(n_221) );
AND2x2_ASAP7_75t_L g265 ( .A(n_178), .B(n_206), .Y(n_265) );
AND2x2_ASAP7_75t_L g286 ( .A(n_178), .B(n_193), .Y(n_286) );
INVx1_ASAP7_75t_L g309 ( .A(n_178), .Y(n_309) );
AND2x4_ASAP7_75t_L g376 ( .A(n_178), .B(n_205), .Y(n_376) );
AND2x2_ASAP7_75t_L g178 ( .A(n_179), .B(n_185), .Y(n_178) );
NOR3xp33_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .C(n_183), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_184), .A2(n_196), .B(n_200), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_184), .B(n_504), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_184), .B(n_506), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_184), .B(n_509), .Y(n_508) );
NOR3xp33_ASAP7_75t_L g511 ( .A(n_184), .B(n_212), .C(n_512), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_184), .A2(n_541), .B(n_542), .Y(n_540) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_190), .A2(n_228), .B(n_236), .Y(n_227) );
AO21x2_ASAP7_75t_L g291 ( .A1(n_190), .A2(n_228), .B(n_236), .Y(n_291) );
AOI21x1_ASAP7_75t_L g548 ( .A1(n_190), .A2(n_549), .B(n_552), .Y(n_548) );
INVx2_ASAP7_75t_SL g190 ( .A(n_191), .Y(n_190) );
OA21x2_ASAP7_75t_L g238 ( .A1(n_191), .A2(n_239), .B(n_243), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_191), .A2(n_575), .B(n_576), .Y(n_574) );
AND2x4_ASAP7_75t_L g392 ( .A(n_192), .B(n_309), .Y(n_392) );
OR2x2_ASAP7_75t_L g433 ( .A(n_192), .B(n_434), .Y(n_433) );
NOR2xp67_ASAP7_75t_SL g452 ( .A(n_192), .B(n_325), .Y(n_452) );
NOR2x1_ASAP7_75t_L g470 ( .A(n_192), .B(n_384), .Y(n_470) );
INVx4_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NOR2x1_ASAP7_75t_SL g270 ( .A(n_193), .B(n_206), .Y(n_270) );
AND2x4_ASAP7_75t_L g308 ( .A(n_193), .B(n_309), .Y(n_308) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_193), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_193), .B(n_268), .Y(n_346) );
INVx2_ASAP7_75t_L g360 ( .A(n_193), .Y(n_360) );
NAND2xp5_ASAP7_75t_SL g382 ( .A(n_193), .B(n_312), .Y(n_382) );
AND2x2_ASAP7_75t_L g474 ( .A(n_193), .B(n_332), .Y(n_474) );
OR2x6_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NOR2x1_ASAP7_75t_L g202 ( .A(n_203), .B(n_222), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_204), .B(n_311), .Y(n_325) );
AND2x2_ASAP7_75t_SL g334 ( .A(n_204), .B(n_314), .Y(n_334) );
AND2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_221), .Y(n_204) );
INVx1_ASAP7_75t_L g312 ( .A(n_205), .Y(n_312) );
INVx3_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g332 ( .A(n_206), .Y(n_332) );
AND2x4_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
OAI21xp5_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_213), .B(n_220), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_212), .B(n_251), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_215), .B1(n_217), .B2(n_218), .Y(n_213) );
INVxp67_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVxp67_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g365 ( .A(n_221), .Y(n_365) );
INVx2_ASAP7_75t_SL g410 ( .A(n_222), .Y(n_410) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_244), .Y(n_224) );
NAND2x1p5_ASAP7_75t_L g319 ( .A(n_225), .B(n_320), .Y(n_319) );
BUFx2_ASAP7_75t_L g356 ( .A(n_225), .Y(n_356) );
AND2x2_ASAP7_75t_L g480 ( .A(n_225), .B(n_305), .Y(n_480) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_237), .Y(n_225) );
AND2x4_ASAP7_75t_L g293 ( .A(n_226), .B(n_275), .Y(n_293) );
INVx1_ASAP7_75t_L g304 ( .A(n_226), .Y(n_304) );
AND2x2_ASAP7_75t_L g335 ( .A(n_226), .B(n_290), .Y(n_335) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_227), .B(n_238), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_227), .B(n_276), .Y(n_367) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_229), .B(n_235), .Y(n_228) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVxp67_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g273 ( .A(n_238), .Y(n_273) );
AND2x4_ASAP7_75t_L g341 ( .A(n_238), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g353 ( .A(n_238), .Y(n_353) );
INVx1_ASAP7_75t_L g395 ( .A(n_238), .Y(n_395) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_238), .Y(n_407) );
AND2x2_ASAP7_75t_L g423 ( .A(n_238), .B(n_246), .Y(n_423) );
BUFx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g370 ( .A(n_245), .B(n_328), .Y(n_370) );
INVx1_ASAP7_75t_SL g372 ( .A(n_245), .Y(n_372) );
AND2x2_ASAP7_75t_L g393 ( .A(n_245), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x4_ASAP7_75t_L g272 ( .A(n_246), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g300 ( .A(n_246), .Y(n_300) );
INVx2_ASAP7_75t_L g306 ( .A(n_246), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_246), .B(n_276), .Y(n_321) );
OR2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_255), .Y(n_246) );
AO21x2_ASAP7_75t_L g276 ( .A1(n_254), .A2(n_277), .B(n_283), .Y(n_276) );
AO21x2_ASAP7_75t_L g290 ( .A1(n_254), .A2(n_277), .B(n_283), .Y(n_290) );
OAI22xp5_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_259), .B1(n_260), .B2(n_261), .Y(n_255) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OAI21xp5_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_266), .B(n_271), .Y(n_262) );
INVx1_ASAP7_75t_L g402 ( .A(n_263), .Y(n_402) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
INVx2_ASAP7_75t_L g322 ( .A(n_265), .Y(n_322) );
AND2x2_ASAP7_75t_L g378 ( .A(n_265), .B(n_314), .Y(n_378) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_270), .Y(n_266) );
INVx1_ASAP7_75t_L g292 ( .A(n_267), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_267), .B(n_308), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_267), .B(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g399 ( .A(n_267), .B(n_392), .Y(n_399) );
AND2x2_ASAP7_75t_L g473 ( .A(n_267), .B(n_474), .Y(n_473) );
INVx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_268), .Y(n_461) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_269), .Y(n_381) );
AND2x2_ASAP7_75t_L g294 ( .A(n_270), .B(n_295), .Y(n_294) );
OAI21xp33_ASAP7_75t_L g482 ( .A1(n_270), .A2(n_483), .B(n_485), .Y(n_482) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
INVx3_ASAP7_75t_L g368 ( .A(n_272), .Y(n_368) );
NAND2x1_ASAP7_75t_SL g412 ( .A(n_272), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g415 ( .A(n_272), .B(n_293), .Y(n_415) );
AND2x2_ASAP7_75t_L g327 ( .A(n_274), .B(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g464 ( .A(n_274), .B(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g475 ( .A(n_274), .B(n_423), .Y(n_475) );
INVx3_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2x1p5_ASAP7_75t_L g351 ( .A(n_275), .B(n_352), .Y(n_351) );
INVx3_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g406 ( .A(n_276), .B(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
OAI21xp5_ASAP7_75t_SL g284 ( .A1(n_285), .A2(n_298), .B(n_301), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_287), .B1(n_293), .B2(n_294), .Y(n_285) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_286), .Y(n_343) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_292), .Y(n_287) );
AND2x2_ASAP7_75t_L g316 ( .A(n_288), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g422 ( .A(n_288), .B(n_423), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_288), .A2(n_441), .B1(n_442), .B2(n_443), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_288), .B(n_449), .Y(n_448) );
AND2x4_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g305 ( .A(n_290), .B(n_306), .Y(n_305) );
NOR2xp67_ASAP7_75t_L g386 ( .A(n_290), .B(n_306), .Y(n_386) );
NOR2x1_ASAP7_75t_L g394 ( .A(n_290), .B(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g342 ( .A(n_291), .Y(n_342) );
AND2x2_ASAP7_75t_L g350 ( .A(n_291), .B(n_306), .Y(n_350) );
INVx1_ASAP7_75t_L g413 ( .A(n_291), .Y(n_413) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2x1_ASAP7_75t_L g331 ( .A(n_296), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g443 ( .A(n_299), .B(n_328), .Y(n_443) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g317 ( .A(n_300), .Y(n_317) );
AND2x2_ASAP7_75t_L g340 ( .A(n_300), .B(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g428 ( .A(n_300), .B(n_335), .Y(n_428) );
AOI22xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_307), .B1(n_313), .B2(n_316), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g436 ( .A(n_303), .B(n_437), .Y(n_436) );
NAND2x1p5_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
AND2x2_ASAP7_75t_L g466 ( .A(n_306), .B(n_353), .Y(n_466) );
AND2x2_ASAP7_75t_SL g307 ( .A(n_308), .B(n_310), .Y(n_307) );
INVx2_ASAP7_75t_L g333 ( .A(n_308), .Y(n_333) );
OAI21xp33_ASAP7_75t_SL g479 ( .A1(n_308), .A2(n_480), .B(n_481), .Y(n_479) );
AND2x4_ASAP7_75t_SL g310 ( .A(n_311), .B(n_312), .Y(n_310) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_311), .Y(n_469) );
AND2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
O2A1O1Ixp33_ASAP7_75t_SL g411 ( .A1(n_314), .A2(n_412), .B(n_414), .C(n_416), .Y(n_411) );
AND2x2_ASAP7_75t_SL g363 ( .A(n_315), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g416 ( .A(n_315), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_315), .B(n_392), .Y(n_456) );
INVx1_ASAP7_75t_SL g323 ( .A(n_316), .Y(n_323) );
AND2x2_ASAP7_75t_L g404 ( .A(n_317), .B(n_341), .Y(n_404) );
INVx1_ASAP7_75t_L g449 ( .A(n_317), .Y(n_449) );
OAI221xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_322), .B1(n_323), .B2(n_324), .C(n_326), .Y(n_318) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_319), .Y(n_438) );
INVx2_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g486 ( .A(n_321), .B(n_329), .Y(n_486) );
OR2x2_ASAP7_75t_L g345 ( .A(n_322), .B(n_346), .Y(n_345) );
NOR2x1_ASAP7_75t_L g358 ( .A(n_322), .B(n_359), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_322), .B(n_446), .Y(n_445) );
OR2x2_ASAP7_75t_L g484 ( .A(n_322), .B(n_381), .Y(n_484) );
BUFx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AOI32xp33_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_330), .A3(n_333), .B1(n_334), .B2(n_335), .Y(n_326) );
INVx1_ASAP7_75t_L g347 ( .A(n_328), .Y(n_347) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_330), .B(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g442 ( .A(n_331), .Y(n_442) );
OAI22xp33_ASAP7_75t_SL g424 ( .A1(n_333), .A2(n_425), .B1(n_427), .B2(n_429), .Y(n_424) );
INVx1_ASAP7_75t_L g455 ( .A(n_334), .Y(n_455) );
AOI211x1_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_343), .B(n_344), .C(n_361), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_340), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_338), .B(n_423), .Y(n_429) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x4_ASAP7_75t_L g385 ( .A(n_341), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g451 ( .A(n_341), .Y(n_451) );
OAI222xp33_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_347), .B1(n_348), .B2(n_354), .C1(n_355), .C2(n_357), .Y(n_344) );
INVxp67_ASAP7_75t_L g441 ( .A(n_345), .Y(n_441) );
OR2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_351), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_349), .B(n_434), .Y(n_481) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g397 ( .A(n_350), .B(n_394), .Y(n_397) );
INVx3_ASAP7_75t_L g437 ( .A(n_352), .Y(n_437) );
BUFx3_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g375 ( .A(n_360), .B(n_376), .Y(n_375) );
OAI221xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_366), .B1(n_369), .B2(n_374), .C(n_377), .Y(n_361) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
OAI21xp5_ASAP7_75t_L g419 ( .A1(n_363), .A2(n_420), .B(n_422), .Y(n_419) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
INVx1_ASAP7_75t_L g373 ( .A(n_367), .Y(n_373) );
OR2x2_ASAP7_75t_L g477 ( .A(n_368), .B(n_413), .Y(n_477) );
NOR2xp67_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_371), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
OAI21xp5_ASAP7_75t_L g471 ( .A1(n_374), .A2(n_403), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OAI21xp5_ASAP7_75t_L g453 ( .A1(n_375), .A2(n_447), .B(n_454), .Y(n_453) );
INVx4_ASAP7_75t_L g384 ( .A(n_376), .Y(n_384) );
OAI31xp33_ASAP7_75t_SL g377 ( .A1(n_378), .A2(n_379), .A3(n_383), .B(n_385), .Y(n_377) );
INVx1_ASAP7_75t_L g435 ( .A(n_379), .Y(n_435) );
NOR2x1_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g409 ( .A(n_384), .Y(n_409) );
AND2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_400), .Y(n_387) );
NAND4xp25_ASAP7_75t_L g488 ( .A(n_388), .B(n_400), .C(n_419), .D(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_398), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_393), .B1(n_396), .B2(n_397), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g460 ( .A(n_392), .B(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_393), .B(n_413), .Y(n_421) );
INVx1_ASAP7_75t_SL g434 ( .A(n_396), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_401), .B(n_411), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B1(n_405), .B2(n_408), .Y(n_401) );
INVx3_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NAND2x1_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_410), .A2(n_473), .B1(n_475), .B2(n_476), .Y(n_472) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NOR3xp33_ASAP7_75t_L g417 ( .A(n_418), .B(n_424), .C(n_430), .Y(n_417) );
INVxp67_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g489 ( .A(n_424), .Y(n_489) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OAI21xp33_ASAP7_75t_L g490 ( .A1(n_430), .A2(n_491), .B(n_492), .Y(n_490) );
INVxp33_ASAP7_75t_L g491 ( .A(n_431), .Y(n_491) );
AND2x2_ASAP7_75t_L g800 ( .A(n_431), .B(n_457), .Y(n_800) );
NOR2xp67_ASAP7_75t_L g431 ( .A(n_432), .B(n_439), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_435), .B1(n_436), .B2(n_438), .Y(n_432) );
OAI21xp5_ASAP7_75t_L g458 ( .A1(n_436), .A2(n_459), .B(n_462), .Y(n_458) );
INVx2_ASAP7_75t_L g446 ( .A(n_437), .Y(n_446) );
NAND3xp33_ASAP7_75t_SL g439 ( .A(n_440), .B(n_444), .C(n_453), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_447), .B1(n_450), .B2(n_452), .Y(n_444) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
INVxp33_ASAP7_75t_SL g492 ( .A(n_457), .Y(n_492) );
NOR3x1_ASAP7_75t_L g457 ( .A(n_458), .B(n_471), .C(n_478), .Y(n_457) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_463), .B(n_467), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_479), .B(n_482), .Y(n_478) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g802 ( .A(n_488), .Y(n_802) );
CKINVDCx11_ASAP7_75t_R g493 ( .A(n_494), .Y(n_493) );
INVx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x4_ASAP7_75t_L g496 ( .A(n_497), .B(n_660), .Y(n_496) );
NOR4xp25_ASAP7_75t_L g497 ( .A(n_498), .B(n_603), .C(n_642), .D(n_649), .Y(n_497) );
OAI221xp5_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_524), .B1(n_561), .B2(n_570), .C(n_589), .Y(n_498) );
OR2x2_ASAP7_75t_L g733 ( .A(n_499), .B(n_595), .Y(n_733) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g648 ( .A(n_500), .B(n_573), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_500), .B(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_SL g713 ( .A(n_500), .B(n_714), .Y(n_713) );
AND2x4_ASAP7_75t_L g500 ( .A(n_501), .B(n_513), .Y(n_500) );
AND2x4_ASAP7_75t_SL g572 ( .A(n_501), .B(n_573), .Y(n_572) );
INVx3_ASAP7_75t_L g594 ( .A(n_501), .Y(n_594) );
AND2x2_ASAP7_75t_L g629 ( .A(n_501), .B(n_602), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_501), .B(n_514), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_501), .B(n_596), .Y(n_681) );
OR2x2_ASAP7_75t_L g759 ( .A(n_501), .B(n_573), .Y(n_759) );
AND2x4_ASAP7_75t_L g501 ( .A(n_502), .B(n_507), .Y(n_501) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g581 ( .A(n_514), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_514), .B(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g607 ( .A(n_514), .Y(n_607) );
OR2x2_ASAP7_75t_L g612 ( .A(n_514), .B(n_596), .Y(n_612) );
AND2x2_ASAP7_75t_L g625 ( .A(n_514), .B(n_583), .Y(n_625) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_514), .Y(n_628) );
INVx1_ASAP7_75t_L g640 ( .A(n_514), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_514), .B(n_594), .Y(n_705) );
INVx3_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_521), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_525), .B(n_534), .Y(n_524) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OR2x2_ASAP7_75t_L g569 ( .A(n_526), .B(n_553), .Y(n_569) );
AND2x4_ASAP7_75t_L g599 ( .A(n_526), .B(n_538), .Y(n_599) );
INVx2_ASAP7_75t_L g633 ( .A(n_526), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_526), .B(n_553), .Y(n_691) );
AND2x2_ASAP7_75t_L g738 ( .A(n_526), .B(n_567), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_532), .Y(n_527) );
AOI222xp33_ASAP7_75t_L g726 ( .A1(n_534), .A2(n_598), .B1(n_641), .B2(n_701), .C1(n_727), .C2(n_729), .Y(n_726) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_546), .Y(n_535) );
AND2x2_ASAP7_75t_L g645 ( .A(n_536), .B(n_565), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_536), .B(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g774 ( .A(n_536), .B(n_614), .Y(n_774) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_537), .A2(n_605), .B(n_609), .Y(n_604) );
AND2x2_ASAP7_75t_L g685 ( .A(n_537), .B(n_568), .Y(n_685) );
OR2x2_ASAP7_75t_L g710 ( .A(n_537), .B(n_569), .Y(n_710) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx5_ASAP7_75t_L g564 ( .A(n_538), .Y(n_564) );
AND2x2_ASAP7_75t_L g651 ( .A(n_538), .B(n_633), .Y(n_651) );
AND2x2_ASAP7_75t_L g677 ( .A(n_538), .B(n_553), .Y(n_677) );
OR2x2_ASAP7_75t_L g680 ( .A(n_538), .B(n_567), .Y(n_680) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_538), .Y(n_698) );
AND2x4_ASAP7_75t_SL g755 ( .A(n_538), .B(n_632), .Y(n_755) );
OR2x2_ASAP7_75t_L g764 ( .A(n_538), .B(n_591), .Y(n_764) );
OR2x6_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
INVx1_ASAP7_75t_L g597 ( .A(n_546), .Y(n_597) );
AOI221xp5_ASAP7_75t_SL g715 ( .A1(n_546), .A2(n_599), .B1(n_716), .B2(n_718), .C(n_719), .Y(n_715) );
AND2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_553), .Y(n_546) );
OR2x2_ASAP7_75t_L g654 ( .A(n_547), .B(n_624), .Y(n_654) );
OR2x2_ASAP7_75t_L g664 ( .A(n_547), .B(n_665), .Y(n_664) );
OR2x2_ASAP7_75t_L g690 ( .A(n_547), .B(n_691), .Y(n_690) );
AND2x4_ASAP7_75t_L g696 ( .A(n_547), .B(n_615), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_547), .B(n_679), .Y(n_708) );
INVx2_ASAP7_75t_L g721 ( .A(n_547), .Y(n_721) );
NAND2xp5_ASAP7_75t_SL g742 ( .A(n_547), .B(n_599), .Y(n_742) );
AND2x2_ASAP7_75t_L g746 ( .A(n_547), .B(n_568), .Y(n_746) );
AND2x2_ASAP7_75t_L g754 ( .A(n_547), .B(n_755), .Y(n_754) );
BUFx6f_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g567 ( .A(n_548), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_553), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g598 ( .A(n_553), .B(n_567), .Y(n_598) );
INVx2_ASAP7_75t_L g615 ( .A(n_553), .Y(n_615) );
AND2x4_ASAP7_75t_L g632 ( .A(n_553), .B(n_633), .Y(n_632) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_553), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_559), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_562), .B(n_565), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OR2x2_ASAP7_75t_L g744 ( .A(n_563), .B(n_566), .Y(n_744) );
AND2x4_ASAP7_75t_L g590 ( .A(n_564), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g631 ( .A(n_564), .B(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g658 ( .A(n_564), .B(n_598), .Y(n_658) );
AND2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_568), .Y(n_565) );
AND2x2_ASAP7_75t_L g762 ( .A(n_566), .B(n_763), .Y(n_762) );
BUFx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g614 ( .A(n_567), .B(n_615), .Y(n_614) );
OAI21xp5_ASAP7_75t_SL g634 ( .A1(n_568), .A2(n_635), .B(n_641), .Y(n_634) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_581), .Y(n_571) );
INVx1_ASAP7_75t_SL g688 ( .A(n_572), .Y(n_688) );
AND2x2_ASAP7_75t_L g718 ( .A(n_572), .B(n_628), .Y(n_718) );
AND2x4_ASAP7_75t_L g729 ( .A(n_572), .B(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_L g595 ( .A(n_573), .B(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g602 ( .A(n_573), .Y(n_602) );
AND2x4_ASAP7_75t_L g608 ( .A(n_573), .B(n_594), .Y(n_608) );
INVx2_ASAP7_75t_L g619 ( .A(n_573), .Y(n_619) );
INVx1_ASAP7_75t_L g668 ( .A(n_573), .Y(n_668) );
OR2x2_ASAP7_75t_L g689 ( .A(n_573), .B(n_673), .Y(n_689) );
OR2x2_ASAP7_75t_L g703 ( .A(n_573), .B(n_583), .Y(n_703) );
HB1xp67_ASAP7_75t_L g769 ( .A(n_573), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_573), .B(n_625), .Y(n_775) );
OR2x6_ASAP7_75t_L g573 ( .A(n_574), .B(n_580), .Y(n_573) );
INVx1_ASAP7_75t_L g620 ( .A(n_581), .Y(n_620) );
AND2x2_ASAP7_75t_L g753 ( .A(n_581), .B(n_619), .Y(n_753) );
AND2x2_ASAP7_75t_L g778 ( .A(n_581), .B(n_608), .Y(n_778) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g596 ( .A(n_583), .Y(n_596) );
BUFx3_ASAP7_75t_L g638 ( .A(n_583), .Y(n_638) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_583), .Y(n_665) );
INVx1_ASAP7_75t_L g674 ( .A(n_583), .Y(n_674) );
AOI33xp33_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_592), .A3(n_597), .B1(n_598), .B2(n_599), .B3(n_600), .Y(n_589) );
AOI21x1_ASAP7_75t_SL g692 ( .A1(n_590), .A2(n_614), .B(n_676), .Y(n_692) );
INVx2_ASAP7_75t_L g722 ( .A(n_590), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_590), .B(n_721), .Y(n_728) );
AND2x2_ASAP7_75t_L g676 ( .A(n_591), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
AND2x2_ASAP7_75t_L g639 ( .A(n_594), .B(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g740 ( .A(n_595), .Y(n_740) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_596), .Y(n_730) );
OAI32xp33_ASAP7_75t_L g779 ( .A1(n_597), .A2(n_599), .A3(n_775), .B1(n_780), .B2(n_782), .Y(n_779) );
AND2x2_ASAP7_75t_L g697 ( .A(n_598), .B(n_698), .Y(n_697) );
INVx2_ASAP7_75t_SL g687 ( .A(n_599), .Y(n_687) );
AND2x2_ASAP7_75t_L g752 ( .A(n_599), .B(n_696), .Y(n_752) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
OAI221xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_613), .B1(n_616), .B2(n_630), .C(n_634), .Y(n_603) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_607), .B(n_674), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_608), .B(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_608), .B(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_608), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g657 ( .A(n_612), .Y(n_657) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NOR3xp33_ASAP7_75t_L g616 ( .A(n_617), .B(n_621), .C(n_626), .Y(n_616) );
INVx1_ASAP7_75t_SL g617 ( .A(n_618), .Y(n_617) );
OAI22xp33_ASAP7_75t_L g719 ( .A1(n_618), .A2(n_680), .B1(n_720), .B2(n_723), .Y(n_719) );
OR2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
INVx1_ASAP7_75t_L g623 ( .A(n_619), .Y(n_623) );
NOR2x1p5_ASAP7_75t_L g637 ( .A(n_619), .B(n_638), .Y(n_637) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_619), .Y(n_659) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
OAI322xp33_ASAP7_75t_L g686 ( .A1(n_622), .A2(n_664), .A3(n_687), .B1(n_688), .B2(n_689), .C1(n_690), .C2(n_692), .Y(n_686) );
OR2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
A2O1A1Ixp33_ASAP7_75t_L g642 ( .A1(n_624), .A2(n_643), .B(n_644), .C(n_646), .Y(n_642) );
OR2x2_ASAP7_75t_L g734 ( .A(n_624), .B(n_688), .Y(n_734) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g641 ( .A(n_625), .B(n_629), .Y(n_641) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g647 ( .A(n_631), .B(n_648), .Y(n_647) );
INVx3_ASAP7_75t_SL g679 ( .A(n_632), .Y(n_679) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_636), .B(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_637), .B(n_639), .Y(n_636) );
INVx1_ASAP7_75t_SL g683 ( .A(n_639), .Y(n_683) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_640), .Y(n_725) );
OR2x6_ASAP7_75t_SL g780 ( .A(n_643), .B(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVxp67_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AOI211xp5_ASAP7_75t_L g770 ( .A1(n_648), .A2(n_771), .B(n_772), .C(n_779), .Y(n_770) );
O2A1O1Ixp33_ASAP7_75t_SL g649 ( .A1(n_650), .A2(n_652), .B(n_655), .C(n_659), .Y(n_649) );
OAI211xp5_ASAP7_75t_SL g661 ( .A1(n_650), .A2(n_662), .B(n_669), .C(n_693), .Y(n_661) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx3_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVxp67_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
NOR3xp33_ASAP7_75t_L g660 ( .A(n_661), .B(n_706), .C(n_750), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_666), .Y(n_662) );
INVx1_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_665), .Y(n_757) );
INVx1_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g712 ( .A(n_668), .Y(n_712) );
NOR3xp33_ASAP7_75t_SL g669 ( .A(n_670), .B(n_682), .C(n_686), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_675), .B1(n_678), .B2(n_681), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g714 ( .A(n_674), .Y(n_714) );
INVxp67_ASAP7_75t_SL g781 ( .A(n_674), .Y(n_781) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OR2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
INVx1_ASAP7_75t_SL g767 ( .A(n_680), .Y(n_767) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
OR2x2_ASAP7_75t_L g717 ( .A(n_683), .B(n_703), .Y(n_717) );
OR2x2_ASAP7_75t_L g768 ( .A(n_683), .B(n_769), .Y(n_768) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g766 ( .A(n_691), .Y(n_766) );
OR2x2_ASAP7_75t_L g782 ( .A(n_691), .B(n_721), .Y(n_782) );
OAI21xp33_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_697), .B(n_699), .Y(n_693) );
OAI31xp33_ASAP7_75t_L g707 ( .A1(n_694), .A2(n_708), .A3(n_709), .B(n_711), .Y(n_707) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_702), .B(n_704), .Y(n_701) );
INVx1_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
AND2x4_ASAP7_75t_L g739 ( .A(n_704), .B(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NAND4xp25_ASAP7_75t_SL g706 ( .A(n_707), .B(n_715), .C(n_726), .D(n_731), .Y(n_706) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
HB1xp67_ASAP7_75t_L g749 ( .A(n_714), .Y(n_749) );
INVx1_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
OR2x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
INVxp67_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
AOI221xp5_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_735), .B1(n_739), .B2(n_741), .C(n_743), .Y(n_731) );
NAND2xp33_ASAP7_75t_SL g732 ( .A(n_733), .B(n_734), .Y(n_732) );
INVx1_ASAP7_75t_L g776 ( .A(n_735), .Y(n_776) );
AND2x2_ASAP7_75t_SL g735 ( .A(n_736), .B(n_738), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
AOI21xp33_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_745), .B(n_747), .Y(n_743) );
INVx1_ASAP7_75t_L g771 ( .A(n_745), .Y(n_771) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
NAND2xp5_ASAP7_75t_SL g750 ( .A(n_751), .B(n_770), .Y(n_750) );
AOI221xp5_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_753), .B1(n_754), .B2(n_756), .C(n_760), .Y(n_751) );
AND2x2_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
INVx1_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
AOI21xp33_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_765), .B(n_768), .Y(n_760) );
INVxp33_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_SL g763 ( .A(n_764), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_773), .A2(n_775), .B1(n_776), .B2(n_777), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
CKINVDCx5p33_ASAP7_75t_R g783 ( .A(n_784), .Y(n_783) );
CKINVDCx20_ASAP7_75t_R g789 ( .A(n_784), .Y(n_789) );
CKINVDCx11_ASAP7_75t_R g784 ( .A(n_785), .Y(n_784) );
CKINVDCx5p33_ASAP7_75t_R g790 ( .A(n_791), .Y(n_790) );
CKINVDCx5p33_ASAP7_75t_R g791 ( .A(n_792), .Y(n_791) );
INVx3_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
OAI22xp33_ASAP7_75t_SL g796 ( .A1(n_797), .A2(n_798), .B1(n_803), .B2(n_804), .Y(n_796) );
INVxp67_ASAP7_75t_SL g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
NAND3x1_ASAP7_75t_L g799 ( .A(n_800), .B(n_801), .C(n_802), .Y(n_799) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
endmodule