module real_jpeg_11205_n_17 (n_301, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_301;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_286;
wire n_288;
wire n_166;
wire n_221;
wire n_176;
wire n_215;
wire n_249;
wire n_292;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_299;
wire n_173;
wire n_243;
wire n_115;
wire n_255;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_167;
wire n_128;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

BUFx24_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_1),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_1),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

AOI21xp33_ASAP7_75t_L g221 ( 
.A1(n_1),
.A2(n_9),
.B(n_32),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_2),
.A2(n_27),
.B1(n_34),
.B2(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_2),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_2),
.A2(n_47),
.B1(n_48),
.B2(n_94),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_2),
.A2(n_63),
.B1(n_66),
.B2(n_94),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_94),
.Y(n_181)
);

BUFx10_ASAP7_75t_L g85 ( 
.A(n_3),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_4),
.Y(n_65)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

BUFx6f_ASAP7_75t_SL g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_8),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_8),
.A2(n_47),
.B1(n_48),
.B2(n_51),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_8),
.A2(n_51),
.B1(n_63),
.B2(n_66),
.Y(n_225)
);

A2O1A1O1Ixp25_ASAP7_75t_L g128 ( 
.A1(n_9),
.A2(n_48),
.B(n_58),
.C(n_129),
.D(n_130),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_9),
.B(n_48),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_9),
.B(n_46),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_9),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_9),
.A2(n_83),
.B(n_148),
.Y(n_165)
);

A2O1A1O1Ixp25_ASAP7_75t_L g178 ( 
.A1(n_9),
.A2(n_31),
.B(n_42),
.C(n_179),
.D(n_180),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_9),
.B(n_31),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_9),
.B(n_117),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_9),
.A2(n_27),
.B1(n_34),
.B2(n_161),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_10),
.A2(n_47),
.B1(n_48),
.B2(n_54),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_10),
.A2(n_54),
.B1(n_63),
.B2(n_66),
.Y(n_107)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_12),
.A2(n_27),
.B1(n_34),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_37),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_12),
.A2(n_37),
.B1(n_47),
.B2(n_48),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_12),
.A2(n_37),
.B1(n_63),
.B2(n_66),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_13),
.A2(n_47),
.B1(n_48),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_13),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_13),
.A2(n_63),
.B1(n_66),
.B2(n_69),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_14),
.A2(n_27),
.B1(n_34),
.B2(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_14),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_14),
.A2(n_63),
.B1(n_66),
.B2(n_115),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_14),
.A2(n_47),
.B1(n_48),
.B2(n_115),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_115),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_15),
.A2(n_27),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_35),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_15),
.A2(n_35),
.B1(n_63),
.B2(n_66),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_15),
.A2(n_35),
.B1(n_47),
.B2(n_48),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_16),
.A2(n_47),
.B1(n_48),
.B2(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_16),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_16),
.A2(n_63),
.B1(n_66),
.B2(n_143),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_16),
.A2(n_31),
.B1(n_32),
.B2(n_143),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_16),
.A2(n_27),
.B1(n_34),
.B2(n_143),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_120),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_118),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_96),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_20),
.B(n_96),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_79),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_71),
.B2(n_72),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_38),
.B2(n_39),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_30),
.B1(n_33),
.B2(n_36),
.Y(n_25)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_26),
.A2(n_114),
.B(n_116),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_26),
.A2(n_30),
.B1(n_114),
.B2(n_247),
.Y(n_267)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_28),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g220 ( 
.A1(n_27),
.A2(n_28),
.B(n_161),
.C(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_30),
.A2(n_33),
.B(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_30),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_L g246 ( 
.A1(n_30),
.A2(n_92),
.B(n_247),
.Y(n_246)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

O2A1O1Ixp33_ASAP7_75t_SL g42 ( 
.A1(n_32),
.A2(n_43),
.B(n_45),
.C(n_46),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_43),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_55),
.B1(n_56),
.B2(n_70),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_40),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_49),
.B1(n_52),
.B2(n_53),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_41),
.A2(n_52),
.B1(n_199),
.B2(n_235),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_41),
.A2(n_235),
.B(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_42),
.A2(n_46),
.B1(n_50),
.B2(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_42),
.A2(n_46),
.B1(n_74),
.B2(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_42),
.B(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_43),
.B(n_48),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_45),
.A2(n_47),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_46),
.Y(n_52)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

O2A1O1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_59),
.B(n_61),
.C(n_62),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_59),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_52),
.B(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_52),
.A2(n_199),
.B(n_200),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_52),
.A2(n_200),
.B(n_265),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_67),
.B(n_68),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_57),
.A2(n_67),
.B1(n_77),
.B2(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_57),
.A2(n_67),
.B1(n_89),
.B2(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_57),
.A2(n_67),
.B1(n_142),
.B2(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_57),
.A2(n_177),
.B(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_57),
.A2(n_67),
.B1(n_109),
.B2(n_232),
.Y(n_255)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_62),
.B1(n_76),
.B2(n_78),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_58),
.B(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_60),
.B1(n_63),
.B2(n_66),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_59),
.B(n_66),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_61),
.A2(n_63),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_63),
.Y(n_66)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_66),
.B(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_66),
.B(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_67),
.B(n_131),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_67),
.A2(n_142),
.B(n_144),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_67),
.B(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_67),
.A2(n_144),
.B(n_232),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_68),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_72),
.A2(n_73),
.B(n_75),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_90),
.B(n_91),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_81),
.B1(n_98),
.B2(n_100),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_88),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_82),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_90),
.B1(n_91),
.B2(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_82),
.A2(n_88),
.B1(n_90),
.B2(n_282),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_86),
.B(n_87),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_83),
.A2(n_86),
.B1(n_87),
.B2(n_107),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_83),
.A2(n_147),
.B(n_148),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_83),
.A2(n_86),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_83),
.A2(n_86),
.B1(n_107),
.B2(n_225),
.Y(n_254)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_84),
.A2(n_85),
.B1(n_153),
.B2(n_155),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_84),
.B(n_149),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_84),
.A2(n_85),
.B1(n_190),
.B2(n_205),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_85),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_85),
.B(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_86),
.A2(n_154),
.B(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_86),
.B(n_161),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_86),
.A2(n_163),
.B(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_88),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_91),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_93),
.B(n_117),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_95),
.A2(n_238),
.B(n_239),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_101),
.C(n_103),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_97),
.A2(n_101),
.B1(n_102),
.B2(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_97),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_98),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_103),
.A2(n_104),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_110),
.C(n_112),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_105),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_108),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_106),
.B(n_108),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_110),
.A2(n_112),
.B1(n_113),
.B2(n_280),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_110),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_111),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_116),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI321xp33_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_275),
.A3(n_288),
.B1(n_294),
.B2(n_299),
.C(n_301),
.Y(n_120)
);

NOR3xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_241),
.C(n_271),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_214),
.B(n_240),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_193),
.B(n_213),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_171),
.B(n_192),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_150),
.B(n_170),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_136),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_127),
.B(n_136),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_132),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_128),
.A2(n_132),
.B1(n_133),
.B2(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_129),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_130),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_131),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_146),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_141),
.C(n_146),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_147),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_158),
.B(n_169),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_156),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_152),
.B(n_156),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_164),
.B(n_168),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_160),
.B(n_162),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_172),
.B(n_173),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_184),
.B2(n_191),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_178),
.B1(n_182),
.B2(n_183),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_176),
.Y(n_183)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_178),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_183),
.C(n_191),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_179),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_180),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_181),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_184),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_188),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_194),
.B(n_195),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_207),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_209),
.C(n_211),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_202),
.B2(n_206),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_203),
.C(n_204),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_202),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_205),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_211),
.B2(n_212),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_208),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_209),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_215),
.B(n_216),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_229),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_218),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_218),
.B(n_228),
.C(n_229),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_222),
.B2(n_223),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_219),
.B(n_223),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_226),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_237),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_233),
.B1(n_234),
.B2(n_236),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_231),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_236),
.C(n_237),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

AOI21xp33_ASAP7_75t_L g295 ( 
.A1(n_242),
.A2(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_257),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_243),
.B(n_257),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_253),
.C(n_256),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_244),
.B(n_274),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_252),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_248),
.B1(n_249),
.B2(n_251),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_246),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_251),
.C(n_252),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_256),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_255),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_269),
.B2(n_270),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_260),
.B(n_261),
.C(n_270),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_266),
.C(n_268),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_264),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_269),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_273),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_284),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_276),
.B(n_284),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_281),
.C(n_283),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_277),
.A2(n_278),
.B1(n_281),
.B2(n_293),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_281),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_289),
.A2(n_295),
.B(n_298),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_290),
.B(n_291),
.Y(n_298)
);


endmodule