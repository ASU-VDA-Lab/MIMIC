module fake_jpeg_7072_n_43 (n_3, n_2, n_1, n_0, n_4, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

AND2x2_ASAP7_75t_SL g10 ( 
.A(n_5),
.B(n_2),
.Y(n_10)
);

BUFx10_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_10),
.B(n_0),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_18),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g15 ( 
.A(n_10),
.B(n_0),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_19),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_13),
.A2(n_4),
.B1(n_0),
.B2(n_1),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_17),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_13),
.A2(n_10),
.B1(n_6),
.B2(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_19),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_1),
.Y(n_21)
);

OA21x2_ASAP7_75t_L g26 ( 
.A1(n_21),
.A2(n_11),
.B(n_12),
.Y(n_26)
);

INVxp67_ASAP7_75t_SL g25 ( 
.A(n_21),
.Y(n_25)
);

INVxp33_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

OA21x2_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_15),
.B(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_28),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_31),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_23),
.A2(n_20),
.B1(n_18),
.B2(n_8),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_25),
.C(n_22),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_35),
.Y(n_38)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

NAND4xp25_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_26),
.C(n_24),
.D(n_9),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_26),
.C(n_9),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_37),
.B(n_9),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_24),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_39),
.B(n_4),
.Y(n_41)
);

A2O1A1O1Ixp25_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_41),
.B(n_39),
.C(n_4),
.D(n_38),
.Y(n_42)
);

AO21x1_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_38),
.B(n_8),
.Y(n_43)
);


endmodule