module real_jpeg_33837_n_11 (n_108, n_8, n_0, n_111, n_2, n_10, n_114, n_9, n_107, n_6, n_106, n_110, n_112, n_7, n_3, n_5, n_4, n_105, n_109, n_1, n_113, n_11);

input n_108;
input n_8;
input n_0;
input n_111;
input n_2;
input n_10;
input n_114;
input n_9;
input n_107;
input n_6;
input n_106;
input n_110;
input n_112;
input n_7;
input n_3;
input n_5;
input n_4;
input n_105;
input n_109;
input n_1;
input n_113;

output n_11;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx1_ASAP7_75t_L g78 ( 
.A(n_0),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_1),
.B(n_40),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_2),
.B(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_4),
.B(n_23),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_4),
.Y(n_101)
);

AOI221xp5_ASAP7_75t_L g61 ( 
.A1(n_5),
.A2(n_10),
.B1(n_62),
.B2(n_67),
.C(n_70),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_5),
.B(n_62),
.C(n_67),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_6),
.B(n_90),
.Y(n_89)
);

HAxp5_ASAP7_75t_SL g95 ( 
.A(n_6),
.B(n_96),
.CON(n_95),
.SN(n_95)
);

OAI22xp5_ASAP7_75t_L g12 ( 
.A1(n_7),
.A2(n_13),
.B1(n_14),
.B2(n_20),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_8),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_9),
.B(n_30),
.Y(n_98)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_10),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_21),
.Y(n_11)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_105),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

HB1xp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_27),
.B(n_99),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_23),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_36),
.B(n_97),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_35),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_89),
.B(n_95),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_48),
.B(n_87),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_47),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_80),
.C(n_81),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_74),
.B(n_79),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_61),
.B1(n_72),
.B2(n_73),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_63),
.B(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_111),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_78),
.Y(n_79)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx24_ASAP7_75t_SL g103 ( 
.A(n_95),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_106),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_107),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_108),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_109),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_110),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_112),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_113),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_114),
.Y(n_91)
);


endmodule