module fake_ariane_464_n_1226 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1226);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1226;

wire n_295;
wire n_356;
wire n_556;
wire n_190;
wire n_698;
wire n_1127;
wire n_1072;
wire n_695;
wire n_913;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_1209;
wire n_1137;
wire n_646;
wire n_1174;
wire n_197;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_176;
wire n_691;
wire n_1214;
wire n_404;
wire n_172;
wire n_943;
wire n_1118;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_423;
wire n_347;
wire n_1042;
wire n_961;
wire n_183;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_1123;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_1169;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_1029;
wire n_341;
wire n_1187;
wire n_985;
wire n_421;
wire n_245;
wire n_1167;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_1180;
wire n_969;
wire n_283;
wire n_1109;
wire n_919;
wire n_187;
wire n_525;
wire n_806;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_643;
wire n_679;
wire n_244;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_261;
wire n_220;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_952;
wire n_864;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_1154;
wire n_1166;
wire n_387;
wire n_1200;
wire n_406;
wire n_826;
wire n_1130;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_756;
wire n_466;
wire n_940;
wire n_1016;
wire n_346;
wire n_1138;
wire n_214;
wire n_1149;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_1196;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_1181;
wire n_379;
wire n_515;
wire n_445;
wire n_807;
wire n_765;
wire n_1131;
wire n_264;
wire n_891;
wire n_1225;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_1217;
wire n_385;
wire n_637;
wire n_917;
wire n_1208;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_1177;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_1170;
wire n_1151;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_905;
wire n_279;
wire n_945;
wire n_702;
wire n_958;
wire n_207;
wire n_790;
wire n_898;
wire n_857;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_194;
wire n_1064;
wire n_633;
wire n_900;
wire n_1133;
wire n_883;
wire n_338;
wire n_1163;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_186;
wire n_801;
wire n_1184;
wire n_202;
wire n_193;
wire n_761;
wire n_733;
wire n_818;
wire n_500;
wire n_665;
wire n_754;
wire n_336;
wire n_779;
wire n_731;
wire n_871;
wire n_315;
wire n_903;
wire n_1073;
wire n_594;
wire n_1173;
wire n_311;
wire n_239;
wire n_402;
wire n_1052;
wire n_1068;
wire n_272;
wire n_829;
wire n_1198;
wire n_1062;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_1117;
wire n_422;
wire n_1106;
wire n_648;
wire n_784;
wire n_597;
wire n_269;
wire n_816;
wire n_1018;
wire n_855;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_1224;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_1125;
wire n_625;
wire n_405;
wire n_557;
wire n_1201;
wire n_1107;
wire n_173;
wire n_858;
wire n_645;
wire n_242;
wire n_989;
wire n_320;
wire n_331;
wire n_309;
wire n_559;
wire n_1134;
wire n_1185;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_1141;
wire n_350;
wire n_291;
wire n_822;
wire n_1143;
wire n_381;
wire n_344;
wire n_840;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_1053;
wire n_795;
wire n_1084;
wire n_398;
wire n_210;
wire n_1090;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_821;
wire n_839;
wire n_1099;
wire n_928;
wire n_271;
wire n_1153;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_569;
wire n_247;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_1145;
wire n_971;
wire n_369;
wire n_240;
wire n_1192;
wire n_224;
wire n_894;
wire n_787;
wire n_1105;
wire n_547;
wire n_1195;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_1172;
wire n_478;
wire n_703;
wire n_222;
wire n_1207;
wire n_748;
wire n_1212;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_1160;
wire n_874;
wire n_188;
wire n_323;
wire n_550;
wire n_1023;
wire n_997;
wire n_635;
wire n_707;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_1116;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1113;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_301;
wire n_248;
wire n_467;
wire n_1085;
wire n_1152;
wire n_432;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_1197;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_1165;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_206;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_192;
wire n_1128;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1122;
wire n_1049;
wire n_1205;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_1132;
wire n_390;
wire n_1156;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_1120;
wire n_440;
wire n_1202;
wire n_627;
wire n_1039;
wire n_1188;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_1150;
wire n_233;
wire n_728;
wire n_957;
wire n_388;
wire n_449;
wire n_333;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_977;
wire n_1216;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_1218;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_321;
wire n_221;
wire n_1136;
wire n_911;
wire n_361;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_623;
wire n_838;
wire n_1213;
wire n_237;
wire n_780;
wire n_861;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_1119;
wire n_734;
wire n_491;
wire n_810;
wire n_181;
wire n_723;
wire n_1142;
wire n_616;
wire n_617;
wire n_705;
wire n_658;
wire n_630;
wire n_1140;
wire n_570;
wire n_1055;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_1121;
wire n_209;
wire n_490;
wire n_262;
wire n_743;
wire n_1194;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_1112;
wire n_700;
wire n_1159;
wire n_910;
wire n_1210;
wire n_290;
wire n_527;
wire n_772;
wire n_741;
wire n_747;
wire n_847;
wire n_939;
wire n_1135;
wire n_371;
wire n_888;
wire n_845;
wire n_199;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_1114;
wire n_676;
wire n_178;
wire n_708;
wire n_551;
wire n_308;
wire n_1223;
wire n_417;
wire n_201;
wire n_1038;
wire n_572;
wire n_343;
wire n_1199;
wire n_865;
wire n_1222;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_860;
wire n_534;
wire n_249;
wire n_1108;
wire n_355;
wire n_444;
wire n_609;
wire n_212;
wire n_278;
wire n_1043;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_1193;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_1179;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_1081;
wire n_182;
wire n_696;
wire n_1040;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_1158;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_774;
wire n_407;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_1168;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_1157;
wire n_555;
wire n_492;
wire n_234;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_252;
wire n_629;
wire n_664;
wire n_215;
wire n_1075;
wire n_454;
wire n_992;
wire n_966;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_1182;
wire n_763;
wire n_655;
wire n_540;
wire n_544;
wire n_216;
wire n_692;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_179;
wire n_812;
wire n_1126;
wire n_395;
wire n_621;
wire n_851;
wire n_1178;
wire n_195;
wire n_606;
wire n_1026;
wire n_951;
wire n_213;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_583;
wire n_509;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_1206;
wire n_378;
wire n_203;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1146;
wire n_1100;
wire n_1171;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_1203;
wire n_619;
wire n_337;
wire n_437;
wire n_697;
wire n_274;
wire n_622;
wire n_967;
wire n_998;
wire n_999;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_174;
wire n_275;
wire n_704;
wire n_1060;
wire n_1175;
wire n_1044;
wire n_1148;
wire n_204;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_1211;
wire n_963;
wire n_873;
wire n_1082;
wire n_1139;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_1221;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_1115;
wire n_824;
wire n_428;
wire n_1002;
wire n_580;
wire n_358;
wire n_1051;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_1101;
wire n_975;
wire n_1102;
wire n_1129;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_1189;
wire n_1124;
wire n_250;
wire n_932;
wire n_1183;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_1110;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_944;
wire n_749;
wire n_1204;
wire n_994;
wire n_548;
wire n_289;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_650;
wire n_258;
wire n_782;
wire n_856;
wire n_425;
wire n_1161;
wire n_431;
wire n_1176;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1155;
wire n_1191;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_767;
wire n_736;
wire n_1025;
wire n_1164;
wire n_1215;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_1011;
wire n_211;
wire n_642;
wire n_978;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_1147;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_1220;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_148),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_92),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_9),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_164),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_79),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_38),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_145),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_32),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_103),
.Y(n_181)
);

BUFx10_ASAP7_75t_L g182 ( 
.A(n_169),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_93),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_121),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_19),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_127),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_69),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_56),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_99),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_150),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_16),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_162),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_86),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_101),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_50),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_9),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_81),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_137),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_120),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_50),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_37),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_12),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_160),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_67),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_14),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_35),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_40),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_168),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_24),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_117),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_135),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_65),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_139),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_163),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_154),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_144),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_153),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_62),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_10),
.Y(n_219)
);

BUFx5_ASAP7_75t_L g220 ( 
.A(n_88),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_132),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_170),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_155),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_104),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_146),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_45),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_0),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_49),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_124),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_45),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_83),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_28),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_152),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_122),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_119),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_156),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_25),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_64),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_90),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_141),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_123),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_54),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_78),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_100),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_91),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_165),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_80),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_138),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_136),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_18),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_63),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_116),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_41),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_161),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_110),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_13),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_27),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_126),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_85),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_167),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_41),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_166),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_158),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_131),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_74),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_24),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_107),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_159),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_142),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_171),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_15),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_57),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_34),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_102),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_46),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_32),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_10),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_17),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_149),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_94),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_96),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_25),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_12),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_115),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_17),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_20),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_0),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_71),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_106),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_38),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_49),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_53),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_261),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_174),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_266),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_261),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_256),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_191),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_217),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_195),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_261),
.Y(n_301)
);

NOR2xp67_ASAP7_75t_L g302 ( 
.A(n_178),
.B(n_1),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_179),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_196),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_261),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_283),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_197),
.B(n_1),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_200),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_202),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_R g310 ( 
.A(n_179),
.B(n_52),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_283),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_283),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_205),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_207),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_283),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_232),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_209),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_185),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_219),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_206),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_237),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_208),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_208),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_226),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_271),
.B(n_2),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_214),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_228),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_259),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_232),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_271),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_243),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_253),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_250),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_214),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_257),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_275),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_238),
.B(n_2),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_R g338 ( 
.A(n_259),
.B(n_55),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_182),
.B(n_3),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_291),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_277),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_273),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_260),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_278),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_276),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_290),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_282),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_292),
.B(n_3),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_291),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_260),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_172),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_173),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_285),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_176),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_287),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_177),
.Y(n_356)
);

NOR2xp67_ASAP7_75t_L g357 ( 
.A(n_251),
.B(n_4),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_267),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_192),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_181),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_190),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_201),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_193),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_183),
.B(n_4),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_189),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_180),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_267),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_194),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_210),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_268),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_198),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_268),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_180),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_213),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_229),
.B(n_5),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_233),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_235),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_236),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_239),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_199),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_252),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_182),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_227),
.Y(n_383)
);

AND3x2_ASAP7_75t_L g384 ( 
.A(n_339),
.B(n_362),
.C(n_307),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_293),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_356),
.B(n_360),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_293),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_326),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_296),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_365),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_296),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_301),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_301),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_305),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_305),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_306),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_306),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_351),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_330),
.B(n_182),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_325),
.B(n_326),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_311),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_311),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_356),
.B(n_263),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_312),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_297),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_352),
.B(n_248),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_365),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_354),
.Y(n_408)
);

AND2x6_ASAP7_75t_L g409 ( 
.A(n_339),
.B(n_175),
.Y(n_409)
);

OR2x2_ASAP7_75t_L g410 ( 
.A(n_330),
.B(n_251),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_312),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_382),
.B(n_184),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_315),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_349),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_315),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_382),
.B(n_184),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_325),
.B(n_279),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_360),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_316),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_368),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_368),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_369),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_369),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_374),
.B(n_186),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_374),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_376),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_376),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_378),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_378),
.B(n_186),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_379),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_334),
.B(n_175),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_379),
.B(n_187),
.Y(n_432)
);

OA21x2_ASAP7_75t_L g433 ( 
.A1(n_375),
.A2(n_188),
.B(n_187),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_381),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_381),
.B(n_188),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_377),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_318),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_334),
.B(n_175),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_329),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_377),
.B(n_246),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_318),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_320),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_320),
.Y(n_443)
);

OAI21x1_ASAP7_75t_L g444 ( 
.A1(n_337),
.A2(n_220),
.B(n_175),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_324),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_324),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_327),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_340),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_327),
.B(n_254),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_332),
.Y(n_450)
);

NAND2xp33_ASAP7_75t_L g451 ( 
.A(n_361),
.B(n_220),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_332),
.Y(n_452)
);

NAND2x1p5_ASAP7_75t_L g453 ( 
.A(n_357),
.B(n_265),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_389),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_398),
.B(n_299),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_385),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_387),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_434),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_434),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_388),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_409),
.A2(n_348),
.B1(n_364),
.B2(n_357),
.Y(n_461)
);

OR2x6_ASAP7_75t_L g462 ( 
.A(n_453),
.B(n_302),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_388),
.B(n_436),
.Y(n_463)
);

AO22x2_ASAP7_75t_L g464 ( 
.A1(n_410),
.A2(n_359),
.B1(n_363),
.B2(n_294),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_387),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_385),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_388),
.B(n_371),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_434),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_391),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_385),
.Y(n_470)
);

AND3x2_ASAP7_75t_L g471 ( 
.A(n_405),
.B(n_383),
.C(n_366),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_394),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_391),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_392),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_392),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_434),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_L g477 ( 
.A1(n_409),
.A2(n_302),
.B1(n_353),
.B2(n_338),
.Y(n_477)
);

OAI22xp33_ASAP7_75t_L g478 ( 
.A1(n_410),
.A2(n_227),
.B1(n_230),
.B2(n_286),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_434),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_436),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g481 ( 
.A(n_408),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_393),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_393),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_394),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_396),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_406),
.B(n_299),
.Y(n_486)
);

AND2x2_ASAP7_75t_SL g487 ( 
.A(n_433),
.B(n_331),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_396),
.Y(n_488)
);

BUFx6f_ASAP7_75t_SL g489 ( 
.A(n_409),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_397),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_436),
.B(n_380),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_436),
.B(n_336),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_394),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_397),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_409),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_412),
.B(n_331),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_401),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_409),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_401),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_409),
.Y(n_500)
);

BUFx10_ASAP7_75t_L g501 ( 
.A(n_409),
.Y(n_501)
);

INVx5_ASAP7_75t_L g502 ( 
.A(n_409),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_419),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_395),
.Y(n_504)
);

INVx6_ASAP7_75t_L g505 ( 
.A(n_431),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_443),
.B(n_336),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_443),
.B(n_341),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_402),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_402),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_435),
.B(n_298),
.Y(n_510)
);

AOI22xp33_ASAP7_75t_L g511 ( 
.A1(n_437),
.A2(n_310),
.B1(n_355),
.B2(n_344),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_395),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_395),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_404),
.Y(n_514)
);

BUFx4f_ASAP7_75t_L g515 ( 
.A(n_433),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_404),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_411),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_413),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_414),
.Y(n_519)
);

OAI22xp33_ASAP7_75t_L g520 ( 
.A1(n_453),
.A2(n_230),
.B1(n_286),
.B2(n_341),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_435),
.B(n_344),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_413),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_411),
.Y(n_523)
);

CKINVDCx11_ASAP7_75t_R g524 ( 
.A(n_450),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_467),
.B(n_511),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_521),
.B(n_400),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_487),
.A2(n_433),
.B1(n_453),
.B2(n_417),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_491),
.B(n_400),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_491),
.B(n_400),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_503),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_457),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_521),
.B(n_400),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_496),
.B(n_486),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_461),
.A2(n_417),
.B1(n_448),
.B2(n_439),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_521),
.B(n_399),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_510),
.B(n_416),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_467),
.B(n_492),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_495),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_457),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_456),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_503),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_511),
.B(n_439),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_495),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_487),
.A2(n_417),
.B1(n_433),
.B2(n_427),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_492),
.B(n_399),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_465),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_477),
.B(n_448),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_481),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_506),
.B(n_440),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_465),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_456),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_481),
.B(n_419),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_469),
.Y(n_553)
);

NAND2xp33_ASAP7_75t_SL g554 ( 
.A(n_519),
.B(n_424),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_456),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g556 ( 
.A(n_462),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_506),
.B(n_440),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_469),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_507),
.B(n_417),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_507),
.B(n_424),
.Y(n_560)
);

OAI22xp33_ASAP7_75t_L g561 ( 
.A1(n_462),
.A2(n_403),
.B1(n_386),
.B2(n_449),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_464),
.B(n_300),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_462),
.B(n_429),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_462),
.B(n_429),
.Y(n_564)
);

BUFx8_ASAP7_75t_L g565 ( 
.A(n_489),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_462),
.B(n_295),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_473),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_487),
.A2(n_433),
.B1(n_426),
.B2(n_427),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_462),
.B(n_432),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_466),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_L g571 ( 
.A1(n_515),
.A2(n_444),
.B(n_451),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_477),
.B(n_432),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_495),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_473),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_520),
.B(n_304),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_463),
.B(n_449),
.Y(n_576)
);

NOR3xp33_ASAP7_75t_L g577 ( 
.A(n_520),
.B(n_443),
.C(n_386),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_463),
.B(n_480),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_455),
.B(n_308),
.Y(n_579)
);

OAI21xp5_ASAP7_75t_L g580 ( 
.A1(n_515),
.A2(n_444),
.B(n_403),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_471),
.Y(n_581)
);

AO221x1_ASAP7_75t_L g582 ( 
.A1(n_478),
.A2(n_384),
.B1(n_443),
.B2(n_270),
.C(n_434),
.Y(n_582)
);

A2O1A1Ixp33_ASAP7_75t_L g583 ( 
.A1(n_515),
.A2(n_444),
.B(n_420),
.C(n_422),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_480),
.B(n_418),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_474),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_505),
.B(n_309),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_478),
.B(n_313),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_480),
.B(n_418),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_464),
.B(n_421),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_466),
.Y(n_590)
);

NAND2xp33_ASAP7_75t_L g591 ( 
.A(n_500),
.B(n_421),
.Y(n_591)
);

NAND2x1p5_ASAP7_75t_L g592 ( 
.A(n_498),
.B(n_431),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_474),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_464),
.B(n_422),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_464),
.B(n_423),
.Y(n_595)
);

NAND2x1_ASAP7_75t_L g596 ( 
.A(n_500),
.B(n_423),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_500),
.B(n_314),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_464),
.B(n_425),
.Y(n_598)
);

BUFx5_ASAP7_75t_L g599 ( 
.A(n_501),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_475),
.B(n_425),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_475),
.B(n_428),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_498),
.B(n_317),
.Y(n_602)
);

BUFx5_ASAP7_75t_L g603 ( 
.A(n_501),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_471),
.B(n_319),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_482),
.B(n_428),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_505),
.B(n_321),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_498),
.A2(n_426),
.B1(n_427),
.B2(n_452),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_505),
.B(n_333),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_501),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_505),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_505),
.A2(n_430),
.B1(n_384),
.B2(n_346),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_460),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_482),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_483),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_483),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_485),
.B(n_430),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_460),
.B(n_335),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_460),
.B(n_342),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_485),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_488),
.B(n_431),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_488),
.B(n_431),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_552),
.B(n_303),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_545),
.B(n_441),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_537),
.A2(n_578),
.B(n_560),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_561),
.B(n_515),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_533),
.B(n_458),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_540),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_576),
.B(n_549),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_551),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_528),
.A2(n_499),
.B1(n_523),
.B2(n_497),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_531),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_561),
.B(n_454),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_557),
.A2(n_459),
.B(n_458),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_530),
.B(n_322),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_525),
.A2(n_372),
.B1(n_370),
.B2(n_323),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_526),
.B(n_502),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_535),
.B(n_441),
.Y(n_637)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_526),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_529),
.A2(n_459),
.B(n_458),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_571),
.A2(n_459),
.B(n_458),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_539),
.Y(n_641)
);

AO21x1_ASAP7_75t_L g642 ( 
.A1(n_580),
.A2(n_572),
.B(n_564),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_581),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_547),
.B(n_459),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_582),
.A2(n_490),
.B1(n_523),
.B2(n_494),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_546),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_538),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_555),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_586),
.B(n_442),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_584),
.A2(n_476),
.B(n_468),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_588),
.A2(n_476),
.B(n_468),
.Y(n_651)
);

OAI21xp5_ASAP7_75t_L g652 ( 
.A1(n_583),
.A2(n_494),
.B(n_490),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_550),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_606),
.B(n_442),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_608),
.B(n_445),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_559),
.A2(n_476),
.B(n_468),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_530),
.B(n_468),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_532),
.B(n_445),
.Y(n_658)
);

AND2x4_ASAP7_75t_L g659 ( 
.A(n_556),
.B(n_502),
.Y(n_659)
);

INVx4_ASAP7_75t_L g660 ( 
.A(n_538),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_563),
.B(n_454),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_577),
.B(n_446),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_577),
.B(n_446),
.Y(n_663)
);

AND2x2_ASAP7_75t_SL g664 ( 
.A(n_527),
.B(n_438),
.Y(n_664)
);

INVx11_ASAP7_75t_L g665 ( 
.A(n_565),
.Y(n_665)
);

OAI22xp5_ASAP7_75t_L g666 ( 
.A1(n_553),
.A2(n_508),
.B1(n_517),
.B2(n_516),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_541),
.B(n_328),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_534),
.B(n_447),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_591),
.A2(n_601),
.B(n_600),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_570),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_542),
.B(n_447),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_605),
.A2(n_479),
.B(n_476),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_538),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_558),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_616),
.A2(n_479),
.B(n_508),
.Y(n_675)
);

OAI22xp5_ASAP7_75t_L g676 ( 
.A1(n_567),
.A2(n_514),
.B1(n_509),
.B2(n_517),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_541),
.B(n_426),
.Y(n_677)
);

O2A1O1Ixp33_ASAP7_75t_L g678 ( 
.A1(n_574),
.A2(n_516),
.B(n_514),
.C(n_509),
.Y(n_678)
);

INVx5_ASAP7_75t_L g679 ( 
.A(n_538),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_536),
.A2(n_350),
.B1(n_358),
.B2(n_367),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_569),
.B(n_454),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_590),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_543),
.B(n_573),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_585),
.Y(n_684)
);

O2A1O1Ixp33_ASAP7_75t_L g685 ( 
.A1(n_593),
.A2(n_479),
.B(n_437),
.C(n_452),
.Y(n_685)
);

NOR3xp33_ASAP7_75t_L g686 ( 
.A(n_554),
.B(n_345),
.C(n_347),
.Y(n_686)
);

BUFx3_ASAP7_75t_L g687 ( 
.A(n_604),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_613),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_596),
.A2(n_479),
.B(n_470),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_614),
.B(n_450),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_615),
.B(n_450),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_619),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_556),
.B(n_450),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_562),
.B(n_610),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_620),
.A2(n_470),
.B(n_466),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_543),
.B(n_454),
.Y(n_696)
);

NOR2xp67_ASAP7_75t_L g697 ( 
.A(n_548),
.B(n_390),
.Y(n_697)
);

AOI21xp5_ASAP7_75t_L g698 ( 
.A1(n_621),
.A2(n_472),
.B(n_470),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_589),
.B(n_450),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_612),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_543),
.B(n_454),
.Y(n_701)
);

OAI21xp33_ASAP7_75t_L g702 ( 
.A1(n_548),
.A2(n_343),
.B(n_437),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_543),
.Y(n_703)
);

INVxp67_ASAP7_75t_L g704 ( 
.A(n_594),
.Y(n_704)
);

NOR3xp33_ASAP7_75t_L g705 ( 
.A(n_579),
.B(n_355),
.C(n_347),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_544),
.A2(n_489),
.B1(n_502),
.B2(n_452),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_565),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_587),
.B(n_373),
.Y(n_708)
);

BUFx4f_ASAP7_75t_L g709 ( 
.A(n_592),
.Y(n_709)
);

INVxp67_ASAP7_75t_L g710 ( 
.A(n_595),
.Y(n_710)
);

HB1xp67_ASAP7_75t_L g711 ( 
.A(n_573),
.Y(n_711)
);

INVx8_ASAP7_75t_L g712 ( 
.A(n_573),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_L g713 ( 
.A1(n_597),
.A2(n_484),
.B(n_472),
.Y(n_713)
);

BUFx2_ASAP7_75t_L g714 ( 
.A(n_611),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_612),
.A2(n_484),
.B(n_472),
.Y(n_715)
);

O2A1O1Ixp33_ASAP7_75t_L g716 ( 
.A1(n_617),
.A2(n_484),
.B(n_522),
.C(n_518),
.Y(n_716)
);

NAND3xp33_ASAP7_75t_L g717 ( 
.A(n_705),
.B(n_575),
.C(n_618),
.Y(n_717)
);

NAND2x2_ASAP7_75t_L g718 ( 
.A(n_707),
.B(n_5),
.Y(n_718)
);

A2O1A1Ixp33_ASAP7_75t_L g719 ( 
.A1(n_628),
.A2(n_544),
.B(n_598),
.C(n_566),
.Y(n_719)
);

AOI21xp5_ASAP7_75t_L g720 ( 
.A1(n_624),
.A2(n_602),
.B(n_609),
.Y(n_720)
);

A2O1A1Ixp33_ASAP7_75t_L g721 ( 
.A1(n_626),
.A2(n_568),
.B(n_607),
.C(n_512),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_626),
.B(n_573),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_631),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_634),
.A2(n_524),
.B1(n_592),
.B2(n_607),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_705),
.B(n_390),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_667),
.B(n_450),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_627),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_680),
.B(n_568),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_673),
.Y(n_729)
);

O2A1O1Ixp33_ASAP7_75t_L g730 ( 
.A1(n_686),
.A2(n_407),
.B(n_390),
.C(n_522),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_714),
.A2(n_489),
.B1(n_438),
.B2(n_504),
.Y(n_731)
);

O2A1O1Ixp5_ASAP7_75t_L g732 ( 
.A1(n_625),
.A2(n_512),
.B(n_493),
.C(n_504),
.Y(n_732)
);

NAND2x1p5_ASAP7_75t_L g733 ( 
.A(n_709),
.B(n_609),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_622),
.B(n_454),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_L g735 ( 
.A1(n_668),
.A2(n_390),
.B1(n_407),
.B2(n_518),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_629),
.Y(n_736)
);

AOI21x1_ASAP7_75t_L g737 ( 
.A1(n_625),
.A2(n_504),
.B(n_493),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_669),
.A2(n_609),
.B(n_502),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_665),
.Y(n_739)
);

OAI21xp5_ASAP7_75t_L g740 ( 
.A1(n_652),
.A2(n_512),
.B(n_493),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_635),
.B(n_454),
.Y(n_741)
);

A2O1A1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_678),
.A2(n_644),
.B(n_663),
.C(n_662),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_649),
.A2(n_609),
.B(n_502),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_641),
.Y(n_744)
);

NOR3xp33_ASAP7_75t_SL g745 ( 
.A(n_657),
.B(n_204),
.C(n_203),
.Y(n_745)
);

INVx4_ASAP7_75t_L g746 ( 
.A(n_709),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_702),
.B(n_513),
.Y(n_747)
);

OAI22xp5_ASAP7_75t_L g748 ( 
.A1(n_658),
.A2(n_407),
.B1(n_518),
.B2(n_513),
.Y(n_748)
);

AOI21x1_ASAP7_75t_L g749 ( 
.A1(n_632),
.A2(n_522),
.B(n_513),
.Y(n_749)
);

OAI22x1_ASAP7_75t_L g750 ( 
.A1(n_708),
.A2(n_407),
.B1(n_438),
.B2(n_281),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_654),
.A2(n_502),
.B(n_599),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_646),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_638),
.B(n_438),
.Y(n_753)
);

AO32x2_ASAP7_75t_L g754 ( 
.A1(n_630),
.A2(n_415),
.A3(n_413),
.B1(n_389),
.B2(n_11),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_636),
.B(n_502),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_686),
.A2(n_489),
.B1(n_599),
.B2(n_603),
.Y(n_756)
);

BUFx4f_ASAP7_75t_L g757 ( 
.A(n_636),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_638),
.B(n_415),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_653),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_637),
.B(n_415),
.Y(n_760)
);

AND2x2_ASAP7_75t_SL g761 ( 
.A(n_664),
.B(n_270),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_643),
.B(n_389),
.Y(n_762)
);

HB1xp67_ASAP7_75t_L g763 ( 
.A(n_700),
.Y(n_763)
);

A2O1A1Ixp33_ASAP7_75t_SL g764 ( 
.A1(n_657),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_764)
);

HB1xp67_ASAP7_75t_L g765 ( 
.A(n_694),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_655),
.A2(n_603),
.B(n_599),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_674),
.B(n_269),
.Y(n_767)
);

OAI21xp33_ASAP7_75t_L g768 ( 
.A1(n_623),
.A2(n_211),
.B(n_212),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_697),
.A2(n_599),
.B1(n_603),
.B2(n_501),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_684),
.B(n_215),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_688),
.B(n_216),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_692),
.B(n_599),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_704),
.B(n_603),
.Y(n_773)
);

HB1xp67_ASAP7_75t_L g774 ( 
.A(n_711),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_679),
.B(n_603),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_677),
.B(n_6),
.Y(n_776)
);

AO32x1_ASAP7_75t_L g777 ( 
.A1(n_666),
.A2(n_389),
.A3(n_8),
.B1(n_11),
.B2(n_13),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_640),
.A2(n_247),
.B(n_289),
.Y(n_778)
);

NOR2xp67_ASAP7_75t_L g779 ( 
.A(n_707),
.B(n_218),
.Y(n_779)
);

OAI21x1_ASAP7_75t_L g780 ( 
.A1(n_713),
.A2(n_220),
.B(n_389),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_761),
.A2(n_664),
.B1(n_676),
.B2(n_645),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_763),
.B(n_687),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_728),
.B(n_704),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_766),
.A2(n_632),
.B(n_696),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_723),
.Y(n_785)
);

BUFx2_ASAP7_75t_L g786 ( 
.A(n_774),
.Y(n_786)
);

OAI21x1_ASAP7_75t_L g787 ( 
.A1(n_780),
.A2(n_642),
.B(n_695),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_734),
.B(n_710),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_744),
.Y(n_789)
);

AO31x2_ASAP7_75t_L g790 ( 
.A1(n_721),
.A2(n_644),
.A3(n_699),
.B(n_706),
.Y(n_790)
);

OAI221xp5_ASAP7_75t_L g791 ( 
.A1(n_717),
.A2(n_645),
.B1(n_671),
.B2(n_685),
.C(n_675),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_SL g792 ( 
.A1(n_742),
.A2(n_719),
.B(n_722),
.Y(n_792)
);

INVxp67_ASAP7_75t_SL g793 ( 
.A(n_722),
.Y(n_793)
);

HB1xp67_ASAP7_75t_SL g794 ( 
.A(n_739),
.Y(n_794)
);

BUFx2_ASAP7_75t_L g795 ( 
.A(n_757),
.Y(n_795)
);

AO31x2_ASAP7_75t_L g796 ( 
.A1(n_773),
.A2(n_698),
.A3(n_715),
.B(n_639),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_752),
.Y(n_797)
);

OAI21xp5_ASAP7_75t_SL g798 ( 
.A1(n_724),
.A2(n_691),
.B(n_690),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_757),
.B(n_710),
.Y(n_799)
);

NOR2xp67_ASAP7_75t_L g800 ( 
.A(n_746),
.B(n_679),
.Y(n_800)
);

OAI21x1_ASAP7_75t_L g801 ( 
.A1(n_737),
.A2(n_681),
.B(n_661),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_746),
.B(n_711),
.Y(n_802)
);

A2O1A1Ixp33_ASAP7_75t_L g803 ( 
.A1(n_725),
.A2(n_716),
.B(n_633),
.C(n_656),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_767),
.B(n_648),
.Y(n_804)
);

OAI21x1_ASAP7_75t_L g805 ( 
.A1(n_749),
.A2(n_681),
.B(n_661),
.Y(n_805)
);

CKINVDCx8_ASAP7_75t_R g806 ( 
.A(n_729),
.Y(n_806)
);

NOR2xp67_ASAP7_75t_L g807 ( 
.A(n_765),
.B(n_679),
.Y(n_807)
);

O2A1O1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_764),
.A2(n_693),
.B(n_672),
.C(n_701),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_772),
.A2(n_651),
.B(n_650),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_729),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_759),
.B(n_670),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_770),
.B(n_659),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_726),
.B(n_682),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_729),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_741),
.B(n_771),
.Y(n_815)
);

BUFx2_ASAP7_75t_L g816 ( 
.A(n_762),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_758),
.B(n_647),
.Y(n_817)
);

OAI21x1_ASAP7_75t_L g818 ( 
.A1(n_720),
.A2(n_689),
.B(n_683),
.Y(n_818)
);

AND2x6_ASAP7_75t_L g819 ( 
.A(n_772),
.B(n_673),
.Y(n_819)
);

OAI21x1_ASAP7_75t_L g820 ( 
.A1(n_732),
.A2(n_683),
.B(n_703),
.Y(n_820)
);

OAI21x1_ASAP7_75t_L g821 ( 
.A1(n_740),
.A2(n_738),
.B(n_773),
.Y(n_821)
);

AOI221xp5_ASAP7_75t_L g822 ( 
.A1(n_750),
.A2(n_703),
.B1(n_647),
.B2(n_389),
.C(n_659),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_751),
.A2(n_679),
.B(n_712),
.Y(n_823)
);

OAI22x1_ASAP7_75t_L g824 ( 
.A1(n_747),
.A2(n_660),
.B1(n_221),
.B2(n_249),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_727),
.Y(n_825)
);

AO21x2_ASAP7_75t_L g826 ( 
.A1(n_740),
.A2(n_673),
.B(n_660),
.Y(n_826)
);

A2O1A1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_776),
.A2(n_712),
.B(n_673),
.C(n_270),
.Y(n_827)
);

A2O1A1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_730),
.A2(n_712),
.B(n_270),
.C(n_284),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_768),
.A2(n_288),
.B1(n_280),
.B2(n_274),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_756),
.B(n_745),
.Y(n_830)
);

AOI221x1_ASAP7_75t_L g831 ( 
.A1(n_735),
.A2(n_220),
.B1(n_14),
.B2(n_15),
.C(n_16),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_736),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_755),
.B(n_58),
.Y(n_833)
);

OAI21x1_ASAP7_75t_SL g834 ( 
.A1(n_760),
.A2(n_7),
.B(n_18),
.Y(n_834)
);

INVx6_ASAP7_75t_L g835 ( 
.A(n_810),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_793),
.B(n_754),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_815),
.A2(n_779),
.B1(n_731),
.B2(n_718),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_786),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_815),
.A2(n_753),
.B1(n_748),
.B2(n_735),
.Y(n_839)
);

INVx3_ASAP7_75t_SL g840 ( 
.A(n_794),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_793),
.Y(n_841)
);

OAI22xp33_ASAP7_75t_L g842 ( 
.A1(n_781),
.A2(n_733),
.B1(n_769),
.B2(n_778),
.Y(n_842)
);

BUFx2_ASAP7_75t_L g843 ( 
.A(n_826),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_783),
.A2(n_733),
.B1(n_748),
.B2(n_743),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_804),
.B(n_19),
.Y(n_845)
);

BUFx2_ASAP7_75t_L g846 ( 
.A(n_826),
.Y(n_846)
);

CKINVDCx11_ASAP7_75t_R g847 ( 
.A(n_806),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_819),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_821),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_821),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_812),
.A2(n_220),
.B1(n_754),
.B2(n_775),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_816),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_805),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_801),
.Y(n_854)
);

BUFx3_ASAP7_75t_L g855 ( 
.A(n_810),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_796),
.Y(n_856)
);

CKINVDCx11_ASAP7_75t_R g857 ( 
.A(n_810),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_SL g858 ( 
.A1(n_799),
.A2(n_754),
.B1(n_777),
.B2(n_220),
.Y(n_858)
);

AND2x4_ASAP7_75t_L g859 ( 
.A(n_814),
.B(n_59),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_822),
.A2(n_220),
.B1(n_777),
.B2(n_264),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_SL g861 ( 
.A1(n_833),
.A2(n_777),
.B1(n_272),
.B2(n_262),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_790),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_796),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_792),
.A2(n_258),
.B1(n_255),
.B2(n_245),
.Y(n_864)
);

OAI22xp33_ASAP7_75t_SL g865 ( 
.A1(n_788),
.A2(n_244),
.B1(n_242),
.B2(n_241),
.Y(n_865)
);

BUFx4_ASAP7_75t_SL g866 ( 
.A(n_814),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_810),
.Y(n_867)
);

INVx4_ASAP7_75t_L g868 ( 
.A(n_819),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_825),
.A2(n_240),
.B1(n_234),
.B2(n_231),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_L g870 ( 
.A1(n_802),
.A2(n_225),
.B1(n_224),
.B2(n_223),
.Y(n_870)
);

BUFx2_ASAP7_75t_L g871 ( 
.A(n_819),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_796),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_796),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_791),
.A2(n_222),
.B1(n_21),
.B2(n_22),
.Y(n_874)
);

INVx5_ASAP7_75t_L g875 ( 
.A(n_819),
.Y(n_875)
);

OAI22xp5_ASAP7_75t_L g876 ( 
.A1(n_830),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_818),
.Y(n_877)
);

AOI22xp5_ASAP7_75t_SL g878 ( 
.A1(n_819),
.A2(n_23),
.B1(n_26),
.B2(n_27),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_818),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_790),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_825),
.A2(n_23),
.B1(n_26),
.B2(n_28),
.Y(n_881)
);

BUFx3_ASAP7_75t_L g882 ( 
.A(n_802),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_830),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_883)
);

INVx6_ASAP7_75t_L g884 ( 
.A(n_833),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_832),
.A2(n_782),
.B1(n_824),
.B2(n_813),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_809),
.A2(n_29),
.B(n_30),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_832),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_790),
.Y(n_888)
);

BUFx2_ASAP7_75t_L g889 ( 
.A(n_790),
.Y(n_889)
);

INVx4_ASAP7_75t_L g890 ( 
.A(n_833),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_787),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_785),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_892)
);

HB1xp67_ASAP7_75t_L g893 ( 
.A(n_849),
.Y(n_893)
);

HB1xp67_ASAP7_75t_L g894 ( 
.A(n_849),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_862),
.Y(n_895)
);

OAI21x1_ASAP7_75t_L g896 ( 
.A1(n_856),
.A2(n_787),
.B(n_784),
.Y(n_896)
);

OAI21x1_ASAP7_75t_L g897 ( 
.A1(n_856),
.A2(n_820),
.B(n_808),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_862),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_863),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_891),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_880),
.Y(n_901)
);

OA21x2_ASAP7_75t_L g902 ( 
.A1(n_863),
.A2(n_803),
.B(n_831),
.Y(n_902)
);

HB1xp67_ASAP7_75t_L g903 ( 
.A(n_850),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_872),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_874),
.A2(n_789),
.B1(n_797),
.B2(n_811),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_880),
.Y(n_906)
);

OAI21x1_ASAP7_75t_L g907 ( 
.A1(n_872),
.A2(n_823),
.B(n_834),
.Y(n_907)
);

BUFx4f_ASAP7_75t_SL g908 ( 
.A(n_840),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_841),
.Y(n_909)
);

HB1xp67_ASAP7_75t_L g910 ( 
.A(n_850),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_872),
.Y(n_911)
);

HB1xp67_ASAP7_75t_L g912 ( 
.A(n_841),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_889),
.B(n_803),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_891),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_873),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_873),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_873),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_888),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_888),
.Y(n_919)
);

AO21x2_ASAP7_75t_L g920 ( 
.A1(n_891),
.A2(n_827),
.B(n_798),
.Y(n_920)
);

OR2x6_ASAP7_75t_L g921 ( 
.A(n_868),
.B(n_827),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_854),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_889),
.B(n_36),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_882),
.B(n_836),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_888),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_854),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_836),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_853),
.Y(n_928)
);

BUFx2_ASAP7_75t_L g929 ( 
.A(n_877),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_927),
.B(n_843),
.Y(n_930)
);

NAND3xp33_ASAP7_75t_L g931 ( 
.A(n_905),
.B(n_878),
.C(n_876),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_912),
.B(n_882),
.Y(n_932)
);

OAI21x1_ASAP7_75t_L g933 ( 
.A1(n_897),
.A2(n_879),
.B(n_877),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_927),
.B(n_924),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_905),
.A2(n_884),
.B1(n_883),
.B2(n_861),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_924),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_927),
.B(n_913),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_923),
.A2(n_878),
.B(n_837),
.C(n_870),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_909),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_899),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_908),
.B(n_840),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_913),
.B(n_843),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_913),
.B(n_875),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_908),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_912),
.B(n_882),
.Y(n_945)
);

AND3x1_ASAP7_75t_L g946 ( 
.A(n_923),
.B(n_838),
.C(n_845),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_923),
.B(n_846),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_909),
.B(n_846),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_909),
.B(n_853),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_902),
.A2(n_886),
.B(n_858),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_895),
.B(n_852),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_921),
.B(n_875),
.Y(n_952)
);

AOI221xp5_ASAP7_75t_L g953 ( 
.A1(n_895),
.A2(n_865),
.B1(n_892),
.B2(n_887),
.C(n_881),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_895),
.B(n_852),
.Y(n_954)
);

AOI22xp5_ASAP7_75t_L g955 ( 
.A1(n_920),
.A2(n_884),
.B1(n_890),
.B2(n_839),
.Y(n_955)
);

OAI21x1_ASAP7_75t_SL g956 ( 
.A1(n_902),
.A2(n_890),
.B(n_868),
.Y(n_956)
);

OR2x2_ASAP7_75t_L g957 ( 
.A(n_898),
.B(n_901),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_921),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_899),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_929),
.B(n_853),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_898),
.B(n_852),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_900),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_921),
.Y(n_963)
);

OR2x2_ASAP7_75t_L g964 ( 
.A(n_898),
.B(n_877),
.Y(n_964)
);

AND2x2_ASAP7_75t_SL g965 ( 
.A(n_902),
.B(n_890),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_901),
.B(n_871),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_926),
.B(n_840),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_929),
.B(n_879),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_901),
.Y(n_969)
);

INVx2_ASAP7_75t_SL g970 ( 
.A(n_962),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_952),
.B(n_962),
.Y(n_971)
);

OR2x6_ASAP7_75t_L g972 ( 
.A(n_952),
.B(n_921),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_937),
.B(n_929),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_969),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_937),
.B(n_900),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_940),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_965),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_934),
.B(n_900),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_962),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_934),
.B(n_900),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_965),
.B(n_900),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_965),
.B(n_968),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_952),
.B(n_900),
.Y(n_983)
);

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_936),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_948),
.B(n_926),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_969),
.Y(n_986)
);

INVx3_ASAP7_75t_L g987 ( 
.A(n_962),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_940),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_948),
.B(n_926),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_968),
.B(n_914),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_960),
.B(n_949),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_957),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_960),
.B(n_914),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_949),
.B(n_914),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_982),
.B(n_947),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_974),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_974),
.Y(n_997)
);

OR2x2_ASAP7_75t_L g998 ( 
.A(n_984),
.B(n_932),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_982),
.B(n_947),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_984),
.B(n_944),
.Y(n_1000)
);

AOI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_977),
.A2(n_931),
.B1(n_946),
.B2(n_938),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_973),
.B(n_932),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_974),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_982),
.B(n_943),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_992),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_986),
.Y(n_1006)
);

OAI211xp5_ASAP7_75t_L g1007 ( 
.A1(n_977),
.A2(n_931),
.B(n_935),
.C(n_967),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_977),
.A2(n_955),
.B(n_935),
.C(n_953),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_976),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_986),
.Y(n_1010)
);

INVx1_ASAP7_75t_SL g1011 ( 
.A(n_985),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_977),
.B(n_981),
.Y(n_1012)
);

OAI22xp33_ASAP7_75t_L g1013 ( 
.A1(n_977),
.A2(n_955),
.B1(n_884),
.B2(n_963),
.Y(n_1013)
);

NOR3xp33_ASAP7_75t_SL g1014 ( 
.A(n_985),
.B(n_941),
.C(n_945),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_976),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_1011),
.B(n_992),
.Y(n_1016)
);

NAND2x1_ASAP7_75t_L g1017 ( 
.A(n_1012),
.B(n_977),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_1009),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_1014),
.B(n_992),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_996),
.Y(n_1020)
);

HB1xp67_ASAP7_75t_L g1021 ( 
.A(n_998),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_998),
.B(n_973),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_1004),
.B(n_995),
.Y(n_1023)
);

INVx1_ASAP7_75t_SL g1024 ( 
.A(n_1000),
.Y(n_1024)
);

OR2x2_ASAP7_75t_L g1025 ( 
.A(n_1005),
.B(n_989),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_996),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_1019),
.B(n_1001),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_1018),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1020),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1026),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_1023),
.B(n_1004),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1021),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_1016),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1032),
.B(n_1001),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_1032),
.B(n_1023),
.Y(n_1035)
);

NAND4xp25_ASAP7_75t_L g1036 ( 
.A(n_1027),
.B(n_1024),
.C(n_1008),
.D(n_1007),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_1031),
.B(n_995),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_1034),
.A2(n_1035),
.B1(n_1037),
.B2(n_1031),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_1036),
.B(n_1033),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1035),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_1034),
.A2(n_946),
.B1(n_977),
.B2(n_1017),
.Y(n_1041)
);

OAI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_1034),
.A2(n_1030),
.B(n_1029),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_1037),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_1034),
.B(n_1030),
.Y(n_1044)
);

NAND4xp75_ASAP7_75t_L g1045 ( 
.A(n_1034),
.B(n_1028),
.C(n_982),
.D(n_950),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_1034),
.B(n_1025),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_1034),
.A2(n_977),
.B1(n_1017),
.B2(n_1012),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_1037),
.B(n_1012),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1044),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1040),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1046),
.Y(n_1051)
);

OR4x1_ASAP7_75t_L g1052 ( 
.A(n_1042),
.B(n_979),
.C(n_970),
.D(n_1006),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_1039),
.B(n_1025),
.Y(n_1053)
);

OAI211xp5_ASAP7_75t_SL g1054 ( 
.A1(n_1038),
.A2(n_1022),
.B(n_1002),
.C(n_997),
.Y(n_1054)
);

OAI32xp33_ASAP7_75t_L g1055 ( 
.A1(n_1041),
.A2(n_1043),
.A3(n_1047),
.B1(n_1045),
.B2(n_1028),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1048),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1048),
.Y(n_1057)
);

INVxp67_ASAP7_75t_L g1058 ( 
.A(n_1039),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_1042),
.B(n_999),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_1043),
.B(n_999),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_1048),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_1042),
.B(n_1012),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1042),
.B(n_997),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_1043),
.B(n_1003),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1050),
.Y(n_1065)
);

AOI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_1058),
.A2(n_977),
.B1(n_1018),
.B2(n_1013),
.Y(n_1066)
);

O2A1O1Ixp5_ASAP7_75t_L g1067 ( 
.A1(n_1055),
.A2(n_1010),
.B(n_1006),
.C(n_1003),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1049),
.Y(n_1068)
);

AOI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_1053),
.A2(n_865),
.B1(n_884),
.B2(n_885),
.Y(n_1069)
);

OAI221xp5_ASAP7_75t_L g1070 ( 
.A1(n_1053),
.A2(n_950),
.B1(n_870),
.B2(n_864),
.C(n_884),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1051),
.Y(n_1071)
);

NAND3x1_ASAP7_75t_L g1072 ( 
.A(n_1061),
.B(n_847),
.C(n_987),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1064),
.Y(n_1073)
);

AOI221xp5_ASAP7_75t_L g1074 ( 
.A1(n_1063),
.A2(n_860),
.B1(n_851),
.B2(n_1010),
.C(n_1015),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1060),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1061),
.B(n_1056),
.Y(n_1076)
);

O2A1O1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_1062),
.A2(n_1054),
.B(n_1059),
.C(n_1057),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1061),
.B(n_986),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1062),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1052),
.B(n_973),
.Y(n_1080)
);

AOI22x1_ASAP7_75t_L g1081 ( 
.A1(n_1052),
.A2(n_970),
.B1(n_979),
.B2(n_987),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1050),
.Y(n_1082)
);

OA21x2_ASAP7_75t_SL g1083 ( 
.A1(n_1062),
.A2(n_971),
.B(n_983),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1076),
.Y(n_1084)
);

NOR3xp33_ASAP7_75t_L g1085 ( 
.A(n_1067),
.B(n_800),
.C(n_857),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_1077),
.A2(n_1015),
.B(n_1009),
.Y(n_1086)
);

OAI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_1079),
.A2(n_981),
.B(n_945),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1075),
.Y(n_1088)
);

NOR2x1p5_ASAP7_75t_SL g1089 ( 
.A(n_1065),
.B(n_957),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_1073),
.B(n_970),
.Y(n_1090)
);

NAND4xp25_ASAP7_75t_L g1091 ( 
.A(n_1083),
.B(n_971),
.C(n_981),
.D(n_987),
.Y(n_1091)
);

AND3x1_ASAP7_75t_L g1092 ( 
.A(n_1071),
.B(n_987),
.C(n_981),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1082),
.A2(n_869),
.B(n_829),
.Y(n_1093)
);

XNOR2xp5_ASAP7_75t_L g1094 ( 
.A(n_1069),
.B(n_795),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_1066),
.A2(n_920),
.B1(n_972),
.B2(n_921),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1068),
.B(n_1078),
.Y(n_1096)
);

NAND4xp25_ASAP7_75t_SL g1097 ( 
.A(n_1080),
.B(n_978),
.C(n_980),
.D(n_989),
.Y(n_1097)
);

AOI322xp5_ASAP7_75t_L g1098 ( 
.A1(n_1078),
.A2(n_942),
.A3(n_973),
.B1(n_991),
.B2(n_930),
.C1(n_975),
.C2(n_980),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_1081),
.B(n_970),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1070),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1084),
.B(n_1074),
.Y(n_1101)
);

AOI211xp5_ASAP7_75t_L g1102 ( 
.A1(n_1088),
.A2(n_1072),
.B(n_859),
.C(n_866),
.Y(n_1102)
);

OAI221xp5_ASAP7_75t_L g1103 ( 
.A1(n_1085),
.A2(n_890),
.B1(n_902),
.B2(n_828),
.C(n_966),
.Y(n_1103)
);

OAI211xp5_ASAP7_75t_SL g1104 ( 
.A1(n_1096),
.A2(n_37),
.B(n_39),
.C(n_40),
.Y(n_1104)
);

A2O1A1O1Ixp25_ASAP7_75t_L g1105 ( 
.A1(n_1086),
.A2(n_39),
.B(n_42),
.C(n_43),
.D(n_44),
.Y(n_1105)
);

AOI222xp33_ASAP7_75t_L g1106 ( 
.A1(n_1089),
.A2(n_942),
.B1(n_988),
.B2(n_976),
.C1(n_842),
.C2(n_828),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_1100),
.A2(n_920),
.B1(n_972),
.B2(n_921),
.Y(n_1107)
);

AOI221xp5_ASAP7_75t_SL g1108 ( 
.A1(n_1090),
.A2(n_987),
.B1(n_980),
.B2(n_978),
.C(n_939),
.Y(n_1108)
);

AOI221xp5_ASAP7_75t_L g1109 ( 
.A1(n_1093),
.A2(n_1092),
.B1(n_1087),
.B2(n_1095),
.C(n_1094),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_1098),
.B(n_978),
.Y(n_1110)
);

AOI211xp5_ASAP7_75t_L g1111 ( 
.A1(n_1097),
.A2(n_859),
.B(n_954),
.C(n_961),
.Y(n_1111)
);

AOI221xp5_ASAP7_75t_L g1112 ( 
.A1(n_1093),
.A2(n_920),
.B1(n_956),
.B2(n_954),
.C(n_961),
.Y(n_1112)
);

NOR2x1_ASAP7_75t_L g1113 ( 
.A(n_1091),
.B(n_859),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_1099),
.A2(n_951),
.B1(n_939),
.B2(n_971),
.Y(n_1114)
);

OAI211xp5_ASAP7_75t_SL g1115 ( 
.A1(n_1084),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_1115)
);

AOI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_1085),
.A2(n_920),
.B1(n_991),
.B2(n_943),
.Y(n_1116)
);

XNOR2x1_ASAP7_75t_L g1117 ( 
.A(n_1094),
.B(n_859),
.Y(n_1117)
);

NAND4xp25_ASAP7_75t_L g1118 ( 
.A(n_1088),
.B(n_971),
.C(n_987),
.D(n_978),
.Y(n_1118)
);

AOI211xp5_ASAP7_75t_L g1119 ( 
.A1(n_1084),
.A2(n_844),
.B(n_975),
.C(n_971),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1096),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1096),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_1084),
.B(n_979),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1084),
.B(n_980),
.Y(n_1123)
);

AOI211xp5_ASAP7_75t_L g1124 ( 
.A1(n_1084),
.A2(n_975),
.B(n_971),
.C(n_48),
.Y(n_1124)
);

AOI322xp5_ASAP7_75t_L g1125 ( 
.A1(n_1101),
.A2(n_991),
.A3(n_930),
.B1(n_975),
.B2(n_958),
.C1(n_993),
.C2(n_966),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1109),
.A2(n_920),
.B1(n_983),
.B2(n_902),
.Y(n_1126)
);

AOI322xp5_ASAP7_75t_L g1127 ( 
.A1(n_1120),
.A2(n_993),
.A3(n_990),
.B1(n_952),
.B2(n_994),
.C1(n_943),
.C2(n_988),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1104),
.Y(n_1128)
);

OAI211xp5_ASAP7_75t_L g1129 ( 
.A1(n_1121),
.A2(n_979),
.B(n_47),
.C(n_48),
.Y(n_1129)
);

AO221x1_ASAP7_75t_L g1130 ( 
.A1(n_1114),
.A2(n_956),
.B1(n_848),
.B2(n_871),
.C(n_51),
.Y(n_1130)
);

AOI221xp5_ASAP7_75t_SL g1131 ( 
.A1(n_1122),
.A2(n_46),
.B1(n_47),
.B2(n_51),
.C(n_993),
.Y(n_1131)
);

OAI22xp33_ASAP7_75t_L g1132 ( 
.A1(n_1105),
.A2(n_921),
.B1(n_902),
.B2(n_972),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1115),
.A2(n_983),
.B(n_922),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_1123),
.B(n_835),
.Y(n_1134)
);

NOR2x1_ASAP7_75t_L g1135 ( 
.A(n_1113),
.B(n_1118),
.Y(n_1135)
);

AND4x1_ASAP7_75t_L g1136 ( 
.A(n_1124),
.B(n_1102),
.C(n_1119),
.D(n_1106),
.Y(n_1136)
);

NAND3xp33_ASAP7_75t_L g1137 ( 
.A(n_1103),
.B(n_855),
.C(n_867),
.Y(n_1137)
);

AOI211xp5_ASAP7_75t_SL g1138 ( 
.A1(n_1111),
.A2(n_922),
.B(n_910),
.C(n_903),
.Y(n_1138)
);

AOI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1116),
.A2(n_983),
.B1(n_902),
.B2(n_943),
.Y(n_1139)
);

O2A1O1Ixp5_ASAP7_75t_L g1140 ( 
.A1(n_1110),
.A2(n_983),
.B(n_988),
.C(n_976),
.Y(n_1140)
);

AOI221xp5_ASAP7_75t_L g1141 ( 
.A1(n_1112),
.A2(n_988),
.B1(n_993),
.B2(n_817),
.C(n_990),
.Y(n_1141)
);

OAI321xp33_ASAP7_75t_L g1142 ( 
.A1(n_1107),
.A2(n_972),
.A3(n_921),
.B1(n_867),
.B2(n_906),
.C(n_964),
.Y(n_1142)
);

AOI21xp33_ASAP7_75t_SL g1143 ( 
.A1(n_1117),
.A2(n_983),
.B(n_61),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1108),
.B(n_990),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1120),
.B(n_994),
.Y(n_1145)
);

OAI211xp5_ASAP7_75t_SL g1146 ( 
.A1(n_1120),
.A2(n_848),
.B(n_903),
.C(n_894),
.Y(n_1146)
);

AOI221xp5_ASAP7_75t_L g1147 ( 
.A1(n_1101),
.A2(n_994),
.B1(n_910),
.B2(n_893),
.C(n_894),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_R g1148 ( 
.A(n_1120),
.B(n_60),
.Y(n_1148)
);

INVxp67_ASAP7_75t_L g1149 ( 
.A(n_1128),
.Y(n_1149)
);

NOR2x1_ASAP7_75t_L g1150 ( 
.A(n_1129),
.B(n_855),
.Y(n_1150)
);

OR2x2_ASAP7_75t_L g1151 ( 
.A(n_1145),
.B(n_893),
.Y(n_1151)
);

XNOR2x1_ASAP7_75t_L g1152 ( 
.A(n_1135),
.B(n_807),
.Y(n_1152)
);

OR2x2_ASAP7_75t_L g1153 ( 
.A(n_1144),
.B(n_964),
.Y(n_1153)
);

NAND4xp75_ASAP7_75t_L g1154 ( 
.A(n_1131),
.B(n_906),
.C(n_928),
.D(n_879),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1130),
.B(n_972),
.Y(n_1155)
);

NOR2x1_ASAP7_75t_L g1156 ( 
.A(n_1134),
.B(n_855),
.Y(n_1156)
);

NOR2x1_ASAP7_75t_L g1157 ( 
.A(n_1132),
.B(n_868),
.Y(n_1157)
);

NOR3xp33_ASAP7_75t_L g1158 ( 
.A(n_1143),
.B(n_868),
.C(n_848),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1136),
.Y(n_1159)
);

NOR3xp33_ASAP7_75t_SL g1160 ( 
.A(n_1146),
.B(n_66),
.C(n_68),
.Y(n_1160)
);

OAI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_1139),
.A2(n_972),
.B1(n_875),
.B2(n_835),
.Y(n_1161)
);

INVx2_ASAP7_75t_SL g1162 ( 
.A(n_1148),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1126),
.Y(n_1163)
);

AOI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1137),
.A2(n_1141),
.B1(n_1147),
.B2(n_1133),
.Y(n_1164)
);

INVxp67_ASAP7_75t_L g1165 ( 
.A(n_1138),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_1142),
.B(n_835),
.Y(n_1166)
);

XNOR2xp5_ASAP7_75t_L g1167 ( 
.A(n_1140),
.B(n_972),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1125),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1127),
.Y(n_1169)
);

OR2x2_ASAP7_75t_L g1170 ( 
.A(n_1129),
.B(n_914),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1159),
.A2(n_972),
.B(n_897),
.Y(n_1171)
);

OR3x2_ASAP7_75t_L g1172 ( 
.A(n_1169),
.B(n_906),
.C(n_72),
.Y(n_1172)
);

NAND3xp33_ASAP7_75t_L g1173 ( 
.A(n_1149),
.B(n_875),
.C(n_848),
.Y(n_1173)
);

AND3x2_ASAP7_75t_L g1174 ( 
.A(n_1165),
.B(n_70),
.C(n_73),
.Y(n_1174)
);

NAND3x1_ASAP7_75t_L g1175 ( 
.A(n_1150),
.B(n_914),
.C(n_835),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1168),
.B(n_835),
.Y(n_1176)
);

NOR2x1_ASAP7_75t_L g1177 ( 
.A(n_1154),
.B(n_75),
.Y(n_1177)
);

OR2x2_ASAP7_75t_L g1178 ( 
.A(n_1170),
.B(n_914),
.Y(n_1178)
);

AOI221xp5_ASAP7_75t_L g1179 ( 
.A1(n_1162),
.A2(n_1163),
.B1(n_1155),
.B2(n_1164),
.C(n_1166),
.Y(n_1179)
);

NAND3xp33_ASAP7_75t_SL g1180 ( 
.A(n_1158),
.B(n_928),
.C(n_959),
.Y(n_1180)
);

AOI222xp33_ASAP7_75t_L g1181 ( 
.A1(n_1163),
.A2(n_928),
.B1(n_915),
.B2(n_917),
.C1(n_907),
.C2(n_959),
.Y(n_1181)
);

A2O1A1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1160),
.A2(n_907),
.B(n_897),
.C(n_933),
.Y(n_1182)
);

NOR3xp33_ASAP7_75t_L g1183 ( 
.A(n_1156),
.B(n_907),
.C(n_77),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_L g1184 ( 
.A(n_1152),
.B(n_76),
.Y(n_1184)
);

NOR2x1_ASAP7_75t_L g1185 ( 
.A(n_1151),
.B(n_82),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1185),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_1172),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1178),
.A2(n_1153),
.B1(n_1157),
.B2(n_1167),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1174),
.B(n_1161),
.Y(n_1189)
);

INVx3_ASAP7_75t_L g1190 ( 
.A(n_1175),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_SL g1191 ( 
.A(n_1176),
.B(n_875),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_SL g1192 ( 
.A1(n_1184),
.A2(n_875),
.B1(n_940),
.B2(n_959),
.Y(n_1192)
);

INVx1_ASAP7_75t_SL g1193 ( 
.A(n_1177),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_1179),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1182),
.Y(n_1195)
);

XNOR2xp5_ASAP7_75t_L g1196 ( 
.A(n_1183),
.B(n_84),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1173),
.A2(n_915),
.B1(n_917),
.B2(n_919),
.Y(n_1197)
);

AOI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1180),
.A2(n_907),
.B1(n_897),
.B2(n_933),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1181),
.Y(n_1199)
);

AO22x1_ASAP7_75t_L g1200 ( 
.A1(n_1171),
.A2(n_87),
.B1(n_89),
.B2(n_95),
.Y(n_1200)
);

AOI211xp5_ASAP7_75t_SL g1201 ( 
.A1(n_1194),
.A2(n_97),
.B(n_98),
.C(n_105),
.Y(n_1201)
);

AO22x2_ASAP7_75t_L g1202 ( 
.A1(n_1193),
.A2(n_917),
.B1(n_915),
.B2(n_918),
.Y(n_1202)
);

AO22x2_ASAP7_75t_L g1203 ( 
.A1(n_1186),
.A2(n_925),
.B1(n_919),
.B2(n_918),
.Y(n_1203)
);

AOI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1188),
.A2(n_925),
.B1(n_919),
.B2(n_918),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1187),
.Y(n_1205)
);

OAI22x1_ASAP7_75t_L g1206 ( 
.A1(n_1195),
.A2(n_925),
.B1(n_916),
.B2(n_911),
.Y(n_1206)
);

AO22x2_ASAP7_75t_L g1207 ( 
.A1(n_1199),
.A2(n_1190),
.B1(n_1189),
.B2(n_1197),
.Y(n_1207)
);

OAI22x1_ASAP7_75t_L g1208 ( 
.A1(n_1190),
.A2(n_916),
.B1(n_911),
.B2(n_904),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_1198),
.B(n_896),
.Y(n_1209)
);

BUFx4f_ASAP7_75t_SL g1210 ( 
.A(n_1196),
.Y(n_1210)
);

NAND3xp33_ASAP7_75t_L g1211 ( 
.A(n_1205),
.B(n_1200),
.C(n_1191),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1207),
.Y(n_1212)
);

AOI21xp33_ASAP7_75t_L g1213 ( 
.A1(n_1204),
.A2(n_1192),
.B(n_109),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1210),
.B(n_108),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_SL g1215 ( 
.A1(n_1201),
.A2(n_1209),
.B1(n_1206),
.B2(n_1208),
.Y(n_1215)
);

XNOR2xp5_ASAP7_75t_L g1216 ( 
.A(n_1202),
.B(n_111),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1212),
.B(n_1203),
.Y(n_1217)
);

OAI22x1_ASAP7_75t_L g1218 ( 
.A1(n_1211),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1214),
.B(n_896),
.Y(n_1219)
);

HB1xp67_ASAP7_75t_L g1220 ( 
.A(n_1216),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1217),
.A2(n_1220),
.B1(n_1215),
.B2(n_1219),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_SL g1222 ( 
.A1(n_1221),
.A2(n_1218),
.B1(n_1213),
.B2(n_128),
.Y(n_1222)
);

AOI21xp33_ASAP7_75t_L g1223 ( 
.A1(n_1222),
.A2(n_118),
.B(n_125),
.Y(n_1223)
);

XNOR2x1_ASAP7_75t_L g1224 ( 
.A(n_1223),
.B(n_129),
.Y(n_1224)
);

AOI221xp5_ASAP7_75t_L g1225 ( 
.A1(n_1224),
.A2(n_130),
.B1(n_133),
.B2(n_134),
.C(n_140),
.Y(n_1225)
);

AOI211xp5_ASAP7_75t_L g1226 ( 
.A1(n_1225),
.A2(n_143),
.B(n_147),
.C(n_151),
.Y(n_1226)
);


endmodule