module fake_jpeg_24423_n_49 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_49);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_49;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx16f_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx8_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx2_ASAP7_75t_SL g13 ( 
.A(n_3),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_2),
.B(n_1),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_9),
.B(n_0),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_17),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_L g16 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_18),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g17 ( 
.A1(n_9),
.A2(n_11),
.B1(n_10),
.B2(n_14),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_11),
.B(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx6p67_ASAP7_75t_R g27 ( 
.A(n_19),
.Y(n_27)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_7),
.Y(n_21)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_20),
.Y(n_28)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_31),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_21),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_23),
.A2(n_16),
.B1(n_19),
.B2(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_32),
.B(n_27),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_34),
.B1(n_22),
.B2(n_27),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_31),
.C(n_29),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_39),
.C(n_40),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_22),
.Y(n_38)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

OAI31xp33_ASAP7_75t_L g40 ( 
.A1(n_35),
.A2(n_31),
.A3(n_25),
.B(n_27),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_25),
.C(n_26),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_25),
.C(n_12),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_45),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_41),
.A2(n_12),
.B1(n_6),
.B2(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_43),
.C(n_7),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_6),
.Y(n_49)
);


endmodule