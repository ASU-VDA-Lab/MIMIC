module fake_jpeg_30988_n_273 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_273);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_273;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx2_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_33),
.B(n_0),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_47),
.B(n_62),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_21),
.B(n_15),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_60),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_33),
.Y(n_57)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_33),
.A2(n_34),
.B1(n_38),
.B2(n_20),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_66),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_0),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_34),
.Y(n_72)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_65),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_35),
.B1(n_39),
.B2(n_38),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_71),
.A2(n_83),
.B1(n_64),
.B2(n_46),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_66),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_58),
.A2(n_39),
.B1(n_30),
.B2(n_25),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_76),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_57),
.A2(n_34),
.B1(n_36),
.B2(n_27),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_81),
.A2(n_89),
.B1(n_90),
.B2(n_95),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_55),
.A2(n_35),
.B1(n_39),
.B2(n_20),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_30),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_3),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_40),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_86),
.B(n_92),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_44),
.B(n_40),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_88),
.B(n_14),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_57),
.A2(n_36),
.B1(n_35),
.B2(n_19),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_41),
.A2(n_36),
.B1(n_32),
.B2(n_31),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_47),
.B(n_21),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_42),
.A2(n_32),
.B1(n_31),
.B2(n_29),
.Y(n_95)
);

OR2x4_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_29),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_85),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_56),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_100),
.A2(n_104),
.B1(n_43),
.B2(n_45),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_51),
.B(n_18),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_9),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_59),
.A2(n_26),
.B1(n_24),
.B2(n_18),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_108),
.B(n_131),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_109),
.A2(n_79),
.B1(n_99),
.B2(n_67),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_110),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_111),
.B(n_112),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_52),
.C(n_54),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_85),
.A2(n_49),
.B1(n_23),
.B2(n_50),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_113),
.A2(n_121),
.B1(n_77),
.B2(n_79),
.Y(n_148)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_114),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_97),
.A2(n_63),
.B1(n_53),
.B2(n_65),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_82),
.B1(n_75),
.B2(n_94),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_87),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_117),
.Y(n_156)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_118),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_119),
.B(n_125),
.Y(n_158)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

INVxp67_ASAP7_75t_SL g141 ( 
.A(n_123),
.Y(n_141)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_74),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_130),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_77),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_84),
.B(n_4),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_127),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_8),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_8),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_134),
.Y(n_164)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_74),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_133),
.Y(n_144)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_136),
.Y(n_145)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_106),
.A2(n_82),
.B1(n_107),
.B2(n_105),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_137),
.A2(n_142),
.B1(n_155),
.B2(n_96),
.Y(n_186)
);

XNOR2x1_ASAP7_75t_SL g143 ( 
.A(n_127),
.B(n_68),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_131),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_75),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_146),
.B(n_150),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_108),
.A2(n_91),
.B(n_67),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_147),
.A2(n_123),
.B(n_120),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_148),
.A2(n_111),
.B1(n_78),
.B2(n_130),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_91),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_135),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_118),
.A2(n_99),
.B1(n_103),
.B2(n_73),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_111),
.A2(n_78),
.B1(n_73),
.B2(n_103),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_163),
.A2(n_128),
.B1(n_121),
.B2(n_112),
.Y(n_171)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_138),
.B(n_126),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_168),
.B(n_173),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_169),
.Y(n_191)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_170),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_171),
.B(n_176),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_158),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_177),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_138),
.B(n_129),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_124),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_187),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_164),
.B(n_134),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_143),
.B(n_10),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_154),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_178),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_159),
.B(n_10),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_179),
.B(n_184),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_180),
.Y(n_206)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

HAxp5_ASAP7_75t_SL g194 ( 
.A(n_181),
.B(n_183),
.CON(n_194),
.SN(n_194)
);

AOI221xp5_ASAP7_75t_L g192 ( 
.A1(n_182),
.A2(n_185),
.B1(n_186),
.B2(n_148),
.C(n_156),
.Y(n_192)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_156),
.A2(n_114),
.B1(n_136),
.B2(n_122),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_151),
.A2(n_96),
.B1(n_11),
.B2(n_12),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_151),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_13),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_159),
.A2(n_11),
.B(n_12),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_189),
.A2(n_157),
.B(n_145),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_192),
.A2(n_161),
.B1(n_181),
.B2(n_162),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_159),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_204),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_203),
.A2(n_168),
.B1(n_179),
.B2(n_187),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_157),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_152),
.C(n_147),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_209),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_208),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_152),
.C(n_162),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_195),
.Y(n_210)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_210),
.Y(n_231)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_195),
.Y(n_211)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_211),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_166),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_216),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_213),
.A2(n_215),
.B1(n_223),
.B2(n_224),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_193),
.A2(n_165),
.B1(n_169),
.B2(n_177),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_198),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_152),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_191),
.C(n_204),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_193),
.A2(n_171),
.B1(n_169),
.B2(n_183),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_222),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_190),
.A2(n_167),
.B1(n_184),
.B2(n_170),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_201),
.B(n_174),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_194),
.A2(n_185),
.B(n_153),
.Y(n_223)
);

OAI22x1_ASAP7_75t_L g224 ( 
.A1(n_191),
.A2(n_142),
.B1(n_163),
.B2(n_141),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_225),
.A2(n_224),
.B1(n_223),
.B2(n_221),
.Y(n_234)
);

XNOR2x1_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_190),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_229),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_209),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_235),
.C(n_238),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_237),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_202),
.C(n_200),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_226),
.B(n_198),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_208),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_230),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_242),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_232),
.C(n_235),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_227),
.C(n_197),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_201),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_233),
.A2(n_225),
.B1(n_221),
.B2(n_218),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_243),
.A2(n_247),
.B1(n_199),
.B2(n_206),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_236),
.A2(n_208),
.B(n_202),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_246),
.A2(n_228),
.B(n_200),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_238),
.A2(n_222),
.B1(n_211),
.B2(n_199),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_219),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_203),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_252),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_196),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_255),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_254),
.C(n_244),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_162),
.Y(n_254)
);

OAI221xp5_ASAP7_75t_L g256 ( 
.A1(n_253),
.A2(n_243),
.B1(n_240),
.B2(n_241),
.C(n_245),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_256),
.B(n_261),
.Y(n_264)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_250),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_261),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_254),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_251),
.A2(n_244),
.B1(n_180),
.B2(n_178),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_263),
.A2(n_264),
.B(n_265),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_260),
.B(n_160),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_262),
.A2(n_259),
.B(n_258),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_268),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_263),
.A2(n_258),
.B(n_161),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_266),
.A2(n_149),
.B(n_160),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_149),
.C(n_180),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_270),
.C(n_13),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_272),
.A2(n_14),
.B(n_230),
.Y(n_273)
);


endmodule