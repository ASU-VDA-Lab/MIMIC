module fake_jpeg_20320_n_142 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_142);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_142;

wire n_117;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx2_ASAP7_75t_SL g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_21),
.Y(n_30)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_9),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_24),
.Y(n_29)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

OR2x4_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_11),
.Y(n_34)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_27),
.A2(n_11),
.B1(n_13),
.B2(n_12),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_23),
.A2(n_18),
.B1(n_11),
.B2(n_17),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_31),
.A2(n_17),
.B1(n_12),
.B2(n_14),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_22),
.Y(n_41)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_41),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_34),
.A2(n_22),
.B1(n_11),
.B2(n_24),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_45),
.B1(n_33),
.B2(n_27),
.Y(n_48)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_18),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_44),
.B(n_46),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_29),
.A2(n_27),
.B1(n_20),
.B2(n_21),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_26),
.B(n_14),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_48),
.A2(n_55),
.B1(n_45),
.B2(n_58),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_52),
.B(n_57),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_36),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_53),
.B(n_56),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_25),
.B1(n_16),
.B2(n_14),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_17),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_40),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_59),
.B(n_63),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_61),
.A2(n_67),
.B(n_48),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_62),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_47),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_50),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_61),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g67 ( 
.A(n_57),
.B(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_80),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_67),
.A2(n_58),
.B1(n_50),
.B2(n_56),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_73),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_49),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_75),
.B(n_76),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_51),
.Y(n_76)
);

MAJx2_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_82),
.C(n_16),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_48),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_78),
.B(n_12),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_79),
.A2(n_60),
.B1(n_25),
.B2(n_19),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_54),
.B(n_51),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_37),
.B1(n_35),
.B2(n_10),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_81),
.A2(n_16),
.B1(n_1),
.B2(n_2),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_66),
.A2(n_12),
.B(n_13),
.Y(n_82)
);

OAI322xp33_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_68),
.A3(n_69),
.B1(n_10),
.B2(n_19),
.C1(n_14),
.C2(n_13),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_83),
.B(n_96),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_79),
.A2(n_60),
.B1(n_10),
.B2(n_19),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_84),
.A2(n_92),
.B1(n_80),
.B2(n_72),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_87),
.Y(n_99)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_78),
.A2(n_19),
.B1(n_10),
.B2(n_13),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_90),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_15),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_91),
.Y(n_104)
);

AOI221xp5_ASAP7_75t_SL g93 ( 
.A1(n_71),
.A2(n_77),
.B1(n_73),
.B2(n_74),
.C(n_81),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_95),
.Y(n_105)
);

NOR3xp33_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_9),
.C(n_8),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_101),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_88),
.A2(n_8),
.B1(n_7),
.B2(n_6),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_98),
.A2(n_87),
.B(n_89),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_16),
.B1(n_8),
.B2(n_6),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g102 ( 
.A1(n_94),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_102),
.A2(n_90),
.B(n_92),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_6),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_107),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_0),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_108),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_111),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_96),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_106),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_105),
.A2(n_86),
.B(n_1),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_114),
.A2(n_3),
.B(n_4),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_0),
.C(n_1),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_115),
.B(n_98),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_0),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_116),
.A2(n_102),
.B(n_100),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_119),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_3),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_104),
.C(n_107),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_123),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_122),
.A2(n_108),
.B(n_116),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_127),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_120),
.A2(n_112),
.B(n_113),
.Y(n_126)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_5),
.C(n_118),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_5),
.C(n_127),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_125),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_128),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_131),
.Y(n_136)
);

INVxp33_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_133),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_135),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_137),
.A2(n_134),
.B(n_5),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_5),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_136),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_138),
.Y(n_142)
);


endmodule