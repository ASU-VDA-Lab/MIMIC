module fake_jpeg_23163_n_32 (n_3, n_2, n_1, n_0, n_4, n_32);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_32;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_5;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g5 ( 
.A(n_1),
.Y(n_5)
);

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_4),
.B(n_0),
.Y(n_6)
);

INVx3_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

INVx2_ASAP7_75t_R g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx11_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_8),
.B(n_3),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_12),
.B(n_13),
.Y(n_23)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx4_ASAP7_75t_SL g14 ( 
.A(n_5),
.Y(n_14)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_8),
.B(n_11),
.Y(n_15)
);

NAND3xp33_ASAP7_75t_L g19 ( 
.A(n_15),
.B(n_18),
.C(n_14),
.Y(n_19)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

XOR2x1_ASAP7_75t_SL g21 ( 
.A(n_16),
.B(n_17),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_7),
.A2(n_9),
.B1(n_6),
.B2(n_5),
.Y(n_17)
);

OR2x4_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_8),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_19),
.Y(n_26)
);

AND2x6_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_18),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_23),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_23),
.B(n_21),
.Y(n_24)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_25),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_29),
.A2(n_30),
.B(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_20),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);


endmodule