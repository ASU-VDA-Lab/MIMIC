module real_jpeg_23380_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_105;
wire n_40;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_1),
.A2(n_55),
.B1(n_56),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_1),
.A2(n_62),
.B1(n_63),
.B2(n_70),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_1),
.A2(n_26),
.B1(n_29),
.B2(n_70),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_1),
.A2(n_42),
.B1(n_43),
.B2(n_70),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_2),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_41)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_2),
.A2(n_26),
.B1(n_29),
.B2(n_45),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_2),
.A2(n_45),
.B1(n_62),
.B2(n_63),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_4),
.A2(n_62),
.B1(n_63),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_4),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_4),
.A2(n_26),
.B1(n_29),
.B2(n_75),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_4),
.A2(n_55),
.B1(n_56),
.B2(n_75),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_4),
.A2(n_42),
.B1(n_43),
.B2(n_75),
.Y(n_156)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_6),
.A2(n_26),
.B1(n_29),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_6),
.A2(n_35),
.B1(n_42),
.B2(n_43),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_6),
.A2(n_35),
.B1(n_62),
.B2(n_63),
.Y(n_83)
);

INVx8_ASAP7_75t_SL g61 ( 
.A(n_7),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_8),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_8),
.A2(n_30),
.B1(n_42),
.B2(n_43),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_9),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_54)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_9),
.A2(n_57),
.B1(n_62),
.B2(n_63),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_9),
.A2(n_42),
.B1(n_43),
.B2(n_57),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_9),
.A2(n_26),
.B1(n_29),
.B2(n_57),
.Y(n_207)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_10),
.Y(n_79)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_11),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_11),
.B(n_68),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_11),
.B(n_26),
.C(n_39),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_11),
.A2(n_42),
.B1(n_43),
.B2(n_105),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_11),
.B(n_84),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_11),
.A2(n_25),
.B1(n_102),
.B2(n_214),
.Y(n_213)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_13),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_13),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_13),
.A2(n_62),
.B1(n_63),
.B2(n_116),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_13),
.A2(n_42),
.B1(n_43),
.B2(n_116),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_13),
.A2(n_26),
.B1(n_29),
.B2(n_116),
.Y(n_214)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_145),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_144),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_121),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_20),
.B(n_121),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_85),
.C(n_96),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_21),
.A2(n_22),
.B1(n_85),
.B2(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_51),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_23),
.B(n_53),
.C(n_71),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_36),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_24),
.B(n_36),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B(n_31),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_25),
.B(n_34),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_25),
.A2(n_28),
.B1(n_100),
.B2(n_102),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_25),
.A2(n_27),
.B(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_25),
.A2(n_89),
.B(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_25),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_25),
.A2(n_33),
.B1(n_207),
.B2(n_214),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g37 ( 
.A1(n_26),
.A2(n_29),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g179 ( 
.A(n_27),
.Y(n_179)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_27),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_29),
.B(n_216),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_32),
.A2(n_91),
.B(n_205),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B(n_46),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_37),
.A2(n_41),
.B1(n_49),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_37),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_37),
.A2(n_49),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_37),
.A2(n_49),
.B1(n_192),
.B2(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_37),
.B(n_105),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_50)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_42),
.A2(n_43),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

NAND3xp33_ASAP7_75t_L g230 ( 
.A(n_42),
.B(n_63),
.C(n_80),
.Y(n_230)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_43),
.B(n_188),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_43),
.A2(n_79),
.B(n_229),
.C(n_230),
.Y(n_228)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_47),
.B(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_48),
.A2(n_129),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_49),
.A2(n_95),
.B(n_128),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_49),
.A2(n_128),
.B(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_49),
.A2(n_251),
.B(n_252),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_71),
.B2(n_72),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_58),
.B1(n_68),
.B2(n_69),
.Y(n_53)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_54),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_55),
.A2(n_60),
.B1(n_61),
.B2(n_66),
.Y(n_65)
);

NAND3xp33_ASAP7_75t_L g107 ( 
.A(n_55),
.B(n_61),
.C(n_62),
.Y(n_107)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_58),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_58),
.A2(n_68),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_65),
.Y(n_58)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_59),
.A2(n_113),
.B1(n_114),
.B2(n_120),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_60),
.A2(n_63),
.B(n_104),
.C(n_107),
.Y(n_103)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_63),
.B1(n_79),
.B2(n_80),
.Y(n_81)
);

INVx5_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

HAxp5_ASAP7_75t_SL g229 ( 
.A(n_63),
.B(n_105),
.CON(n_229),
.SN(n_229)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_68),
.B(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_69),
.Y(n_135)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_76),
.B(n_82),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_74),
.B(n_84),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_76),
.A2(n_109),
.B(n_111),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_76),
.A2(n_78),
.B1(n_172),
.B2(n_174),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_77),
.B(n_83),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_77),
.A2(n_84),
.B1(n_110),
.B2(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_77),
.A2(n_84),
.B1(n_173),
.B2(n_229),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_78),
.A2(n_139),
.B(n_140),
.Y(n_138)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_85),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_93),
.B2(n_94),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_86),
.B(n_94),
.Y(n_141)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_92),
.Y(n_87)
);

INVxp33_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_91),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_92),
.A2(n_101),
.B(n_179),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_96),
.B(n_265),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_108),
.C(n_112),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_97),
.A2(n_98),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_99),
.B(n_103),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

OAI21xp33_ASAP7_75t_L g160 ( 
.A1(n_104),
.A2(n_105),
.B(n_117),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_105),
.B(n_217),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_108),
.B(n_112),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_113),
.A2(n_135),
.B(n_136),
.Y(n_134)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_114),
.Y(n_161)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_143),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_131),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_127),
.B2(n_130),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_127),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_129),
.B(n_156),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_141),
.B2(n_142),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_138),
.Y(n_133)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_180),
.B(n_262),
.C(n_267),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_165),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_147),
.B(n_165),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_162),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_149),
.B(n_152),
.C(n_162),
.Y(n_263)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_157),
.C(n_159),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_153),
.A2(n_154),
.B1(n_157),
.B2(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_158),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_159),
.B(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.C(n_170),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_166),
.B(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_169),
.B(n_170),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_175),
.C(n_177),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_171),
.B(n_246),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_179),
.A2(n_205),
.B1(n_206),
.B2(n_208),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_261),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_256),
.B(n_260),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_241),
.B(n_255),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_225),
.B(n_240),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_202),
.B(n_224),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_193),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_186),
.B(n_193),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_187),
.A2(n_189),
.B1(n_190),
.B2(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_187),
.Y(n_210)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_200),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_195),
.B(n_198),
.C(n_200),
.Y(n_239)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_199),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_201),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_211),
.B(n_223),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_209),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_209),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_219),
.B(n_222),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_220),
.B(n_221),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_239),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_239),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_234),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_235),
.C(n_238),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_228),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_233),
.Y(n_249)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_231),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_238),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_237),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_242),
.B(n_243),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_247),
.B2(n_248),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_250),
.C(n_253),
.Y(n_259)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_253),
.B2(n_254),
.Y(n_248)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_249),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_250),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_259),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_257),
.B(n_259),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_264),
.Y(n_267)
);


endmodule