module fake_jpeg_28451_n_426 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_426);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_426;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_18),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_42),
.B(n_45),
.Y(n_96)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_17),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_19),
.B(n_16),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_54),
.B(n_55),
.Y(n_128)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_57),
.Y(n_133)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_19),
.B(n_15),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_66),
.B(n_71),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_39),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_35),
.B(n_15),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_32),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_17),
.Y(n_81)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_35),
.B1(n_21),
.B2(n_32),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_89),
.A2(n_126),
.B1(n_136),
.B2(n_22),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_55),
.A2(n_21),
.B1(n_40),
.B2(n_27),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_90),
.A2(n_21),
.B1(n_67),
.B2(n_40),
.Y(n_139)
);

BUFx2_ASAP7_75t_SL g98 ( 
.A(n_42),
.Y(n_98)
);

INVx11_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

AOI21xp33_ASAP7_75t_L g102 ( 
.A1(n_48),
.A2(n_36),
.B(n_31),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_102),
.B(n_36),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_108),
.B(n_111),
.Y(n_172)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_50),
.B(n_31),
.C(n_21),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_112),
.B(n_38),
.C(n_29),
.Y(n_165)
);

INVx6_ASAP7_75t_SL g115 ( 
.A(n_72),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_115),
.Y(n_158)
);

NAND2xp33_ASAP7_75t_SL g118 ( 
.A(n_58),
.B(n_36),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_118),
.B(n_38),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_43),
.Y(n_122)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_74),
.A2(n_82),
.B1(n_77),
.B2(n_56),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_59),
.A2(n_40),
.B1(n_27),
.B2(n_29),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_51),
.Y(n_137)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_137),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_139),
.A2(n_151),
.B1(n_90),
.B2(n_136),
.Y(n_176)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_141),
.Y(n_177)
);

NAND3xp33_ASAP7_75t_L g192 ( 
.A(n_142),
.B(n_148),
.C(n_166),
.Y(n_192)
);

BUFx10_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

INVx6_ASAP7_75t_SL g186 ( 
.A(n_143),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_105),
.B(n_22),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_170),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_134),
.B(n_13),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_150),
.A2(n_173),
.B1(n_125),
.B2(n_127),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_95),
.A2(n_83),
.B1(n_64),
.B2(n_62),
.Y(n_151)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_132),
.A2(n_80),
.B1(n_78),
.B2(n_40),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_155),
.Y(n_175)
);

INVx11_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_132),
.A2(n_40),
.B1(n_27),
.B2(n_67),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_157),
.A2(n_163),
.B1(n_167),
.B2(n_168),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_110),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g182 ( 
.A(n_159),
.Y(n_182)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_88),
.Y(n_160)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_160),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_96),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_162),
.Y(n_178)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_169),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_134),
.B(n_15),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_123),
.Y(n_167)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_107),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_128),
.B(n_38),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_94),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_174),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_125),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_99),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_176),
.A2(n_183),
.B1(n_188),
.B2(n_150),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_L g183 ( 
.A1(n_146),
.A2(n_121),
.B1(n_87),
.B2(n_97),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_142),
.B(n_113),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_193),
.B(n_179),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_96),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_128),
.C(n_152),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_178),
.A2(n_162),
.B1(n_158),
.B2(n_149),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_197),
.A2(n_203),
.B1(n_205),
.B2(n_206),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_180),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_207),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_202),
.Y(n_219)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_200),
.Y(n_226)
);

BUFx4f_ASAP7_75t_SL g201 ( 
.A(n_186),
.Y(n_201)
);

INVxp33_ASAP7_75t_L g220 ( 
.A(n_201),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_179),
.B(n_170),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_172),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_208),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_181),
.A2(n_169),
.B1(n_165),
.B2(n_97),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_176),
.A2(n_158),
.B1(n_171),
.B2(n_153),
.Y(n_206)
);

NOR2x1p5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_143),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_166),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_184),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_209),
.B(n_143),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_211),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_152),
.Y(n_211)
);

MAJx2_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_144),
.C(n_148),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_120),
.Y(n_233)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_213),
.Y(n_227)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_177),
.Y(n_214)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_214),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_175),
.Y(n_215)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_181),
.A2(n_100),
.B1(n_127),
.B2(n_92),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_161),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_186),
.A2(n_119),
.B1(n_168),
.B2(n_135),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_217),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_183),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_229),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_204),
.B(n_13),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_225),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_207),
.B(n_185),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_230),
.A2(n_236),
.B(n_201),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_212),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_208),
.B(n_195),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_237),
.Y(n_259)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_235),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_207),
.A2(n_184),
.B(n_175),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g237 ( 
.A(n_200),
.B(n_144),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_213),
.Y(n_238)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_238),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_224),
.A2(n_203),
.B1(n_206),
.B2(n_199),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_239),
.A2(n_240),
.B1(n_247),
.B2(n_248),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_224),
.A2(n_205),
.B1(n_210),
.B2(n_202),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_211),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_231),
.C(n_233),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_243),
.B(n_242),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_222),
.A2(n_216),
.B1(n_212),
.B2(n_191),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_244),
.A2(n_257),
.B1(n_258),
.B2(n_229),
.Y(n_270)
);

NOR2x1_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_201),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_237),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_218),
.A2(n_191),
.B1(n_189),
.B2(n_159),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_226),
.A2(n_189),
.B1(n_145),
.B2(n_167),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_237),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_255),
.Y(n_264)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_220),
.Y(n_251)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_251),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_252),
.A2(n_253),
.B(n_255),
.Y(n_278)
);

AND2x4_ASAP7_75t_SL g253 ( 
.A(n_230),
.B(n_201),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_230),
.A2(n_164),
.B(n_214),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_227),
.Y(n_256)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_256),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_222),
.A2(n_173),
.B1(n_100),
.B2(n_92),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_226),
.A2(n_187),
.B1(n_190),
.B2(n_177),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_260),
.A2(n_264),
.B(n_268),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_239),
.A2(n_223),
.B1(n_236),
.B2(n_218),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_262),
.A2(n_263),
.B1(n_258),
.B2(n_228),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_241),
.A2(n_223),
.B1(n_236),
.B2(n_235),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_246),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_267),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_219),
.Y(n_266)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_266),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_244),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_245),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_268),
.B(n_277),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_249),
.B(n_225),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_269),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_270),
.A2(n_273),
.B1(n_247),
.B2(n_277),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_219),
.Y(n_271)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_271),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_241),
.A2(n_252),
.B1(n_245),
.B2(n_257),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_256),
.C(n_254),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_218),
.Y(n_276)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_276),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_259),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_278),
.A2(n_253),
.B(n_240),
.Y(n_284)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_254),
.Y(n_279)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_279),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_231),
.Y(n_286)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_282),
.Y(n_305)
);

INVx5_ASAP7_75t_L g283 ( 
.A(n_269),
.Y(n_283)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_283),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_288),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_243),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_285),
.B(n_289),
.C(n_294),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_286),
.B(n_261),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_266),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_287),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_273),
.A2(n_253),
.B1(n_248),
.B2(n_233),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_276),
.B(n_221),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_292),
.B(n_275),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_221),
.Y(n_293)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_293),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_232),
.C(n_253),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_270),
.A2(n_251),
.B1(n_238),
.B2(n_227),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_297),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_261),
.A2(n_251),
.B1(n_232),
.B2(n_228),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_300),
.A2(n_261),
.B1(n_263),
.B2(n_262),
.Y(n_317)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_301),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_260),
.B(n_143),
.Y(n_303)
);

OAI21xp33_ASAP7_75t_L g309 ( 
.A1(n_303),
.A2(n_264),
.B(n_278),
.Y(n_309)
);

INVxp33_ASAP7_75t_L g307 ( 
.A(n_302),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_307),
.B(n_316),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_309),
.B(n_315),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_283),
.B(n_279),
.Y(n_312)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_312),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_286),
.C(n_285),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_313),
.B(n_314),
.C(n_323),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_294),
.B(n_274),
.C(n_280),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_317),
.A2(n_291),
.B1(n_299),
.B2(n_182),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_301),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_318),
.B(n_321),
.Y(n_343)
);

NAND2x1_ASAP7_75t_SL g320 ( 
.A(n_303),
.B(n_278),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_320),
.Y(n_335)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_302),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_284),
.B(n_262),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_324),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_288),
.B(n_275),
.C(n_272),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_282),
.B(n_272),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_299),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_326),
.B(n_327),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_298),
.B(n_190),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_313),
.B(n_297),
.C(n_281),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_330),
.B(n_341),
.C(n_342),
.Y(n_354)
);

FAx1_ASAP7_75t_SL g332 ( 
.A(n_315),
.B(n_281),
.CI(n_295),
.CON(n_332),
.SN(n_332)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_332),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_314),
.B(n_296),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g366 ( 
.A(n_333),
.B(n_340),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_310),
.A2(n_290),
.B(n_295),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_334),
.A2(n_337),
.B(n_312),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_306),
.A2(n_290),
.B(n_291),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_339),
.B(n_320),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_311),
.B(n_164),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_311),
.B(n_187),
.C(n_140),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_323),
.B(n_140),
.C(n_174),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_319),
.A2(n_160),
.B1(n_101),
.B2(n_85),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_344),
.A2(n_325),
.B1(n_305),
.B2(n_182),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_322),
.B(n_141),
.C(n_155),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_345),
.B(n_349),
.C(n_305),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_306),
.B(n_138),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_346),
.B(n_348),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_324),
.B(n_93),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_310),
.B(n_163),
.C(n_106),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_350),
.B(n_353),
.Y(n_378)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_336),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_355),
.B(n_328),
.Y(n_371)
);

OAI321xp33_ASAP7_75t_L g356 ( 
.A1(n_343),
.A2(n_304),
.A3(n_307),
.B1(n_325),
.B2(n_308),
.C(n_317),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_356),
.A2(n_363),
.B1(n_349),
.B2(n_345),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_333),
.B(n_308),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_357),
.B(n_358),
.Y(n_372)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_338),
.Y(n_358)
);

XNOR2x1_ASAP7_75t_L g374 ( 
.A(n_359),
.B(n_147),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_360),
.B(n_361),
.Y(n_380)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_347),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_335),
.A2(n_182),
.B(n_156),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_362),
.A2(n_367),
.B(n_133),
.Y(n_381)
);

OAI321xp33_ASAP7_75t_L g363 ( 
.A1(n_332),
.A2(n_182),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_330),
.A2(n_131),
.B1(n_104),
.B2(n_114),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_364),
.B(n_365),
.Y(n_375)
);

XOR2x2_ASAP7_75t_L g365 ( 
.A(n_328),
.B(n_147),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_329),
.B(n_124),
.C(n_103),
.Y(n_367)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_368),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_351),
.A2(n_342),
.B1(n_341),
.B2(n_329),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_369),
.B(n_370),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_359),
.A2(n_331),
.B1(n_346),
.B2(n_348),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_371),
.B(n_374),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_362),
.A2(n_331),
.B1(n_340),
.B2(n_119),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_373),
.A2(n_354),
.B1(n_366),
.B2(n_116),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_366),
.B(n_22),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_376),
.B(n_377),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_357),
.B(n_352),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_352),
.B(n_29),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_379),
.B(n_381),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_378),
.B(n_367),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_385),
.B(n_389),
.Y(n_400)
);

NAND2xp33_ASAP7_75t_SL g386 ( 
.A(n_371),
.B(n_365),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g399 ( 
.A(n_386),
.B(n_390),
.Y(n_399)
);

XNOR2x1_ASAP7_75t_L g402 ( 
.A(n_387),
.B(n_0),
.Y(n_402)
);

NAND2x1_ASAP7_75t_SL g388 ( 
.A(n_373),
.B(n_354),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_388),
.A2(n_375),
.B(n_2),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_372),
.B(n_23),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_377),
.B(n_23),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_380),
.B(n_91),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_391),
.B(n_0),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_393),
.B(n_379),
.Y(n_394)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_394),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_383),
.B(n_374),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_395),
.B(n_397),
.Y(n_410)
);

OAI21xp33_ASAP7_75t_SL g407 ( 
.A1(n_396),
.A2(n_402),
.B(n_0),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_392),
.B(n_23),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_388),
.A2(n_69),
.B(n_34),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_398),
.A2(n_404),
.B(n_2),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_382),
.B(n_34),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_401),
.B(n_3),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_403),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_391),
.B(n_27),
.C(n_2),
.Y(n_404)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g406 ( 
.A1(n_399),
.A2(n_386),
.B(n_394),
.C(n_392),
.D(n_384),
.Y(n_406)
);

AO21x2_ASAP7_75t_L g417 ( 
.A1(n_406),
.A2(n_407),
.B(n_4),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_408),
.B(n_3),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_411),
.B(n_12),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_400),
.A2(n_403),
.B(n_4),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_412),
.A2(n_12),
.B(n_5),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_413),
.B(n_415),
.C(n_409),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_405),
.B(n_3),
.C(n_4),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_414),
.A2(n_417),
.B(n_410),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_416),
.B(n_5),
.C(n_6),
.Y(n_420)
);

NOR4xp25_ASAP7_75t_L g422 ( 
.A(n_418),
.B(n_419),
.C(n_420),
.D(n_7),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_419),
.A2(n_417),
.B(n_8),
.Y(n_421)
);

A2O1A1O1Ixp25_ASAP7_75t_L g423 ( 
.A1(n_421),
.A2(n_422),
.B(n_8),
.C(n_9),
.D(n_10),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_423),
.B(n_11),
.C(n_8),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_424),
.B(n_10),
.Y(n_425)
);

A2O1A1Ixp33_ASAP7_75t_SL g426 ( 
.A1(n_425),
.A2(n_10),
.B(n_11),
.C(n_419),
.Y(n_426)
);


endmodule