module fake_jpeg_9889_n_248 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_248);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_248;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_22),
.B(n_7),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_39),
.Y(n_46)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_19),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_40),
.B1(n_20),
.B2(n_17),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_25),
.Y(n_58)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_49),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_20),
.B1(n_17),
.B2(n_30),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_47),
.A2(n_52),
.B1(n_55),
.B2(n_56),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_48),
.A2(n_22),
.B1(n_16),
.B2(n_19),
.Y(n_84)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_26),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_62),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_20),
.B1(n_25),
.B2(n_21),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_35),
.A2(n_20),
.B1(n_25),
.B2(n_30),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_33),
.A2(n_25),
.B1(n_30),
.B2(n_16),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_23),
.Y(n_59)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_36),
.A2(n_16),
.B1(n_22),
.B2(n_27),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_60),
.A2(n_66),
.B1(n_24),
.B2(n_31),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_23),
.Y(n_61)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_36),
.B(n_18),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_63),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_41),
.A2(n_23),
.B1(n_18),
.B2(n_21),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

AO22x1_ASAP7_75t_L g68 ( 
.A1(n_64),
.A2(n_42),
.B1(n_32),
.B2(n_26),
.Y(n_68)
);

AO21x1_ASAP7_75t_L g94 ( 
.A1(n_68),
.A2(n_88),
.B(n_49),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_52),
.A2(n_18),
.B1(n_21),
.B2(n_31),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_75),
.A2(n_81),
.B(n_76),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_59),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_78),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_80),
.Y(n_99)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_60),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_85),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_84),
.A2(n_54),
.B1(n_64),
.B2(n_65),
.Y(n_96)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_86),
.A2(n_24),
.B1(n_28),
.B2(n_45),
.Y(n_111)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_64),
.A2(n_42),
.B1(n_32),
.B2(n_38),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_62),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_91),
.Y(n_116)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_90),
.B(n_100),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_46),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_98),
.B1(n_105),
.B2(n_88),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_46),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_104),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_96),
.A2(n_108),
.B1(n_78),
.B2(n_69),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_50),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_86),
.C(n_72),
.Y(n_123)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_85),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_87),
.A2(n_48),
.B1(n_54),
.B2(n_63),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_102),
.A2(n_111),
.B1(n_69),
.B2(n_88),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_82),
.A2(n_54),
.B1(n_65),
.B2(n_27),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_83),
.Y(n_104)
);

AO21x1_ASAP7_75t_SL g105 ( 
.A1(n_84),
.A2(n_56),
.B(n_32),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_83),
.A2(n_65),
.B1(n_44),
.B2(n_57),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_56),
.B1(n_45),
.B2(n_19),
.Y(n_108)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_112),
.B(n_72),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_128),
.Y(n_152)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_114),
.B(n_117),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_115),
.A2(n_122),
.B1(n_109),
.B2(n_105),
.Y(n_146)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_120),
.B(n_121),
.Y(n_143)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_94),
.Y(n_156)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_124),
.B(n_126),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_125),
.A2(n_102),
.B1(n_109),
.B2(n_112),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_95),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_129),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_91),
.B(n_70),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_70),
.C(n_88),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_132),
.C(n_108),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_98),
.B(n_45),
.C(n_68),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_111),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_28),
.C(n_53),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_156),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_137),
.A2(n_147),
.B1(n_121),
.B2(n_120),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_135),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_138),
.B(n_149),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_127),
.A2(n_99),
.B(n_105),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_141),
.B(n_142),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_129),
.A2(n_126),
.B(n_119),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_119),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_148),
.Y(n_168)
);

OA22x2_ASAP7_75t_L g167 ( 
.A1(n_146),
.A2(n_157),
.B1(n_53),
.B2(n_29),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_113),
.A2(n_109),
.B1(n_99),
.B2(n_92),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_135),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_123),
.A2(n_94),
.B1(n_90),
.B2(n_100),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_150),
.A2(n_145),
.B1(n_149),
.B2(n_137),
.Y(n_165)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_122),
.Y(n_154)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_110),
.Y(n_155)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_155),
.Y(n_172)
);

OA22x2_ASAP7_75t_L g157 ( 
.A1(n_134),
.A2(n_68),
.B1(n_101),
.B2(n_28),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_29),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_148),
.A2(n_131),
.B1(n_117),
.B2(n_114),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_160),
.A2(n_138),
.B(n_158),
.Y(n_181)
);

OAI321xp33_ASAP7_75t_L g161 ( 
.A1(n_142),
.A2(n_133),
.A3(n_124),
.B1(n_125),
.B2(n_130),
.C(n_132),
.Y(n_161)
);

AOI221xp5_ASAP7_75t_L g186 ( 
.A1(n_161),
.A2(n_162),
.B1(n_167),
.B2(n_157),
.C(n_139),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_165),
.A2(n_174),
.B(n_169),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_150),
.A2(n_53),
.B1(n_29),
.B2(n_2),
.Y(n_166)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_166),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_169),
.B(n_152),
.Y(n_183)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_175),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_53),
.B1(n_29),
.B2(n_2),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_178),
.C(n_136),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_153),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_179),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_29),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_184),
.C(n_197),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_181),
.A2(n_167),
.B1(n_8),
.B2(n_9),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_168),
.Y(n_182)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_182),
.Y(n_206)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_183),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_151),
.C(n_152),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_159),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_188),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_186),
.B(n_193),
.Y(n_208)
);

FAx1_ASAP7_75t_SL g188 ( 
.A(n_164),
.B(n_157),
.CI(n_139),
.CON(n_188),
.SN(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_172),
.B(n_157),
.Y(n_189)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_191),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_170),
.B(n_0),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_164),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_176),
.Y(n_200)
);

OA21x2_ASAP7_75t_SL g193 ( 
.A1(n_165),
.A2(n_7),
.B(n_14),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_171),
.B(n_0),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_174),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_0),
.C(n_1),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_204),
.C(n_205),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_209),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_160),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_166),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_167),
.C(n_2),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_15),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_195),
.A2(n_8),
.B1(n_14),
.B2(n_12),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_211),
.A2(n_194),
.B1(n_191),
.B2(n_196),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_206),
.A2(n_195),
.B1(n_185),
.B2(n_193),
.Y(n_212)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_212),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_199),
.B(n_187),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_213),
.B(n_215),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_207),
.A2(n_183),
.B1(n_182),
.B2(n_190),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_214),
.A2(n_217),
.B1(n_219),
.B2(n_209),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_198),
.B(n_187),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_207),
.A2(n_181),
.B1(n_188),
.B2(n_189),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_218),
.A2(n_222),
.B1(n_6),
.B2(n_15),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_208),
.A2(n_188),
.B1(n_197),
.B2(n_9),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_10),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_204),
.B(n_5),
.Y(n_222)
);

OAI221xp5_ASAP7_75t_L g223 ( 
.A1(n_214),
.A2(n_208),
.B1(n_202),
.B2(n_203),
.C(n_205),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_225),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_224),
.A2(n_228),
.B(n_220),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_5),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_220),
.A2(n_203),
.B(n_202),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_229),
.A2(n_226),
.B1(n_222),
.B2(n_10),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_216),
.A2(n_200),
.B(n_6),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_230),
.B(n_221),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_233),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_235),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_217),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_12),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_5),
.Y(n_238)
);

A2O1A1Ixp33_ASAP7_75t_L g242 ( 
.A1(n_238),
.A2(n_12),
.B(n_15),
.C(n_3),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_233),
.A2(n_4),
.B(n_10),
.Y(n_240)
);

OAI21x1_ASAP7_75t_SL g243 ( 
.A1(n_240),
.A2(n_241),
.B(n_1),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_242),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_244),
.C(n_237),
.Y(n_246)
);

OAI21x1_ASAP7_75t_L g244 ( 
.A1(n_239),
.A2(n_2),
.B(n_3),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_246),
.A2(n_245),
.B(n_241),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_3),
.Y(n_248)
);


endmodule