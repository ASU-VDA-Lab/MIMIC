module fake_ariane_3104_n_1810 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1810);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1810;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_197;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_236;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_19),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_26),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_155),
.Y(n_158)
);

INVx4_ASAP7_75t_R g159 ( 
.A(n_16),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_55),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_146),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_39),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_99),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_124),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_56),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_116),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_125),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_5),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_11),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_30),
.Y(n_171)
);

BUFx10_ASAP7_75t_L g172 ( 
.A(n_80),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_38),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_46),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_71),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_29),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_74),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_34),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_56),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_72),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_113),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_64),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_17),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_114),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_77),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_39),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_81),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_83),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_98),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_106),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_69),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_1),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_144),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_131),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_73),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_31),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_111),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_40),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_49),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_121),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_87),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_55),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_84),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_115),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_8),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_123),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_76),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_129),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_57),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_35),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_79),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_152),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_53),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_40),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_96),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_35),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_49),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_107),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_154),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_88),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_42),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_3),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_97),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_38),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_78),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_46),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_60),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_50),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_15),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_33),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_15),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_68),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_126),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_137),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_29),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_18),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_104),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_120),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_136),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_23),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_127),
.Y(n_243)
);

INVxp33_ASAP7_75t_SL g244 ( 
.A(n_58),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_54),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_70),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_102),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_89),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_143),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_109),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_53),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_149),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_91),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_122),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_134),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_133),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_23),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_19),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_33),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_30),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_135),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_4),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_27),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_14),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_85),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_32),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_61),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_8),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_24),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_32),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_48),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_45),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_130),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_117),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_2),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_54),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_94),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_10),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_31),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_5),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_57),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_6),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_139),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_119),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_142),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_118),
.Y(n_286)
);

BUFx2_ASAP7_75t_SL g287 ( 
.A(n_128),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_67),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_37),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_48),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_14),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_92),
.Y(n_292)
);

BUFx10_ASAP7_75t_L g293 ( 
.A(n_2),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_43),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_34),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_112),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_62),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_58),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_17),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_3),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_59),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_26),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_151),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_50),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_44),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_140),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_10),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_95),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_1),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_148),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_193),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_179),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_176),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_158),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_221),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_227),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_251),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_166),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_283),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_283),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_158),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_166),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_264),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_264),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_216),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_301),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_301),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_244),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_167),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_167),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_156),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_177),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_214),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_160),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_298),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_177),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_279),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_184),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_184),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_171),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_185),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_206),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_206),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_220),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_188),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_200),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_201),
.Y(n_347)
);

INVxp33_ASAP7_75t_SL g348 ( 
.A(n_207),
.Y(n_348)
);

BUFx6f_ASAP7_75t_SL g349 ( 
.A(n_172),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_220),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_298),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_211),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_222),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_214),
.B(n_0),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_212),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_222),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_247),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_247),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_292),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_249),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_249),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_164),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_250),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_250),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_215),
.Y(n_365)
);

BUFx10_ASAP7_75t_L g366 ( 
.A(n_205),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_265),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_218),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_254),
.B(n_0),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_228),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_230),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_265),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_273),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_254),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_231),
.Y(n_375)
);

INVxp33_ASAP7_75t_L g376 ( 
.A(n_157),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_238),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_172),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_242),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_157),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_274),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_362),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_362),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_323),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_314),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_362),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_314),
.B(n_274),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_362),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_362),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_362),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_330),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_330),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_321),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_321),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_329),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_329),
.B(n_273),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_332),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_332),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_336),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_336),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_338),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_338),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_339),
.Y(n_403)
);

INVx4_ASAP7_75t_L g404 ( 
.A(n_366),
.Y(n_404)
);

AND2x2_ASAP7_75t_SL g405 ( 
.A(n_378),
.B(n_164),
.Y(n_405)
);

NAND2xp33_ASAP7_75t_L g406 ( 
.A(n_354),
.B(n_205),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_339),
.Y(n_407)
);

AND3x2_ASAP7_75t_L g408 ( 
.A(n_369),
.B(n_279),
.C(n_196),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_342),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_342),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_343),
.B(n_344),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_343),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_333),
.A2(n_275),
.B1(n_224),
.B2(n_194),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_344),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_350),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g416 ( 
.A(n_324),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_350),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_353),
.B(n_284),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_353),
.B(n_284),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_356),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_356),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_357),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_357),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_358),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_358),
.B(n_288),
.Y(n_425)
);

OA21x2_ASAP7_75t_L g426 ( 
.A1(n_360),
.A2(n_288),
.B(n_186),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_360),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_361),
.B(n_161),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_361),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_367),
.Y(n_430)
);

OA21x2_ASAP7_75t_L g431 ( 
.A1(n_367),
.A2(n_186),
.B(n_164),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_372),
.B(n_161),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_363),
.A2(n_275),
.B1(n_237),
.B2(n_233),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_337),
.Y(n_434)
);

AND3x2_ASAP7_75t_L g435 ( 
.A(n_312),
.B(n_196),
.C(n_163),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_372),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_373),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_373),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_335),
.Y(n_439)
);

AND2x6_ASAP7_75t_L g440 ( 
.A(n_374),
.B(n_186),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_351),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_366),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_380),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_366),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_366),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_374),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_395),
.Y(n_447)
);

OR2x6_ASAP7_75t_L g448 ( 
.A(n_446),
.B(n_232),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g449 ( 
.A(n_434),
.B(n_319),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_446),
.B(n_374),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_391),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_446),
.B(n_439),
.Y(n_452)
);

BUFx10_ASAP7_75t_L g453 ( 
.A(n_405),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_391),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_405),
.B(n_319),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_395),
.Y(n_456)
);

OR2x2_ASAP7_75t_L g457 ( 
.A(n_434),
.B(n_320),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_405),
.B(n_378),
.Y(n_458)
);

BUFx2_ASAP7_75t_L g459 ( 
.A(n_384),
.Y(n_459)
);

NAND3xp33_ASAP7_75t_L g460 ( 
.A(n_393),
.B(n_219),
.C(n_163),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_405),
.A2(n_349),
.B1(n_381),
.B2(n_364),
.Y(n_461)
);

AOI22xp33_ASAP7_75t_L g462 ( 
.A1(n_440),
.A2(n_349),
.B1(n_376),
.B2(n_325),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_L g463 ( 
.A1(n_440),
.A2(n_349),
.B1(n_232),
.B2(n_269),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_L g464 ( 
.A1(n_440),
.A2(n_349),
.B1(n_163),
.B2(n_272),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_385),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_439),
.B(n_359),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_413),
.A2(n_320),
.B1(n_263),
.B2(n_294),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_442),
.B(n_359),
.Y(n_468)
);

INVx4_ASAP7_75t_L g469 ( 
.A(n_395),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_395),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_384),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_391),
.Y(n_472)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_395),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_442),
.B(n_444),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_395),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_439),
.B(n_348),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_391),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_442),
.B(n_331),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_441),
.B(n_334),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_395),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_391),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_443),
.B(n_340),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_395),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_441),
.B(n_341),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_391),
.Y(n_485)
);

AO22x2_ASAP7_75t_L g486 ( 
.A1(n_446),
.A2(n_387),
.B1(n_441),
.B2(n_433),
.Y(n_486)
);

INVx2_ASAP7_75t_SL g487 ( 
.A(n_444),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_440),
.A2(n_219),
.B1(n_269),
.B2(n_272),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_384),
.B(n_311),
.Y(n_489)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_395),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_416),
.B(n_315),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_442),
.B(n_444),
.Y(n_492)
);

BUFx6f_ASAP7_75t_SL g493 ( 
.A(n_440),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_442),
.B(n_345),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_443),
.B(n_346),
.Y(n_495)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_385),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_391),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_L g498 ( 
.A1(n_440),
.A2(n_385),
.B1(n_426),
.B2(n_413),
.Y(n_498)
);

OAI22xp33_ASAP7_75t_SL g499 ( 
.A1(n_428),
.A2(n_326),
.B1(n_327),
.B2(n_328),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_444),
.B(n_347),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_445),
.B(n_352),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_415),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_391),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_445),
.B(n_355),
.Y(n_504)
);

CKINVDCx16_ASAP7_75t_R g505 ( 
.A(n_416),
.Y(n_505)
);

INVxp33_ASAP7_75t_L g506 ( 
.A(n_433),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_445),
.B(n_404),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_415),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_443),
.B(n_298),
.Y(n_509)
);

INVx4_ASAP7_75t_L g510 ( 
.A(n_415),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_416),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_445),
.B(n_365),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_415),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_391),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_415),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_415),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_415),
.Y(n_517)
);

OR2x2_ASAP7_75t_L g518 ( 
.A(n_387),
.B(n_316),
.Y(n_518)
);

NAND3xp33_ASAP7_75t_L g519 ( 
.A(n_393),
.B(n_269),
.C(n_219),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_415),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_440),
.B(n_385),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_415),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_420),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_404),
.B(n_368),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g525 ( 
.A1(n_440),
.A2(n_426),
.B1(n_431),
.B2(n_428),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_420),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_420),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_420),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_420),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_420),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_432),
.Y(n_531)
);

NAND3xp33_ASAP7_75t_L g532 ( 
.A(n_393),
.B(n_276),
.C(n_272),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_408),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_420),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_404),
.B(n_370),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_408),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_440),
.A2(n_426),
.B1(n_431),
.B2(n_432),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_404),
.B(n_371),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_404),
.B(n_375),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_420),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_420),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_404),
.B(n_377),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_397),
.B(n_379),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_399),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_440),
.A2(n_276),
.B1(n_281),
.B2(n_304),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_421),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_421),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_411),
.B(n_293),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_411),
.B(n_397),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_383),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_421),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_421),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_398),
.B(n_313),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_421),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_421),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_421),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_398),
.B(n_322),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_440),
.A2(n_276),
.B1(n_309),
.B2(n_281),
.Y(n_558)
);

INVx1_ASAP7_75t_SL g559 ( 
.A(n_435),
.Y(n_559)
);

BUFx6f_ASAP7_75t_SL g560 ( 
.A(n_424),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_399),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_426),
.A2(n_281),
.B1(n_309),
.B2(n_304),
.Y(n_562)
);

INVx4_ASAP7_75t_L g563 ( 
.A(n_421),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_421),
.Y(n_564)
);

BUFx4f_ASAP7_75t_L g565 ( 
.A(n_426),
.Y(n_565)
);

NAND2xp33_ASAP7_75t_L g566 ( 
.A(n_394),
.B(n_304),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_383),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_394),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_383),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_399),
.B(n_293),
.Y(n_570)
);

INVxp67_ASAP7_75t_SL g571 ( 
.A(n_399),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_394),
.Y(n_572)
);

INVxp67_ASAP7_75t_SL g573 ( 
.A(n_399),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_410),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_410),
.B(n_175),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_410),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_401),
.Y(n_577)
);

OR2x2_ASAP7_75t_L g578 ( 
.A(n_396),
.B(n_418),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_426),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_410),
.B(n_293),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_383),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_383),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_424),
.B(n_293),
.Y(n_583)
);

NAND3xp33_ASAP7_75t_L g584 ( 
.A(n_401),
.B(n_309),
.C(n_170),
.Y(n_584)
);

INVx4_ASAP7_75t_L g585 ( 
.A(n_410),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_401),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_396),
.B(n_169),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_431),
.A2(n_194),
.B1(n_305),
.B2(n_300),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_422),
.B(n_175),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_422),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_422),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_422),
.B(n_191),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_422),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_402),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_568),
.Y(n_595)
);

INVxp67_ASAP7_75t_L g596 ( 
.A(n_459),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_568),
.Y(n_597)
);

NAND2xp33_ASAP7_75t_L g598 ( 
.A(n_524),
.B(n_402),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_572),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_453),
.B(n_402),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_504),
.B(n_403),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_494),
.B(n_403),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_578),
.B(n_403),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_572),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_465),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_583),
.B(n_427),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_578),
.B(n_409),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_479),
.B(n_409),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_471),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_531),
.B(n_406),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_465),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_548),
.A2(n_406),
.B1(n_429),
.B2(n_430),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_484),
.B(n_409),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_577),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_548),
.B(n_414),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_577),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_586),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_586),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_486),
.A2(n_431),
.B1(n_392),
.B2(n_436),
.Y(n_619)
);

INVxp67_ASAP7_75t_L g620 ( 
.A(n_459),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_594),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_594),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_549),
.B(n_414),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_453),
.B(n_414),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_453),
.B(n_417),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_452),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_455),
.B(n_458),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_549),
.B(n_417),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_511),
.B(n_318),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_543),
.B(n_417),
.Y(n_630)
);

OR2x2_ASAP7_75t_L g631 ( 
.A(n_505),
.B(n_418),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_452),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_452),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_452),
.Y(n_634)
);

INVxp67_ASAP7_75t_SL g635 ( 
.A(n_465),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_507),
.A2(n_425),
.B(n_419),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_590),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_476),
.B(n_437),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_590),
.Y(n_639)
);

NOR3xp33_ASAP7_75t_L g640 ( 
.A(n_505),
.B(n_170),
.C(n_169),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_590),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_511),
.B(n_317),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_590),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_591),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_458),
.B(n_437),
.Y(n_645)
);

A2O1A1Ixp33_ASAP7_75t_L g646 ( 
.A1(n_506),
.A2(n_437),
.B(n_438),
.C(n_436),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_453),
.B(n_565),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_565),
.B(n_427),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_535),
.B(n_429),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_591),
.Y(n_650)
);

O2A1O1Ixp33_ASAP7_75t_L g651 ( 
.A1(n_587),
.A2(n_430),
.B(n_436),
.C(n_400),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_466),
.B(n_400),
.Y(n_652)
);

INVx4_ASAP7_75t_L g653 ( 
.A(n_521),
.Y(n_653)
);

OAI22xp33_ASAP7_75t_L g654 ( 
.A1(n_467),
.A2(n_425),
.B1(n_419),
.B2(n_400),
.Y(n_654)
);

AND2x2_ASAP7_75t_SL g655 ( 
.A(n_498),
.B(n_431),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_591),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_449),
.B(n_400),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_486),
.A2(n_431),
.B1(n_392),
.B2(n_436),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_591),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_544),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_SL g661 ( 
.A1(n_467),
.A2(n_245),
.B1(n_258),
.B2(n_259),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_544),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_583),
.B(n_407),
.Y(n_663)
);

INVx8_ASAP7_75t_L g664 ( 
.A(n_560),
.Y(n_664)
);

OAI22xp5_ASAP7_75t_L g665 ( 
.A1(n_500),
.A2(n_438),
.B1(n_423),
.B2(n_412),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_544),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_501),
.B(n_407),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_561),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_478),
.B(n_407),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_496),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_565),
.B(n_407),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_533),
.B(n_536),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_486),
.A2(n_392),
.B1(n_438),
.B2(n_423),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_561),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_561),
.Y(n_675)
);

AND2x6_ASAP7_75t_L g676 ( 
.A(n_521),
.B(n_496),
.Y(n_676)
);

BUFx12f_ASAP7_75t_SL g677 ( 
.A(n_495),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_585),
.B(n_412),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_585),
.B(n_412),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_574),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_496),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_450),
.B(n_412),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_450),
.B(n_423),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_585),
.B(n_423),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_585),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_574),
.Y(n_686)
);

O2A1O1Ixp33_ASAP7_75t_L g687 ( 
.A1(n_587),
.A2(n_438),
.B(n_267),
.C(n_266),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_521),
.B(n_383),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_450),
.B(n_435),
.Y(n_689)
);

NOR3xp33_ASAP7_75t_L g690 ( 
.A(n_499),
.B(n_174),
.C(n_173),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_449),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_457),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_518),
.B(n_260),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_574),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_521),
.Y(n_695)
);

NOR2xp67_ASAP7_75t_L g696 ( 
.A(n_518),
.B(n_382),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_576),
.Y(n_697)
);

AOI21xp5_ASAP7_75t_L g698 ( 
.A1(n_474),
.A2(n_382),
.B(n_388),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_495),
.A2(n_195),
.B1(n_191),
.B2(n_286),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_468),
.B(n_262),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_576),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_450),
.B(n_382),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_457),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_571),
.B(n_195),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_487),
.B(n_576),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_487),
.B(n_383),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_533),
.B(n_173),
.Y(n_707)
);

HB1xp67_ASAP7_75t_L g708 ( 
.A(n_557),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_593),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_560),
.A2(n_286),
.B1(n_213),
.B2(n_287),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_573),
.B(n_388),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_593),
.Y(n_712)
);

OAI21xp5_ASAP7_75t_L g713 ( 
.A1(n_579),
.A2(n_388),
.B(n_234),
.Y(n_713)
);

A2O1A1Ixp33_ASAP7_75t_L g714 ( 
.A1(n_492),
.A2(n_278),
.B(n_198),
.C(n_204),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_575),
.B(n_589),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_593),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_566),
.Y(n_717)
);

AND2x4_ASAP7_75t_SL g718 ( 
.A(n_461),
.B(n_172),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_592),
.B(n_538),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_525),
.B(n_383),
.Y(n_720)
);

NAND2xp33_ASAP7_75t_SL g721 ( 
.A(n_560),
.B(n_268),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_482),
.B(n_271),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_537),
.B(n_383),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_493),
.Y(n_724)
);

BUFx3_ASAP7_75t_L g725 ( 
.A(n_485),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_579),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_536),
.A2(n_213),
.B1(n_287),
.B2(n_310),
.Y(n_727)
);

OR2x2_ASAP7_75t_L g728 ( 
.A(n_553),
.B(n_174),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_512),
.B(n_388),
.Y(n_729)
);

O2A1O1Ixp33_ASAP7_75t_L g730 ( 
.A1(n_570),
.A2(n_198),
.B(n_204),
.C(n_223),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_580),
.B(n_280),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_509),
.B(n_180),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_509),
.B(n_180),
.Y(n_733)
);

NOR3xp33_ASAP7_75t_L g734 ( 
.A(n_499),
.B(n_237),
.C(n_257),
.Y(n_734)
);

HB1xp67_ASAP7_75t_L g735 ( 
.A(n_559),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_516),
.Y(n_736)
);

OR2x2_ASAP7_75t_L g737 ( 
.A(n_509),
.B(n_223),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_509),
.B(n_224),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_539),
.B(n_226),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_516),
.Y(n_740)
);

NAND2xp33_ASAP7_75t_L g741 ( 
.A(n_542),
.B(n_386),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_584),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_584),
.Y(n_743)
);

NOR3xp33_ASAP7_75t_L g744 ( 
.A(n_469),
.B(n_257),
.C(n_266),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_462),
.B(n_226),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_523),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_486),
.B(n_229),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_588),
.B(n_229),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_460),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_448),
.B(n_233),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_448),
.A2(n_178),
.B1(n_181),
.B2(n_182),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_523),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_485),
.B(n_386),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_448),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_460),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_519),
.Y(n_756)
);

INVx4_ASAP7_75t_L g757 ( 
.A(n_493),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_489),
.B(n_267),
.Y(n_758)
);

INVx8_ASAP7_75t_L g759 ( 
.A(n_493),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_448),
.B(n_270),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_448),
.B(n_270),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_SL g762 ( 
.A1(n_491),
.A2(n_299),
.B1(n_290),
.B2(n_307),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_562),
.A2(n_289),
.B1(n_278),
.B2(n_300),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_469),
.B(n_282),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_502),
.B(n_289),
.Y(n_765)
);

INVxp67_ASAP7_75t_SL g766 ( 
.A(n_485),
.Y(n_766)
);

CKINVDCx6p67_ASAP7_75t_R g767 ( 
.A(n_664),
.Y(n_767)
);

OAI21xp5_ASAP7_75t_L g768 ( 
.A1(n_671),
.A2(n_456),
.B(n_447),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_719),
.A2(n_456),
.B(n_447),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_638),
.B(n_463),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_645),
.B(n_464),
.Y(n_771)
);

OAI22xp33_ASAP7_75t_L g772 ( 
.A1(n_708),
.A2(n_302),
.B1(n_291),
.B2(n_295),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_677),
.B(n_469),
.Y(n_773)
);

OAI22xp5_ASAP7_75t_L g774 ( 
.A1(n_608),
.A2(n_473),
.B1(n_490),
.B2(n_469),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_645),
.B(n_473),
.Y(n_775)
);

OAI21xp5_ASAP7_75t_L g776 ( 
.A1(n_671),
.A2(n_475),
.B(n_470),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_604),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_627),
.B(n_672),
.Y(n_778)
);

A2O1A1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_693),
.A2(n_532),
.B(n_519),
.C(n_305),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_627),
.B(n_473),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_614),
.Y(n_781)
);

OAI21xp5_ASAP7_75t_L g782 ( 
.A1(n_648),
.A2(n_475),
.B(n_470),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_595),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_630),
.B(n_473),
.Y(n_784)
);

OR2x6_ASAP7_75t_L g785 ( 
.A(n_664),
.B(n_532),
.Y(n_785)
);

O2A1O1Ixp33_ASAP7_75t_L g786 ( 
.A1(n_693),
.A2(n_520),
.B(n_483),
.C(n_508),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_602),
.A2(n_483),
.B(n_480),
.Y(n_787)
);

AOI21x1_ASAP7_75t_L g788 ( 
.A1(n_720),
.A2(n_723),
.B(n_648),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_603),
.B(n_490),
.Y(n_789)
);

BUFx3_ASAP7_75t_L g790 ( 
.A(n_695),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_695),
.B(n_485),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_607),
.B(n_490),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_613),
.B(n_606),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_601),
.A2(n_508),
.B(n_480),
.Y(n_794)
);

AND2x4_ASAP7_75t_SL g795 ( 
.A(n_672),
.B(n_172),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_715),
.A2(n_515),
.B(n_513),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_606),
.B(n_490),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_606),
.B(n_510),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_L g799 ( 
.A1(n_623),
.A2(n_510),
.B1(n_563),
.B2(n_529),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_595),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_615),
.B(n_510),
.Y(n_801)
);

A2O1A1Ixp33_ASAP7_75t_L g802 ( 
.A1(n_628),
.A2(n_488),
.B(n_558),
.C(n_545),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_618),
.Y(n_803)
);

AOI21x1_ASAP7_75t_L g804 ( 
.A1(n_720),
.A2(n_515),
.B(n_513),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_598),
.A2(n_522),
.B(n_534),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_609),
.B(n_297),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_SL g807 ( 
.A(n_664),
.B(n_162),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_622),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_669),
.A2(n_522),
.B(n_534),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_636),
.A2(n_540),
.B(n_530),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_653),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_696),
.B(n_510),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_642),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_695),
.B(n_485),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_672),
.B(n_563),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_653),
.B(n_563),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_597),
.Y(n_817)
);

O2A1O1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_714),
.A2(n_527),
.B(n_517),
.C(n_520),
.Y(n_818)
);

AOI21x1_ASAP7_75t_L g819 ( 
.A1(n_723),
.A2(n_527),
.B(n_526),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_678),
.A2(n_530),
.B(n_517),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_678),
.A2(n_540),
.B(n_526),
.Y(n_821)
);

OAI21xp5_ASAP7_75t_L g822 ( 
.A1(n_679),
.A2(n_551),
.B(n_556),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_631),
.B(n_691),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_597),
.Y(n_824)
);

BUFx3_ASAP7_75t_L g825 ( 
.A(n_695),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_685),
.B(n_497),
.Y(n_826)
);

HB1xp67_ASAP7_75t_L g827 ( 
.A(n_596),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_679),
.A2(n_556),
.B(n_551),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_700),
.B(n_563),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_629),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_684),
.A2(n_528),
.B(n_541),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_685),
.B(n_497),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_599),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_692),
.B(n_564),
.Y(n_834)
);

A2O1A1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_646),
.A2(n_651),
.B(n_610),
.C(n_616),
.Y(n_835)
);

OAI21xp5_ASAP7_75t_L g836 ( 
.A1(n_684),
.A2(n_528),
.B(n_541),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_766),
.A2(n_547),
.B(n_555),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_655),
.A2(n_308),
.B1(n_187),
.B2(n_234),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_620),
.Y(n_839)
);

AND2x4_ASAP7_75t_L g840 ( 
.A(n_626),
.B(n_502),
.Y(n_840)
);

A2O1A1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_646),
.A2(n_564),
.B(n_554),
.C(n_555),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_599),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_616),
.Y(n_843)
);

CKINVDCx6p67_ASAP7_75t_R g844 ( 
.A(n_758),
.Y(n_844)
);

OAI21xp5_ASAP7_75t_L g845 ( 
.A1(n_667),
.A2(n_554),
.B(n_547),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_661),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_617),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_617),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_703),
.B(n_564),
.Y(n_849)
);

INVx3_ASAP7_75t_L g850 ( 
.A(n_676),
.Y(n_850)
);

AND2x4_ASAP7_75t_SL g851 ( 
.A(n_735),
.B(n_497),
.Y(n_851)
);

INVx4_ASAP7_75t_L g852 ( 
.A(n_676),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_667),
.A2(n_639),
.B(n_637),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_621),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_728),
.B(n_502),
.Y(n_855)
);

BUFx2_ASAP7_75t_L g856 ( 
.A(n_754),
.Y(n_856)
);

AO21x1_ASAP7_75t_L g857 ( 
.A1(n_649),
.A2(n_187),
.B(n_306),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_621),
.Y(n_858)
);

OAI21xp5_ASAP7_75t_L g859 ( 
.A1(n_643),
.A2(n_454),
.B(n_472),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_676),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_657),
.Y(n_861)
);

INVx3_ASAP7_75t_L g862 ( 
.A(n_676),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_711),
.A2(n_582),
.B(n_581),
.Y(n_863)
);

NOR2x1_ASAP7_75t_L g864 ( 
.A(n_704),
.B(n_502),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_700),
.B(n_529),
.Y(n_865)
);

A2O1A1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_610),
.A2(n_552),
.B(n_546),
.C(n_529),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_L g867 ( 
.A1(n_652),
.A2(n_663),
.B1(n_632),
.B2(n_634),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_654),
.B(n_529),
.Y(n_868)
);

AO21x1_ASAP7_75t_L g869 ( 
.A1(n_665),
.A2(n_234),
.B(n_187),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_736),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_709),
.B(n_497),
.Y(n_871)
);

OAI21xp33_ASAP7_75t_L g872 ( 
.A1(n_722),
.A2(n_546),
.B(n_552),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_633),
.A2(n_546),
.B1(n_552),
.B2(n_497),
.Y(n_873)
);

O2A1O1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_714),
.A2(n_546),
.B(n_552),
.C(n_481),
.Y(n_874)
);

AO21x1_ASAP7_75t_L g875 ( 
.A1(n_647),
.A2(n_713),
.B(n_624),
.Y(n_875)
);

OR2x2_ASAP7_75t_L g876 ( 
.A(n_707),
.B(n_451),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_641),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_753),
.A2(n_582),
.B(n_581),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_753),
.A2(n_582),
.B(n_581),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_706),
.A2(n_569),
.B(n_451),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_736),
.Y(n_881)
);

O2A1O1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_687),
.A2(n_503),
.B(n_481),
.C(n_451),
.Y(n_882)
);

INVx1_ASAP7_75t_SL g883 ( 
.A(n_762),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_740),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_706),
.A2(n_705),
.B(n_698),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_705),
.A2(n_569),
.B(n_481),
.Y(n_886)
);

AO21x1_ASAP7_75t_L g887 ( 
.A1(n_647),
.A2(n_306),
.B(n_308),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_707),
.B(n_503),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_709),
.B(n_550),
.Y(n_889)
);

OAI22xp5_ASAP7_75t_L g890 ( 
.A1(n_668),
.A2(n_503),
.B1(n_454),
.B2(n_477),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_740),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_641),
.A2(n_569),
.B(n_477),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_644),
.A2(n_514),
.B(n_472),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_650),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_707),
.B(n_640),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_689),
.B(n_718),
.Y(n_896)
);

NOR2xp67_ASAP7_75t_L g897 ( 
.A(n_699),
.B(n_514),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_718),
.B(n_722),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_650),
.A2(n_567),
.B(n_550),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_612),
.B(n_550),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_656),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_676),
.Y(n_902)
);

AOI21x1_ASAP7_75t_L g903 ( 
.A1(n_600),
.A2(n_308),
.B(n_306),
.Y(n_903)
);

OAI22xp5_ASAP7_75t_L g904 ( 
.A1(n_668),
.A2(n_567),
.B1(n_550),
.B2(n_390),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_725),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_674),
.A2(n_567),
.B1(n_550),
.B2(n_390),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_656),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_L g908 ( 
.A1(n_655),
.A2(n_390),
.B1(n_389),
.B2(n_386),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_765),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_742),
.B(n_567),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_746),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_635),
.A2(n_567),
.B(n_390),
.Y(n_912)
);

AOI21xp33_ASAP7_75t_L g913 ( 
.A1(n_731),
.A2(n_236),
.B(n_165),
.Y(n_913)
);

O2A1O1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_739),
.A2(n_159),
.B(n_6),
.C(n_7),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_688),
.B(n_4),
.Y(n_915)
);

AOI21x1_ASAP7_75t_L g916 ( 
.A1(n_600),
.A2(n_390),
.B(n_389),
.Y(n_916)
);

OAI21xp5_ASAP7_75t_L g917 ( 
.A1(n_659),
.A2(n_239),
.B(n_168),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_746),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_741),
.A2(n_390),
.B(n_389),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_752),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_R g921 ( 
.A(n_759),
.B(n_183),
.Y(n_921)
);

A2O1A1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_743),
.A2(n_390),
.B(n_389),
.C(n_386),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_605),
.B(n_386),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_702),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_732),
.B(n_386),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_674),
.A2(n_390),
.B1(n_389),
.B2(n_386),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_688),
.B(n_7),
.Y(n_927)
);

O2A1O1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_744),
.A2(n_159),
.B(n_11),
.C(n_12),
.Y(n_928)
);

OAI321xp33_ASAP7_75t_L g929 ( 
.A1(n_763),
.A2(n_390),
.A3(n_389),
.B1(n_386),
.B2(n_16),
.C(n_18),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_733),
.B(n_386),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_752),
.A2(n_726),
.B(n_686),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_660),
.B(n_9),
.Y(n_932)
);

AO21x1_ASAP7_75t_L g933 ( 
.A1(n_624),
.A2(n_389),
.B(n_105),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_726),
.A2(n_389),
.B(n_303),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_709),
.B(n_716),
.Y(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_737),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_682),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_675),
.A2(n_389),
.B(n_296),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_675),
.A2(n_285),
.B(n_277),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_738),
.B(n_189),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_725),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_763),
.B(n_261),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_764),
.B(n_256),
.Y(n_943)
);

O2A1O1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_662),
.A2(n_9),
.B(n_12),
.C(n_13),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_680),
.A2(n_255),
.B(n_253),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_680),
.A2(n_252),
.B1(n_248),
.B2(n_246),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_686),
.Y(n_947)
);

INVx4_ASAP7_75t_L g948 ( 
.A(n_759),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_666),
.B(n_13),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_764),
.B(n_243),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_683),
.Y(n_951)
);

O2A1O1Ixp5_ASAP7_75t_L g952 ( 
.A1(n_731),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_952)
);

OAI21xp5_ASAP7_75t_L g953 ( 
.A1(n_694),
.A2(n_241),
.B(n_240),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_750),
.B(n_235),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_L g955 ( 
.A1(n_709),
.A2(n_225),
.B1(n_217),
.B2(n_210),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_936),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_915),
.A2(n_734),
.B(n_690),
.C(n_730),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_777),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_829),
.A2(n_670),
.B(n_625),
.Y(n_959)
);

INVx5_ASAP7_75t_L g960 ( 
.A(n_860),
.Y(n_960)
);

BUFx2_ASAP7_75t_L g961 ( 
.A(n_813),
.Y(n_961)
);

OAI21xp33_ASAP7_75t_SL g962 ( 
.A1(n_838),
.A2(n_793),
.B(n_915),
.Y(n_962)
);

A2O1A1Ixp33_ASAP7_75t_SL g963 ( 
.A1(n_786),
.A2(n_712),
.B(n_701),
.C(n_697),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_775),
.A2(n_670),
.B(n_625),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_838),
.A2(n_605),
.B1(n_716),
.B2(n_611),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_783),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_780),
.B(n_611),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_767),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_921),
.Y(n_969)
);

HB1xp67_ASAP7_75t_L g970 ( 
.A(n_861),
.Y(n_970)
);

O2A1O1Ixp33_ASAP7_75t_SL g971 ( 
.A1(n_866),
.A2(n_729),
.B(n_747),
.C(n_756),
.Y(n_971)
);

INVx4_ASAP7_75t_L g972 ( 
.A(n_860),
.Y(n_972)
);

O2A1O1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_772),
.A2(n_761),
.B(n_760),
.C(n_745),
.Y(n_973)
);

BUFx2_ASAP7_75t_L g974 ( 
.A(n_813),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_784),
.A2(n_681),
.B(n_611),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_781),
.Y(n_976)
);

INVx4_ASAP7_75t_L g977 ( 
.A(n_860),
.Y(n_977)
);

INVx4_ASAP7_75t_L g978 ( 
.A(n_860),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_865),
.A2(n_681),
.B(n_611),
.Y(n_979)
);

NAND2xp33_ASAP7_75t_L g980 ( 
.A(n_811),
.B(n_716),
.Y(n_980)
);

INVx2_ASAP7_75t_SL g981 ( 
.A(n_844),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_778),
.B(n_710),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_927),
.A2(n_717),
.B(n_727),
.C(n_749),
.Y(n_983)
);

INVxp67_ASAP7_75t_L g984 ( 
.A(n_827),
.Y(n_984)
);

INVx3_ASAP7_75t_SL g985 ( 
.A(n_830),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_780),
.B(n_681),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_943),
.A2(n_716),
.B1(n_681),
.B2(n_751),
.Y(n_987)
);

O2A1O1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_913),
.A2(n_748),
.B(n_755),
.C(n_673),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_778),
.B(n_673),
.Y(n_989)
);

OR2x6_ASAP7_75t_L g990 ( 
.A(n_852),
.B(n_759),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_950),
.A2(n_619),
.B1(n_658),
.B2(n_757),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_823),
.B(n_619),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_852),
.B(n_658),
.Y(n_993)
);

OAI21xp33_ASAP7_75t_SL g994 ( 
.A1(n_927),
.A2(n_757),
.B(n_724),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_867),
.A2(n_724),
.B(n_721),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_928),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_996)
);

OAI21x1_ASAP7_75t_L g997 ( 
.A1(n_788),
.A2(n_819),
.B(n_804),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_803),
.Y(n_998)
);

AOI22xp5_ASAP7_75t_L g999 ( 
.A1(n_846),
.A2(n_199),
.B1(n_208),
.B2(n_203),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_830),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_868),
.A2(n_209),
.B(n_202),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_783),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_800),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_895),
.B(n_24),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_898),
.B(n_896),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_845),
.A2(n_197),
.B(n_192),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_808),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_896),
.B(n_25),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_948),
.B(n_25),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_817),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_800),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_SL g1012 ( 
.A(n_839),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_924),
.B(n_27),
.Y(n_1013)
);

INVx2_ASAP7_75t_SL g1014 ( 
.A(n_856),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_824),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_795),
.B(n_28),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_824),
.Y(n_1017)
);

CKINVDCx6p67_ASAP7_75t_R g1018 ( 
.A(n_846),
.Y(n_1018)
);

INVx2_ASAP7_75t_SL g1019 ( 
.A(n_921),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_842),
.Y(n_1020)
);

O2A1O1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_835),
.A2(n_28),
.B(n_36),
.C(n_37),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_795),
.B(n_36),
.Y(n_1022)
);

NAND3xp33_ASAP7_75t_SL g1023 ( 
.A(n_883),
.B(n_944),
.C(n_914),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_R g1024 ( 
.A(n_807),
.B(n_850),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_863),
.A2(n_190),
.B(n_75),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_806),
.B(n_41),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_790),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_773),
.B(n_41),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_834),
.B(n_42),
.Y(n_1029)
);

OAI22x1_ASAP7_75t_L g1030 ( 
.A1(n_932),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_1030)
);

INVxp67_ASAP7_75t_L g1031 ( 
.A(n_932),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_797),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_937),
.B(n_47),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_842),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_951),
.B(n_855),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_847),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_847),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_773),
.B(n_51),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_815),
.B(n_52),
.Y(n_1039)
);

CKINVDCx8_ASAP7_75t_R g1040 ( 
.A(n_785),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_815),
.B(n_59),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_769),
.A2(n_93),
.B(n_145),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_798),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_1043)
);

AOI22xp33_ASAP7_75t_L g1044 ( 
.A1(n_771),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_876),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_909),
.B(n_82),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_858),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_858),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_833),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_R g1050 ( 
.A(n_850),
.B(n_86),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_849),
.B(n_790),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_870),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_870),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_851),
.B(n_147),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_787),
.A2(n_90),
.B(n_100),
.Y(n_1055)
);

OR2x6_ASAP7_75t_SL g1056 ( 
.A(n_942),
.B(n_101),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_835),
.A2(n_103),
.B(n_108),
.C(n_110),
.Y(n_1057)
);

OA21x2_ASAP7_75t_L g1058 ( 
.A1(n_922),
.A2(n_132),
.B(n_141),
.Y(n_1058)
);

INVxp67_ASAP7_75t_L g1059 ( 
.A(n_949),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_789),
.A2(n_792),
.B(n_885),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_881),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_825),
.B(n_843),
.Y(n_1062)
);

NOR2x1_ASAP7_75t_L g1063 ( 
.A(n_825),
.B(n_811),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_881),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_848),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_854),
.B(n_851),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_794),
.A2(n_810),
.B(n_796),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_809),
.A2(n_801),
.B(n_886),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_899),
.A2(n_812),
.B(n_878),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_948),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_879),
.A2(n_912),
.B(n_872),
.Y(n_1071)
);

INVx4_ASAP7_75t_L g1072 ( 
.A(n_852),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_954),
.B(n_840),
.Y(n_1073)
);

AOI221xp5_ASAP7_75t_L g1074 ( 
.A1(n_929),
.A2(n_779),
.B1(n_949),
.B2(n_952),
.C(n_770),
.Y(n_1074)
);

CKINVDCx14_ASAP7_75t_R g1075 ( 
.A(n_948),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_840),
.B(n_877),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_816),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_888),
.B(n_840),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_905),
.B(n_941),
.Y(n_1079)
);

AOI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_850),
.A2(n_862),
.B1(n_902),
.B2(n_897),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_837),
.A2(n_880),
.B(n_853),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_R g1082 ( 
.A(n_862),
.B(n_902),
.Y(n_1082)
);

AOI22xp33_ASAP7_75t_L g1083 ( 
.A1(n_884),
.A2(n_911),
.B1(n_891),
.B2(n_920),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_785),
.B(n_894),
.Y(n_1084)
);

BUFx3_ASAP7_75t_L g1085 ( 
.A(n_905),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_901),
.B(n_907),
.Y(n_1086)
);

OAI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_816),
.A2(n_866),
.B1(n_873),
.B2(n_940),
.Y(n_1087)
);

BUFx3_ASAP7_75t_L g1088 ( 
.A(n_905),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_884),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_816),
.A2(n_900),
.B1(n_941),
.B2(n_802),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_779),
.A2(n_874),
.B(n_841),
.C(n_818),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_923),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_941),
.B(n_875),
.Y(n_1093)
);

AOI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_785),
.A2(n_955),
.B1(n_946),
.B2(n_791),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_802),
.A2(n_953),
.B1(n_917),
.B2(n_910),
.Y(n_1095)
);

BUFx2_ASAP7_75t_L g1096 ( 
.A(n_923),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_947),
.B(n_918),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_923),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_826),
.A2(n_832),
.B(n_831),
.Y(n_1099)
);

O2A1O1Ixp5_ASAP7_75t_L g1100 ( 
.A1(n_869),
.A2(n_857),
.B(n_933),
.C(n_922),
.Y(n_1100)
);

INVxp33_ASAP7_75t_SL g1101 ( 
.A(n_935),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_947),
.B(n_920),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_SL g1103 ( 
.A1(n_891),
.A2(n_918),
.B1(n_911),
.B2(n_774),
.Y(n_1103)
);

AOI221xp5_ASAP7_75t_SL g1104 ( 
.A1(n_1021),
.A2(n_882),
.B1(n_841),
.B2(n_799),
.C(n_945),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1060),
.A2(n_904),
.B(n_906),
.Y(n_1105)
);

O2A1O1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_1031),
.A2(n_791),
.B(n_814),
.C(n_832),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_970),
.B(n_814),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_989),
.B(n_992),
.Y(n_1108)
);

BUFx3_ASAP7_75t_L g1109 ( 
.A(n_968),
.Y(n_1109)
);

INVxp33_ASAP7_75t_L g1110 ( 
.A(n_1012),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_958),
.Y(n_1111)
);

AOI21xp33_ASAP7_75t_L g1112 ( 
.A1(n_962),
.A2(n_890),
.B(n_887),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_970),
.B(n_908),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_1069),
.A2(n_1071),
.B(n_1067),
.Y(n_1114)
);

AO31x2_ASAP7_75t_L g1115 ( 
.A1(n_1095),
.A2(n_931),
.A3(n_934),
.B(n_938),
.Y(n_1115)
);

O2A1O1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_1059),
.A2(n_826),
.B(n_871),
.C(n_935),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1068),
.A2(n_889),
.B(n_871),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_976),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1081),
.A2(n_889),
.B(n_805),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_967),
.A2(n_986),
.B(n_1087),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_SL g1121 ( 
.A1(n_1030),
.A2(n_908),
.B1(n_864),
.B2(n_782),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_1039),
.A2(n_925),
.B1(n_930),
.B2(n_768),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_997),
.A2(n_916),
.B(n_903),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_998),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_967),
.A2(n_859),
.B(n_893),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1007),
.Y(n_1126)
);

O2A1O1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_957),
.A2(n_939),
.B(n_776),
.C(n_822),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_1028),
.B(n_836),
.Y(n_1128)
);

INVx2_ASAP7_75t_SL g1129 ( 
.A(n_981),
.Y(n_1129)
);

NAND2xp33_ASAP7_75t_SL g1130 ( 
.A(n_1024),
.B(n_926),
.Y(n_1130)
);

AO21x1_ASAP7_75t_L g1131 ( 
.A1(n_1008),
.A2(n_820),
.B(n_821),
.Y(n_1131)
);

BUFx2_ASAP7_75t_L g1132 ( 
.A(n_961),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1099),
.A2(n_919),
.B(n_892),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_974),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_956),
.B(n_828),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_1005),
.B(n_1004),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_956),
.B(n_1045),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1010),
.Y(n_1138)
);

CKINVDCx11_ASAP7_75t_R g1139 ( 
.A(n_985),
.Y(n_1139)
);

BUFx2_ASAP7_75t_L g1140 ( 
.A(n_1000),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_985),
.Y(n_1141)
);

OAI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1091),
.A2(n_1074),
.B(n_983),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1003),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1049),
.Y(n_1144)
);

AOI221xp5_ASAP7_75t_L g1145 ( 
.A1(n_1004),
.A2(n_1023),
.B1(n_957),
.B2(n_996),
.C(n_983),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1100),
.A2(n_979),
.B(n_1093),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1073),
.B(n_1035),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_969),
.Y(n_1148)
);

AO21x2_ASAP7_75t_L g1149 ( 
.A1(n_1093),
.A2(n_993),
.B(n_971),
.Y(n_1149)
);

AOI21x1_ASAP7_75t_L g1150 ( 
.A1(n_986),
.A2(n_1090),
.B(n_959),
.Y(n_1150)
);

AO32x2_ASAP7_75t_L g1151 ( 
.A1(n_991),
.A2(n_1043),
.A3(n_1032),
.B1(n_987),
.B2(n_965),
.Y(n_1151)
);

O2A1O1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_1028),
.A2(n_1039),
.B(n_984),
.C(n_1038),
.Y(n_1152)
);

AO31x2_ASAP7_75t_L g1153 ( 
.A1(n_1091),
.A2(n_1015),
.A3(n_1011),
.B(n_1017),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_964),
.A2(n_971),
.B(n_975),
.Y(n_1154)
);

INVx4_ASAP7_75t_L g1155 ( 
.A(n_1070),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1065),
.Y(n_1156)
);

OA21x2_ASAP7_75t_L g1157 ( 
.A1(n_993),
.A2(n_1025),
.B(n_995),
.Y(n_1157)
);

O2A1O1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_1016),
.A2(n_1022),
.B(n_1041),
.C(n_1013),
.Y(n_1158)
);

INVx3_ASAP7_75t_L g1159 ( 
.A(n_960),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1073),
.B(n_1078),
.Y(n_1160)
);

AO31x2_ASAP7_75t_L g1161 ( 
.A1(n_966),
.A2(n_1047),
.A3(n_1011),
.B(n_1015),
.Y(n_1161)
);

OR2x2_ASAP7_75t_L g1162 ( 
.A(n_1014),
.B(n_1045),
.Y(n_1162)
);

AO31x2_ASAP7_75t_L g1163 ( 
.A1(n_966),
.A2(n_1047),
.A3(n_1017),
.B(n_1064),
.Y(n_1163)
);

NAND3xp33_ASAP7_75t_SL g1164 ( 
.A(n_999),
.B(n_1026),
.C(n_1040),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1020),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_980),
.A2(n_994),
.B(n_1055),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_982),
.B(n_1076),
.Y(n_1167)
);

NAND2xp33_ASAP7_75t_SL g1168 ( 
.A(n_1024),
.B(n_1077),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1009),
.A2(n_1033),
.B1(n_1094),
.B2(n_1077),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1042),
.A2(n_1079),
.B(n_1046),
.Y(n_1170)
);

INVx3_ASAP7_75t_L g1171 ( 
.A(n_960),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1079),
.A2(n_963),
.B(n_1057),
.Y(n_1172)
);

OA21x2_ASAP7_75t_L g1173 ( 
.A1(n_1083),
.A2(n_1097),
.B(n_1102),
.Y(n_1173)
);

OR2x2_ASAP7_75t_L g1174 ( 
.A(n_1029),
.B(n_1018),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1034),
.Y(n_1175)
);

INVx5_ASAP7_75t_L g1176 ( 
.A(n_1077),
.Y(n_1176)
);

NOR2xp67_ASAP7_75t_SL g1177 ( 
.A(n_1019),
.B(n_960),
.Y(n_1177)
);

AOI221x1_ASAP7_75t_L g1178 ( 
.A1(n_1006),
.A2(n_1001),
.B1(n_1076),
.B2(n_1051),
.C(n_1066),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_1101),
.B(n_1075),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_1096),
.A2(n_1048),
.B1(n_1037),
.B2(n_1036),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_1027),
.Y(n_1181)
);

A2O1A1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_973),
.A2(n_988),
.B(n_1086),
.C(n_1044),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1089),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_L g1184 ( 
.A(n_1075),
.B(n_1077),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1103),
.A2(n_963),
.B(n_1044),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_960),
.B(n_1009),
.Y(n_1186)
);

INVx1_ASAP7_75t_SL g1187 ( 
.A(n_1092),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1072),
.A2(n_1058),
.B(n_990),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1072),
.A2(n_1058),
.B(n_990),
.Y(n_1189)
);

O2A1O1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1084),
.A2(n_1088),
.B(n_1085),
.C(n_1062),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1086),
.B(n_1098),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1052),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1058),
.A2(n_1083),
.B(n_1080),
.Y(n_1193)
);

BUFx2_ASAP7_75t_L g1194 ( 
.A(n_1092),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_990),
.A2(n_1088),
.B(n_1085),
.Y(n_1195)
);

AO31x2_ASAP7_75t_L g1196 ( 
.A1(n_1052),
.A2(n_1061),
.A3(n_1064),
.B(n_1053),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_1092),
.B(n_1098),
.Y(n_1197)
);

OAI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1056),
.A2(n_1098),
.B1(n_977),
.B2(n_978),
.Y(n_1198)
);

NOR2x1_ASAP7_75t_R g1199 ( 
.A(n_1070),
.B(n_972),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1063),
.A2(n_1054),
.B(n_1061),
.C(n_1053),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1070),
.A2(n_972),
.B1(n_977),
.B2(n_978),
.Y(n_1201)
);

BUFx2_ASAP7_75t_SL g1202 ( 
.A(n_1070),
.Y(n_1202)
);

INVxp67_ASAP7_75t_L g1203 ( 
.A(n_1082),
.Y(n_1203)
);

OAI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1050),
.A2(n_1031),
.B1(n_1059),
.B2(n_1039),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1050),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_1082),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_989),
.B(n_778),
.Y(n_1207)
);

BUFx2_ASAP7_75t_L g1208 ( 
.A(n_961),
.Y(n_1208)
);

AO31x2_ASAP7_75t_L g1209 ( 
.A1(n_1095),
.A2(n_857),
.A3(n_887),
.B(n_875),
.Y(n_1209)
);

AO31x2_ASAP7_75t_L g1210 ( 
.A1(n_1095),
.A2(n_857),
.A3(n_887),
.B(n_875),
.Y(n_1210)
);

A2O1A1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_962),
.A2(n_1031),
.B(n_1059),
.C(n_983),
.Y(n_1211)
);

AO22x2_ASAP7_75t_L g1212 ( 
.A1(n_1023),
.A2(n_1095),
.B1(n_992),
.B2(n_898),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_968),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1069),
.A2(n_1071),
.B(n_1067),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1060),
.A2(n_602),
.B(n_1067),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_1077),
.B(n_790),
.Y(n_1216)
);

INVx2_ASAP7_75t_SL g1217 ( 
.A(n_981),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_1005),
.B(n_505),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_1077),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_970),
.B(n_823),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_958),
.Y(n_1221)
);

O2A1O1Ixp33_ASAP7_75t_SL g1222 ( 
.A1(n_963),
.A2(n_793),
.B(n_1059),
.C(n_1031),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1060),
.A2(n_602),
.B(n_1067),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1002),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1060),
.A2(n_602),
.B(n_1067),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_958),
.Y(n_1226)
);

AO32x2_ASAP7_75t_L g1227 ( 
.A1(n_1090),
.A2(n_1095),
.A3(n_991),
.B1(n_1087),
.B2(n_1043),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1060),
.A2(n_602),
.B(n_1067),
.Y(n_1228)
);

NAND3xp33_ASAP7_75t_SL g1229 ( 
.A(n_999),
.B(n_491),
.C(n_489),
.Y(n_1229)
);

A2O1A1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_962),
.A2(n_1031),
.B(n_1059),
.C(n_983),
.Y(n_1230)
);

INVx8_ASAP7_75t_L g1231 ( 
.A(n_960),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1060),
.A2(n_602),
.B(n_1067),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_958),
.Y(n_1233)
);

AND2x4_ASAP7_75t_L g1234 ( 
.A(n_1077),
.B(n_790),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1060),
.A2(n_602),
.B(n_1067),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1069),
.A2(n_1071),
.B(n_1067),
.Y(n_1236)
);

INVx3_ASAP7_75t_SL g1237 ( 
.A(n_968),
.Y(n_1237)
);

AND2x4_ASAP7_75t_L g1238 ( 
.A(n_1077),
.B(n_790),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1069),
.A2(n_1071),
.B(n_1067),
.Y(n_1239)
);

OAI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_962),
.A2(n_835),
.B(n_866),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_962),
.A2(n_835),
.B(n_866),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_989),
.B(n_778),
.Y(n_1242)
);

AO31x2_ASAP7_75t_L g1243 ( 
.A1(n_1095),
.A2(n_857),
.A3(n_887),
.B(n_875),
.Y(n_1243)
);

AOI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1004),
.A2(n_505),
.B1(n_846),
.B2(n_471),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1069),
.A2(n_1071),
.B(n_1067),
.Y(n_1245)
);

OA21x2_ASAP7_75t_L g1246 ( 
.A1(n_1100),
.A2(n_1071),
.B(n_1067),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_970),
.B(n_708),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_958),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1077),
.B(n_790),
.Y(n_1249)
);

NAND3xp33_ASAP7_75t_SL g1250 ( 
.A(n_999),
.B(n_491),
.C(n_489),
.Y(n_1250)
);

OA21x2_ASAP7_75t_L g1251 ( 
.A1(n_1100),
.A2(n_1071),
.B(n_1067),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1111),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1136),
.B(n_1167),
.Y(n_1253)
);

OAI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1244),
.A2(n_1229),
.B1(n_1250),
.B2(n_1204),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_1139),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1118),
.Y(n_1256)
);

BUFx3_ASAP7_75t_L g1257 ( 
.A(n_1181),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1124),
.Y(n_1258)
);

CKINVDCx6p67_ASAP7_75t_R g1259 ( 
.A(n_1237),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1167),
.B(n_1147),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1126),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1221),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1145),
.A2(n_1164),
.B1(n_1218),
.B2(n_1212),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_1141),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1212),
.A2(n_1142),
.B1(n_1113),
.B2(n_1108),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1142),
.A2(n_1108),
.B1(n_1204),
.B2(n_1169),
.Y(n_1266)
);

CKINVDCx20_ASAP7_75t_R g1267 ( 
.A(n_1148),
.Y(n_1267)
);

INVx6_ASAP7_75t_L g1268 ( 
.A(n_1176),
.Y(n_1268)
);

CKINVDCx20_ASAP7_75t_R g1269 ( 
.A(n_1109),
.Y(n_1269)
);

INVx1_ASAP7_75t_SL g1270 ( 
.A(n_1132),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1169),
.A2(n_1121),
.B1(n_1185),
.B2(n_1207),
.Y(n_1271)
);

INVx6_ASAP7_75t_L g1272 ( 
.A(n_1176),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1121),
.A2(n_1185),
.B1(n_1207),
.B2(n_1242),
.Y(n_1273)
);

BUFx2_ASAP7_75t_L g1274 ( 
.A(n_1134),
.Y(n_1274)
);

BUFx3_ASAP7_75t_L g1275 ( 
.A(n_1206),
.Y(n_1275)
);

OAI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1152),
.A2(n_1211),
.B1(n_1230),
.B2(n_1247),
.Y(n_1276)
);

OAI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1147),
.A2(n_1242),
.B1(n_1174),
.B2(n_1110),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1226),
.Y(n_1278)
);

OAI21xp33_ASAP7_75t_SL g1279 ( 
.A1(n_1128),
.A2(n_1186),
.B(n_1241),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_1140),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1233),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1220),
.B(n_1160),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_1208),
.Y(n_1283)
);

INVx1_ASAP7_75t_SL g1284 ( 
.A(n_1162),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1182),
.A2(n_1158),
.B1(n_1160),
.B2(n_1203),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1168),
.A2(n_1175),
.B1(n_1183),
.B2(n_1130),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1137),
.B(n_1191),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1248),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1240),
.A2(n_1241),
.B1(n_1179),
.B2(n_1205),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_1231),
.Y(n_1290)
);

CKINVDCx11_ASAP7_75t_R g1291 ( 
.A(n_1213),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_SL g1292 ( 
.A1(n_1240),
.A2(n_1149),
.B1(n_1193),
.B2(n_1191),
.Y(n_1292)
);

OR2x2_ASAP7_75t_L g1293 ( 
.A(n_1107),
.B(n_1153),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1219),
.Y(n_1294)
);

INVx4_ASAP7_75t_L g1295 ( 
.A(n_1231),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1138),
.Y(n_1296)
);

HB1xp67_ASAP7_75t_L g1297 ( 
.A(n_1144),
.Y(n_1297)
);

CKINVDCx11_ASAP7_75t_R g1298 ( 
.A(n_1219),
.Y(n_1298)
);

BUFx4f_ASAP7_75t_SL g1299 ( 
.A(n_1129),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1156),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_SL g1301 ( 
.A1(n_1198),
.A2(n_1120),
.B(n_1127),
.Y(n_1301)
);

OAI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1217),
.A2(n_1178),
.B1(n_1135),
.B2(n_1176),
.Y(n_1302)
);

INVxp67_ASAP7_75t_L g1303 ( 
.A(n_1197),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1166),
.A2(n_1225),
.B(n_1223),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1122),
.A2(n_1172),
.B1(n_1106),
.B2(n_1116),
.Y(n_1305)
);

BUFx12f_ASAP7_75t_L g1306 ( 
.A(n_1219),
.Y(n_1306)
);

INVx3_ASAP7_75t_L g1307 ( 
.A(n_1150),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1143),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1165),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1180),
.A2(n_1224),
.B1(n_1192),
.B2(n_1149),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1163),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_SL g1312 ( 
.A1(n_1157),
.A2(n_1122),
.B1(n_1184),
.B2(n_1227),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1163),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1196),
.Y(n_1314)
);

AND2x4_ASAP7_75t_L g1315 ( 
.A(n_1187),
.B(n_1249),
.Y(n_1315)
);

INVx3_ASAP7_75t_L g1316 ( 
.A(n_1159),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1159),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1196),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_SL g1319 ( 
.A1(n_1157),
.A2(n_1227),
.B1(n_1231),
.B2(n_1151),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1173),
.A2(n_1112),
.B1(n_1249),
.B2(n_1238),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1153),
.Y(n_1321)
);

CKINVDCx11_ASAP7_75t_R g1322 ( 
.A(n_1155),
.Y(n_1322)
);

OAI22xp33_ASAP7_75t_SL g1323 ( 
.A1(n_1187),
.A2(n_1194),
.B1(n_1216),
.B2(n_1238),
.Y(n_1323)
);

OAI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1112),
.A2(n_1227),
.B1(n_1195),
.B2(n_1155),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1153),
.Y(n_1325)
);

BUFx6f_ASAP7_75t_L g1326 ( 
.A(n_1216),
.Y(n_1326)
);

OAI21xp5_ASAP7_75t_SL g1327 ( 
.A1(n_1188),
.A2(n_1189),
.B(n_1170),
.Y(n_1327)
);

AOI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1177),
.A2(n_1234),
.B1(n_1222),
.B2(n_1201),
.Y(n_1328)
);

BUFx6f_ASAP7_75t_L g1329 ( 
.A(n_1234),
.Y(n_1329)
);

CKINVDCx11_ASAP7_75t_R g1330 ( 
.A(n_1201),
.Y(n_1330)
);

INVx3_ASAP7_75t_L g1331 ( 
.A(n_1171),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_SL g1332 ( 
.A1(n_1151),
.A2(n_1173),
.B1(n_1202),
.B2(n_1171),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1190),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_SL g1334 ( 
.A1(n_1151),
.A2(n_1154),
.B1(n_1246),
.B2(n_1251),
.Y(n_1334)
);

INVx2_ASAP7_75t_SL g1335 ( 
.A(n_1146),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1199),
.B(n_1200),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1105),
.A2(n_1125),
.B1(n_1154),
.B2(n_1235),
.Y(n_1337)
);

CKINVDCx20_ASAP7_75t_R g1338 ( 
.A(n_1131),
.Y(n_1338)
);

CKINVDCx11_ASAP7_75t_R g1339 ( 
.A(n_1104),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1209),
.Y(n_1340)
);

BUFx12f_ASAP7_75t_L g1341 ( 
.A(n_1104),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1246),
.A2(n_1251),
.B1(n_1117),
.B2(n_1119),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1215),
.A2(n_1232),
.B1(n_1228),
.B2(n_1123),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1133),
.A2(n_1114),
.B1(n_1245),
.B2(n_1239),
.Y(n_1344)
);

CKINVDCx11_ASAP7_75t_R g1345 ( 
.A(n_1209),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1214),
.A2(n_1236),
.B1(n_1209),
.B2(n_1210),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1210),
.A2(n_718),
.B1(n_506),
.B2(n_1229),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1243),
.Y(n_1348)
);

NAND2x1p5_ASAP7_75t_L g1349 ( 
.A(n_1115),
.B(n_1210),
.Y(n_1349)
);

INVx4_ASAP7_75t_L g1350 ( 
.A(n_1243),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_SL g1351 ( 
.A1(n_1243),
.A2(n_718),
.B1(n_317),
.B2(n_433),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1115),
.A2(n_718),
.B1(n_506),
.B2(n_1229),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1229),
.A2(n_718),
.B1(n_506),
.B2(n_1250),
.Y(n_1353)
);

BUFx6f_ASAP7_75t_L g1354 ( 
.A(n_1231),
.Y(n_1354)
);

INVx1_ASAP7_75t_SL g1355 ( 
.A(n_1141),
.Y(n_1355)
);

CKINVDCx20_ASAP7_75t_R g1356 ( 
.A(n_1139),
.Y(n_1356)
);

INVx3_ASAP7_75t_L g1357 ( 
.A(n_1150),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_1181),
.Y(n_1358)
);

BUFx3_ASAP7_75t_L g1359 ( 
.A(n_1181),
.Y(n_1359)
);

CKINVDCx20_ASAP7_75t_R g1360 ( 
.A(n_1139),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1161),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1229),
.A2(n_718),
.B1(n_506),
.B2(n_1250),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1229),
.A2(n_718),
.B1(n_506),
.B2(n_1250),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1111),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1111),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1148),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1111),
.Y(n_1367)
);

CKINVDCx6p67_ASAP7_75t_R g1368 ( 
.A(n_1237),
.Y(n_1368)
);

BUFx2_ASAP7_75t_L g1369 ( 
.A(n_1181),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1161),
.Y(n_1370)
);

OAI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1244),
.A2(n_489),
.B1(n_491),
.B2(n_467),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_SL g1372 ( 
.A1(n_1136),
.A2(n_718),
.B1(n_317),
.B2(n_433),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_1148),
.Y(n_1373)
);

NAND2x1p5_ASAP7_75t_L g1374 ( 
.A(n_1176),
.B(n_960),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1229),
.A2(n_718),
.B1(n_506),
.B2(n_1250),
.Y(n_1375)
);

AOI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1244),
.A2(n_846),
.B1(n_1136),
.B2(n_491),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1229),
.A2(n_718),
.B1(n_506),
.B2(n_1250),
.Y(n_1377)
);

INVx4_ASAP7_75t_L g1378 ( 
.A(n_1231),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1229),
.A2(n_718),
.B1(n_506),
.B2(n_1250),
.Y(n_1379)
);

INVx6_ASAP7_75t_L g1380 ( 
.A(n_1176),
.Y(n_1380)
);

INVx8_ASAP7_75t_L g1381 ( 
.A(n_1231),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1204),
.A2(n_1244),
.B1(n_1145),
.B2(n_1059),
.Y(n_1382)
);

INVx6_ASAP7_75t_L g1383 ( 
.A(n_1176),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1293),
.B(n_1287),
.Y(n_1384)
);

BUFx8_ASAP7_75t_SL g1385 ( 
.A(n_1255),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1293),
.Y(n_1386)
);

AOI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1304),
.A2(n_1337),
.B(n_1305),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1297),
.B(n_1252),
.Y(n_1388)
);

OA21x2_ASAP7_75t_L g1389 ( 
.A1(n_1327),
.A2(n_1342),
.B(n_1346),
.Y(n_1389)
);

NOR2xp33_ASAP7_75t_L g1390 ( 
.A(n_1253),
.B(n_1366),
.Y(n_1390)
);

OAI22xp33_ASAP7_75t_SL g1391 ( 
.A1(n_1382),
.A2(n_1276),
.B1(n_1376),
.B2(n_1285),
.Y(n_1391)
);

NAND2x1p5_ASAP7_75t_L g1392 ( 
.A(n_1333),
.B(n_1328),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1338),
.Y(n_1393)
);

OAI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1301),
.A2(n_1254),
.B(n_1371),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1321),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1256),
.B(n_1258),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1311),
.Y(n_1397)
);

OR2x6_ASAP7_75t_L g1398 ( 
.A(n_1350),
.B(n_1325),
.Y(n_1398)
);

INVx3_ASAP7_75t_L g1399 ( 
.A(n_1307),
.Y(n_1399)
);

OAI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1279),
.A2(n_1271),
.B(n_1273),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1261),
.B(n_1262),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1313),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1257),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1314),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1344),
.A2(n_1343),
.B(n_1357),
.Y(n_1405)
);

NOR2xp33_ASAP7_75t_L g1406 ( 
.A(n_1366),
.B(n_1373),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1278),
.B(n_1281),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1318),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1257),
.Y(n_1409)
);

INVx2_ASAP7_75t_SL g1410 ( 
.A(n_1358),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1260),
.B(n_1282),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1358),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1307),
.A2(n_1357),
.B(n_1349),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_SL g1414 ( 
.A(n_1269),
.B(n_1267),
.Y(n_1414)
);

INVx3_ASAP7_75t_L g1415 ( 
.A(n_1307),
.Y(n_1415)
);

NOR2x1_ASAP7_75t_SL g1416 ( 
.A(n_1341),
.B(n_1289),
.Y(n_1416)
);

INVxp67_ASAP7_75t_L g1417 ( 
.A(n_1274),
.Y(n_1417)
);

OAI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1263),
.A2(n_1302),
.B(n_1266),
.Y(n_1418)
);

BUFx2_ASAP7_75t_SL g1419 ( 
.A(n_1275),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1288),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1296),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1357),
.A2(n_1349),
.B(n_1340),
.Y(n_1422)
);

BUFx2_ASAP7_75t_L g1423 ( 
.A(n_1338),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1300),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1265),
.B(n_1284),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1364),
.Y(n_1426)
);

OR2x6_ASAP7_75t_L g1427 ( 
.A(n_1350),
.B(n_1348),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1365),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1367),
.Y(n_1429)
);

INVx2_ASAP7_75t_SL g1430 ( 
.A(n_1359),
.Y(n_1430)
);

BUFx2_ASAP7_75t_L g1431 ( 
.A(n_1335),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1312),
.B(n_1319),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_1373),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_SL g1434 ( 
.A1(n_1351),
.A2(n_1372),
.B1(n_1336),
.B2(n_1350),
.Y(n_1434)
);

OA21x2_ASAP7_75t_L g1435 ( 
.A1(n_1320),
.A2(n_1361),
.B(n_1370),
.Y(n_1435)
);

INVx4_ASAP7_75t_L g1436 ( 
.A(n_1330),
.Y(n_1436)
);

CKINVDCx20_ASAP7_75t_R g1437 ( 
.A(n_1255),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1316),
.A2(n_1331),
.B(n_1317),
.Y(n_1438)
);

BUFx2_ASAP7_75t_L g1439 ( 
.A(n_1335),
.Y(n_1439)
);

INVx4_ASAP7_75t_L g1440 ( 
.A(n_1330),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_1290),
.Y(n_1441)
);

O2A1O1Ixp33_ASAP7_75t_L g1442 ( 
.A1(n_1277),
.A2(n_1377),
.B(n_1363),
.C(n_1353),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1292),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1359),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1316),
.A2(n_1317),
.B(n_1331),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1308),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1309),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1334),
.B(n_1339),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1324),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1345),
.Y(n_1450)
);

AO21x2_ASAP7_75t_L g1451 ( 
.A1(n_1315),
.A2(n_1332),
.B(n_1303),
.Y(n_1451)
);

INVxp67_ASAP7_75t_L g1452 ( 
.A(n_1283),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1315),
.Y(n_1453)
);

INVx1_ASAP7_75t_SL g1454 ( 
.A(n_1299),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1316),
.A2(n_1317),
.B(n_1331),
.Y(n_1455)
);

NOR2xp33_ASAP7_75t_L g1456 ( 
.A(n_1267),
.B(n_1275),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_1291),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1310),
.Y(n_1458)
);

BUFx2_ASAP7_75t_SL g1459 ( 
.A(n_1264),
.Y(n_1459)
);

INVx3_ASAP7_75t_L g1460 ( 
.A(n_1295),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1294),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1369),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1270),
.B(n_1280),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1264),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1355),
.B(n_1269),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1323),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1352),
.B(n_1326),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1306),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1286),
.Y(n_1469)
);

BUFx6f_ASAP7_75t_L g1470 ( 
.A(n_1290),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1329),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1329),
.B(n_1347),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1329),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1380),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1420),
.Y(n_1475)
);

O2A1O1Ixp33_ASAP7_75t_L g1476 ( 
.A1(n_1391),
.A2(n_1362),
.B(n_1379),
.C(n_1375),
.Y(n_1476)
);

A2O1A1Ixp33_ASAP7_75t_L g1477 ( 
.A1(n_1394),
.A2(n_1400),
.B(n_1442),
.C(n_1418),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1403),
.B(n_1259),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1434),
.A2(n_1259),
.B1(n_1368),
.B2(n_1360),
.Y(n_1479)
);

OA21x2_ASAP7_75t_L g1480 ( 
.A1(n_1405),
.A2(n_1322),
.B(n_1298),
.Y(n_1480)
);

CKINVDCx11_ASAP7_75t_R g1481 ( 
.A(n_1437),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1384),
.B(n_1368),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1384),
.B(n_1298),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1388),
.B(n_1354),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1420),
.Y(n_1485)
);

BUFx3_ASAP7_75t_L g1486 ( 
.A(n_1385),
.Y(n_1486)
);

AOI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1391),
.A2(n_1383),
.B1(n_1380),
.B2(n_1268),
.Y(n_1487)
);

BUFx12f_ASAP7_75t_L g1488 ( 
.A(n_1457),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1409),
.B(n_1291),
.Y(n_1489)
);

AOI221xp5_ASAP7_75t_L g1490 ( 
.A1(n_1449),
.A2(n_1356),
.B1(n_1360),
.B2(n_1354),
.C(n_1381),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1412),
.B(n_1322),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1444),
.B(n_1356),
.Y(n_1492)
);

OR2x6_ASAP7_75t_L g1493 ( 
.A(n_1436),
.B(n_1440),
.Y(n_1493)
);

OAI221xp5_ASAP7_75t_L g1494 ( 
.A1(n_1392),
.A2(n_1295),
.B1(n_1378),
.B2(n_1383),
.C(n_1380),
.Y(n_1494)
);

AOI21xp33_ASAP7_75t_L g1495 ( 
.A1(n_1443),
.A2(n_1354),
.B(n_1295),
.Y(n_1495)
);

OAI211xp5_ASAP7_75t_SL g1496 ( 
.A1(n_1417),
.A2(n_1381),
.B(n_1378),
.C(n_1272),
.Y(n_1496)
);

CKINVDCx20_ASAP7_75t_R g1497 ( 
.A(n_1433),
.Y(n_1497)
);

O2A1O1Ixp33_ASAP7_75t_L g1498 ( 
.A1(n_1392),
.A2(n_1374),
.B(n_1381),
.C(n_1380),
.Y(n_1498)
);

NAND4xp25_ASAP7_75t_L g1499 ( 
.A(n_1390),
.B(n_1268),
.C(n_1272),
.D(n_1452),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1464),
.B(n_1410),
.Y(n_1500)
);

NOR2xp33_ASAP7_75t_L g1501 ( 
.A(n_1436),
.B(n_1440),
.Y(n_1501)
);

AND2x4_ASAP7_75t_L g1502 ( 
.A(n_1453),
.B(n_1430),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_L g1503 ( 
.A(n_1436),
.B(n_1440),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1436),
.B(n_1440),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1386),
.B(n_1388),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1462),
.B(n_1421),
.Y(n_1506)
);

AND2x2_ASAP7_75t_SL g1507 ( 
.A(n_1432),
.B(n_1393),
.Y(n_1507)
);

OAI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1392),
.A2(n_1387),
.B(n_1448),
.Y(n_1508)
);

A2O1A1Ixp33_ASAP7_75t_L g1509 ( 
.A1(n_1432),
.A2(n_1448),
.B(n_1393),
.C(n_1423),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1396),
.B(n_1401),
.Y(n_1510)
);

CKINVDCx10_ASAP7_75t_R g1511 ( 
.A(n_1414),
.Y(n_1511)
);

OAI211xp5_ASAP7_75t_SL g1512 ( 
.A1(n_1463),
.A2(n_1454),
.B(n_1465),
.C(n_1456),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1386),
.B(n_1411),
.Y(n_1513)
);

OR2x6_ASAP7_75t_L g1514 ( 
.A(n_1419),
.B(n_1459),
.Y(n_1514)
);

A2O1A1Ixp33_ASAP7_75t_L g1515 ( 
.A1(n_1423),
.A2(n_1443),
.B(n_1469),
.C(n_1450),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1459),
.B(n_1419),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1424),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1396),
.B(n_1401),
.Y(n_1518)
);

AOI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1469),
.A2(n_1472),
.B1(n_1451),
.B2(n_1466),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1407),
.B(n_1461),
.Y(n_1520)
);

O2A1O1Ixp33_ASAP7_75t_L g1521 ( 
.A1(n_1458),
.A2(n_1461),
.B(n_1468),
.C(n_1389),
.Y(n_1521)
);

OAI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1387),
.A2(n_1455),
.B(n_1445),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1424),
.Y(n_1523)
);

AOI221xp5_ASAP7_75t_L g1524 ( 
.A1(n_1458),
.A2(n_1429),
.B1(n_1426),
.B2(n_1428),
.C(n_1466),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1431),
.Y(n_1525)
);

NAND4xp25_ASAP7_75t_L g1526 ( 
.A(n_1406),
.B(n_1429),
.C(n_1428),
.D(n_1426),
.Y(n_1526)
);

OR2x6_ASAP7_75t_L g1527 ( 
.A(n_1427),
.B(n_1398),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1447),
.Y(n_1528)
);

INVx3_ASAP7_75t_L g1529 ( 
.A(n_1438),
.Y(n_1529)
);

AOI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1389),
.A2(n_1416),
.B(n_1413),
.Y(n_1530)
);

INVx3_ASAP7_75t_L g1531 ( 
.A(n_1438),
.Y(n_1531)
);

OA21x2_ASAP7_75t_L g1532 ( 
.A1(n_1413),
.A2(n_1422),
.B(n_1439),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1471),
.B(n_1473),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1475),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1485),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1529),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1507),
.A2(n_1425),
.B1(n_1467),
.B2(n_1451),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1517),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_L g1539 ( 
.A(n_1481),
.B(n_1460),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_SL g1540 ( 
.A1(n_1507),
.A2(n_1479),
.B1(n_1508),
.B2(n_1416),
.Y(n_1540)
);

BUFx3_ASAP7_75t_L g1541 ( 
.A(n_1514),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1529),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1505),
.B(n_1510),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1513),
.B(n_1389),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1513),
.B(n_1389),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1523),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1518),
.B(n_1431),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1528),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1520),
.B(n_1439),
.Y(n_1549)
);

INVxp67_ASAP7_75t_SL g1550 ( 
.A(n_1525),
.Y(n_1550)
);

AOI21xp33_ASAP7_75t_L g1551 ( 
.A1(n_1521),
.A2(n_1425),
.B(n_1397),
.Y(n_1551)
);

NOR2x1_ASAP7_75t_L g1552 ( 
.A(n_1514),
.B(n_1474),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1527),
.B(n_1399),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1525),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1505),
.B(n_1402),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1506),
.Y(n_1556)
);

INVx2_ASAP7_75t_SL g1557 ( 
.A(n_1500),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1533),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1477),
.A2(n_1460),
.B1(n_1467),
.B2(n_1441),
.Y(n_1559)
);

INVxp67_ASAP7_75t_L g1560 ( 
.A(n_1482),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1502),
.B(n_1415),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1531),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1524),
.B(n_1408),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1524),
.B(n_1526),
.Y(n_1564)
);

NOR2x1_ASAP7_75t_L g1565 ( 
.A(n_1514),
.B(n_1474),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1519),
.A2(n_1446),
.B1(n_1435),
.B2(n_1398),
.Y(n_1566)
);

INVx3_ASAP7_75t_L g1567 ( 
.A(n_1531),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1483),
.B(n_1408),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1534),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1536),
.B(n_1522),
.Y(n_1570)
);

INVx5_ASAP7_75t_SL g1571 ( 
.A(n_1553),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1534),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1544),
.B(n_1480),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1544),
.B(n_1521),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1535),
.Y(n_1575)
);

OAI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1564),
.A2(n_1476),
.B(n_1515),
.Y(n_1576)
);

BUFx2_ASAP7_75t_L g1577 ( 
.A(n_1567),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_SL g1578 ( 
.A(n_1552),
.B(n_1516),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1542),
.B(n_1480),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1554),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1542),
.B(n_1530),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1542),
.Y(n_1582)
);

NAND3xp33_ASAP7_75t_L g1583 ( 
.A(n_1564),
.B(n_1476),
.C(n_1509),
.Y(n_1583)
);

AOI221x1_ASAP7_75t_SL g1584 ( 
.A1(n_1559),
.A2(n_1499),
.B1(n_1503),
.B2(n_1501),
.C(n_1504),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1553),
.B(n_1530),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1562),
.B(n_1532),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1554),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1547),
.B(n_1532),
.Y(n_1588)
);

NAND4xp25_ASAP7_75t_L g1589 ( 
.A(n_1540),
.B(n_1504),
.C(n_1503),
.D(n_1501),
.Y(n_1589)
);

OAI31xp33_ASAP7_75t_L g1590 ( 
.A1(n_1559),
.A2(n_1512),
.A3(n_1494),
.B(n_1495),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1562),
.Y(n_1591)
);

AO21x2_ASAP7_75t_L g1592 ( 
.A1(n_1551),
.A2(n_1404),
.B(n_1395),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1550),
.Y(n_1593)
);

INVx5_ASAP7_75t_L g1594 ( 
.A(n_1553),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1545),
.B(n_1484),
.Y(n_1595)
);

OR2x2_ASAP7_75t_SL g1596 ( 
.A(n_1563),
.B(n_1470),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1545),
.B(n_1516),
.Y(n_1597)
);

INVx3_ASAP7_75t_L g1598 ( 
.A(n_1567),
.Y(n_1598)
);

AOI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1551),
.A2(n_1498),
.B(n_1494),
.Y(n_1599)
);

AND2x2_ASAP7_75t_SL g1600 ( 
.A(n_1563),
.B(n_1490),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1556),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1580),
.B(n_1538),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1588),
.B(n_1558),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1588),
.B(n_1549),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1588),
.B(n_1579),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1594),
.B(n_1541),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1569),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1580),
.B(n_1546),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1573),
.B(n_1555),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1597),
.B(n_1543),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1579),
.B(n_1549),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1579),
.B(n_1557),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1579),
.B(n_1557),
.Y(n_1613)
);

NOR2x1_ASAP7_75t_L g1614 ( 
.A(n_1589),
.B(n_1493),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1570),
.B(n_1567),
.Y(n_1615)
);

NAND3xp33_ASAP7_75t_SL g1616 ( 
.A(n_1576),
.B(n_1490),
.C(n_1537),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1570),
.B(n_1560),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1570),
.B(n_1561),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1570),
.B(n_1561),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1586),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1587),
.B(n_1546),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1587),
.B(n_1548),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1573),
.B(n_1555),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1594),
.B(n_1585),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1586),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1569),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1586),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1569),
.B(n_1548),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1572),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_L g1630 ( 
.A(n_1583),
.B(n_1486),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1572),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1572),
.B(n_1543),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1573),
.B(n_1568),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1575),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1574),
.B(n_1568),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1575),
.Y(n_1636)
);

INVx1_ASAP7_75t_SL g1637 ( 
.A(n_1635),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1607),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1635),
.B(n_1574),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1635),
.B(n_1576),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1617),
.Y(n_1641)
);

NAND3xp33_ASAP7_75t_L g1642 ( 
.A(n_1614),
.B(n_1583),
.C(n_1590),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1617),
.B(n_1571),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1620),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1607),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1626),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1617),
.B(n_1614),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1626),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1610),
.B(n_1601),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_SL g1650 ( 
.A1(n_1605),
.A2(n_1600),
.B1(n_1592),
.B2(n_1599),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1624),
.B(n_1594),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1620),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1610),
.B(n_1600),
.Y(n_1653)
);

AOI322xp5_ASAP7_75t_L g1654 ( 
.A1(n_1616),
.A2(n_1600),
.A3(n_1566),
.B1(n_1597),
.B2(n_1586),
.C1(n_1581),
.C2(n_1601),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1629),
.Y(n_1655)
);

OAI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1616),
.A2(n_1599),
.B1(n_1589),
.B2(n_1600),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1629),
.Y(n_1657)
);

AO221x1_ASAP7_75t_L g1658 ( 
.A1(n_1620),
.A2(n_1598),
.B1(n_1577),
.B2(n_1584),
.C(n_1596),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_L g1659 ( 
.A(n_1630),
.B(n_1512),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1633),
.B(n_1595),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1624),
.B(n_1594),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1633),
.B(n_1584),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1633),
.B(n_1595),
.Y(n_1663)
);

HB1xp67_ASAP7_75t_L g1664 ( 
.A(n_1602),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1632),
.B(n_1593),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1631),
.Y(n_1666)
);

AOI22xp33_ASAP7_75t_SL g1667 ( 
.A1(n_1605),
.A2(n_1592),
.B1(n_1585),
.B2(n_1581),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1632),
.B(n_1595),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1609),
.B(n_1593),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1631),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1634),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1618),
.B(n_1571),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1634),
.Y(n_1673)
);

NAND2x1p5_ASAP7_75t_L g1674 ( 
.A(n_1606),
.B(n_1552),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1636),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1636),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1618),
.B(n_1571),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1628),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1643),
.B(n_1618),
.Y(n_1679)
);

OAI21xp33_ASAP7_75t_L g1680 ( 
.A1(n_1650),
.A2(n_1605),
.B(n_1627),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1638),
.Y(n_1681)
);

CKINVDCx16_ASAP7_75t_R g1682 ( 
.A(n_1659),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1645),
.Y(n_1683)
);

NAND2x1p5_ASAP7_75t_L g1684 ( 
.A(n_1643),
.B(n_1565),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1672),
.B(n_1619),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1640),
.B(n_1656),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1639),
.B(n_1609),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1659),
.B(n_1497),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1639),
.B(n_1609),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1646),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1672),
.B(n_1619),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1648),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1655),
.Y(n_1693)
);

OAI322xp33_ASAP7_75t_L g1694 ( 
.A1(n_1662),
.A2(n_1623),
.A3(n_1625),
.B1(n_1627),
.B2(n_1608),
.C1(n_1602),
.C2(n_1622),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1637),
.B(n_1664),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1657),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1658),
.B(n_1624),
.Y(n_1697)
);

NOR2x1_ASAP7_75t_L g1698 ( 
.A(n_1642),
.B(n_1606),
.Y(n_1698)
);

BUFx2_ASAP7_75t_L g1699 ( 
.A(n_1641),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1677),
.B(n_1619),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1677),
.B(n_1604),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1658),
.B(n_1604),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1647),
.B(n_1604),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1647),
.B(n_1611),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1666),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1651),
.B(n_1611),
.Y(n_1706)
);

AND2x4_ASAP7_75t_L g1707 ( 
.A(n_1651),
.B(n_1624),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1670),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1651),
.B(n_1611),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1671),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1644),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1673),
.Y(n_1712)
);

BUFx2_ASAP7_75t_L g1713 ( 
.A(n_1649),
.Y(n_1713)
);

HB1xp67_ASAP7_75t_L g1714 ( 
.A(n_1713),
.Y(n_1714)
);

INVxp67_ASAP7_75t_L g1715 ( 
.A(n_1688),
.Y(n_1715)
);

INVx1_ASAP7_75t_SL g1716 ( 
.A(n_1713),
.Y(n_1716)
);

INVxp33_ASAP7_75t_L g1717 ( 
.A(n_1688),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1681),
.Y(n_1718)
);

NAND3xp33_ASAP7_75t_L g1719 ( 
.A(n_1682),
.B(n_1654),
.C(n_1667),
.Y(n_1719)
);

AOI32xp33_ASAP7_75t_L g1720 ( 
.A1(n_1680),
.A2(n_1653),
.A3(n_1627),
.B1(n_1625),
.B2(n_1669),
.Y(n_1720)
);

OAI21xp5_ASAP7_75t_SL g1721 ( 
.A1(n_1698),
.A2(n_1590),
.B(n_1661),
.Y(n_1721)
);

A2O1A1Ixp33_ASAP7_75t_L g1722 ( 
.A1(n_1680),
.A2(n_1625),
.B(n_1663),
.C(n_1660),
.Y(n_1722)
);

OAI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1698),
.A2(n_1649),
.B(n_1665),
.Y(n_1723)
);

AOI21xp33_ASAP7_75t_L g1724 ( 
.A1(n_1686),
.A2(n_1644),
.B(n_1652),
.Y(n_1724)
);

NAND2xp33_ASAP7_75t_L g1725 ( 
.A(n_1697),
.B(n_1674),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1681),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1687),
.B(n_1689),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1683),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1682),
.B(n_1678),
.Y(n_1729)
);

OAI31xp33_ASAP7_75t_L g1730 ( 
.A1(n_1686),
.A2(n_1660),
.A3(n_1663),
.B(n_1674),
.Y(n_1730)
);

AOI22xp5_ASAP7_75t_SL g1731 ( 
.A1(n_1702),
.A2(n_1661),
.B1(n_1492),
.B2(n_1624),
.Y(n_1731)
);

AOI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1702),
.A2(n_1592),
.B1(n_1652),
.B2(n_1585),
.Y(n_1732)
);

OAI22xp5_ASAP7_75t_SL g1733 ( 
.A1(n_1695),
.A2(n_1699),
.B1(n_1684),
.B2(n_1488),
.Y(n_1733)
);

A2O1A1Ixp33_ASAP7_75t_L g1734 ( 
.A1(n_1697),
.A2(n_1687),
.B(n_1689),
.C(n_1695),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1683),
.Y(n_1735)
);

OAI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1697),
.A2(n_1623),
.B1(n_1668),
.B2(n_1487),
.Y(n_1736)
);

NOR2x1p5_ASAP7_75t_L g1737 ( 
.A(n_1707),
.B(n_1661),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1679),
.Y(n_1738)
);

HB1xp67_ASAP7_75t_L g1739 ( 
.A(n_1714),
.Y(n_1739)
);

NOR4xp25_ASAP7_75t_L g1740 ( 
.A(n_1734),
.B(n_1716),
.C(n_1719),
.D(n_1715),
.Y(n_1740)
);

OAI33xp33_ASAP7_75t_L g1741 ( 
.A1(n_1736),
.A2(n_1729),
.A3(n_1727),
.B1(n_1733),
.B2(n_1726),
.B3(n_1735),
.Y(n_1741)
);

NOR3xp33_ASAP7_75t_L g1742 ( 
.A(n_1734),
.B(n_1694),
.C(n_1699),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1738),
.B(n_1704),
.Y(n_1743)
);

INVxp33_ASAP7_75t_L g1744 ( 
.A(n_1717),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1738),
.B(n_1679),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_L g1746 ( 
.A(n_1721),
.B(n_1694),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1722),
.B(n_1668),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1737),
.B(n_1685),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1718),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1728),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1724),
.B(n_1704),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1723),
.B(n_1684),
.Y(n_1752)
);

O2A1O1Ixp33_ASAP7_75t_L g1753 ( 
.A1(n_1722),
.A2(n_1712),
.B(n_1690),
.C(n_1710),
.Y(n_1753)
);

OAI322xp33_ASAP7_75t_L g1754 ( 
.A1(n_1736),
.A2(n_1712),
.A3(n_1690),
.B1(n_1710),
.B2(n_1692),
.C1(n_1708),
.C2(n_1693),
.Y(n_1754)
);

AOI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1732),
.A2(n_1711),
.B1(n_1703),
.B2(n_1592),
.Y(n_1755)
);

AOI222xp33_ASAP7_75t_L g1756 ( 
.A1(n_1725),
.A2(n_1711),
.B1(n_1692),
.B2(n_1708),
.C1(n_1693),
.C2(n_1696),
.Y(n_1756)
);

INVx1_ASAP7_75t_SL g1757 ( 
.A(n_1731),
.Y(n_1757)
);

AOI211xp5_ASAP7_75t_L g1758 ( 
.A1(n_1740),
.A2(n_1730),
.B(n_1703),
.C(n_1705),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1746),
.B(n_1684),
.Y(n_1759)
);

NOR3xp33_ASAP7_75t_L g1760 ( 
.A(n_1741),
.B(n_1746),
.C(n_1742),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1739),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1739),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1745),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_SL g1764 ( 
.A(n_1744),
.B(n_1720),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1743),
.Y(n_1765)
);

O2A1O1Ixp33_ASAP7_75t_L g1766 ( 
.A1(n_1754),
.A2(n_1705),
.B(n_1696),
.C(n_1711),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1748),
.Y(n_1767)
);

AOI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1757),
.A2(n_1592),
.B1(n_1691),
.B2(n_1685),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1751),
.B(n_1691),
.Y(n_1769)
);

NAND3xp33_ASAP7_75t_SL g1770 ( 
.A(n_1760),
.B(n_1758),
.C(n_1759),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1761),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1763),
.B(n_1747),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1762),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1769),
.B(n_1749),
.Y(n_1774)
);

AND3x2_ASAP7_75t_L g1775 ( 
.A(n_1760),
.B(n_1752),
.C(n_1750),
.Y(n_1775)
);

NAND5xp2_ASAP7_75t_L g1776 ( 
.A(n_1759),
.B(n_1756),
.C(n_1752),
.D(n_1753),
.E(n_1755),
.Y(n_1776)
);

HB1xp67_ASAP7_75t_L g1777 ( 
.A(n_1767),
.Y(n_1777)
);

NAND3xp33_ASAP7_75t_L g1778 ( 
.A(n_1764),
.B(n_1700),
.C(n_1701),
.Y(n_1778)
);

NOR2xp67_ASAP7_75t_L g1779 ( 
.A(n_1778),
.B(n_1765),
.Y(n_1779)
);

O2A1O1Ixp5_ASAP7_75t_L g1780 ( 
.A1(n_1772),
.A2(n_1707),
.B(n_1766),
.C(n_1709),
.Y(n_1780)
);

OAI211xp5_ASAP7_75t_L g1781 ( 
.A1(n_1770),
.A2(n_1768),
.B(n_1700),
.C(n_1709),
.Y(n_1781)
);

AOI221xp5_ASAP7_75t_L g1782 ( 
.A1(n_1776),
.A2(n_1707),
.B1(n_1706),
.B2(n_1701),
.C(n_1676),
.Y(n_1782)
);

INVxp67_ASAP7_75t_SL g1783 ( 
.A(n_1772),
.Y(n_1783)
);

NAND3xp33_ASAP7_75t_SL g1784 ( 
.A(n_1780),
.B(n_1777),
.C(n_1771),
.Y(n_1784)
);

A2O1A1Ixp33_ASAP7_75t_L g1785 ( 
.A1(n_1783),
.A2(n_1773),
.B(n_1774),
.C(n_1775),
.Y(n_1785)
);

OAI211xp5_ASAP7_75t_SL g1786 ( 
.A1(n_1781),
.A2(n_1623),
.B(n_1578),
.C(n_1675),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1782),
.Y(n_1787)
);

AOI322xp5_ASAP7_75t_L g1788 ( 
.A1(n_1779),
.A2(n_1707),
.A3(n_1706),
.B1(n_1603),
.B2(n_1613),
.C1(n_1612),
.C2(n_1615),
.Y(n_1788)
);

BUFx2_ASAP7_75t_L g1789 ( 
.A(n_1783),
.Y(n_1789)
);

CKINVDCx12_ASAP7_75t_R g1790 ( 
.A(n_1787),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1789),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1784),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1785),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1788),
.B(n_1615),
.Y(n_1794)
);

NOR3xp33_ASAP7_75t_L g1795 ( 
.A(n_1792),
.B(n_1786),
.C(n_1489),
.Y(n_1795)
);

NAND4xp75_ASAP7_75t_L g1796 ( 
.A(n_1791),
.B(n_1578),
.C(n_1478),
.D(n_1565),
.Y(n_1796)
);

AOI22x1_ASAP7_75t_L g1797 ( 
.A1(n_1793),
.A2(n_1790),
.B1(n_1794),
.B2(n_1577),
.Y(n_1797)
);

OAI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1797),
.A2(n_1793),
.B1(n_1608),
.B2(n_1622),
.Y(n_1798)
);

AOI22x1_ASAP7_75t_SL g1799 ( 
.A1(n_1798),
.A2(n_1795),
.B1(n_1796),
.B2(n_1511),
.Y(n_1799)
);

OA21x2_ASAP7_75t_L g1800 ( 
.A1(n_1799),
.A2(n_1621),
.B(n_1603),
.Y(n_1800)
);

BUFx2_ASAP7_75t_L g1801 ( 
.A(n_1800),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1801),
.B(n_1800),
.Y(n_1802)
);

AOI22xp33_ASAP7_75t_L g1803 ( 
.A1(n_1802),
.A2(n_1606),
.B1(n_1582),
.B2(n_1591),
.Y(n_1803)
);

AOI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1802),
.A2(n_1621),
.B(n_1603),
.Y(n_1804)
);

OA21x2_ASAP7_75t_L g1805 ( 
.A1(n_1804),
.A2(n_1539),
.B(n_1612),
.Y(n_1805)
);

AOI21x1_ASAP7_75t_L g1806 ( 
.A1(n_1803),
.A2(n_1612),
.B(n_1613),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1805),
.Y(n_1807)
);

AOI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1806),
.A2(n_1613),
.B(n_1628),
.Y(n_1808)
);

OAI221xp5_ASAP7_75t_R g1809 ( 
.A1(n_1807),
.A2(n_1808),
.B1(n_1615),
.B2(n_1606),
.C(n_1577),
.Y(n_1809)
);

AOI211xp5_ASAP7_75t_L g1810 ( 
.A1(n_1809),
.A2(n_1491),
.B(n_1606),
.C(n_1496),
.Y(n_1810)
);


endmodule