module fake_ariane_2341_n_1710 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1710);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1710;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_1083;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_10),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_82),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_72),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_126),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_58),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_114),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_91),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_98),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_1),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_146),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_25),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_11),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_30),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_30),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g173 ( 
.A(n_120),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_76),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_67),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_10),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_128),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_93),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_9),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_20),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_83),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_107),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_144),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_23),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_84),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_17),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_13),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_4),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_33),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_80),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_102),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_8),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_124),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_117),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_96),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_29),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_99),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_150),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_89),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_112),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_12),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_110),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_46),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_149),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_14),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_43),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_61),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_155),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_121),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_6),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_32),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_2),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_29),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_154),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_88),
.Y(n_215)
);

BUFx5_ASAP7_75t_L g216 ( 
.A(n_113),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_111),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_15),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_56),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_59),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_148),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_130),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_56),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_4),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_101),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_77),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_37),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_15),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_16),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_52),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_140),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_73),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_60),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_125),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_86),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_27),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_1),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_127),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_2),
.Y(n_239)
);

BUFx5_ASAP7_75t_L g240 ( 
.A(n_85),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_69),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_100),
.Y(n_242)
);

BUFx5_ASAP7_75t_L g243 ( 
.A(n_138),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_143),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_49),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_129),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_64),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_36),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_118),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_108),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_105),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_39),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_37),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_44),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_62),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_65),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_0),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_42),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_28),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_132),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_151),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_50),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_81),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_47),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_0),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_26),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_11),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_36),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_145),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_119),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_123),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_55),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_135),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_52),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_142),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_21),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_90),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_74),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_33),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_54),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_63),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_157),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_94),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_40),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_24),
.Y(n_285)
);

BUFx8_ASAP7_75t_SL g286 ( 
.A(n_109),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_116),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_147),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_104),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_95),
.Y(n_290)
);

BUFx10_ASAP7_75t_L g291 ( 
.A(n_17),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_6),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_79),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_3),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_78),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_131),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_31),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_141),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_106),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_57),
.Y(n_300)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_48),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_115),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_39),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_136),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_34),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_40),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_54),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_55),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_7),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_23),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_161),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_247),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_301),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_3),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_164),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_164),
.Y(n_316)
);

INVxp67_ASAP7_75t_SL g317 ( 
.A(n_188),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_172),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_180),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_201),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_160),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_205),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_166),
.Y(n_323)
);

INVxp33_ASAP7_75t_SL g324 ( 
.A(n_259),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_210),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_175),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_188),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_166),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_248),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_252),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_291),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_253),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_238),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_272),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_162),
.B(n_5),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_174),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_241),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_174),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_163),
.B(n_5),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_280),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_282),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_282),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_188),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_165),
.B(n_9),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_285),
.Y(n_345)
);

NOR2xp67_ASAP7_75t_L g346 ( 
.A(n_186),
.B(n_12),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_269),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_288),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_288),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_283),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_293),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_302),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_289),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_158),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_177),
.B(n_14),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_303),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_307),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_309),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_188),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_190),
.B(n_204),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_186),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_191),
.Y(n_362)
);

NAND2xp33_ASAP7_75t_R g363 ( 
.A(n_289),
.B(n_66),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_228),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_228),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_290),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_286),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_245),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_245),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_215),
.B(n_16),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_232),
.B(n_242),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_292),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_290),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_178),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_295),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_217),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_295),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_167),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_292),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_298),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_298),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_188),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_299),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_299),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_191),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_291),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_304),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_304),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_291),
.Y(n_389)
);

BUFx6f_ASAP7_75t_SL g390 ( 
.A(n_281),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_236),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_281),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_167),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_236),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_179),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_184),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_170),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_343),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_325),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_343),
.Y(n_400)
);

BUFx8_ASAP7_75t_L g401 ( 
.A(n_325),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_362),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_315),
.B(n_193),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_317),
.B(n_249),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_327),
.B(n_359),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_315),
.B(n_260),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_374),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_343),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_382),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_376),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_321),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_391),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_394),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_316),
.B(n_273),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_316),
.B(n_323),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_323),
.B(n_193),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_354),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_326),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_313),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_328),
.B(n_225),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_333),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_337),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_318),
.Y(n_423)
);

INVx5_ASAP7_75t_L g424 ( 
.A(n_390),
.Y(n_424)
);

NOR2x1_ASAP7_75t_L g425 ( 
.A(n_360),
.B(n_168),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_319),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_385),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_347),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_378),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_361),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_350),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_351),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_320),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_352),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_367),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_322),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_390),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_329),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_395),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_364),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_392),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_314),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_365),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_336),
.Y(n_444)
);

AND2x6_ASAP7_75t_L g445 ( 
.A(n_339),
.B(n_159),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_368),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_369),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_372),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_330),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_336),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_332),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_371),
.B(n_236),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_379),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_338),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_334),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_338),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_341),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_311),
.Y(n_458)
);

NAND2xp33_ASAP7_75t_R g459 ( 
.A(n_311),
.B(n_171),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_335),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_340),
.Y(n_461)
);

BUFx10_ASAP7_75t_L g462 ( 
.A(n_341),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_345),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_342),
.B(n_287),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_356),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_342),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_348),
.B(n_225),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_357),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_358),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_468),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_468),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_415),
.B(n_348),
.Y(n_472)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_399),
.B(n_397),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_398),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_398),
.Y(n_475)
);

AND2x4_ASAP7_75t_L g476 ( 
.A(n_402),
.B(n_331),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_408),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_469),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g479 ( 
.A(n_402),
.B(n_386),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_408),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_420),
.B(n_349),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_419),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_405),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_461),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_409),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_467),
.B(n_353),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_460),
.B(n_353),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_442),
.B(n_366),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_406),
.B(n_366),
.Y(n_489)
);

BUFx10_ASAP7_75t_L g490 ( 
.A(n_444),
.Y(n_490)
);

BUFx8_ASAP7_75t_SL g491 ( 
.A(n_458),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_409),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_461),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_414),
.B(n_373),
.Y(n_494)
);

BUFx10_ASAP7_75t_L g495 ( 
.A(n_444),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_461),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_399),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_412),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_460),
.B(n_373),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_460),
.B(n_375),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_400),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_460),
.B(n_375),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_400),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_461),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_461),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_460),
.B(n_377),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_463),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_464),
.B(n_380),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_441),
.Y(n_509)
);

INVx5_ASAP7_75t_L g510 ( 
.A(n_424),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_400),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_452),
.B(n_381),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_462),
.B(n_381),
.Y(n_513)
);

AND2x6_ASAP7_75t_L g514 ( 
.A(n_425),
.B(n_159),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_403),
.B(n_383),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_452),
.B(n_395),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_463),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_463),
.Y(n_518)
);

OR2x6_ASAP7_75t_L g519 ( 
.A(n_427),
.B(n_346),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_445),
.B(n_383),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_412),
.Y(n_521)
);

INVx6_ASAP7_75t_L g522 ( 
.A(n_424),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_423),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_412),
.Y(n_524)
);

INVx4_ASAP7_75t_L g525 ( 
.A(n_424),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_412),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_412),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_413),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_411),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_L g530 ( 
.A1(n_445),
.A2(n_324),
.B1(n_355),
.B2(n_344),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_426),
.B(n_389),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_433),
.Y(n_532)
);

AND2x6_ASAP7_75t_L g533 ( 
.A(n_436),
.B(n_182),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_440),
.Y(n_534)
);

AND2x6_ASAP7_75t_L g535 ( 
.A(n_438),
.B(n_182),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_462),
.B(n_384),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_416),
.B(n_384),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_430),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_445),
.B(n_387),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_429),
.B(n_387),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_424),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_424),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_430),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_440),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_430),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_445),
.B(n_388),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_449),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_443),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_451),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_404),
.B(n_312),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_455),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_443),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_462),
.B(n_450),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_424),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_448),
.Y(n_555)
);

BUFx2_ASAP7_75t_L g556 ( 
.A(n_450),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_448),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_454),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_446),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_445),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_454),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_446),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_445),
.B(n_312),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_465),
.B(n_393),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_447),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_447),
.Y(n_566)
);

BUFx6f_ASAP7_75t_SL g567 ( 
.A(n_427),
.Y(n_567)
);

INVx4_ASAP7_75t_L g568 ( 
.A(n_445),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_466),
.B(n_396),
.Y(n_569)
);

BUFx10_ASAP7_75t_L g570 ( 
.A(n_456),
.Y(n_570)
);

INVx6_ASAP7_75t_L g571 ( 
.A(n_437),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_453),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_456),
.A2(n_294),
.B1(n_310),
.B2(n_308),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_453),
.Y(n_574)
);

INVx4_ASAP7_75t_L g575 ( 
.A(n_457),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_401),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_439),
.B(n_396),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_466),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_457),
.A2(n_370),
.B1(n_390),
.B2(n_169),
.Y(n_579)
);

BUFx2_ASAP7_75t_L g580 ( 
.A(n_401),
.Y(n_580)
);

OR2x6_ASAP7_75t_L g581 ( 
.A(n_401),
.B(n_250),
.Y(n_581)
);

AOI22x1_ASAP7_75t_L g582 ( 
.A1(n_459),
.A2(n_176),
.B1(n_310),
.B2(n_308),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_421),
.Y(n_583)
);

INVx4_ASAP7_75t_L g584 ( 
.A(n_407),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_434),
.Y(n_585)
);

OR2x2_ASAP7_75t_L g586 ( 
.A(n_428),
.B(n_192),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_418),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_417),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_418),
.Y(n_589)
);

OAI221xp5_ASAP7_75t_L g590 ( 
.A1(n_410),
.A2(n_176),
.B1(n_171),
.B2(n_284),
.C(n_294),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_422),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_410),
.B(n_256),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_422),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_431),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_431),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_432),
.Y(n_596)
);

AND3x2_ASAP7_75t_L g597 ( 
.A(n_435),
.B(n_255),
.C(n_194),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_468),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_468),
.Y(n_599)
);

AND2x2_ASAP7_75t_SL g600 ( 
.A(n_437),
.B(n_194),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_402),
.B(n_284),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_468),
.Y(n_602)
);

AND2x6_ASAP7_75t_L g603 ( 
.A(n_425),
.B(n_255),
.Y(n_603)
);

INVx1_ASAP7_75t_SL g604 ( 
.A(n_441),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_460),
.B(n_296),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_559),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_474),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_560),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_481),
.B(n_270),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_560),
.B(n_568),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_486),
.B(n_187),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_474),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_477),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_550),
.A2(n_363),
.B1(n_277),
.B2(n_250),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_497),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_571),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_483),
.B(n_189),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_489),
.B(n_196),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_477),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_560),
.B(n_277),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_556),
.Y(n_621)
);

INVx4_ASAP7_75t_L g622 ( 
.A(n_571),
.Y(n_622)
);

AO221x1_ASAP7_75t_L g623 ( 
.A1(n_573),
.A2(n_236),
.B1(n_300),
.B2(n_263),
.C(n_275),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_571),
.Y(n_624)
);

AND2x6_ASAP7_75t_SL g625 ( 
.A(n_569),
.B(n_297),
.Y(n_625)
);

AND2x2_ASAP7_75t_SL g626 ( 
.A(n_600),
.B(n_263),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_575),
.B(n_297),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_494),
.B(n_203),
.Y(n_628)
);

OR2x2_ASAP7_75t_L g629 ( 
.A(n_473),
.B(n_604),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_499),
.B(n_206),
.Y(n_630)
);

OR2x6_ASAP7_75t_L g631 ( 
.A(n_580),
.B(n_275),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_472),
.B(n_211),
.Y(n_632)
);

BUFx8_ASAP7_75t_L g633 ( 
.A(n_588),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_488),
.B(n_212),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_500),
.B(n_213),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_508),
.B(n_218),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_568),
.B(n_173),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_480),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_568),
.B(n_173),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_520),
.B(n_173),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_571),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_563),
.A2(n_214),
.B1(n_222),
.B2(n_221),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_480),
.Y(n_643)
);

NAND3xp33_ASAP7_75t_L g644 ( 
.A(n_540),
.B(n_306),
.C(n_305),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_559),
.B(n_219),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_556),
.B(n_577),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_539),
.B(n_173),
.Y(n_647)
);

OR2x6_ASAP7_75t_L g648 ( 
.A(n_580),
.B(n_236),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_546),
.B(n_173),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_485),
.Y(n_650)
);

OAI21xp5_ASAP7_75t_L g651 ( 
.A1(n_605),
.A2(n_207),
.B(n_278),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_533),
.A2(n_279),
.B1(n_276),
.B2(n_274),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_485),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_528),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_508),
.B(n_223),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_572),
.B(n_538),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_487),
.B(n_224),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_528),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_566),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_492),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_492),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_572),
.B(n_227),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_566),
.B(n_173),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_538),
.B(n_229),
.Y(n_664)
);

OAI22xp33_ASAP7_75t_L g665 ( 
.A1(n_558),
.A2(n_268),
.B1(n_267),
.B2(n_266),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_487),
.B(n_502),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_502),
.B(n_230),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_543),
.Y(n_668)
);

OR2x6_ASAP7_75t_L g669 ( 
.A(n_576),
.B(n_237),
.Y(n_669)
);

A2O1A1Ixp33_ASAP7_75t_L g670 ( 
.A1(n_515),
.A2(n_265),
.B(n_264),
.C(n_262),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_543),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_SL g672 ( 
.A(n_584),
.B(n_239),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_588),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_545),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_586),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_490),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_501),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_577),
.B(n_254),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_501),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_566),
.B(n_173),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_503),
.Y(n_681)
);

OAI221xp5_ASAP7_75t_L g682 ( 
.A1(n_530),
.A2(n_257),
.B1(n_258),
.B2(n_271),
.C(n_261),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_506),
.B(n_18),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_562),
.B(n_181),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_566),
.B(n_173),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_565),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_574),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_516),
.B(n_183),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_516),
.B(n_185),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_511),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_523),
.B(n_195),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_511),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_532),
.B(n_197),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_475),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_506),
.B(n_18),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_561),
.B(n_198),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_475),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_557),
.Y(n_698)
);

BUFx6f_ASAP7_75t_SL g699 ( 
.A(n_576),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_473),
.B(n_19),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_561),
.B(n_216),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_547),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_549),
.B(n_199),
.Y(n_703)
);

OAI22xp33_ASAP7_75t_L g704 ( 
.A1(n_512),
.A2(n_251),
.B1(n_246),
.B2(n_244),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_537),
.B(n_19),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_578),
.B(n_243),
.Y(n_706)
);

AOI21xp5_ASAP7_75t_L g707 ( 
.A1(n_605),
.A2(n_220),
.B(n_202),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_513),
.B(n_21),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_601),
.B(n_243),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_475),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_581),
.B(n_22),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_551),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_490),
.B(n_22),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_470),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_491),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_601),
.B(n_484),
.Y(n_716)
);

A2O1A1Ixp33_ASAP7_75t_L g717 ( 
.A1(n_471),
.A2(n_200),
.B(n_208),
.C(n_209),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_548),
.B(n_231),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_476),
.B(n_226),
.Y(n_719)
);

HB1xp67_ASAP7_75t_L g720 ( 
.A(n_509),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_548),
.Y(n_721)
);

HB1xp67_ASAP7_75t_L g722 ( 
.A(n_509),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_513),
.B(n_24),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_586),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_478),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_476),
.B(n_233),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_598),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_533),
.A2(n_243),
.B1(n_240),
.B2(n_216),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_583),
.Y(n_729)
);

BUFx6f_ASAP7_75t_SL g730 ( 
.A(n_583),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_599),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_476),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_602),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_491),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_548),
.B(n_235),
.Y(n_735)
);

NOR3xp33_ASAP7_75t_L g736 ( 
.A(n_553),
.B(n_234),
.C(n_26),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_533),
.A2(n_243),
.B1(n_240),
.B2(n_216),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_552),
.B(n_243),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_552),
.B(n_243),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_552),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_482),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_603),
.B(n_243),
.Y(n_742)
);

AO221x1_ASAP7_75t_L g743 ( 
.A1(n_591),
.A2(n_25),
.B1(n_27),
.B2(n_31),
.C(n_34),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_603),
.B(n_243),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_536),
.B(n_35),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_495),
.B(n_35),
.Y(n_746)
);

INVxp67_ASAP7_75t_L g747 ( 
.A(n_585),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_603),
.B(n_240),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_603),
.B(n_240),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_536),
.B(n_38),
.Y(n_750)
);

OAI22xp5_ASAP7_75t_L g751 ( 
.A1(n_609),
.A2(n_553),
.B1(n_564),
.B2(n_601),
.Y(n_751)
);

OR2x6_ASAP7_75t_L g752 ( 
.A(n_669),
.B(n_581),
.Y(n_752)
);

NOR2x1_ASAP7_75t_L g753 ( 
.A(n_622),
.B(n_616),
.Y(n_753)
);

INVx4_ASAP7_75t_L g754 ( 
.A(n_622),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_637),
.A2(n_505),
.B(n_518),
.Y(n_755)
);

INVx5_ASAP7_75t_L g756 ( 
.A(n_608),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_702),
.Y(n_757)
);

OAI21xp5_ASAP7_75t_L g758 ( 
.A1(n_637),
.A2(n_504),
.B(n_507),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_705),
.B(n_564),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_639),
.A2(n_496),
.B(n_517),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_607),
.Y(n_761)
);

A2O1A1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_705),
.A2(n_531),
.B(n_579),
.C(n_591),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_L g763 ( 
.A1(n_639),
.A2(n_493),
.B(n_531),
.Y(n_763)
);

INVx1_ASAP7_75t_SL g764 ( 
.A(n_629),
.Y(n_764)
);

AO21x1_ASAP7_75t_L g765 ( 
.A1(n_683),
.A2(n_524),
.B(n_526),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_640),
.A2(n_531),
.B(n_498),
.Y(n_766)
);

INVx4_ASAP7_75t_L g767 ( 
.A(n_616),
.Y(n_767)
);

NAND2xp33_ASAP7_75t_L g768 ( 
.A(n_608),
.B(n_533),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_672),
.B(n_495),
.Y(n_769)
);

O2A1O1Ixp33_ASAP7_75t_L g770 ( 
.A1(n_611),
.A2(n_618),
.B(n_628),
.C(n_632),
.Y(n_770)
);

OAI21x1_ASAP7_75t_L g771 ( 
.A1(n_640),
.A2(n_526),
.B(n_527),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_610),
.A2(n_525),
.B(n_554),
.Y(n_772)
);

NAND2x1p5_ASAP7_75t_L g773 ( 
.A(n_659),
.B(n_534),
.Y(n_773)
);

O2A1O1Ixp33_ASAP7_75t_L g774 ( 
.A1(n_708),
.A2(n_590),
.B(n_593),
.C(n_591),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_610),
.A2(n_525),
.B(n_554),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_630),
.B(n_635),
.Y(n_776)
);

OAI21xp5_ASAP7_75t_L g777 ( 
.A1(n_606),
.A2(n_498),
.B(n_527),
.Y(n_777)
);

O2A1O1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_708),
.A2(n_593),
.B(n_592),
.C(n_596),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_646),
.B(n_495),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_621),
.B(n_529),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_614),
.A2(n_570),
.B1(n_587),
.B2(n_595),
.Y(n_781)
);

O2A1O1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_723),
.A2(n_750),
.B(n_745),
.C(n_695),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_701),
.A2(n_525),
.B(n_542),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_659),
.Y(n_784)
);

OAI22xp5_ASAP7_75t_L g785 ( 
.A1(n_666),
.A2(n_584),
.B1(n_582),
.B2(n_593),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_633),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_732),
.B(n_570),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_712),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_701),
.A2(n_541),
.B(n_542),
.Y(n_789)
);

NOR2x1_ASAP7_75t_L g790 ( 
.A(n_676),
.B(n_584),
.Y(n_790)
);

A2O1A1Ixp33_ASAP7_75t_L g791 ( 
.A1(n_683),
.A2(n_695),
.B(n_745),
.C(n_723),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_620),
.A2(n_541),
.B(n_510),
.Y(n_792)
);

OAI21xp33_ASAP7_75t_L g793 ( 
.A1(n_636),
.A2(n_529),
.B(n_589),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_657),
.B(n_603),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_612),
.Y(n_795)
);

NOR2xp67_ASAP7_75t_SL g796 ( 
.A(n_676),
.B(n_589),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_647),
.A2(n_498),
.B(n_521),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_657),
.B(n_603),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_L g799 ( 
.A1(n_686),
.A2(n_595),
.B1(n_594),
.B2(n_587),
.Y(n_799)
);

CKINVDCx10_ASAP7_75t_R g800 ( 
.A(n_730),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_741),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_667),
.B(n_514),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_612),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_647),
.A2(n_479),
.B(n_484),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_687),
.A2(n_479),
.B1(n_557),
.B2(n_555),
.Y(n_805)
);

NOR2x1p5_ASAP7_75t_SL g806 ( 
.A(n_668),
.B(n_216),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_667),
.B(n_514),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_626),
.B(n_585),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_636),
.B(n_514),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_626),
.B(n_519),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_R g811 ( 
.A(n_734),
.B(n_567),
.Y(n_811)
);

AOI21x1_ASAP7_75t_L g812 ( 
.A1(n_649),
.A2(n_519),
.B(n_581),
.Y(n_812)
);

INVx1_ASAP7_75t_SL g813 ( 
.A(n_615),
.Y(n_813)
);

NAND3xp33_ASAP7_75t_L g814 ( 
.A(n_655),
.B(n_557),
.C(n_534),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_654),
.Y(n_815)
);

AND2x2_ASAP7_75t_SL g816 ( 
.A(n_711),
.B(n_581),
.Y(n_816)
);

BUFx2_ASAP7_75t_SL g817 ( 
.A(n_699),
.Y(n_817)
);

BUFx4f_ASAP7_75t_L g818 ( 
.A(n_669),
.Y(n_818)
);

NOR3xp33_ASAP7_75t_L g819 ( 
.A(n_665),
.B(n_597),
.C(n_567),
.Y(n_819)
);

OR2x6_ASAP7_75t_SL g820 ( 
.A(n_700),
.B(n_567),
.Y(n_820)
);

A2O1A1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_655),
.A2(n_555),
.B(n_544),
.C(n_534),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_678),
.B(n_519),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_649),
.A2(n_484),
.B(n_544),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_673),
.B(n_519),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_634),
.B(n_617),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_662),
.B(n_535),
.Y(n_826)
);

BUFx2_ASAP7_75t_L g827 ( 
.A(n_633),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_658),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_613),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_675),
.B(n_535),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_688),
.B(n_535),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_706),
.A2(n_510),
.B(n_533),
.Y(n_832)
);

NOR2x1_ASAP7_75t_R g833 ( 
.A(n_711),
.B(n_216),
.Y(n_833)
);

CKINVDCx10_ASAP7_75t_R g834 ( 
.A(n_730),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_706),
.A2(n_510),
.B(n_533),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_677),
.A2(n_510),
.B(n_535),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_689),
.B(n_535),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_620),
.A2(n_510),
.B(n_522),
.Y(n_838)
);

NOR2xp67_ASAP7_75t_L g839 ( 
.A(n_624),
.B(n_103),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_714),
.B(n_41),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_679),
.A2(n_522),
.B(n_240),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_681),
.A2(n_216),
.B(n_42),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_681),
.A2(n_216),
.B(n_97),
.Y(n_843)
);

AOI22x1_ASAP7_75t_L g844 ( 
.A1(n_694),
.A2(n_216),
.B1(n_44),
.B2(n_45),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_619),
.Y(n_845)
);

NAND2x1_ASAP7_75t_L g846 ( 
.A(n_698),
.B(n_156),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_L g847 ( 
.A1(n_645),
.A2(n_41),
.B1(n_45),
.B2(n_48),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_674),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_690),
.A2(n_122),
.B(n_153),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_690),
.A2(n_92),
.B(n_152),
.Y(n_850)
);

BUFx12f_ASAP7_75t_L g851 ( 
.A(n_669),
.Y(n_851)
);

O2A1O1Ixp33_ASAP7_75t_SL g852 ( 
.A1(n_696),
.A2(n_50),
.B(n_51),
.C(n_53),
.Y(n_852)
);

O2A1O1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_682),
.A2(n_51),
.B(n_53),
.C(n_68),
.Y(n_853)
);

AOI21x1_ASAP7_75t_L g854 ( 
.A1(n_663),
.A2(n_70),
.B(n_71),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_720),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_724),
.B(n_722),
.Y(n_856)
);

OAI21xp5_ASAP7_75t_L g857 ( 
.A1(n_668),
.A2(n_75),
.B(n_87),
.Y(n_857)
);

OAI321xp33_ASAP7_75t_L g858 ( 
.A1(n_652),
.A2(n_651),
.A3(n_737),
.B1(n_728),
.B2(n_670),
.C(n_644),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_664),
.A2(n_133),
.B1(n_134),
.B2(n_139),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_725),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_638),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_727),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_692),
.A2(n_671),
.B(n_697),
.Y(n_863)
);

NOR2xp67_ASAP7_75t_L g864 ( 
.A(n_641),
.B(n_729),
.Y(n_864)
);

BUFx2_ASAP7_75t_L g865 ( 
.A(n_648),
.Y(n_865)
);

BUFx4f_ASAP7_75t_L g866 ( 
.A(n_648),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_L g867 ( 
.A1(n_721),
.A2(n_740),
.B1(n_652),
.B2(n_697),
.Y(n_867)
);

OAI21x1_ASAP7_75t_L g868 ( 
.A1(n_738),
.A2(n_739),
.B(n_685),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_631),
.B(n_648),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_731),
.B(n_733),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_716),
.B(n_693),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_692),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_694),
.A2(n_710),
.B(n_740),
.Y(n_873)
);

OR2x6_ASAP7_75t_L g874 ( 
.A(n_631),
.B(n_747),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_631),
.B(n_713),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_710),
.A2(n_721),
.B(n_680),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_638),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_680),
.A2(n_684),
.B(n_709),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_709),
.A2(n_735),
.B(n_718),
.Y(n_879)
);

INVxp67_ASAP7_75t_L g880 ( 
.A(n_691),
.Y(n_880)
);

O2A1O1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_736),
.A2(n_627),
.B(n_717),
.C(n_703),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_704),
.B(n_746),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_719),
.B(n_726),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_650),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_650),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_643),
.A2(n_653),
.B(n_660),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_653),
.A2(n_661),
.B(n_749),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_742),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_L g889 ( 
.A1(n_642),
.A2(n_737),
.B1(n_728),
.B2(n_748),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_744),
.A2(n_707),
.B(n_623),
.Y(n_890)
);

NAND2x1_ASAP7_75t_L g891 ( 
.A(n_743),
.B(n_699),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_625),
.B(n_715),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_656),
.A2(n_639),
.B(n_637),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_702),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_705),
.A2(n_609),
.B1(n_486),
.B2(n_481),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_609),
.B(n_481),
.Y(n_896)
);

OAI21xp33_ASAP7_75t_L g897 ( 
.A1(n_705),
.A2(n_486),
.B(n_481),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_609),
.B(n_481),
.Y(n_898)
);

AO21x1_ASAP7_75t_L g899 ( 
.A1(n_705),
.A2(n_695),
.B(n_683),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_616),
.B(n_622),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_702),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_609),
.B(n_481),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_776),
.A2(n_897),
.B(n_791),
.Y(n_903)
);

BUFx2_ASAP7_75t_L g904 ( 
.A(n_813),
.Y(n_904)
);

OAI21x1_ASAP7_75t_SL g905 ( 
.A1(n_782),
.A2(n_899),
.B(n_871),
.Y(n_905)
);

AOI21xp33_ASAP7_75t_L g906 ( 
.A1(n_895),
.A2(n_759),
.B(n_774),
.Y(n_906)
);

AND2x4_ASAP7_75t_L g907 ( 
.A(n_900),
.B(n_874),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_825),
.A2(n_768),
.B(n_770),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_764),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_761),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_898),
.B(n_902),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_901),
.Y(n_912)
);

INVx4_ASAP7_75t_L g913 ( 
.A(n_900),
.Y(n_913)
);

AO31x2_ASAP7_75t_L g914 ( 
.A1(n_765),
.A2(n_821),
.A3(n_879),
.B(n_887),
.Y(n_914)
);

INVx5_ASAP7_75t_L g915 ( 
.A(n_754),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_754),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_767),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_757),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_893),
.A2(n_873),
.B(n_878),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_751),
.B(n_810),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_788),
.Y(n_921)
);

OAI22x1_ASAP7_75t_L g922 ( 
.A1(n_808),
.A2(n_781),
.B1(n_824),
.B2(n_869),
.Y(n_922)
);

INVx5_ASAP7_75t_L g923 ( 
.A(n_767),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_873),
.A2(n_878),
.B(n_876),
.Y(n_924)
);

OR2x6_ASAP7_75t_L g925 ( 
.A(n_817),
.B(n_851),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_874),
.B(n_752),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_762),
.A2(n_870),
.B1(n_801),
.B2(n_894),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_860),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_880),
.B(n_793),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_780),
.B(n_862),
.Y(n_930)
);

A2O1A1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_778),
.A2(n_881),
.B(n_858),
.C(n_809),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_856),
.B(n_822),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_799),
.B(n_816),
.Y(n_933)
);

INVx8_ASAP7_75t_L g934 ( 
.A(n_752),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_840),
.A2(n_882),
.B1(n_866),
.B2(n_798),
.Y(n_935)
);

OAI21x1_ASAP7_75t_L g936 ( 
.A1(n_886),
.A2(n_823),
.B(n_863),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_890),
.A2(n_867),
.B(n_797),
.Y(n_937)
);

BUFx12f_ASAP7_75t_L g938 ( 
.A(n_827),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_875),
.B(n_874),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_818),
.B(n_855),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_866),
.B(n_818),
.Y(n_941)
);

OAI21x1_ASAP7_75t_L g942 ( 
.A1(n_755),
.A2(n_760),
.B(n_836),
.Y(n_942)
);

OAI21x1_ASAP7_75t_L g943 ( 
.A1(n_755),
.A2(n_760),
.B(n_836),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_766),
.A2(n_763),
.B(n_777),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_884),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_883),
.B(n_769),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_830),
.B(n_865),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_815),
.B(n_828),
.Y(n_948)
);

A2O1A1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_794),
.A2(n_802),
.B(n_807),
.C(n_853),
.Y(n_949)
);

AND2x2_ASAP7_75t_SL g950 ( 
.A(n_819),
.B(n_892),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_786),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_848),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_831),
.A2(n_837),
.B(n_826),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_872),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_756),
.B(n_811),
.Y(n_955)
);

OAI21x1_ASAP7_75t_L g956 ( 
.A1(n_758),
.A2(n_783),
.B(n_775),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_796),
.B(n_790),
.Y(n_957)
);

OAI21x1_ASAP7_75t_L g958 ( 
.A1(n_772),
.A2(n_789),
.B(n_804),
.Y(n_958)
);

INVxp67_ASAP7_75t_L g959 ( 
.A(n_833),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_779),
.B(n_805),
.Y(n_960)
);

INVx3_ASAP7_75t_L g961 ( 
.A(n_756),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_885),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_795),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_784),
.B(n_864),
.Y(n_964)
);

OAI21xp5_ASAP7_75t_L g965 ( 
.A1(n_842),
.A2(n_889),
.B(n_832),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_842),
.A2(n_832),
.B(n_835),
.Y(n_966)
);

OAI21x1_ASAP7_75t_SL g967 ( 
.A1(n_812),
.A2(n_844),
.B(n_857),
.Y(n_967)
);

INVx2_ASAP7_75t_SL g968 ( 
.A(n_800),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_803),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_756),
.A2(n_841),
.B(n_792),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_784),
.B(n_845),
.Y(n_971)
);

AOI21xp33_ASAP7_75t_L g972 ( 
.A1(n_847),
.A2(n_888),
.B(n_814),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_829),
.Y(n_973)
);

AO22x1_ASAP7_75t_L g974 ( 
.A1(n_753),
.A2(n_752),
.B1(n_820),
.B2(n_834),
.Y(n_974)
);

OAI21x1_ASAP7_75t_L g975 ( 
.A1(n_835),
.A2(n_854),
.B(n_838),
.Y(n_975)
);

OAI21x1_ASAP7_75t_L g976 ( 
.A1(n_843),
.A2(n_846),
.B(n_773),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_861),
.Y(n_977)
);

O2A1O1Ixp5_ASAP7_75t_L g978 ( 
.A1(n_787),
.A2(n_859),
.B(n_891),
.C(n_849),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_884),
.B(n_839),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_877),
.B(n_884),
.Y(n_980)
);

OAI21x1_ASAP7_75t_L g981 ( 
.A1(n_850),
.A2(n_806),
.B(n_852),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_896),
.B(n_898),
.Y(n_982)
);

INVxp67_ASAP7_75t_L g983 ( 
.A(n_764),
.Y(n_983)
);

OR2x6_ASAP7_75t_L g984 ( 
.A(n_817),
.B(n_851),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_764),
.B(n_646),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_761),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_764),
.B(n_646),
.Y(n_987)
);

NAND2x1p5_ASAP7_75t_L g988 ( 
.A(n_900),
.B(n_754),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_900),
.Y(n_989)
);

NAND2x1p5_ASAP7_75t_L g990 ( 
.A(n_900),
.B(n_754),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_757),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_776),
.A2(n_897),
.B(n_791),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_L g993 ( 
.A1(n_791),
.A2(n_782),
.B(n_893),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_757),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_896),
.B(n_898),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_896),
.B(n_898),
.Y(n_996)
);

AOI21xp33_ASAP7_75t_L g997 ( 
.A1(n_782),
.A2(n_791),
.B(n_776),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_896),
.B(n_898),
.Y(n_998)
);

AOI21xp33_ASAP7_75t_L g999 ( 
.A1(n_782),
.A2(n_791),
.B(n_776),
.Y(n_999)
);

NOR2x1_ASAP7_75t_L g1000 ( 
.A(n_817),
.B(n_583),
.Y(n_1000)
);

AOI21xp33_ASAP7_75t_L g1001 ( 
.A1(n_782),
.A2(n_791),
.B(n_776),
.Y(n_1001)
);

NOR3xp33_ASAP7_75t_L g1002 ( 
.A(n_897),
.B(n_793),
.C(n_569),
.Y(n_1002)
);

OAI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_791),
.A2(n_782),
.B(n_893),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_813),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_813),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_754),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_791),
.A2(n_782),
.B(n_893),
.Y(n_1007)
);

OAI21x1_ASAP7_75t_L g1008 ( 
.A1(n_771),
.A2(n_887),
.B(n_868),
.Y(n_1008)
);

NAND2x1p5_ASAP7_75t_L g1009 ( 
.A(n_900),
.B(n_754),
.Y(n_1009)
);

O2A1O1Ixp5_ASAP7_75t_L g1010 ( 
.A1(n_776),
.A2(n_899),
.B(n_791),
.C(n_705),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_896),
.B(n_898),
.Y(n_1011)
);

AOI221x1_ASAP7_75t_L g1012 ( 
.A1(n_791),
.A2(n_897),
.B1(n_776),
.B2(n_705),
.C(n_762),
.Y(n_1012)
);

BUFx12f_ASAP7_75t_L g1013 ( 
.A(n_827),
.Y(n_1013)
);

AOI21x1_ASAP7_75t_SL g1014 ( 
.A1(n_776),
.A2(n_898),
.B(n_896),
.Y(n_1014)
);

AO31x2_ASAP7_75t_L g1015 ( 
.A1(n_765),
.A2(n_899),
.A3(n_791),
.B(n_821),
.Y(n_1015)
);

INVx1_ASAP7_75t_SL g1016 ( 
.A(n_813),
.Y(n_1016)
);

OAI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_791),
.A2(n_782),
.B(n_893),
.Y(n_1017)
);

NAND2x1p5_ASAP7_75t_L g1018 ( 
.A(n_900),
.B(n_754),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_776),
.A2(n_897),
.B(n_791),
.Y(n_1019)
);

AND3x2_ASAP7_75t_L g1020 ( 
.A(n_827),
.B(n_580),
.C(n_588),
.Y(n_1020)
);

BUFx5_ASAP7_75t_L g1021 ( 
.A(n_888),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_776),
.A2(n_897),
.B(n_791),
.Y(n_1022)
);

OAI21xp33_ASAP7_75t_L g1023 ( 
.A1(n_897),
.A2(n_895),
.B(n_776),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_895),
.A2(n_791),
.B1(n_776),
.B2(n_759),
.Y(n_1024)
);

AO31x2_ASAP7_75t_L g1025 ( 
.A1(n_765),
.A2(n_899),
.A3(n_791),
.B(n_821),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_761),
.Y(n_1026)
);

AOI21x1_ASAP7_75t_L g1027 ( 
.A1(n_765),
.A2(n_879),
.B(n_823),
.Y(n_1027)
);

NAND2x1p5_ASAP7_75t_L g1028 ( 
.A(n_900),
.B(n_754),
.Y(n_1028)
);

BUFx10_ASAP7_75t_L g1029 ( 
.A(n_968),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_1023),
.B(n_1002),
.Y(n_1030)
);

OAI21xp33_ASAP7_75t_L g1031 ( 
.A1(n_1024),
.A2(n_911),
.B(n_997),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_913),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_912),
.Y(n_1033)
);

NAND3xp33_ASAP7_75t_L g1034 ( 
.A(n_1012),
.B(n_1010),
.C(n_992),
.Y(n_1034)
);

INVx2_ASAP7_75t_SL g1035 ( 
.A(n_904),
.Y(n_1035)
);

BUFx12f_ASAP7_75t_L g1036 ( 
.A(n_938),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_989),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_918),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_921),
.Y(n_1039)
);

BUFx10_ASAP7_75t_L g1040 ( 
.A(n_1020),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_989),
.Y(n_1041)
);

AOI22xp33_ASAP7_75t_L g1042 ( 
.A1(n_920),
.A2(n_987),
.B1(n_985),
.B2(n_1024),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_SL g1043 ( 
.A1(n_935),
.A2(n_927),
.B(n_908),
.Y(n_1043)
);

BUFx4f_ASAP7_75t_SL g1044 ( 
.A(n_1013),
.Y(n_1044)
);

INVx1_ASAP7_75t_SL g1045 ( 
.A(n_1016),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_910),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_982),
.B(n_995),
.Y(n_1047)
);

OR2x6_ASAP7_75t_L g1048 ( 
.A(n_934),
.B(n_974),
.Y(n_1048)
);

INVx4_ASAP7_75t_L g1049 ( 
.A(n_915),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_928),
.Y(n_1050)
);

AOI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_933),
.A2(n_909),
.B1(n_1011),
.B2(n_996),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_930),
.B(n_929),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_925),
.Y(n_1053)
);

OAI21xp33_ASAP7_75t_L g1054 ( 
.A1(n_997),
.A2(n_1001),
.B(n_999),
.Y(n_1054)
);

INVx1_ASAP7_75t_SL g1055 ( 
.A(n_1016),
.Y(n_1055)
);

OA21x2_ASAP7_75t_L g1056 ( 
.A1(n_965),
.A2(n_919),
.B(n_937),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_998),
.B(n_1019),
.Y(n_1057)
);

NOR2x1_ASAP7_75t_L g1058 ( 
.A(n_955),
.B(n_913),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_1022),
.B(n_999),
.Y(n_1059)
);

INVxp67_ASAP7_75t_SL g1060 ( 
.A(n_1004),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_1005),
.Y(n_1061)
);

INVx1_ASAP7_75t_SL g1062 ( 
.A(n_940),
.Y(n_1062)
);

INVx2_ASAP7_75t_SL g1063 ( 
.A(n_925),
.Y(n_1063)
);

O2A1O1Ixp5_ASAP7_75t_L g1064 ( 
.A1(n_993),
.A2(n_1017),
.B(n_1003),
.C(n_1007),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_965),
.A2(n_1017),
.B(n_993),
.Y(n_1065)
);

BUFx4f_ASAP7_75t_L g1066 ( 
.A(n_925),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_983),
.B(n_932),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_963),
.Y(n_1068)
);

OR2x2_ASAP7_75t_L g1069 ( 
.A(n_939),
.B(n_926),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_977),
.Y(n_1070)
);

AOI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_927),
.A2(n_935),
.B1(n_922),
.B2(n_950),
.Y(n_1071)
);

OR2x6_ASAP7_75t_L g1072 ( 
.A(n_934),
.B(n_926),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_986),
.Y(n_1073)
);

INVx3_ASAP7_75t_L g1074 ( 
.A(n_915),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_946),
.B(n_907),
.Y(n_1075)
);

BUFx3_ASAP7_75t_L g1076 ( 
.A(n_951),
.Y(n_1076)
);

OR2x2_ASAP7_75t_L g1077 ( 
.A(n_991),
.B(n_994),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_959),
.B(n_989),
.Y(n_1078)
);

AO31x2_ASAP7_75t_L g1079 ( 
.A1(n_931),
.A2(n_949),
.A3(n_953),
.B(n_970),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_906),
.A2(n_948),
.B1(n_960),
.B2(n_952),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_944),
.A2(n_906),
.B(n_966),
.Y(n_1081)
);

BUFx12f_ASAP7_75t_L g1082 ( 
.A(n_984),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_966),
.A2(n_919),
.B(n_924),
.Y(n_1083)
);

OR2x6_ASAP7_75t_SL g1084 ( 
.A(n_957),
.B(n_964),
.Y(n_1084)
);

AND2x4_ASAP7_75t_L g1085 ( 
.A(n_941),
.B(n_915),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_984),
.B(n_954),
.Y(n_1086)
);

OAI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_988),
.A2(n_1028),
.B1(n_1018),
.B2(n_1009),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_984),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_917),
.Y(n_1089)
);

INVxp67_ASAP7_75t_L g1090 ( 
.A(n_1000),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_945),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_945),
.Y(n_1092)
);

AOI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_947),
.A2(n_1021),
.B1(n_962),
.B2(n_934),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_1026),
.Y(n_1094)
);

AND2x4_ASAP7_75t_L g1095 ( 
.A(n_923),
.B(n_917),
.Y(n_1095)
);

OAI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_972),
.A2(n_978),
.B(n_942),
.Y(n_1096)
);

INVx2_ASAP7_75t_SL g1097 ( 
.A(n_917),
.Y(n_1097)
);

INVx3_ASAP7_75t_L g1098 ( 
.A(n_945),
.Y(n_1098)
);

NOR2xp67_ASAP7_75t_L g1099 ( 
.A(n_961),
.B(n_923),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_905),
.B(n_969),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_923),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_973),
.Y(n_1102)
);

INVx3_ASAP7_75t_SL g1103 ( 
.A(n_923),
.Y(n_1103)
);

NAND3xp33_ASAP7_75t_SL g1104 ( 
.A(n_988),
.B(n_1018),
.C(n_1009),
.Y(n_1104)
);

HB1xp67_ASAP7_75t_L g1105 ( 
.A(n_971),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_980),
.Y(n_1106)
);

NAND2x1_ASAP7_75t_L g1107 ( 
.A(n_961),
.B(n_916),
.Y(n_1107)
);

INVx2_ASAP7_75t_SL g1108 ( 
.A(n_990),
.Y(n_1108)
);

CKINVDCx11_ASAP7_75t_R g1109 ( 
.A(n_1021),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1021),
.Y(n_1110)
);

INVx3_ASAP7_75t_SL g1111 ( 
.A(n_916),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_990),
.B(n_1028),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1006),
.B(n_1021),
.Y(n_1113)
);

BUFx3_ASAP7_75t_L g1114 ( 
.A(n_1006),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1015),
.B(n_1025),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1015),
.B(n_1025),
.Y(n_1116)
);

OR2x6_ASAP7_75t_L g1117 ( 
.A(n_979),
.B(n_976),
.Y(n_1117)
);

INVx2_ASAP7_75t_SL g1118 ( 
.A(n_914),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_981),
.A2(n_943),
.B(n_975),
.C(n_956),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_958),
.B(n_914),
.Y(n_1120)
);

AND2x4_ASAP7_75t_L g1121 ( 
.A(n_936),
.B(n_1027),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_1008),
.Y(n_1122)
);

AOI221x1_ASAP7_75t_L g1123 ( 
.A1(n_1014),
.A2(n_791),
.B1(n_897),
.B2(n_1023),
.C(n_999),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_904),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_985),
.B(n_987),
.Y(n_1125)
);

INVx5_ASAP7_75t_L g1126 ( 
.A(n_925),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_912),
.Y(n_1127)
);

INVxp67_ASAP7_75t_SL g1128 ( 
.A(n_904),
.Y(n_1128)
);

AOI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_911),
.A2(n_705),
.B1(n_895),
.B2(n_897),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_911),
.B(n_982),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_1024),
.A2(n_895),
.B1(n_759),
.B2(n_791),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_912),
.Y(n_1132)
);

NAND3xp33_ASAP7_75t_L g1133 ( 
.A(n_1012),
.B(n_895),
.C(n_897),
.Y(n_1133)
);

INVxp67_ASAP7_75t_SL g1134 ( 
.A(n_904),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1023),
.B(n_1024),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_910),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_910),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_912),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_910),
.Y(n_1139)
);

OR2x2_ASAP7_75t_L g1140 ( 
.A(n_985),
.B(n_764),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_989),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_903),
.A2(n_776),
.B(n_791),
.Y(n_1142)
);

CKINVDCx11_ASAP7_75t_R g1143 ( 
.A(n_938),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_1023),
.A2(n_782),
.B(n_897),
.C(n_776),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_968),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_1023),
.B(n_776),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1023),
.B(n_1024),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_985),
.B(n_987),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_907),
.B(n_913),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_910),
.Y(n_1150)
);

INVx2_ASAP7_75t_SL g1151 ( 
.A(n_904),
.Y(n_1151)
);

CKINVDCx20_ASAP7_75t_R g1152 ( 
.A(n_968),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_911),
.B(n_982),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1023),
.A2(n_782),
.B(n_897),
.C(n_776),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_985),
.B(n_987),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_910),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_904),
.Y(n_1157)
);

BUFx6f_ASAP7_75t_L g1158 ( 
.A(n_989),
.Y(n_1158)
);

AO32x1_ASAP7_75t_L g1159 ( 
.A1(n_1024),
.A2(n_927),
.A3(n_935),
.B1(n_847),
.B2(n_785),
.Y(n_1159)
);

A2O1A1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_1023),
.A2(n_782),
.B(n_897),
.C(n_776),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_912),
.Y(n_1161)
);

OR2x2_ASAP7_75t_L g1162 ( 
.A(n_985),
.B(n_764),
.Y(n_1162)
);

INVx3_ASAP7_75t_SL g1163 ( 
.A(n_968),
.Y(n_1163)
);

NAND2x1p5_ASAP7_75t_L g1164 ( 
.A(n_1093),
.B(n_1049),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_SL g1165 ( 
.A1(n_1131),
.A2(n_1080),
.B1(n_1133),
.B2(n_1135),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1033),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1038),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_L g1168 ( 
.A1(n_1031),
.A2(n_1129),
.B1(n_1071),
.B2(n_1131),
.Y(n_1168)
);

AOI22xp33_ASAP7_75t_L g1169 ( 
.A1(n_1031),
.A2(n_1129),
.B1(n_1071),
.B2(n_1148),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_1076),
.Y(n_1170)
);

OAI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_1130),
.A2(n_1153),
.B1(n_1047),
.B2(n_1147),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1039),
.Y(n_1172)
);

CKINVDCx11_ASAP7_75t_R g1173 ( 
.A(n_1152),
.Y(n_1173)
);

OR2x2_ASAP7_75t_L g1174 ( 
.A(n_1116),
.B(n_1115),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1050),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1127),
.Y(n_1176)
);

INVx3_ASAP7_75t_L g1177 ( 
.A(n_1109),
.Y(n_1177)
);

AOI22xp33_ASAP7_75t_SL g1178 ( 
.A1(n_1080),
.A2(n_1133),
.B1(n_1147),
.B2(n_1135),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1125),
.B(n_1155),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_1042),
.A2(n_1162),
.B1(n_1140),
.B2(n_1051),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_1072),
.B(n_1149),
.Y(n_1181)
);

INVx4_ASAP7_75t_L g1182 ( 
.A(n_1101),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1132),
.Y(n_1183)
);

BUFx4f_ASAP7_75t_SL g1184 ( 
.A(n_1036),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1138),
.Y(n_1185)
);

HB1xp67_ASAP7_75t_L g1186 ( 
.A(n_1157),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1067),
.B(n_1075),
.Y(n_1187)
);

INVx2_ASAP7_75t_SL g1188 ( 
.A(n_1126),
.Y(n_1188)
);

OAI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1060),
.A2(n_1128),
.B1(n_1134),
.B2(n_1124),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_1061),
.Y(n_1190)
);

BUFx2_ASAP7_75t_L g1191 ( 
.A(n_1120),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1161),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1064),
.B(n_1065),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1102),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1046),
.Y(n_1195)
);

BUFx2_ASAP7_75t_R g1196 ( 
.A(n_1145),
.Y(n_1196)
);

INVx4_ASAP7_75t_L g1197 ( 
.A(n_1101),
.Y(n_1197)
);

OAI22xp33_ASAP7_75t_R g1198 ( 
.A1(n_1144),
.A2(n_1160),
.B1(n_1154),
.B2(n_1030),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1045),
.B(n_1055),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1068),
.Y(n_1200)
);

BUFx2_ASAP7_75t_L g1201 ( 
.A(n_1120),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1070),
.A2(n_1136),
.B1(n_1094),
.B2(n_1139),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1073),
.A2(n_1137),
.B1(n_1156),
.B2(n_1150),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1105),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1062),
.A2(n_1146),
.B1(n_1106),
.B2(n_1055),
.Y(n_1205)
);

AOI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1052),
.A2(n_1151),
.B1(n_1035),
.B2(n_1086),
.Y(n_1206)
);

CKINVDCx11_ASAP7_75t_R g1207 ( 
.A(n_1163),
.Y(n_1207)
);

BUFx2_ASAP7_75t_L g1208 ( 
.A(n_1056),
.Y(n_1208)
);

INVx2_ASAP7_75t_SL g1209 ( 
.A(n_1126),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1142),
.A2(n_1054),
.B(n_1043),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1096),
.A2(n_1083),
.B(n_1081),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1100),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1100),
.Y(n_1213)
);

OR2x2_ASAP7_75t_L g1214 ( 
.A(n_1056),
.B(n_1045),
.Y(n_1214)
);

NAND2x1p5_ASAP7_75t_L g1215 ( 
.A(n_1093),
.B(n_1049),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_1101),
.Y(n_1216)
);

INVx4_ASAP7_75t_L g1217 ( 
.A(n_1103),
.Y(n_1217)
);

INVx4_ASAP7_75t_L g1218 ( 
.A(n_1066),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1057),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1118),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1054),
.A2(n_1034),
.B1(n_1059),
.B2(n_1057),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1062),
.A2(n_1048),
.B1(n_1066),
.B2(n_1040),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1069),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1110),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_1037),
.Y(n_1225)
);

INVx3_ASAP7_75t_L g1226 ( 
.A(n_1117),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1091),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1059),
.B(n_1092),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1092),
.Y(n_1229)
);

CKINVDCx11_ASAP7_75t_R g1230 ( 
.A(n_1143),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1098),
.Y(n_1231)
);

AO21x1_ASAP7_75t_L g1232 ( 
.A1(n_1113),
.A2(n_1159),
.B(n_1121),
.Y(n_1232)
);

HB1xp67_ASAP7_75t_L g1233 ( 
.A(n_1089),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1098),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1112),
.Y(n_1235)
);

INVx4_ASAP7_75t_L g1236 ( 
.A(n_1126),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1037),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1037),
.Y(n_1238)
);

BUFx2_ASAP7_75t_L g1239 ( 
.A(n_1121),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1041),
.Y(n_1240)
);

BUFx3_ASAP7_75t_L g1241 ( 
.A(n_1041),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1141),
.Y(n_1242)
);

OA21x2_ASAP7_75t_L g1243 ( 
.A1(n_1119),
.A2(n_1034),
.B(n_1123),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1149),
.B(n_1084),
.Y(n_1244)
);

INVx4_ASAP7_75t_L g1245 ( 
.A(n_1095),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1111),
.A2(n_1032),
.B1(n_1114),
.B2(n_1088),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1048),
.A2(n_1040),
.B1(n_1082),
.B2(n_1072),
.Y(n_1247)
);

BUFx2_ASAP7_75t_L g1248 ( 
.A(n_1079),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1048),
.A2(n_1072),
.B1(n_1085),
.B2(n_1104),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1141),
.B(n_1158),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1141),
.Y(n_1251)
);

CKINVDCx11_ASAP7_75t_R g1252 ( 
.A(n_1029),
.Y(n_1252)
);

AOI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1099),
.A2(n_1107),
.B(n_1087),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1078),
.A2(n_1063),
.B1(n_1158),
.B2(n_1090),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1032),
.B(n_1097),
.Y(n_1255)
);

INVx1_ASAP7_75t_SL g1256 ( 
.A(n_1053),
.Y(n_1256)
);

AOI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1099),
.A2(n_1087),
.B(n_1058),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1108),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1074),
.A2(n_1122),
.B(n_1159),
.Y(n_1259)
);

CKINVDCx11_ASAP7_75t_R g1260 ( 
.A(n_1029),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1095),
.Y(n_1261)
);

INVx8_ASAP7_75t_L g1262 ( 
.A(n_1044),
.Y(n_1262)
);

INVx1_ASAP7_75t_SL g1263 ( 
.A(n_1159),
.Y(n_1263)
);

OAI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1129),
.A2(n_895),
.B1(n_1071),
.B2(n_776),
.Y(n_1264)
);

AO21x1_ASAP7_75t_L g1265 ( 
.A1(n_1080),
.A2(n_782),
.B(n_1131),
.Y(n_1265)
);

AO21x1_ASAP7_75t_L g1266 ( 
.A1(n_1080),
.A2(n_782),
.B(n_1131),
.Y(n_1266)
);

AND2x4_ASAP7_75t_L g1267 ( 
.A(n_1072),
.B(n_926),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1031),
.A2(n_626),
.B1(n_418),
.B2(n_422),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1077),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_SL g1270 ( 
.A1(n_1131),
.A2(n_626),
.B1(n_321),
.B2(n_333),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1064),
.B(n_1071),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1077),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1157),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1031),
.A2(n_626),
.B1(n_418),
.B2(n_422),
.Y(n_1274)
);

BUFx3_ASAP7_75t_L g1275 ( 
.A(n_1076),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1077),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1077),
.Y(n_1277)
);

INVx3_ASAP7_75t_L g1278 ( 
.A(n_1109),
.Y(n_1278)
);

BUFx2_ASAP7_75t_SL g1279 ( 
.A(n_1126),
.Y(n_1279)
);

INVxp33_ASAP7_75t_L g1280 ( 
.A(n_1125),
.Y(n_1280)
);

OAI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1129),
.A2(n_895),
.B1(n_1071),
.B2(n_776),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1031),
.A2(n_626),
.B1(n_418),
.B2(n_422),
.Y(n_1282)
);

AO21x2_ASAP7_75t_L g1283 ( 
.A1(n_1096),
.A2(n_967),
.B(n_966),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1177),
.Y(n_1284)
);

HB1xp67_ASAP7_75t_L g1285 ( 
.A(n_1208),
.Y(n_1285)
);

INVx3_ASAP7_75t_L g1286 ( 
.A(n_1259),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1271),
.B(n_1193),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1271),
.B(n_1193),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1219),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1174),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1174),
.Y(n_1291)
);

AO21x1_ASAP7_75t_SL g1292 ( 
.A1(n_1210),
.A2(n_1168),
.B(n_1169),
.Y(n_1292)
);

AND2x2_ASAP7_75t_SL g1293 ( 
.A(n_1248),
.B(n_1191),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1201),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1201),
.B(n_1214),
.Y(n_1295)
);

OR2x6_ASAP7_75t_L g1296 ( 
.A(n_1164),
.B(n_1215),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1171),
.B(n_1178),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1214),
.B(n_1228),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1190),
.B(n_1256),
.Y(n_1299)
);

BUFx4f_ASAP7_75t_L g1300 ( 
.A(n_1181),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1270),
.A2(n_1265),
.B1(n_1266),
.B2(n_1282),
.Y(n_1301)
);

INVx3_ASAP7_75t_L g1302 ( 
.A(n_1259),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1221),
.B(n_1165),
.Y(n_1303)
);

BUFx2_ASAP7_75t_L g1304 ( 
.A(n_1239),
.Y(n_1304)
);

HB1xp67_ASAP7_75t_L g1305 ( 
.A(n_1212),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1213),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1228),
.Y(n_1307)
);

NOR2x1_ASAP7_75t_R g1308 ( 
.A(n_1230),
.B(n_1207),
.Y(n_1308)
);

AND2x4_ASAP7_75t_SL g1309 ( 
.A(n_1177),
.B(n_1278),
.Y(n_1309)
);

HB1xp67_ASAP7_75t_L g1310 ( 
.A(n_1248),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1220),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1224),
.Y(n_1312)
);

BUFx2_ASAP7_75t_SL g1313 ( 
.A(n_1217),
.Y(n_1313)
);

BUFx3_ASAP7_75t_L g1314 ( 
.A(n_1278),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1239),
.B(n_1211),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1166),
.B(n_1167),
.Y(n_1316)
);

NOR2x1_ASAP7_75t_SL g1317 ( 
.A(n_1279),
.B(n_1253),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1265),
.B(n_1266),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1283),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1172),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_1278),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_1283),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1175),
.B(n_1176),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1183),
.B(n_1185),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1243),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1268),
.A2(n_1274),
.B1(n_1264),
.B2(n_1281),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1198),
.A2(n_1180),
.B1(n_1280),
.B2(n_1195),
.Y(n_1327)
);

OA21x2_ASAP7_75t_L g1328 ( 
.A1(n_1232),
.A2(n_1263),
.B(n_1194),
.Y(n_1328)
);

BUFx3_ASAP7_75t_L g1329 ( 
.A(n_1215),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1192),
.Y(n_1330)
);

INVx4_ASAP7_75t_L g1331 ( 
.A(n_1215),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1226),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1280),
.B(n_1226),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1243),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1226),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1232),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1235),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1204),
.Y(n_1338)
);

BUFx2_ASAP7_75t_SL g1339 ( 
.A(n_1217),
.Y(n_1339)
);

HB1xp67_ASAP7_75t_L g1340 ( 
.A(n_1186),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1200),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_1244),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1273),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1269),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1272),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1276),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1277),
.Y(n_1347)
);

AO21x2_ASAP7_75t_L g1348 ( 
.A1(n_1257),
.A2(n_1199),
.B(n_1258),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1198),
.A2(n_1189),
.B(n_1205),
.Y(n_1349)
);

AO21x2_ASAP7_75t_L g1350 ( 
.A1(n_1227),
.A2(n_1234),
.B(n_1231),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1229),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1181),
.B(n_1245),
.Y(n_1352)
);

OAI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1246),
.A2(n_1206),
.B(n_1187),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1179),
.B(n_1223),
.Y(n_1354)
);

INVx3_ASAP7_75t_L g1355 ( 
.A(n_1217),
.Y(n_1355)
);

OAI221xp5_ASAP7_75t_L g1356 ( 
.A1(n_1301),
.A2(n_1254),
.B1(n_1222),
.B2(n_1247),
.C(n_1249),
.Y(n_1356)
);

AND2x4_ASAP7_75t_SL g1357 ( 
.A(n_1352),
.B(n_1296),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1287),
.B(n_1233),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1340),
.Y(n_1359)
);

INVx2_ASAP7_75t_SL g1360 ( 
.A(n_1284),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1312),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1288),
.B(n_1250),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1288),
.B(n_1250),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1298),
.B(n_1237),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1307),
.B(n_1238),
.Y(n_1365)
);

INVxp67_ASAP7_75t_L g1366 ( 
.A(n_1340),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1315),
.B(n_1240),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1343),
.B(n_1170),
.Y(n_1368)
);

INVxp67_ASAP7_75t_L g1369 ( 
.A(n_1343),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1315),
.B(n_1242),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1290),
.B(n_1170),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1296),
.B(n_1331),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1290),
.B(n_1275),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1303),
.A2(n_1261),
.B1(n_1203),
.B2(n_1202),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1295),
.B(n_1251),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1305),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1295),
.B(n_1275),
.Y(n_1377)
);

INVx4_ASAP7_75t_L g1378 ( 
.A(n_1300),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1306),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1306),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1303),
.A2(n_1218),
.B1(n_1230),
.B2(n_1267),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1320),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1297),
.A2(n_1218),
.B1(n_1267),
.B2(n_1209),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1291),
.B(n_1225),
.Y(n_1384)
);

AO21x2_ASAP7_75t_L g1385 ( 
.A1(n_1325),
.A2(n_1255),
.B(n_1267),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1291),
.B(n_1225),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1320),
.Y(n_1387)
);

NOR2x1_ASAP7_75t_L g1388 ( 
.A(n_1348),
.B(n_1182),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1294),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1318),
.B(n_1241),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1286),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1293),
.B(n_1216),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1305),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1354),
.B(n_1241),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1293),
.B(n_1216),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1326),
.A2(n_1218),
.B1(n_1184),
.B2(n_1196),
.Y(n_1396)
);

OAI211xp5_ASAP7_75t_L g1397 ( 
.A1(n_1297),
.A2(n_1260),
.B(n_1252),
.C(n_1207),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1286),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1293),
.B(n_1182),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1333),
.B(n_1197),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_SL g1401 ( 
.A1(n_1349),
.A2(n_1279),
.B1(n_1236),
.B2(n_1188),
.Y(n_1401)
);

BUFx2_ASAP7_75t_L g1402 ( 
.A(n_1285),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_SL g1403 ( 
.A(n_1401),
.B(n_1349),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1362),
.B(n_1363),
.Y(n_1404)
);

NOR3xp33_ASAP7_75t_L g1405 ( 
.A(n_1396),
.B(n_1336),
.C(n_1353),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1376),
.B(n_1336),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1362),
.B(n_1285),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_SL g1408 ( 
.A1(n_1356),
.A2(n_1353),
.B1(n_1342),
.B2(n_1328),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1393),
.B(n_1359),
.Y(n_1409)
);

AND2x2_ASAP7_75t_SL g1410 ( 
.A(n_1357),
.B(n_1304),
.Y(n_1410)
);

NAND3xp33_ASAP7_75t_L g1411 ( 
.A(n_1390),
.B(n_1338),
.C(n_1322),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1366),
.B(n_1338),
.Y(n_1412)
);

AOI21xp33_ASAP7_75t_L g1413 ( 
.A1(n_1388),
.A2(n_1348),
.B(n_1328),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1369),
.B(n_1328),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1402),
.B(n_1328),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1402),
.B(n_1389),
.Y(n_1416)
);

NAND3xp33_ASAP7_75t_L g1417 ( 
.A(n_1384),
.B(n_1319),
.C(n_1322),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1389),
.B(n_1328),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1358),
.B(n_1316),
.Y(n_1419)
);

OAI21xp5_ASAP7_75t_SL g1420 ( 
.A1(n_1397),
.A2(n_1309),
.B(n_1327),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1364),
.B(n_1323),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_SL g1422 ( 
.A1(n_1357),
.A2(n_1342),
.B1(n_1329),
.B2(n_1310),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1377),
.B(n_1286),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1361),
.Y(n_1424)
);

AOI221x1_ASAP7_75t_L g1425 ( 
.A1(n_1368),
.A2(n_1335),
.B1(n_1332),
.B2(n_1299),
.C(n_1337),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1377),
.B(n_1302),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1382),
.Y(n_1427)
);

OAI221xp5_ASAP7_75t_L g1428 ( 
.A1(n_1381),
.A2(n_1345),
.B1(n_1347),
.B2(n_1346),
.C(n_1337),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1388),
.A2(n_1317),
.B(n_1319),
.Y(n_1429)
);

OAI21xp5_ASAP7_75t_SL g1430 ( 
.A1(n_1383),
.A2(n_1309),
.B(n_1308),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1379),
.B(n_1323),
.Y(n_1431)
);

OAI221xp5_ASAP7_75t_L g1432 ( 
.A1(n_1371),
.A2(n_1345),
.B1(n_1346),
.B2(n_1347),
.C(n_1330),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1375),
.B(n_1302),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1379),
.B(n_1324),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1365),
.B(n_1324),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1374),
.A2(n_1292),
.B1(n_1348),
.B2(n_1341),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1375),
.B(n_1302),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1367),
.B(n_1302),
.Y(n_1438)
);

HB1xp67_ASAP7_75t_L g1439 ( 
.A(n_1373),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1370),
.B(n_1350),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1370),
.B(n_1350),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1372),
.A2(n_1292),
.B1(n_1348),
.B2(n_1341),
.Y(n_1442)
);

NAND3xp33_ASAP7_75t_L g1443 ( 
.A(n_1386),
.B(n_1351),
.C(n_1289),
.Y(n_1443)
);

OAI221xp5_ASAP7_75t_SL g1444 ( 
.A1(n_1386),
.A2(n_1330),
.B1(n_1334),
.B2(n_1325),
.C(n_1311),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1394),
.B(n_1308),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1404),
.B(n_1391),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1424),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1414),
.B(n_1380),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1427),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1427),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1410),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1409),
.B(n_1416),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1424),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1406),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1440),
.B(n_1398),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1441),
.B(n_1433),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1414),
.B(n_1380),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1441),
.B(n_1398),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1406),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1424),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1412),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1412),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1437),
.B(n_1438),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1409),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1443),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1407),
.B(n_1400),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1443),
.Y(n_1467)
);

INVx4_ASAP7_75t_L g1468 ( 
.A(n_1410),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1415),
.B(n_1382),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1431),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1415),
.B(n_1387),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1418),
.B(n_1411),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1418),
.B(n_1411),
.Y(n_1473)
);

INVx5_ASAP7_75t_L g1474 ( 
.A(n_1438),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1425),
.B(n_1431),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1434),
.Y(n_1476)
);

AND4x1_ASAP7_75t_L g1477 ( 
.A(n_1405),
.B(n_1399),
.C(n_1395),
.D(n_1392),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1434),
.Y(n_1478)
);

CKINVDCx20_ASAP7_75t_R g1479 ( 
.A(n_1439),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1425),
.B(n_1387),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1408),
.A2(n_1385),
.B1(n_1372),
.B2(n_1344),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1416),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1432),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1423),
.B(n_1360),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1451),
.B(n_1468),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1449),
.Y(n_1486)
);

NAND2x1p5_ASAP7_75t_L g1487 ( 
.A(n_1468),
.B(n_1410),
.Y(n_1487)
);

NOR2xp33_ASAP7_75t_L g1488 ( 
.A(n_1483),
.B(n_1252),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1483),
.B(n_1260),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1451),
.B(n_1468),
.Y(n_1490)
);

NAND2x1p5_ASAP7_75t_L g1491 ( 
.A(n_1468),
.B(n_1378),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1447),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1449),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1447),
.Y(n_1494)
);

BUFx2_ASAP7_75t_L g1495 ( 
.A(n_1465),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1474),
.B(n_1423),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1450),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1450),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1461),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1474),
.B(n_1417),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1465),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1474),
.B(n_1426),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_L g1503 ( 
.A(n_1479),
.B(n_1173),
.Y(n_1503)
);

INVx2_ASAP7_75t_SL g1504 ( 
.A(n_1474),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1461),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1467),
.B(n_1435),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1462),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1447),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1467),
.B(n_1421),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_L g1510 ( 
.A(n_1477),
.B(n_1173),
.Y(n_1510)
);

NAND2x1p5_ASAP7_75t_L g1511 ( 
.A(n_1474),
.B(n_1378),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_1477),
.B(n_1445),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1462),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1464),
.B(n_1482),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1470),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1453),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1470),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1464),
.B(n_1482),
.Y(n_1518)
);

OAI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1472),
.A2(n_1403),
.B(n_1417),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1476),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1474),
.B(n_1426),
.Y(n_1521)
);

INVx1_ASAP7_75t_SL g1522 ( 
.A(n_1452),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_SL g1523 ( 
.A(n_1474),
.B(n_1422),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1452),
.B(n_1419),
.Y(n_1524)
);

INVxp33_ASAP7_75t_L g1525 ( 
.A(n_1466),
.Y(n_1525)
);

AOI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1488),
.A2(n_1481),
.B1(n_1436),
.B2(n_1475),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1516),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1519),
.A2(n_1475),
.B1(n_1473),
.B2(n_1472),
.Y(n_1528)
);

INVx3_ASAP7_75t_L g1529 ( 
.A(n_1500),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1486),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1495),
.B(n_1454),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1486),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1495),
.B(n_1454),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1485),
.B(n_1456),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1493),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1516),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1522),
.B(n_1459),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1493),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1497),
.Y(n_1539)
);

NOR2x1_ASAP7_75t_L g1540 ( 
.A(n_1510),
.B(n_1420),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1497),
.Y(n_1541)
);

NOR2x1_ASAP7_75t_L g1542 ( 
.A(n_1489),
.B(n_1420),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1498),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1516),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1492),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1498),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1492),
.Y(n_1547)
);

INVx2_ASAP7_75t_SL g1548 ( 
.A(n_1485),
.Y(n_1548)
);

NAND2x2_ASAP7_75t_L g1549 ( 
.A(n_1504),
.B(n_1314),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1501),
.Y(n_1550)
);

INVx1_ASAP7_75t_SL g1551 ( 
.A(n_1503),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1499),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1506),
.B(n_1459),
.Y(n_1553)
);

AND2x4_ASAP7_75t_SL g1554 ( 
.A(n_1490),
.B(n_1484),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1524),
.B(n_1476),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1524),
.B(n_1478),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1509),
.B(n_1478),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1514),
.B(n_1473),
.Y(n_1558)
);

A2O1A1Ixp33_ASAP7_75t_L g1559 ( 
.A1(n_1512),
.A2(n_1480),
.B(n_1523),
.C(n_1500),
.Y(n_1559)
);

INVxp67_ASAP7_75t_L g1560 ( 
.A(n_1499),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1505),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1505),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1518),
.B(n_1480),
.Y(n_1563)
);

INVx2_ASAP7_75t_SL g1564 ( 
.A(n_1490),
.Y(n_1564)
);

NAND2x1p5_ASAP7_75t_L g1565 ( 
.A(n_1500),
.B(n_1378),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1507),
.B(n_1456),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1525),
.B(n_1446),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1507),
.Y(n_1568)
);

INVxp67_ASAP7_75t_L g1569 ( 
.A(n_1551),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1554),
.B(n_1500),
.Y(n_1570)
);

INVx1_ASAP7_75t_SL g1571 ( 
.A(n_1550),
.Y(n_1571)
);

AO22x1_ASAP7_75t_L g1572 ( 
.A1(n_1542),
.A2(n_1504),
.B1(n_1521),
.B2(n_1496),
.Y(n_1572)
);

NOR2x1p5_ASAP7_75t_L g1573 ( 
.A(n_1529),
.B(n_1314),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1530),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1528),
.B(n_1513),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1527),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1554),
.B(n_1496),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1532),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1535),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1538),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1527),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1528),
.B(n_1513),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1529),
.B(n_1502),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1529),
.B(n_1502),
.Y(n_1584)
);

CKINVDCx16_ASAP7_75t_R g1585 ( 
.A(n_1540),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_L g1586 ( 
.A1(n_1526),
.A2(n_1442),
.B1(n_1413),
.B2(n_1494),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1539),
.Y(n_1587)
);

INVx1_ASAP7_75t_SL g1588 ( 
.A(n_1548),
.Y(n_1588)
);

AOI222xp33_ASAP7_75t_L g1589 ( 
.A1(n_1559),
.A2(n_1560),
.B1(n_1533),
.B2(n_1531),
.C1(n_1537),
.C2(n_1568),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1548),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1534),
.B(n_1565),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1541),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1536),
.Y(n_1593)
);

INVx1_ASAP7_75t_SL g1594 ( 
.A(n_1564),
.Y(n_1594)
);

AO21x2_ASAP7_75t_L g1595 ( 
.A1(n_1559),
.A2(n_1544),
.B(n_1536),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1560),
.Y(n_1596)
);

INVx1_ASAP7_75t_SL g1597 ( 
.A(n_1564),
.Y(n_1597)
);

INVx2_ASAP7_75t_SL g1598 ( 
.A(n_1565),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1544),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1534),
.B(n_1521),
.Y(n_1600)
);

NOR2x1_ASAP7_75t_L g1601 ( 
.A(n_1552),
.B(n_1430),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1561),
.B(n_1515),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1543),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1567),
.B(n_1487),
.Y(n_1604)
);

AOI22x1_ASAP7_75t_L g1605 ( 
.A1(n_1585),
.A2(n_1491),
.B1(n_1487),
.B2(n_1511),
.Y(n_1605)
);

AOI221x1_ASAP7_75t_L g1606 ( 
.A1(n_1575),
.A2(n_1562),
.B1(n_1546),
.B2(n_1547),
.C(n_1545),
.Y(n_1606)
);

NAND4xp25_ASAP7_75t_L g1607 ( 
.A(n_1589),
.B(n_1558),
.C(n_1563),
.D(n_1566),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1603),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1569),
.B(n_1553),
.Y(n_1609)
);

AOI322xp5_ASAP7_75t_L g1610 ( 
.A1(n_1585),
.A2(n_1547),
.A3(n_1545),
.B1(n_1456),
.B2(n_1457),
.C1(n_1448),
.C2(n_1469),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1569),
.B(n_1557),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1588),
.B(n_1555),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1603),
.Y(n_1613)
);

OAI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1601),
.A2(n_1582),
.B1(n_1575),
.B2(n_1586),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1582),
.A2(n_1595),
.B1(n_1589),
.B2(n_1601),
.Y(n_1615)
);

OAI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1596),
.A2(n_1487),
.B(n_1430),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1596),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1591),
.B(n_1556),
.Y(n_1618)
);

NAND3xp33_ASAP7_75t_L g1619 ( 
.A(n_1590),
.B(n_1517),
.C(n_1515),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1574),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1574),
.Y(n_1621)
);

AND2x4_ASAP7_75t_SL g1622 ( 
.A(n_1591),
.B(n_1484),
.Y(n_1622)
);

A2O1A1Ixp33_ASAP7_75t_L g1623 ( 
.A1(n_1604),
.A2(n_1444),
.B(n_1413),
.C(n_1457),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1588),
.B(n_1517),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1594),
.B(n_1520),
.Y(n_1625)
);

AOI221xp5_ASAP7_75t_L g1626 ( 
.A1(n_1595),
.A2(n_1448),
.B1(n_1469),
.B2(n_1471),
.C(n_1428),
.Y(n_1626)
);

AOI321xp33_ASAP7_75t_L g1627 ( 
.A1(n_1604),
.A2(n_1591),
.A3(n_1593),
.B1(n_1599),
.B2(n_1581),
.C(n_1576),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1600),
.Y(n_1628)
);

OAI21xp33_ASAP7_75t_SL g1629 ( 
.A1(n_1570),
.A2(n_1520),
.B(n_1463),
.Y(n_1629)
);

NAND2x1_ASAP7_75t_L g1630 ( 
.A(n_1570),
.B(n_1577),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1578),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1628),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1615),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1611),
.B(n_1571),
.Y(n_1634)
);

BUFx2_ASAP7_75t_L g1635 ( 
.A(n_1617),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1618),
.B(n_1594),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1622),
.B(n_1597),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1627),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1630),
.B(n_1597),
.Y(n_1639)
);

INVx1_ASAP7_75t_SL g1640 ( 
.A(n_1609),
.Y(n_1640)
);

NAND3xp33_ASAP7_75t_L g1641 ( 
.A(n_1614),
.B(n_1572),
.C(n_1578),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1616),
.B(n_1604),
.Y(n_1642)
);

INVxp67_ASAP7_75t_L g1643 ( 
.A(n_1612),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1614),
.B(n_1571),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1607),
.B(n_1602),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1606),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1607),
.B(n_1602),
.Y(n_1647)
);

INVxp67_ASAP7_75t_SL g1648 ( 
.A(n_1608),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1613),
.B(n_1572),
.Y(n_1649)
);

HB1xp67_ASAP7_75t_L g1650 ( 
.A(n_1624),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1620),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1626),
.B(n_1579),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1616),
.B(n_1600),
.Y(n_1653)
);

NAND3xp33_ASAP7_75t_L g1654 ( 
.A(n_1644),
.B(n_1623),
.C(n_1610),
.Y(n_1654)
);

OAI221xp5_ASAP7_75t_L g1655 ( 
.A1(n_1638),
.A2(n_1646),
.B1(n_1641),
.B2(n_1645),
.C(n_1647),
.Y(n_1655)
);

NAND3xp33_ASAP7_75t_SL g1656 ( 
.A(n_1638),
.B(n_1625),
.C(n_1570),
.Y(n_1656)
);

NOR2x1_ASAP7_75t_L g1657 ( 
.A(n_1646),
.B(n_1635),
.Y(n_1657)
);

AOI222xp33_ASAP7_75t_L g1658 ( 
.A1(n_1633),
.A2(n_1619),
.B1(n_1631),
.B2(n_1621),
.C1(n_1599),
.C2(n_1581),
.Y(n_1658)
);

OAI21xp5_ASAP7_75t_SL g1659 ( 
.A1(n_1645),
.A2(n_1598),
.B(n_1584),
.Y(n_1659)
);

AOI221xp5_ASAP7_75t_L g1660 ( 
.A1(n_1652),
.A2(n_1633),
.B1(n_1647),
.B2(n_1634),
.C(n_1640),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1639),
.Y(n_1661)
);

NAND4xp25_ASAP7_75t_L g1662 ( 
.A(n_1636),
.B(n_1584),
.C(n_1583),
.D(n_1577),
.Y(n_1662)
);

AOI21xp5_ASAP7_75t_L g1663 ( 
.A1(n_1649),
.A2(n_1595),
.B(n_1598),
.Y(n_1663)
);

O2A1O1Ixp33_ASAP7_75t_SL g1664 ( 
.A1(n_1643),
.A2(n_1598),
.B(n_1579),
.C(n_1587),
.Y(n_1664)
);

O2A1O1Ixp33_ASAP7_75t_L g1665 ( 
.A1(n_1648),
.A2(n_1595),
.B(n_1629),
.C(n_1580),
.Y(n_1665)
);

O2A1O1Ixp33_ASAP7_75t_L g1666 ( 
.A1(n_1635),
.A2(n_1580),
.B(n_1587),
.C(n_1592),
.Y(n_1666)
);

AND5x1_ASAP7_75t_L g1667 ( 
.A(n_1660),
.B(n_1653),
.C(n_1642),
.D(n_1639),
.E(n_1650),
.Y(n_1667)
);

NOR2xp67_ASAP7_75t_L g1668 ( 
.A(n_1662),
.B(n_1632),
.Y(n_1668)
);

NOR3x1_ASAP7_75t_L g1669 ( 
.A(n_1656),
.B(n_1651),
.C(n_1592),
.Y(n_1669)
);

NAND3x1_ASAP7_75t_SL g1670 ( 
.A(n_1657),
.B(n_1642),
.C(n_1653),
.Y(n_1670)
);

NOR3xp33_ASAP7_75t_L g1671 ( 
.A(n_1655),
.B(n_1632),
.C(n_1637),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_SL g1672 ( 
.A(n_1661),
.B(n_1637),
.Y(n_1672)
);

OA22x2_ASAP7_75t_SL g1673 ( 
.A1(n_1659),
.A2(n_1605),
.B1(n_1573),
.B2(n_1584),
.Y(n_1673)
);

OAI21xp33_ASAP7_75t_L g1674 ( 
.A1(n_1654),
.A2(n_1658),
.B(n_1663),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1666),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1664),
.Y(n_1676)
);

NAND4xp25_ASAP7_75t_L g1677 ( 
.A(n_1669),
.B(n_1665),
.C(n_1583),
.D(n_1577),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1668),
.B(n_1600),
.Y(n_1678)
);

NAND4xp25_ASAP7_75t_SL g1679 ( 
.A(n_1671),
.B(n_1583),
.C(n_1262),
.D(n_1593),
.Y(n_1679)
);

AOI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1674),
.A2(n_1581),
.B(n_1576),
.Y(n_1680)
);

NOR3xp33_ASAP7_75t_L g1681 ( 
.A(n_1670),
.B(n_1593),
.C(n_1576),
.Y(n_1681)
);

NOR3xp33_ASAP7_75t_L g1682 ( 
.A(n_1675),
.B(n_1599),
.C(n_1262),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1678),
.Y(n_1683)
);

AOI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1681),
.A2(n_1672),
.B1(n_1676),
.B2(n_1667),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1680),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1682),
.B(n_1573),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_SL g1687 ( 
.A(n_1679),
.B(n_1673),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_SL g1688 ( 
.A(n_1677),
.B(n_1262),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1678),
.Y(n_1689)
);

AOI21xp5_ASAP7_75t_L g1690 ( 
.A1(n_1687),
.A2(n_1262),
.B(n_1471),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1685),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1684),
.B(n_1463),
.Y(n_1692)
);

OR3x1_ASAP7_75t_L g1693 ( 
.A(n_1683),
.B(n_1549),
.C(n_1491),
.Y(n_1693)
);

NAND3xp33_ASAP7_75t_L g1694 ( 
.A(n_1689),
.B(n_1508),
.C(n_1494),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_R g1695 ( 
.A(n_1686),
.B(n_1355),
.Y(n_1695)
);

XNOR2xp5_ASAP7_75t_L g1696 ( 
.A(n_1692),
.B(n_1688),
.Y(n_1696)
);

XOR2x1_ASAP7_75t_L g1697 ( 
.A(n_1691),
.B(n_1491),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1694),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1698),
.Y(n_1699)
);

NAND5xp2_ASAP7_75t_L g1700 ( 
.A(n_1699),
.B(n_1690),
.C(n_1697),
.D(n_1696),
.E(n_1695),
.Y(n_1700)
);

AOI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1700),
.A2(n_1693),
.B1(n_1549),
.B2(n_1508),
.Y(n_1701)
);

AOI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1700),
.A2(n_1460),
.B1(n_1453),
.B2(n_1511),
.Y(n_1702)
);

OR2x6_ASAP7_75t_L g1703 ( 
.A(n_1701),
.B(n_1702),
.Y(n_1703)
);

INVxp33_ASAP7_75t_SL g1704 ( 
.A(n_1701),
.Y(n_1704)
);

OAI21xp33_ASAP7_75t_L g1705 ( 
.A1(n_1704),
.A2(n_1511),
.B(n_1309),
.Y(n_1705)
);

OR2x6_ASAP7_75t_L g1706 ( 
.A(n_1703),
.B(n_1313),
.Y(n_1706)
);

AOI222xp33_ASAP7_75t_L g1707 ( 
.A1(n_1705),
.A2(n_1460),
.B1(n_1453),
.B2(n_1354),
.C1(n_1458),
.C2(n_1455),
.Y(n_1707)
);

AOI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1707),
.A2(n_1706),
.B1(n_1313),
.B2(n_1339),
.Y(n_1708)
);

AOI221xp5_ASAP7_75t_L g1709 ( 
.A1(n_1708),
.A2(n_1339),
.B1(n_1429),
.B2(n_1458),
.C(n_1455),
.Y(n_1709)
);

AOI211xp5_ASAP7_75t_L g1710 ( 
.A1(n_1709),
.A2(n_1321),
.B(n_1314),
.C(n_1355),
.Y(n_1710)
);


endmodule