module fake_jpeg_9646_n_341 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_37),
.B(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_36),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_32),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_44),
.Y(n_52)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_0),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_23),
.Y(n_49)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_23),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_50),
.B(n_57),
.Y(n_95)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_44),
.B(n_28),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_46),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_63),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_30),
.Y(n_63)
);

AO22x1_ASAP7_75t_SL g66 ( 
.A1(n_40),
.A2(n_19),
.B1(n_35),
.B2(n_33),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_66),
.A2(n_41),
.B1(n_39),
.B2(n_42),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_30),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_21),
.Y(n_74)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_72),
.B(n_84),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_44),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_77),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_74),
.B(n_75),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_26),
.Y(n_75)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g125 ( 
.A(n_76),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_52),
.Y(n_77)
);

NAND2xp33_ASAP7_75t_SL g113 ( 
.A(n_78),
.B(n_94),
.Y(n_113)
);

CKINVDCx9p33_ASAP7_75t_R g79 ( 
.A(n_66),
.Y(n_79)
);

INVxp67_ASAP7_75t_SL g110 ( 
.A(n_79),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_66),
.A2(n_17),
.B1(n_47),
.B2(n_41),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_42),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_86),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_83),
.B1(n_56),
.B2(n_57),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_52),
.B1(n_43),
.B2(n_56),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

CKINVDCx12_ASAP7_75t_R g85 ( 
.A(n_51),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_43),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_91),
.Y(n_124)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_65),
.Y(n_93)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_26),
.Y(n_94)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_65),
.Y(n_97)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_56),
.A2(n_17),
.B1(n_31),
.B2(n_24),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_98),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_122)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_58),
.B(n_21),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_31),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_107),
.B1(n_122),
.B2(n_73),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_46),
.C(n_40),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_45),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_79),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_129),
.Y(n_137)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_88),
.A2(n_45),
.B1(n_48),
.B2(n_39),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_112),
.A2(n_76),
.B1(n_87),
.B2(n_99),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_126),
.B(n_94),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_78),
.A2(n_34),
.B1(n_25),
.B2(n_27),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_128),
.A2(n_70),
.B1(n_28),
.B2(n_34),
.Y(n_144)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_130),
.A2(n_135),
.B1(n_39),
.B2(n_101),
.Y(n_161)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_132),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_126),
.Y(n_132)
);

OAI21xp33_ASAP7_75t_L g133 ( 
.A1(n_110),
.A2(n_78),
.B(n_95),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_133),
.A2(n_128),
.B(n_122),
.Y(n_173)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_136),
.B(n_138),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_125),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_86),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_139),
.A2(n_147),
.B(n_158),
.Y(n_188)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_141),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_127),
.Y(n_141)
);

BUFx12_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_142),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_143),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_144),
.A2(n_132),
.B1(n_141),
.B2(n_115),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_112),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_146),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_104),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_106),
.B(n_75),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_149),
.Y(n_163)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_106),
.B(n_92),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_159),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_111),
.B(n_69),
.Y(n_152)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_152),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_104),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_153),
.Y(n_160)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_155),
.Y(n_162)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_102),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_156),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_129),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_157),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_115),
.A2(n_29),
.B(n_89),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_103),
.B(n_91),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_161),
.A2(n_39),
.B1(n_58),
.B2(n_64),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_189),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_103),
.C(n_111),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_180),
.C(n_181),
.Y(n_206)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_175),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_173),
.A2(n_185),
.B(n_29),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_113),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_174),
.A2(n_48),
.B(n_45),
.Y(n_224)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_159),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_184),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_135),
.A2(n_109),
.B1(n_112),
.B2(n_124),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_178),
.A2(n_147),
.B1(n_154),
.B2(n_90),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_139),
.B(n_121),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_144),
.A2(n_120),
.B1(n_71),
.B2(n_114),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_182),
.A2(n_193),
.B1(n_58),
.B2(n_156),
.Y(n_203)
);

XNOR2x1_ASAP7_75t_SL g183 ( 
.A(n_139),
.B(n_45),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_45),
.Y(n_207)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_138),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_158),
.A2(n_123),
.B(n_121),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_146),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_148),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_35),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_151),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_168),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_131),
.A2(n_71),
.B1(n_123),
.B2(n_116),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_167),
.B(n_69),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_194),
.B(n_196),
.Y(n_243)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_176),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_162),
.A2(n_140),
.B1(n_136),
.B2(n_134),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_197),
.A2(n_211),
.B1(n_217),
.B2(n_222),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_198),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_155),
.Y(n_199)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_199),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_134),
.Y(n_200)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_179),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_202),
.B(n_210),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_203),
.A2(n_214),
.B(n_220),
.Y(n_239)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_208),
.Y(n_237)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_212),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_207),
.B(n_224),
.Y(n_232)
);

INVx13_ASAP7_75t_L g208 ( 
.A(n_168),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_166),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_172),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_183),
.A2(n_163),
.B1(n_177),
.B2(n_165),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_213),
.A2(n_169),
.B1(n_186),
.B2(n_160),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_193),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_215),
.B(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_163),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_169),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_178),
.A2(n_154),
.B1(n_91),
.B2(n_61),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_170),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_185),
.C(n_171),
.Y(n_236)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_174),
.A2(n_173),
.B(n_188),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_190),
.A2(n_61),
.B1(n_22),
.B2(n_18),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_142),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_223),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_180),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_228),
.B(n_236),
.C(n_45),
.Y(n_262)
);

XNOR2x1_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_188),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_231),
.B(n_235),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_216),
.A2(n_175),
.B1(n_184),
.B2(n_182),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_233),
.A2(n_195),
.B1(n_205),
.B2(n_212),
.Y(n_251)
);

XNOR2x1_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_174),
.Y(n_235)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_240),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_209),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_244),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_242),
.B(n_33),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_209),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_201),
.B(n_35),
.Y(n_245)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_245),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_201),
.B(n_35),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_249),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_33),
.Y(n_249)
);

HAxp5_ASAP7_75t_L g250 ( 
.A(n_211),
.B(n_142),
.CON(n_250),
.SN(n_250)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_250),
.A2(n_214),
.B(n_208),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_251),
.A2(n_254),
.B1(n_266),
.B2(n_269),
.Y(n_274)
);

MAJx2_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_206),
.C(n_218),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_256),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_250),
.A2(n_203),
.B1(n_196),
.B2(n_204),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_250),
.A2(n_217),
.B1(n_222),
.B2(n_224),
.Y(n_255)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_255),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_207),
.Y(n_256)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_243),
.Y(n_258)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_258),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_252),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_227),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_264),
.B(n_265),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_64),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_225),
.A2(n_33),
.B1(n_22),
.B2(n_2),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_225),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_234),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_268),
.A2(n_240),
.B1(n_246),
.B2(n_245),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_242),
.A2(n_22),
.B1(n_36),
.B2(n_2),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_234),
.B(n_0),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_271),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_229),
.B(n_230),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_236),
.C(n_226),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_277),
.C(n_278),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_275),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_282),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_231),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_239),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_239),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_287),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_233),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_286),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_267),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_259),
.B(n_226),
.C(n_232),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_288),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_251),
.B(n_249),
.Y(n_289)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_289),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_273),
.A2(n_263),
.B1(n_266),
.B2(n_260),
.Y(n_290)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_290),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_284),
.A2(n_247),
.B1(n_248),
.B2(n_261),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_301),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_261),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_298),
.Y(n_306)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_281),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_302),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_283),
.A2(n_252),
.B1(n_253),
.B2(n_232),
.Y(n_301)
);

INVx11_ASAP7_75t_L g302 ( 
.A(n_276),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_274),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_303),
.A2(n_280),
.B(n_2),
.Y(n_310)
);

AO221x1_ASAP7_75t_L g304 ( 
.A1(n_288),
.A2(n_48),
.B1(n_22),
.B2(n_3),
.C(n_5),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_304),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_299),
.B(n_272),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_305),
.B(n_307),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_295),
.B(n_277),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_285),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_309),
.B(n_297),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_310),
.A2(n_313),
.B(n_304),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_300),
.A2(n_280),
.B(n_3),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_302),
.A2(n_36),
.B1(n_5),
.B2(n_6),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_316),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_303),
.A2(n_1),
.B1(n_6),
.B2(n_7),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_312),
.A2(n_294),
.B(n_295),
.Y(n_317)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_317),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_312),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_319),
.Y(n_331)
);

FAx1_ASAP7_75t_SL g320 ( 
.A(n_314),
.B(n_298),
.CI(n_291),
.CON(n_320),
.SN(n_320)
);

AOI31xp67_ASAP7_75t_L g326 ( 
.A1(n_320),
.A2(n_325),
.A3(n_311),
.B(n_6),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_321),
.A2(n_1),
.B1(n_8),
.B2(n_9),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_308),
.A2(n_292),
.B(n_293),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_324),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_297),
.C(n_290),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_326),
.B(n_327),
.Y(n_332)
);

AOI21x1_ASAP7_75t_L g328 ( 
.A1(n_319),
.A2(n_8),
.B(n_9),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_318),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_331),
.B(n_320),
.Y(n_333)
);

O2A1O1Ixp33_ASAP7_75t_SL g335 ( 
.A1(n_333),
.A2(n_334),
.B(n_326),
.C(n_329),
.Y(n_335)
);

AOI322xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_330),
.A3(n_332),
.B1(n_322),
.B2(n_15),
.C1(n_10),
.C2(n_14),
.Y(n_336)
);

AO21x1_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_322),
.B(n_12),
.Y(n_337)
);

AOI322xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_10),
.A3(n_12),
.B1(n_14),
.B2(n_15),
.C1(n_16),
.C2(n_48),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_16),
.B(n_48),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_16),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_48),
.Y(n_341)
);


endmodule