module fake_jpeg_247_n_44 (n_3, n_2, n_1, n_0, n_4, n_5, n_44);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_4),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

AND2x2_ASAP7_75t_SL g9 ( 
.A(n_2),
.B(n_0),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

OAI22xp33_ASAP7_75t_SL g15 ( 
.A1(n_12),
.A2(n_3),
.B1(n_5),
.B2(n_2),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_15),
.A2(n_7),
.B1(n_6),
.B2(n_11),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g16 ( 
.A(n_13),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_16),
.A2(n_17),
.B1(n_18),
.B2(n_20),
.Y(n_23)
);

CKINVDCx12_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

OR2x2_ASAP7_75t_SL g19 ( 
.A(n_9),
.B(n_12),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_SL g25 ( 
.A(n_19),
.B(n_9),
.Y(n_25)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_19),
.B(n_9),
.C(n_8),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_24),
.C(n_25),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_8),
.B(n_9),
.Y(n_24)
);

AO21x2_ASAP7_75t_L g27 ( 
.A1(n_26),
.A2(n_16),
.B(n_6),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_30),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_24),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_17),
.C(n_18),
.Y(n_30)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_28),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_35),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_23),
.B(n_26),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_32),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_39),
.B1(n_11),
.B2(n_14),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_36),
.A2(n_33),
.B1(n_7),
.B2(n_22),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_5),
.B(n_1),
.Y(n_40)
);

AOI322xp5_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_41),
.A3(n_14),
.B1(n_39),
.B2(n_2),
.C1(n_0),
.C2(n_1),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_0),
.C(n_1),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_0),
.B(n_1),
.Y(n_44)
);


endmodule