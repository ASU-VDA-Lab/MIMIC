module real_aes_2810_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_357;
wire n_287;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_456;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
INVx1_ASAP7_75t_L g174 ( .A(n_0), .Y(n_174) );
AOI22xp33_ASAP7_75t_L g165 ( .A1(n_1), .A2(n_43), .B1(n_166), .B2(n_168), .Y(n_165) );
AO22x2_ASAP7_75t_L g106 ( .A1(n_2), .A2(n_54), .B1(n_96), .B2(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_3), .B(n_225), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_4), .B(n_251), .Y(n_263) );
INVx1_ASAP7_75t_L g197 ( .A(n_5), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g89 ( .A(n_6), .B(n_90), .Y(n_89) );
AOI22xp5_ASAP7_75t_L g175 ( .A1(n_7), .A2(n_176), .B1(n_177), .B2(n_183), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_7), .Y(n_176) );
AO22x2_ASAP7_75t_L g103 ( .A1(n_8), .A2(n_18), .B1(n_96), .B2(n_104), .Y(n_103) );
AND2x2_ASAP7_75t_L g254 ( .A(n_9), .B(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g265 ( .A(n_10), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g214 ( .A(n_11), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_12), .B(n_251), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g157 ( .A1(n_13), .A2(n_69), .B1(n_158), .B2(n_161), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_14), .B(n_225), .Y(n_305) );
AOI22xp5_ASAP7_75t_L g149 ( .A1(n_15), .A2(n_72), .B1(n_150), .B2(n_153), .Y(n_149) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_16), .A2(n_71), .B1(n_218), .B2(n_225), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g121 ( .A1(n_17), .A2(n_30), .B1(n_122), .B2(n_127), .Y(n_121) );
OAI221xp5_ASAP7_75t_L g189 ( .A1(n_18), .A2(n_54), .B1(n_58), .B2(n_190), .C(n_192), .Y(n_189) );
OR2x2_ASAP7_75t_L g215 ( .A(n_19), .B(n_70), .Y(n_215) );
OA21x2_ASAP7_75t_L g244 ( .A1(n_19), .A2(n_70), .B(n_214), .Y(n_244) );
INVx3_ASAP7_75t_L g96 ( .A(n_20), .Y(n_96) );
AO21x2_ASAP7_75t_L g315 ( .A1(n_21), .A2(n_255), .B(n_316), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_22), .A2(n_233), .B(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_23), .B(n_251), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_23), .A2(n_86), .B1(n_172), .B2(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_23), .Y(n_522) );
INVx1_ASAP7_75t_SL g97 ( .A(n_24), .Y(n_97) );
AOI22xp5_ASAP7_75t_SL g142 ( .A1(n_25), .A2(n_62), .B1(n_143), .B2(n_146), .Y(n_142) );
INVx1_ASAP7_75t_L g199 ( .A(n_26), .Y(n_199) );
AND2x2_ASAP7_75t_L g223 ( .A(n_26), .B(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g231 ( .A(n_26), .B(n_197), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_27), .B(n_225), .Y(n_264) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_28), .A2(n_86), .B1(n_172), .B2(n_530), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_28), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_29), .B(n_251), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_31), .B(n_225), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_32), .A2(n_233), .B(n_247), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_33), .A2(n_36), .B1(n_180), .B2(n_181), .Y(n_179) );
INVx1_ASAP7_75t_L g181 ( .A(n_33), .Y(n_181) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_34), .A2(n_58), .B1(n_96), .B2(n_100), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_35), .B(n_249), .Y(n_277) );
INVx1_ASAP7_75t_L g180 ( .A(n_36), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g317 ( .A(n_37), .B(n_225), .Y(n_317) );
INVx1_ASAP7_75t_L g221 ( .A(n_38), .Y(n_221) );
INVx1_ASAP7_75t_L g228 ( .A(n_38), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_39), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g285 ( .A(n_40), .B(n_212), .Y(n_285) );
INVx1_ASAP7_75t_L g98 ( .A(n_41), .Y(n_98) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_42), .B(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_44), .B(n_249), .Y(n_299) );
INVx1_ASAP7_75t_L g539 ( .A(n_44), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_45), .B(n_225), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g131 ( .A1(n_46), .A2(n_53), .B1(n_132), .B2(n_138), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_47), .B(n_225), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_48), .A2(n_233), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g311 ( .A(n_49), .B(n_213), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_50), .B(n_249), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_51), .B(n_249), .Y(n_321) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_52), .A2(n_73), .B1(n_233), .B2(n_235), .Y(n_232) );
INVxp33_ASAP7_75t_L g194 ( .A(n_54), .Y(n_194) );
INVx1_ASAP7_75t_L g84 ( .A(n_55), .Y(n_84) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_55), .B(n_251), .Y(n_308) );
INVx1_ASAP7_75t_L g224 ( .A(n_56), .Y(n_224) );
INVx1_ASAP7_75t_L g230 ( .A(n_56), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_57), .B(n_249), .Y(n_262) );
INVxp67_ASAP7_75t_L g193 ( .A(n_58), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g108 ( .A1(n_59), .A2(n_67), .B1(n_109), .B2(n_115), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_60), .A2(n_233), .B(n_289), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_61), .A2(n_233), .B(n_275), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_63), .A2(n_233), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g302 ( .A(n_64), .B(n_213), .Y(n_302) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_65), .B(n_212), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_66), .A2(n_178), .B1(n_179), .B2(n_182), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_66), .Y(n_178) );
AND2x2_ASAP7_75t_L g278 ( .A(n_68), .B(n_266), .Y(n_278) );
OAI22xp5_ASAP7_75t_L g82 ( .A1(n_73), .A2(n_83), .B1(n_84), .B2(n_85), .Y(n_82) );
INVx1_ASAP7_75t_L g85 ( .A(n_73), .Y(n_85) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_74), .A2(n_233), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_75), .B(n_251), .Y(n_276) );
BUFx2_ASAP7_75t_L g310 ( .A(n_76), .Y(n_310) );
BUFx2_ASAP7_75t_SL g191 ( .A(n_77), .Y(n_191) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_186), .B1(n_200), .B2(n_517), .C(n_520), .Y(n_78) );
XOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_173), .Y(n_79) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_81), .A2(n_82), .B1(n_86), .B2(n_172), .Y(n_80) );
CKINVDCx16_ASAP7_75t_R g81 ( .A(n_82), .Y(n_81) );
INVx1_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
CKINVDCx16_ASAP7_75t_R g172 ( .A(n_86), .Y(n_172) );
HB1xp67_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
NOR2x1_ASAP7_75t_L g87 ( .A(n_88), .B(n_141), .Y(n_87) );
NAND4xp25_ASAP7_75t_L g88 ( .A(n_89), .B(n_108), .C(n_121), .D(n_131), .Y(n_88) );
INVx3_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx6_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
AND2x2_ASAP7_75t_L g92 ( .A(n_93), .B(n_101), .Y(n_92) );
AND2x4_ASAP7_75t_L g117 ( .A(n_93), .B(n_118), .Y(n_117) );
AND2x4_ASAP7_75t_L g155 ( .A(n_93), .B(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_L g93 ( .A(n_94), .B(n_99), .Y(n_93) );
INVx2_ASAP7_75t_L g114 ( .A(n_94), .Y(n_114) );
AND2x2_ASAP7_75t_L g130 ( .A(n_94), .B(n_125), .Y(n_130) );
HB1xp67_ASAP7_75t_L g164 ( .A(n_94), .Y(n_164) );
OAI22x1_ASAP7_75t_L g94 ( .A1(n_95), .A2(n_96), .B1(n_97), .B2(n_98), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
INVx1_ASAP7_75t_L g100 ( .A(n_96), .Y(n_100) );
INVx2_ASAP7_75t_L g104 ( .A(n_96), .Y(n_104) );
INVx1_ASAP7_75t_L g107 ( .A(n_96), .Y(n_107) );
AND2x2_ASAP7_75t_L g113 ( .A(n_99), .B(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g125 ( .A(n_99), .Y(n_125) );
BUFx2_ASAP7_75t_L g140 ( .A(n_99), .Y(n_140) );
AND2x4_ASAP7_75t_L g129 ( .A(n_101), .B(n_130), .Y(n_129) );
AND2x4_ASAP7_75t_L g148 ( .A(n_101), .B(n_124), .Y(n_148) );
AND2x2_ASAP7_75t_L g167 ( .A(n_101), .B(n_113), .Y(n_167) );
AND2x4_ASAP7_75t_L g101 ( .A(n_102), .B(n_105), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x4_ASAP7_75t_L g112 ( .A(n_103), .B(n_105), .Y(n_112) );
INVx1_ASAP7_75t_L g120 ( .A(n_103), .Y(n_120) );
AND2x2_ASAP7_75t_L g126 ( .A(n_103), .B(n_106), .Y(n_126) );
INVxp67_ASAP7_75t_L g156 ( .A(n_105), .Y(n_156) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_L g137 ( .A(n_106), .B(n_120), .Y(n_137) );
BUFx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
AND2x4_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
AND2x2_ASAP7_75t_L g160 ( .A(n_112), .B(n_130), .Y(n_160) );
AND2x4_ASAP7_75t_L g171 ( .A(n_112), .B(n_124), .Y(n_171) );
AND2x2_ASAP7_75t_L g136 ( .A(n_113), .B(n_137), .Y(n_136) );
AND2x4_ASAP7_75t_L g124 ( .A(n_114), .B(n_125), .Y(n_124) );
BUFx6f_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
BUFx3_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_SL g122 ( .A(n_123), .Y(n_122) );
AND2x4_ASAP7_75t_L g123 ( .A(n_124), .B(n_126), .Y(n_123) );
AND2x4_ASAP7_75t_L g145 ( .A(n_124), .B(n_137), .Y(n_145) );
AND2x4_ASAP7_75t_L g139 ( .A(n_126), .B(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g163 ( .A(n_126), .B(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx6_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g152 ( .A(n_130), .B(n_137), .Y(n_152) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
NAND4xp25_ASAP7_75t_L g141 ( .A(n_142), .B(n_149), .C(n_157), .D(n_165), .Y(n_141) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx8_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx8_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx6f_ASAP7_75t_SL g150 ( .A(n_151), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx6_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
BUFx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
BUFx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
BUFx12f_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
BUFx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
HB1xp67_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B1(n_184), .B2(n_185), .Y(n_173) );
INVx1_ASAP7_75t_L g184 ( .A(n_174), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_175), .Y(n_185) );
CKINVDCx16_ASAP7_75t_R g183 ( .A(n_177), .Y(n_183) );
INVx1_ASAP7_75t_L g182 ( .A(n_179), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_187), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g187 ( .A(n_188), .Y(n_187) );
AND3x1_ASAP7_75t_SL g188 ( .A(n_189), .B(n_195), .C(n_198), .Y(n_188) );
INVxp67_ASAP7_75t_L g528 ( .A(n_189), .Y(n_528) );
CKINVDCx8_ASAP7_75t_R g190 ( .A(n_191), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_193), .B(n_194), .Y(n_192) );
CKINVDCx16_ASAP7_75t_R g526 ( .A(n_195), .Y(n_526) );
AOI21xp33_ASAP7_75t_L g535 ( .A1(n_195), .A2(n_536), .B(n_537), .Y(n_535) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g219 ( .A(n_196), .B(n_220), .Y(n_219) );
OR2x2_ASAP7_75t_SL g533 ( .A(n_196), .B(n_198), .Y(n_533) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g234 ( .A(n_197), .B(n_221), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_198), .B(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NOR2x1p5_ASAP7_75t_L g236 ( .A(n_199), .B(n_237), .Y(n_236) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
OR2x6_ASAP7_75t_L g201 ( .A(n_202), .B(n_454), .Y(n_201) );
NAND3xp33_ASAP7_75t_L g202 ( .A(n_203), .B(n_370), .C(n_407), .Y(n_202) );
NOR3xp33_ASAP7_75t_L g203 ( .A(n_204), .B(n_338), .C(n_353), .Y(n_203) );
OAI221xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_282), .B1(n_312), .B2(n_324), .C(n_325), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_207), .B(n_267), .Y(n_206) );
OAI22xp33_ASAP7_75t_SL g398 ( .A1(n_207), .A2(n_362), .B1(n_399), .B2(n_402), .Y(n_398) );
OR2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_239), .Y(n_207) );
OAI21xp33_ASAP7_75t_SL g408 ( .A1(n_208), .A2(n_409), .B(n_415), .Y(n_408) );
OR2x2_ASAP7_75t_L g437 ( .A(n_208), .B(n_269), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_208), .B(n_357), .Y(n_438) );
INVx2_ASAP7_75t_L g469 ( .A(n_208), .Y(n_469) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_209), .B(n_329), .Y(n_450) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
OR2x2_ASAP7_75t_L g324 ( .A(n_210), .B(n_242), .Y(n_324) );
BUFx3_ASAP7_75t_L g350 ( .A(n_210), .Y(n_350) );
AND2x2_ASAP7_75t_L g486 ( .A(n_210), .B(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g509 ( .A(n_210), .B(n_270), .Y(n_509) );
AND2x4_ASAP7_75t_L g210 ( .A(n_211), .B(n_216), .Y(n_210) );
AND2x4_ASAP7_75t_L g281 ( .A(n_211), .B(n_216), .Y(n_281) );
AO21x2_ASAP7_75t_L g216 ( .A1(n_212), .A2(n_217), .B(n_232), .Y(n_216) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_212), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_212), .A2(n_273), .B(n_274), .Y(n_272) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_SL g213 ( .A(n_214), .B(n_215), .Y(n_213) );
AND2x4_ASAP7_75t_L g292 ( .A(n_214), .B(n_215), .Y(n_292) );
INVx1_ASAP7_75t_L g519 ( .A(n_218), .Y(n_519) );
AND2x4_ASAP7_75t_L g218 ( .A(n_219), .B(n_222), .Y(n_218) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_220), .Y(n_536) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AND2x4_ASAP7_75t_L g251 ( .A(n_221), .B(n_229), .Y(n_251) );
INVx1_ASAP7_75t_L g538 ( .A(n_222), .Y(n_538) );
BUFx3_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x6_ASAP7_75t_L g233 ( .A(n_223), .B(n_234), .Y(n_233) );
INVx2_ASAP7_75t_L g238 ( .A(n_224), .Y(n_238) );
AND2x6_ASAP7_75t_L g249 ( .A(n_224), .B(n_227), .Y(n_249) );
AND2x4_ASAP7_75t_L g225 ( .A(n_226), .B(n_231), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_227), .B(n_229), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx5_ASAP7_75t_L g252 ( .A(n_231), .Y(n_252) );
AND2x4_ASAP7_75t_L g235 ( .A(n_234), .B(n_236), .Y(n_235) );
INVx3_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_SL g239 ( .A(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_240), .B(n_270), .Y(n_429) );
INVx1_ASAP7_75t_L g466 ( .A(n_240), .Y(n_466) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_256), .Y(n_240) );
AND2x2_ASAP7_75t_L g280 ( .A(n_241), .B(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g487 ( .A(n_241), .Y(n_487) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g330 ( .A(n_242), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_242), .B(n_256), .Y(n_331) );
AND2x2_ASAP7_75t_L g352 ( .A(n_242), .B(n_271), .Y(n_352) );
AND2x2_ASAP7_75t_L g434 ( .A(n_242), .B(n_257), .Y(n_434) );
AO21x2_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_245), .B(n_254), .Y(n_242) );
INVx4_ASAP7_75t_L g255 ( .A(n_243), .Y(n_255) );
INVx3_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
BUFx4f_ASAP7_75t_L g266 ( .A(n_244), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_253), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_250), .B(n_252), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_249), .B(n_310), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_252), .A2(n_262), .B(n_263), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_252), .A2(n_276), .B(n_277), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_252), .A2(n_290), .B(n_291), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g298 ( .A1(n_252), .A2(n_299), .B(n_300), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_252), .A2(n_308), .B(n_309), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g319 ( .A1(n_252), .A2(n_320), .B(n_321), .Y(n_319) );
INVx3_ASAP7_75t_L g295 ( .A(n_255), .Y(n_295) );
AND2x4_ASAP7_75t_SL g327 ( .A(n_256), .B(n_271), .Y(n_327) );
INVx1_ASAP7_75t_L g358 ( .A(n_256), .Y(n_358) );
INVx2_ASAP7_75t_L g366 ( .A(n_256), .Y(n_366) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_256), .Y(n_390) );
INVx3_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_257), .Y(n_279) );
AOI21x1_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_259), .B(n_265), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_264), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_266), .A2(n_305), .B(n_306), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_280), .Y(n_267) );
AND2x2_ASAP7_75t_L g505 ( .A(n_268), .B(n_368), .Y(n_505) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_279), .Y(n_269) );
NAND2x1p5_ASAP7_75t_L g364 ( .A(n_270), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g416 ( .A(n_270), .B(n_331), .Y(n_416) );
AND2x2_ASAP7_75t_L g433 ( .A(n_270), .B(n_434), .Y(n_433) );
INVx4_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x4_ASAP7_75t_L g357 ( .A(n_271), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g373 ( .A(n_271), .Y(n_373) );
AND2x2_ASAP7_75t_L g417 ( .A(n_271), .B(n_418), .Y(n_417) );
OR2x2_ASAP7_75t_L g424 ( .A(n_271), .B(n_425), .Y(n_424) );
NOR2x1_ASAP7_75t_L g439 ( .A(n_271), .B(n_330), .Y(n_439) );
BUFx2_ASAP7_75t_L g449 ( .A(n_271), .Y(n_449) );
AND2x2_ASAP7_75t_L g474 ( .A(n_271), .B(n_434), .Y(n_474) );
AND2x2_ASAP7_75t_L g495 ( .A(n_271), .B(n_496), .Y(n_495) );
OR2x6_ASAP7_75t_L g271 ( .A(n_272), .B(n_278), .Y(n_271) );
INVx1_ASAP7_75t_L g426 ( .A(n_279), .Y(n_426) );
NAND2xp5_ASAP7_75t_SL g372 ( .A(n_280), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g456 ( .A(n_280), .B(n_327), .Y(n_456) );
INVx3_ASAP7_75t_L g363 ( .A(n_281), .Y(n_363) );
AND2x2_ASAP7_75t_L g496 ( .A(n_281), .B(n_418), .Y(n_496) );
INVx1_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
AOI22xp5_ASAP7_75t_L g325 ( .A1(n_283), .A2(n_326), .B1(n_331), .B2(n_332), .Y(n_325) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_293), .Y(n_283) );
INVx4_ASAP7_75t_L g323 ( .A(n_284), .Y(n_323) );
INVx2_ASAP7_75t_L g360 ( .A(n_284), .Y(n_360) );
NAND2x1_ASAP7_75t_L g386 ( .A(n_284), .B(n_303), .Y(n_386) );
OR2x2_ASAP7_75t_L g401 ( .A(n_284), .B(n_336), .Y(n_401) );
OR2x2_ASAP7_75t_SL g428 ( .A(n_284), .B(n_400), .Y(n_428) );
AND2x2_ASAP7_75t_L g441 ( .A(n_284), .B(n_315), .Y(n_441) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_284), .Y(n_462) );
OR2x6_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
AOI21xp5_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_288), .B(n_292), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_292), .A2(n_317), .B(n_318), .Y(n_316) );
INVx2_ASAP7_75t_L g341 ( .A(n_293), .Y(n_341) );
AND2x2_ASAP7_75t_L g473 ( .A(n_293), .B(n_447), .Y(n_473) );
NOR2x1_ASAP7_75t_SL g293 ( .A(n_294), .B(n_303), .Y(n_293) );
AND2x2_ASAP7_75t_L g314 ( .A(n_294), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g490 ( .A(n_294), .B(n_413), .Y(n_490) );
AO21x1_ASAP7_75t_SL g294 ( .A1(n_295), .A2(n_296), .B(n_302), .Y(n_294) );
AO21x2_ASAP7_75t_L g337 ( .A1(n_295), .A2(n_296), .B(n_302), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_301), .Y(n_296) );
OR2x2_ASAP7_75t_L g322 ( .A(n_303), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g333 ( .A(n_303), .B(n_323), .Y(n_333) );
AND2x2_ASAP7_75t_L g379 ( .A(n_303), .B(n_336), .Y(n_379) );
OR2x2_ASAP7_75t_L g400 ( .A(n_303), .B(n_315), .Y(n_400) );
INVx2_ASAP7_75t_SL g406 ( .A(n_303), .Y(n_406) );
AND2x2_ASAP7_75t_L g412 ( .A(n_303), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g422 ( .A(n_303), .B(n_405), .Y(n_422) );
BUFx2_ASAP7_75t_L g444 ( .A(n_303), .Y(n_444) );
OR2x6_ASAP7_75t_L g303 ( .A(n_304), .B(n_311), .Y(n_303) );
INVx2_ASAP7_75t_L g491 ( .A(n_312), .Y(n_491) );
OR2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_322), .Y(n_312) );
OR2x2_ASAP7_75t_L g516 ( .A(n_313), .B(n_360), .Y(n_516) );
INVx2_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_314), .B(n_323), .Y(n_382) );
AND2x2_ASAP7_75t_L g453 ( .A(n_314), .B(n_333), .Y(n_453) );
INVx1_ASAP7_75t_L g335 ( .A(n_315), .Y(n_335) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_315), .Y(n_344) );
INVx1_ASAP7_75t_L g377 ( .A(n_315), .Y(n_377) );
INVx2_ASAP7_75t_L g413 ( .A(n_315), .Y(n_413) );
NOR2xp67_ASAP7_75t_L g343 ( .A(n_323), .B(n_344), .Y(n_343) );
BUFx2_ASAP7_75t_L g403 ( .A(n_323), .Y(n_403) );
INVx2_ASAP7_75t_SL g479 ( .A(n_324), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_326), .A2(n_381), .B1(n_383), .B2(n_387), .Y(n_380) );
AND2x2_ASAP7_75t_SL g326 ( .A(n_327), .B(n_328), .Y(n_326) );
AND2x2_ASAP7_75t_L g507 ( .A(n_327), .B(n_363), .Y(n_507) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_329), .B(n_373), .Y(n_452) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g418 ( .A(n_330), .B(n_366), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_331), .B(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g361 ( .A(n_332), .Y(n_361) );
AOI221xp5_ASAP7_75t_L g475 ( .A1(n_332), .A2(n_476), .B1(n_480), .B2(n_482), .C(n_484), .Y(n_475) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
AND2x2_ASAP7_75t_L g345 ( .A(n_333), .B(n_346), .Y(n_345) );
INVxp67_ASAP7_75t_SL g369 ( .A(n_333), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_333), .B(n_376), .Y(n_431) );
INVx1_ASAP7_75t_SL g427 ( .A(n_334), .Y(n_427) );
AOI221xp5_ASAP7_75t_SL g455 ( .A1(n_334), .A2(n_345), .B1(n_456), .B2(n_457), .C(n_460), .Y(n_455) );
AOI322xp5_ASAP7_75t_L g488 ( .A1(n_334), .A2(n_406), .A3(n_433), .B1(n_489), .B2(n_491), .C1(n_492), .C2(n_495), .Y(n_488) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
BUFx2_ASAP7_75t_L g355 ( .A(n_335), .Y(n_355) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_336), .Y(n_347) );
INVx2_ASAP7_75t_L g405 ( .A(n_336), .Y(n_405) );
AND2x2_ASAP7_75t_L g446 ( .A(n_336), .B(n_447), .Y(n_446) );
INVx3_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OA21x2_ASAP7_75t_SL g338 ( .A1(n_339), .A2(n_345), .B(n_348), .Y(n_338) );
AOI211xp5_ASAP7_75t_L g508 ( .A1(n_339), .A2(n_509), .B(n_510), .C(n_514), .Y(n_508) );
INVx1_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
OR2x2_ASAP7_75t_L g397 ( .A(n_341), .B(n_359), .Y(n_397) );
OR2x2_ASAP7_75t_L g481 ( .A(n_341), .B(n_376), .Y(n_481) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g421 ( .A(n_343), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g499 ( .A(n_346), .Y(n_499) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g385 ( .A(n_347), .Y(n_385) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
OR2x2_ASAP7_75t_L g354 ( .A(n_350), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g389 ( .A(n_352), .B(n_390), .Y(n_389) );
OAI322xp33_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_356), .A3(n_359), .B1(n_361), .B2(n_362), .C1(n_367), .C2(n_369), .Y(n_353) );
INVx1_ASAP7_75t_L g395 ( .A(n_354), .Y(n_395) );
OR2x2_ASAP7_75t_L g367 ( .A(n_356), .B(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_356), .B(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g378 ( .A(n_360), .B(n_379), .Y(n_378) );
OAI32xp33_ASAP7_75t_L g423 ( .A1(n_360), .A2(n_424), .A3(n_427), .B1(n_428), .B2(n_429), .Y(n_423) );
OR2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
INVx2_ASAP7_75t_L g368 ( .A(n_363), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_363), .B(n_426), .Y(n_425) );
NOR2x1_ASAP7_75t_L g465 ( .A(n_363), .B(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g489 ( .A(n_363), .B(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g410 ( .A(n_364), .Y(n_410) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_368), .B(n_434), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_371), .B(n_391), .Y(n_370) );
OAI21xp33_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_374), .B(n_380), .Y(n_371) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x4_ASAP7_75t_SL g375 ( .A(n_376), .B(n_378), .Y(n_375) );
INVx3_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g440 ( .A(n_379), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g503 ( .A1(n_382), .A2(n_402), .B1(n_504), .B2(n_506), .Y(n_503) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
A2O1A1Ixp33_ASAP7_75t_L g430 ( .A1(n_384), .A2(n_431), .B(n_432), .C(n_435), .Y(n_430) );
OR2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
INVx3_ASAP7_75t_L g512 ( .A(n_386), .Y(n_512) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g393 ( .A(n_390), .Y(n_393) );
AO21x1_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_394), .B(n_398), .Y(n_391) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g458 ( .A(n_393), .Y(n_458) );
AND2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_399), .B(n_485), .Y(n_484) );
OR2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_401), .Y(n_399) );
INVx1_ASAP7_75t_L g414 ( .A(n_401), .Y(n_414) );
OR2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVx1_ASAP7_75t_L g471 ( .A(n_404), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
NOR3xp33_ASAP7_75t_L g407 ( .A(n_408), .B(n_430), .C(n_442), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
OAI21xp5_ASAP7_75t_SL g472 ( .A1(n_411), .A2(n_473), .B(n_474), .Y(n_472) );
AND2x4_ASAP7_75t_L g411 ( .A(n_412), .B(n_414), .Y(n_411) );
INVx1_ASAP7_75t_L g447 ( .A(n_413), .Y(n_447) );
O2A1O1Ixp5_ASAP7_75t_SL g415 ( .A1(n_416), .A2(n_417), .B(n_419), .C(n_423), .Y(n_415) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_425), .Y(n_515) );
INVx2_ASAP7_75t_L g500 ( .A(n_428), .Y(n_500) );
AOI21xp33_ASAP7_75t_L g514 ( .A1(n_429), .A2(n_515), .B(n_516), .Y(n_514) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g494 ( .A(n_434), .Y(n_494) );
OAI31xp33_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_438), .A3(n_439), .B(n_440), .Y(n_435) );
INVx1_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g513 ( .A(n_441), .Y(n_513) );
OAI21xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_448), .B(n_451), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
BUFx2_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g463 ( .A(n_446), .Y(n_463) );
AOI21xp33_ASAP7_75t_SL g510 ( .A1(n_448), .A2(n_511), .B(n_513), .Y(n_510) );
OR2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
INVx2_ASAP7_75t_L g478 ( .A(n_449), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_449), .B(n_469), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_449), .B(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g459 ( .A(n_450), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
NAND5xp2_ASAP7_75t_L g454 ( .A(n_455), .B(n_475), .C(n_488), .D(n_497), .E(n_508), .Y(n_454) );
AND2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
OAI221xp5_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_464), .B1(n_467), .B2(n_470), .C(n_472), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVxp67_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVxp67_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_501), .B(n_503), .Y(n_497) );
AND2x4_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
INVx1_ASAP7_75t_SL g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
INVxp67_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_518), .Y(n_517) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
OAI222xp33_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_523), .B1(n_529), .B2(n_531), .C1(n_534), .C2(n_539), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_524), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_525), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
INVxp67_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
endmodule