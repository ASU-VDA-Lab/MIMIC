module real_aes_8993_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_182;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_502;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_741;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_359;
wire n_156;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g109 ( .A(n_0), .Y(n_109) );
A2O1A1Ixp33_ASAP7_75t_L g245 ( .A1(n_1), .A2(n_163), .B(n_166), .C(n_246), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_2), .A2(n_192), .B(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g493 ( .A(n_3), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_4), .B(n_222), .Y(n_221) );
AOI21xp33_ASAP7_75t_L g476 ( .A1(n_5), .A2(n_192), .B(n_477), .Y(n_476) );
AND2x6_ASAP7_75t_L g163 ( .A(n_6), .B(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g259 ( .A(n_7), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_8), .B(n_115), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_8), .B(n_42), .Y(n_128) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_9), .A2(n_191), .B(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_10), .B(n_175), .Y(n_248) );
INVx1_ASAP7_75t_L g481 ( .A(n_11), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_12), .B(n_216), .Y(n_516) );
INVx1_ASAP7_75t_L g155 ( .A(n_13), .Y(n_155) );
INVx1_ASAP7_75t_L g528 ( .A(n_14), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g135 ( .A1(n_15), .A2(n_79), .B1(n_136), .B2(n_137), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_15), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g280 ( .A1(n_16), .A2(n_200), .B(n_281), .C(n_283), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_17), .B(n_222), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_18), .B(n_459), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_19), .B(n_192), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_20), .B(n_206), .Y(n_205) );
A2O1A1Ixp33_ASAP7_75t_L g266 ( .A1(n_21), .A2(n_216), .B(n_267), .C(n_269), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_22), .B(n_222), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_23), .B(n_175), .Y(n_174) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_24), .A2(n_202), .B(n_283), .C(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_25), .B(n_175), .Y(n_230) );
CKINVDCx16_ASAP7_75t_R g157 ( .A(n_26), .Y(n_157) );
INVx1_ASAP7_75t_L g229 ( .A(n_27), .Y(n_229) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_28), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g244 ( .A(n_29), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_30), .B(n_175), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_31), .A2(n_104), .B1(n_116), .B2(n_747), .Y(n_103) );
INVx1_ASAP7_75t_L g198 ( .A(n_32), .Y(n_198) );
INVx1_ASAP7_75t_L g471 ( .A(n_33), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g132 ( .A1(n_34), .A2(n_133), .B1(n_134), .B2(n_135), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_34), .Y(n_133) );
INVx2_ASAP7_75t_L g161 ( .A(n_35), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g250 ( .A(n_36), .Y(n_250) );
A2O1A1Ixp33_ASAP7_75t_L g215 ( .A1(n_37), .A2(n_216), .B(n_217), .C(n_219), .Y(n_215) );
INVxp67_ASAP7_75t_L g201 ( .A(n_38), .Y(n_201) );
CKINVDCx14_ASAP7_75t_R g214 ( .A(n_39), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_40), .A2(n_166), .B(n_228), .C(n_232), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g503 ( .A1(n_41), .A2(n_163), .B(n_166), .C(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g115 ( .A(n_42), .Y(n_115) );
INVx1_ASAP7_75t_L g470 ( .A(n_43), .Y(n_470) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_44), .A2(n_177), .B(n_257), .C(n_258), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_45), .B(n_175), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g234 ( .A(n_46), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_47), .Y(n_194) );
INVx1_ASAP7_75t_L g265 ( .A(n_48), .Y(n_265) );
CKINVDCx16_ASAP7_75t_R g472 ( .A(n_49), .Y(n_472) );
OAI22xp5_ASAP7_75t_SL g741 ( .A1(n_50), .A2(n_59), .B1(n_742), .B2(n_743), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_50), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_51), .B(n_192), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g468 ( .A1(n_52), .A2(n_166), .B1(n_269), .B2(n_469), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_53), .Y(n_508) );
CKINVDCx16_ASAP7_75t_R g490 ( .A(n_54), .Y(n_490) );
CKINVDCx14_ASAP7_75t_R g255 ( .A(n_55), .Y(n_255) );
A2O1A1Ixp33_ASAP7_75t_L g479 ( .A1(n_56), .A2(n_219), .B(n_257), .C(n_480), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_57), .Y(n_540) );
INVx1_ASAP7_75t_L g478 ( .A(n_58), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_59), .Y(n_743) );
INVx1_ASAP7_75t_L g164 ( .A(n_60), .Y(n_164) );
INVx1_ASAP7_75t_L g154 ( .A(n_61), .Y(n_154) );
INVx1_ASAP7_75t_SL g218 ( .A(n_62), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_63), .Y(n_122) );
OAI22xp5_ASAP7_75t_SL g740 ( .A1(n_64), .A2(n_741), .B1(n_744), .B2(n_745), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_64), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_65), .B(n_222), .Y(n_271) );
INVx1_ASAP7_75t_L g170 ( .A(n_66), .Y(n_170) );
AOI222xp33_ASAP7_75t_SL g130 ( .A1(n_67), .A2(n_131), .B1(n_132), .B2(n_138), .C1(n_732), .C2(n_734), .Y(n_130) );
A2O1A1Ixp33_ASAP7_75t_SL g458 ( .A1(n_68), .A2(n_219), .B(n_459), .C(n_460), .Y(n_458) );
INVxp67_ASAP7_75t_L g461 ( .A(n_69), .Y(n_461) );
INVx1_ASAP7_75t_L g112 ( .A(n_70), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_71), .A2(n_192), .B(n_254), .Y(n_253) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_72), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_73), .A2(n_192), .B(n_278), .Y(n_277) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_74), .Y(n_474) );
INVx1_ASAP7_75t_L g534 ( .A(n_75), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_76), .A2(n_191), .B(n_193), .Y(n_190) );
CKINVDCx16_ASAP7_75t_R g226 ( .A(n_77), .Y(n_226) );
INVx1_ASAP7_75t_L g279 ( .A(n_78), .Y(n_279) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_79), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_80), .A2(n_163), .B(n_166), .C(n_536), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_81), .A2(n_192), .B(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g282 ( .A(n_82), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_83), .B(n_199), .Y(n_505) );
INVx2_ASAP7_75t_L g152 ( .A(n_84), .Y(n_152) );
INVx1_ASAP7_75t_L g247 ( .A(n_85), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_86), .B(n_459), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_87), .A2(n_163), .B(n_166), .C(n_492), .Y(n_491) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_88), .B(n_109), .C(n_110), .Y(n_108) );
OR2x2_ASAP7_75t_L g125 ( .A(n_88), .B(n_126), .Y(n_125) );
OR2x2_ASAP7_75t_L g445 ( .A(n_88), .B(n_127), .Y(n_445) );
INVx2_ASAP7_75t_L g731 ( .A(n_88), .Y(n_731) );
A2O1A1Ixp33_ASAP7_75t_L g165 ( .A1(n_89), .A2(n_166), .B(n_169), .C(n_179), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_90), .B(n_184), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_91), .Y(n_497) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_92), .A2(n_163), .B(n_166), .C(n_514), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_93), .Y(n_520) );
INVx1_ASAP7_75t_L g457 ( .A(n_94), .Y(n_457) );
CKINVDCx16_ASAP7_75t_R g525 ( .A(n_95), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_96), .B(n_199), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_97), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_98), .B(n_150), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_99), .B(n_150), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_100), .B(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g268 ( .A(n_101), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_102), .A2(n_192), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_SL g749 ( .A(n_106), .Y(n_749) );
AND2x2_ASAP7_75t_SL g106 ( .A(n_107), .B(n_113), .Y(n_106) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g127 ( .A(n_109), .B(n_128), .Y(n_127) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
INVxp67_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AOI22xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_130), .B1(n_737), .B2(n_738), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g118 ( .A(n_119), .B(n_123), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_SL g737 ( .A(n_121), .Y(n_737) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AOI21xp5_ASAP7_75t_L g738 ( .A1(n_123), .A2(n_739), .B(n_746), .Y(n_738) );
NOR2xp33_ASAP7_75t_SL g123 ( .A(n_124), .B(n_129), .Y(n_123) );
HB1xp67_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_125), .Y(n_746) );
NOR2x2_ASAP7_75t_L g736 ( .A(n_126), .B(n_731), .Y(n_736) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OR2x2_ASAP7_75t_L g730 ( .A(n_127), .B(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OAI22xp5_ASAP7_75t_SL g138 ( .A1(n_139), .A2(n_445), .B1(n_446), .B2(n_728), .Y(n_138) );
INVx2_ASAP7_75t_L g733 ( .A(n_139), .Y(n_733) );
XOR2xp5_ASAP7_75t_L g739 ( .A(n_139), .B(n_740), .Y(n_739) );
OR2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_379), .Y(n_139) );
NAND5xp2_ASAP7_75t_L g140 ( .A(n_141), .B(n_308), .C(n_338), .D(n_359), .E(n_365), .Y(n_140) );
AOI221xp5_ASAP7_75t_SL g141 ( .A1(n_142), .A2(n_238), .B1(n_272), .B2(n_274), .C(n_285), .Y(n_141) );
INVxp67_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_144), .B(n_235), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g144 ( .A(n_145), .B(n_207), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
A2O1A1Ixp33_ASAP7_75t_SL g359 ( .A1(n_146), .A2(n_223), .B(n_360), .C(n_363), .Y(n_359) );
AND2x2_ASAP7_75t_L g429 ( .A(n_146), .B(n_224), .Y(n_429) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_185), .Y(n_146) );
AND2x2_ASAP7_75t_L g287 ( .A(n_147), .B(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g291 ( .A(n_147), .B(n_288), .Y(n_291) );
OR2x2_ASAP7_75t_L g317 ( .A(n_147), .B(n_224), .Y(n_317) );
AND2x2_ASAP7_75t_L g319 ( .A(n_147), .B(n_210), .Y(n_319) );
AND2x2_ASAP7_75t_L g337 ( .A(n_147), .B(n_209), .Y(n_337) );
INVx1_ASAP7_75t_L g370 ( .A(n_147), .Y(n_370) );
INVx2_ASAP7_75t_SL g147 ( .A(n_148), .Y(n_147) );
BUFx2_ASAP7_75t_L g237 ( .A(n_148), .Y(n_237) );
AND2x2_ASAP7_75t_L g273 ( .A(n_148), .B(n_210), .Y(n_273) );
AND2x2_ASAP7_75t_L g426 ( .A(n_148), .B(n_224), .Y(n_426) );
AO21x2_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_156), .B(n_181), .Y(n_148) );
INVx3_ASAP7_75t_L g222 ( .A(n_149), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_149), .B(n_234), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_149), .B(n_250), .Y(n_249) );
NOR2xp33_ASAP7_75t_SL g507 ( .A(n_149), .B(n_508), .Y(n_507) );
INVx4_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
HB1xp67_ASAP7_75t_L g211 ( .A(n_150), .Y(n_211) );
OA21x2_ASAP7_75t_L g454 ( .A1(n_150), .A2(n_455), .B(n_462), .Y(n_454) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g188 ( .A(n_151), .Y(n_188) );
AND2x2_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
AND2x2_ASAP7_75t_SL g184 ( .A(n_152), .B(n_153), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
OAI21xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_158), .B(n_165), .Y(n_156) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_158), .A2(n_184), .B(n_226), .C(n_227), .Y(n_225) );
OAI21xp5_ASAP7_75t_L g243 ( .A1(n_158), .A2(n_244), .B(n_245), .Y(n_243) );
OAI22xp33_ASAP7_75t_L g467 ( .A1(n_158), .A2(n_180), .B1(n_468), .B2(n_472), .Y(n_467) );
OAI21xp5_ASAP7_75t_L g489 ( .A1(n_158), .A2(n_490), .B(n_491), .Y(n_489) );
OAI21xp5_ASAP7_75t_L g533 ( .A1(n_158), .A2(n_534), .B(n_535), .Y(n_533) );
NAND2x1p5_ASAP7_75t_L g158 ( .A(n_159), .B(n_163), .Y(n_158) );
AND2x4_ASAP7_75t_L g192 ( .A(n_159), .B(n_163), .Y(n_192) );
AND2x2_ASAP7_75t_L g159 ( .A(n_160), .B(n_162), .Y(n_159) );
INVx1_ASAP7_75t_L g203 ( .A(n_160), .Y(n_203) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g167 ( .A(n_161), .Y(n_167) );
INVx1_ASAP7_75t_L g270 ( .A(n_161), .Y(n_270) );
INVx1_ASAP7_75t_L g168 ( .A(n_162), .Y(n_168) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_162), .Y(n_173) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_162), .Y(n_175) );
INVx3_ASAP7_75t_L g200 ( .A(n_162), .Y(n_200) );
INVx1_ASAP7_75t_L g459 ( .A(n_162), .Y(n_459) );
INVx4_ASAP7_75t_SL g180 ( .A(n_163), .Y(n_180) );
BUFx3_ASAP7_75t_L g232 ( .A(n_163), .Y(n_232) );
INVx5_ASAP7_75t_L g195 ( .A(n_166), .Y(n_195) );
AND2x6_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
BUFx3_ASAP7_75t_L g178 ( .A(n_167), .Y(n_178) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_167), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_174), .C(n_176), .Y(n_169) );
O2A1O1Ixp5_ASAP7_75t_L g246 ( .A1(n_171), .A2(n_176), .B(n_247), .C(n_248), .Y(n_246) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
OAI22xp5_ASAP7_75t_SL g469 ( .A1(n_172), .A2(n_173), .B1(n_470), .B2(n_471), .Y(n_469) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx4_ASAP7_75t_L g202 ( .A(n_173), .Y(n_202) );
INVx4_ASAP7_75t_L g216 ( .A(n_175), .Y(n_216) );
INVx2_ASAP7_75t_L g257 ( .A(n_175), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_176), .A2(n_505), .B(n_506), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_176), .A2(n_537), .B(n_538), .Y(n_536) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g283 ( .A(n_178), .Y(n_283) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
O2A1O1Ixp33_ASAP7_75t_SL g193 ( .A1(n_180), .A2(n_194), .B(n_195), .C(n_196), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_L g213 ( .A1(n_180), .A2(n_195), .B(n_214), .C(n_215), .Y(n_213) );
O2A1O1Ixp33_ASAP7_75t_SL g254 ( .A1(n_180), .A2(n_195), .B(n_255), .C(n_256), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_SL g264 ( .A1(n_180), .A2(n_195), .B(n_265), .C(n_266), .Y(n_264) );
O2A1O1Ixp33_ASAP7_75t_SL g278 ( .A1(n_180), .A2(n_195), .B(n_279), .C(n_280), .Y(n_278) );
O2A1O1Ixp33_ASAP7_75t_L g456 ( .A1(n_180), .A2(n_195), .B(n_457), .C(n_458), .Y(n_456) );
O2A1O1Ixp33_ASAP7_75t_L g477 ( .A1(n_180), .A2(n_195), .B(n_478), .C(n_479), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_L g524 ( .A1(n_180), .A2(n_195), .B(n_525), .C(n_526), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_182), .B(n_183), .Y(n_181) );
INVx1_ASAP7_75t_L g206 ( .A(n_183), .Y(n_206) );
AO21x2_ASAP7_75t_L g511 ( .A1(n_183), .A2(n_512), .B(n_519), .Y(n_511) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g242 ( .A(n_184), .Y(n_242) );
OA21x2_ASAP7_75t_L g252 ( .A1(n_184), .A2(n_253), .B(n_260), .Y(n_252) );
OA21x2_ASAP7_75t_L g522 ( .A1(n_184), .A2(n_523), .B(n_529), .Y(n_522) );
AND2x2_ASAP7_75t_L g307 ( .A(n_185), .B(n_208), .Y(n_307) );
OR2x2_ASAP7_75t_L g311 ( .A(n_185), .B(n_224), .Y(n_311) );
AND2x2_ASAP7_75t_L g336 ( .A(n_185), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_SL g383 ( .A(n_185), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_185), .B(n_345), .Y(n_431) );
AO21x2_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_189), .B(n_204), .Y(n_185) );
INVx1_ASAP7_75t_L g289 ( .A(n_186), .Y(n_289) );
AO21x2_ASAP7_75t_L g532 ( .A1(n_186), .A2(n_533), .B(n_539), .Y(n_532) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AOI21xp5_ASAP7_75t_SL g501 ( .A1(n_187), .A2(n_502), .B(n_503), .Y(n_501) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AO21x2_ASAP7_75t_L g466 ( .A1(n_188), .A2(n_467), .B(n_473), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_188), .B(n_474), .Y(n_473) );
AO21x2_ASAP7_75t_L g488 ( .A1(n_188), .A2(n_489), .B(n_496), .Y(n_488) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
OA21x2_ASAP7_75t_L g288 ( .A1(n_190), .A2(n_205), .B(n_289), .Y(n_288) );
BUFx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_197), .B(n_203), .Y(n_196) );
OAI22xp33_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B1(n_201), .B2(n_202), .Y(n_197) );
O2A1O1Ixp33_ASAP7_75t_L g228 ( .A1(n_199), .A2(n_229), .B(n_230), .C(n_231), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_L g492 ( .A1(n_199), .A2(n_493), .B(n_494), .C(n_495), .Y(n_492) );
INVx5_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_200), .B(n_259), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_200), .B(n_461), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_200), .B(n_481), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_202), .B(n_268), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_202), .B(n_282), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_202), .B(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g231 ( .A(n_203), .Y(n_231) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
OAI322xp33_ASAP7_75t_L g432 ( .A1(n_207), .A2(n_368), .A3(n_391), .B1(n_412), .B2(n_433), .C1(n_435), .C2(n_436), .Y(n_432) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_208), .B(n_288), .Y(n_435) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_223), .Y(n_208) );
AND2x2_ASAP7_75t_L g236 ( .A(n_209), .B(n_237), .Y(n_236) );
AND2x4_ASAP7_75t_L g304 ( .A(n_209), .B(n_224), .Y(n_304) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g345 ( .A(n_210), .B(n_224), .Y(n_345) );
AND2x2_ASAP7_75t_L g389 ( .A(n_210), .B(n_223), .Y(n_389) );
OA21x2_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_221), .Y(n_210) );
OA21x2_ASAP7_75t_L g262 ( .A1(n_211), .A2(n_263), .B(n_271), .Y(n_262) );
OA21x2_ASAP7_75t_L g276 ( .A1(n_211), .A2(n_277), .B(n_284), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_216), .B(n_218), .Y(n_217) );
INVx3_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_220), .Y(n_517) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_222), .A2(n_476), .B(n_482), .Y(n_475) );
AND2x2_ASAP7_75t_L g272 ( .A(n_223), .B(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g290 ( .A(n_223), .B(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_223), .B(n_319), .Y(n_443) );
INVx3_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g235 ( .A(n_224), .B(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_224), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g357 ( .A(n_224), .B(n_288), .Y(n_357) );
AND2x2_ASAP7_75t_L g384 ( .A(n_224), .B(n_319), .Y(n_384) );
OR2x2_ASAP7_75t_L g440 ( .A(n_224), .B(n_291), .Y(n_440) );
OR2x6_ASAP7_75t_L g224 ( .A(n_225), .B(n_233), .Y(n_224) );
INVx1_ASAP7_75t_SL g326 ( .A(n_235), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_236), .B(n_357), .Y(n_358) );
AND2x2_ASAP7_75t_L g392 ( .A(n_236), .B(n_382), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_236), .B(n_315), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_236), .B(n_437), .Y(n_436) );
OAI31xp33_ASAP7_75t_L g410 ( .A1(n_238), .A2(n_272), .A3(n_411), .B(n_413), .Y(n_410) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_251), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g377 ( .A(n_239), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g393 ( .A(n_239), .B(n_328), .Y(n_393) );
OR2x2_ASAP7_75t_L g400 ( .A(n_239), .B(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g412 ( .A(n_239), .B(n_301), .Y(n_412) );
CKINVDCx16_ASAP7_75t_R g239 ( .A(n_240), .Y(n_239) );
OR2x2_ASAP7_75t_L g346 ( .A(n_240), .B(n_347), .Y(n_346) );
BUFx3_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g274 ( .A(n_241), .B(n_275), .Y(n_274) );
INVx4_ASAP7_75t_L g295 ( .A(n_241), .Y(n_295) );
AND2x2_ASAP7_75t_L g332 ( .A(n_241), .B(n_276), .Y(n_332) );
AO21x2_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_243), .B(n_249), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_242), .B(n_497), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_242), .B(n_520), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_242), .B(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g331 ( .A(n_251), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_SL g401 ( .A(n_251), .Y(n_401) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_261), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_252), .B(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g301 ( .A(n_252), .B(n_262), .Y(n_301) );
INVx2_ASAP7_75t_L g321 ( .A(n_252), .Y(n_321) );
AND2x2_ASAP7_75t_L g335 ( .A(n_252), .B(n_262), .Y(n_335) );
AND2x2_ASAP7_75t_L g342 ( .A(n_252), .B(n_298), .Y(n_342) );
BUFx3_ASAP7_75t_L g352 ( .A(n_252), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_252), .B(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g297 ( .A(n_261), .Y(n_297) );
AND2x2_ASAP7_75t_L g305 ( .A(n_261), .B(n_295), .Y(n_305) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g275 ( .A(n_262), .B(n_276), .Y(n_275) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_262), .Y(n_329) );
INVx2_ASAP7_75t_L g495 ( .A(n_269), .Y(n_495) );
INVx3_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx2_ASAP7_75t_SL g312 ( .A(n_273), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_273), .B(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_273), .B(n_382), .Y(n_403) );
NAND2xp5_ASAP7_75t_SL g405 ( .A(n_274), .B(n_352), .Y(n_405) );
INVx1_ASAP7_75t_SL g439 ( .A(n_274), .Y(n_439) );
INVx1_ASAP7_75t_SL g347 ( .A(n_275), .Y(n_347) );
INVx1_ASAP7_75t_SL g298 ( .A(n_276), .Y(n_298) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_276), .Y(n_309) );
OR2x2_ASAP7_75t_L g320 ( .A(n_276), .B(n_295), .Y(n_320) );
AND2x2_ASAP7_75t_L g334 ( .A(n_276), .B(n_295), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_276), .B(n_324), .Y(n_386) );
A2O1A1Ixp33_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_290), .B(n_292), .C(n_303), .Y(n_285) );
AOI31xp33_ASAP7_75t_L g402 ( .A1(n_286), .A2(n_403), .A3(n_404), .B(n_405), .Y(n_402) );
AND2x2_ASAP7_75t_L g375 ( .A(n_287), .B(n_304), .Y(n_375) );
BUFx3_ASAP7_75t_L g315 ( .A(n_288), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_288), .B(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g351 ( .A(n_288), .B(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_288), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_SL g306 ( .A(n_291), .Y(n_306) );
OAI222xp33_ASAP7_75t_L g415 ( .A1(n_291), .A2(n_416), .B1(n_419), .B2(n_420), .C1(n_421), .C2(n_422), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_293), .B(n_299), .Y(n_292) );
INVx1_ASAP7_75t_L g421 ( .A(n_293), .Y(n_421) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_296), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_295), .B(n_298), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_295), .B(n_321), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_295), .B(n_296), .Y(n_391) );
INVx1_ASAP7_75t_L g442 ( .A(n_295), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g372 ( .A(n_296), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g444 ( .A(n_296), .Y(n_444) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
INVx2_ASAP7_75t_L g324 ( .A(n_297), .Y(n_324) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_298), .Y(n_367) );
AOI32xp33_ASAP7_75t_L g303 ( .A1(n_299), .A2(n_304), .A3(n_305), .B1(n_306), .B2(n_307), .Y(n_303) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_301), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g378 ( .A(n_301), .Y(n_378) );
OR2x2_ASAP7_75t_L g419 ( .A(n_301), .B(n_320), .Y(n_419) );
INVx1_ASAP7_75t_L g355 ( .A(n_302), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_304), .B(n_315), .Y(n_340) );
INVx3_ASAP7_75t_L g349 ( .A(n_304), .Y(n_349) );
AOI322xp5_ASAP7_75t_L g365 ( .A1(n_304), .A2(n_349), .A3(n_366), .B1(n_368), .B2(n_371), .C1(n_375), .C2(n_376), .Y(n_365) );
AND2x2_ASAP7_75t_L g341 ( .A(n_305), .B(n_342), .Y(n_341) );
INVxp67_ASAP7_75t_L g418 ( .A(n_305), .Y(n_418) );
A2O1A1O1Ixp25_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_310), .B(n_313), .C(n_321), .D(n_322), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_309), .B(n_352), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
OAI221xp5_ASAP7_75t_L g322 ( .A1(n_311), .A2(n_323), .B1(n_326), .B2(n_327), .C(n_330), .Y(n_322) );
INVx1_ASAP7_75t_SL g437 ( .A(n_311), .Y(n_437) );
AOI21xp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_318), .B(n_320), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g425 ( .A(n_315), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OAI221xp5_ASAP7_75t_SL g407 ( .A1(n_317), .A2(n_401), .B1(n_408), .B2(n_409), .C(n_410), .Y(n_407) );
OAI222xp33_ASAP7_75t_L g438 ( .A1(n_318), .A2(n_439), .B1(n_440), .B2(n_441), .C1(n_443), .C2(n_444), .Y(n_438) );
AND2x2_ASAP7_75t_L g396 ( .A(n_319), .B(n_382), .Y(n_396) );
AOI21xp5_ASAP7_75t_L g408 ( .A1(n_319), .A2(n_334), .B(n_381), .Y(n_408) );
INVx1_ASAP7_75t_L g422 ( .A(n_319), .Y(n_422) );
INVx2_ASAP7_75t_SL g325 ( .A(n_320), .Y(n_325) );
AND2x2_ASAP7_75t_L g328 ( .A(n_321), .B(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx1_ASAP7_75t_SL g362 ( .A(n_324), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_324), .B(n_334), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_325), .B(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_325), .B(n_335), .Y(n_364) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OAI21xp5_ASAP7_75t_SL g330 ( .A1(n_331), .A2(n_333), .B(n_336), .Y(n_330) );
INVx1_ASAP7_75t_SL g348 ( .A(n_332), .Y(n_348) );
AND2x2_ASAP7_75t_L g395 ( .A(n_332), .B(n_378), .Y(n_395) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
AND2x2_ASAP7_75t_L g434 ( .A(n_334), .B(n_352), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_335), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_SL g420 ( .A(n_336), .Y(n_420) );
AOI221xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_341), .B1(n_343), .B2(n_350), .C(n_353), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
OAI22xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_346), .B1(n_348), .B2(n_349), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OAI22xp33_ASAP7_75t_L g353 ( .A1(n_347), .A2(n_354), .B1(n_356), .B2(n_358), .Y(n_353) );
OR2x2_ASAP7_75t_L g424 ( .A(n_348), .B(n_352), .Y(n_424) );
OR2x2_ASAP7_75t_L g427 ( .A(n_348), .B(n_362), .Y(n_427) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OAI221xp5_ASAP7_75t_L g423 ( .A1(n_369), .A2(n_424), .B1(n_425), .B2(n_427), .C(n_428), .Y(n_423) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVxp67_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND3xp33_ASAP7_75t_SL g379 ( .A(n_380), .B(n_394), .C(n_406), .Y(n_379) );
AOI222xp33_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_385), .B1(n_387), .B2(n_390), .C1(n_392), .C2(n_393), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_384), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_382), .B(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g404 ( .A(n_384), .Y(n_404) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVxp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AOI221xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B1(n_397), .B2(n_399), .C(n_402), .Y(n_394) );
INVx1_ASAP7_75t_L g409 ( .A(n_395), .Y(n_409) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
OAI21xp33_ASAP7_75t_L g428 ( .A1(n_399), .A2(n_429), .B(n_430), .Y(n_428) );
INVx1_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
NOR5xp2_ASAP7_75t_L g406 ( .A(n_407), .B(n_415), .C(n_423), .D(n_432), .E(n_438), .Y(n_406) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
INVxp67_ASAP7_75t_SL g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OAI22xp5_ASAP7_75t_SL g732 ( .A1(n_445), .A2(n_447), .B1(n_728), .B2(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_SL g447 ( .A(n_448), .B(n_665), .Y(n_447) );
NOR4xp25_ASAP7_75t_L g448 ( .A(n_449), .B(n_595), .C(n_626), .D(n_645), .Y(n_448) );
NAND4xp25_ASAP7_75t_L g449 ( .A(n_450), .B(n_553), .C(n_568), .D(n_586), .Y(n_449) );
AOI222xp33_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_498), .B1(n_530), .B2(n_541), .C1(n_546), .C2(n_548), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_483), .Y(n_451) );
INVx1_ASAP7_75t_L g609 ( .A(n_452), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_463), .Y(n_452) );
AND2x2_ASAP7_75t_L g484 ( .A(n_453), .B(n_475), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_453), .B(n_487), .Y(n_638) );
INVx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g545 ( .A(n_454), .B(n_465), .Y(n_545) );
AND2x2_ASAP7_75t_L g554 ( .A(n_454), .B(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g580 ( .A(n_454), .Y(n_580) );
AND2x2_ASAP7_75t_L g601 ( .A(n_454), .B(n_465), .Y(n_601) );
BUFx2_ASAP7_75t_L g624 ( .A(n_454), .Y(n_624) );
AND2x2_ASAP7_75t_L g648 ( .A(n_454), .B(n_466), .Y(n_648) );
AND2x2_ASAP7_75t_L g712 ( .A(n_454), .B(n_475), .Y(n_712) );
AND2x2_ASAP7_75t_L g613 ( .A(n_463), .B(n_544), .Y(n_613) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_464), .B(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_475), .Y(n_464) );
OR2x2_ASAP7_75t_L g573 ( .A(n_465), .B(n_488), .Y(n_573) );
AND2x2_ASAP7_75t_L g585 ( .A(n_465), .B(n_544), .Y(n_585) );
BUFx2_ASAP7_75t_L g717 ( .A(n_465), .Y(n_717) );
INVx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OR2x2_ASAP7_75t_L g486 ( .A(n_466), .B(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g567 ( .A(n_466), .B(n_488), .Y(n_567) );
AND2x2_ASAP7_75t_L g620 ( .A(n_466), .B(n_475), .Y(n_620) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_466), .Y(n_656) );
AND2x2_ASAP7_75t_L g543 ( .A(n_475), .B(n_544), .Y(n_543) );
INVx1_ASAP7_75t_SL g555 ( .A(n_475), .Y(n_555) );
INVx2_ASAP7_75t_L g566 ( .A(n_475), .Y(n_566) );
BUFx2_ASAP7_75t_L g590 ( .A(n_475), .Y(n_590) );
AND2x2_ASAP7_75t_SL g647 ( .A(n_475), .B(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
AOI332xp33_ASAP7_75t_L g568 ( .A1(n_484), .A2(n_569), .A3(n_573), .B1(n_574), .B2(n_578), .B3(n_581), .C1(n_582), .C2(n_584), .Y(n_568) );
NAND2x1_ASAP7_75t_L g653 ( .A(n_484), .B(n_544), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_484), .B(n_558), .Y(n_704) );
A2O1A1Ixp33_ASAP7_75t_SL g586 ( .A1(n_485), .A2(n_587), .B(n_590), .C(n_591), .Y(n_586) );
AND2x2_ASAP7_75t_L g725 ( .A(n_485), .B(n_566), .Y(n_725) );
INVx3_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
OR2x2_ASAP7_75t_L g622 ( .A(n_486), .B(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g627 ( .A(n_486), .B(n_624), .Y(n_627) );
INVx1_ASAP7_75t_L g558 ( .A(n_487), .Y(n_558) );
AND2x2_ASAP7_75t_L g661 ( .A(n_487), .B(n_620), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_487), .B(n_601), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_487), .B(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_487), .B(n_579), .Y(n_687) );
INVx3_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx3_ASAP7_75t_L g544 ( .A(n_488), .Y(n_544) );
OAI31xp33_ASAP7_75t_L g726 ( .A1(n_498), .A2(n_647), .A3(n_654), .B(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_509), .Y(n_498) );
AND2x2_ASAP7_75t_L g530 ( .A(n_499), .B(n_531), .Y(n_530) );
NAND2x1_ASAP7_75t_SL g549 ( .A(n_499), .B(n_550), .Y(n_549) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_499), .Y(n_636) );
AND2x2_ASAP7_75t_L g641 ( .A(n_499), .B(n_552), .Y(n_641) );
INVx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g553 ( .A1(n_500), .A2(n_554), .B(n_556), .C(n_559), .Y(n_553) );
OR2x2_ASAP7_75t_L g570 ( .A(n_500), .B(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g583 ( .A(n_500), .Y(n_583) );
AND2x2_ASAP7_75t_L g589 ( .A(n_500), .B(n_532), .Y(n_589) );
INVx2_ASAP7_75t_L g607 ( .A(n_500), .Y(n_607) );
AND2x2_ASAP7_75t_L g618 ( .A(n_500), .B(n_572), .Y(n_618) );
AND2x2_ASAP7_75t_L g650 ( .A(n_500), .B(n_608), .Y(n_650) );
AND2x2_ASAP7_75t_L g654 ( .A(n_500), .B(n_577), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_500), .B(n_509), .Y(n_659) );
AND2x2_ASAP7_75t_L g693 ( .A(n_500), .B(n_694), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_500), .B(n_596), .Y(n_727) );
OR2x6_ASAP7_75t_L g500 ( .A(n_501), .B(n_507), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_509), .B(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g635 ( .A(n_509), .Y(n_635) );
AND2x2_ASAP7_75t_L g697 ( .A(n_509), .B(n_618), .Y(n_697) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_521), .Y(n_509) );
OR2x2_ASAP7_75t_L g551 ( .A(n_510), .B(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g561 ( .A(n_510), .B(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_510), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g669 ( .A(n_510), .Y(n_669) );
AND2x2_ASAP7_75t_L g686 ( .A(n_510), .B(n_532), .Y(n_686) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g577 ( .A(n_511), .B(n_521), .Y(n_577) );
AND2x2_ASAP7_75t_L g606 ( .A(n_511), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g617 ( .A(n_511), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_511), .B(n_572), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_518), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B(n_517), .Y(n_514) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g531 ( .A(n_522), .B(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g552 ( .A(n_522), .Y(n_552) );
AND2x2_ASAP7_75t_L g608 ( .A(n_522), .B(n_572), .Y(n_608) );
INVx1_ASAP7_75t_L g710 ( .A(n_530), .Y(n_710) );
INVx1_ASAP7_75t_L g714 ( .A(n_531), .Y(n_714) );
INVx2_ASAP7_75t_L g572 ( .A(n_532), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_542), .B(n_545), .Y(n_541) );
INVx1_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_543), .B(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_543), .B(n_648), .Y(n_706) );
OR2x2_ASAP7_75t_L g547 ( .A(n_544), .B(n_545), .Y(n_547) );
INVx1_ASAP7_75t_SL g599 ( .A(n_544), .Y(n_599) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AOI221xp5_ASAP7_75t_L g602 ( .A1(n_550), .A2(n_603), .B1(n_605), .B2(n_609), .C(n_610), .Y(n_602) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
OR2x2_ASAP7_75t_L g630 ( .A(n_551), .B(n_594), .Y(n_630) );
INVx2_ASAP7_75t_L g562 ( .A(n_552), .Y(n_562) );
INVx1_ASAP7_75t_L g588 ( .A(n_552), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_552), .B(n_572), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_552), .B(n_575), .Y(n_682) );
INVx1_ASAP7_75t_L g690 ( .A(n_552), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_554), .B(n_558), .Y(n_604) );
AND2x4_ASAP7_75t_L g579 ( .A(n_555), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g692 ( .A(n_558), .B(n_648), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_560), .B(n_563), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_561), .B(n_593), .Y(n_592) );
INVxp67_ASAP7_75t_L g700 ( .A(n_562), .Y(n_700) );
INVxp67_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_567), .Y(n_564) );
INVx1_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g600 ( .A(n_566), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g672 ( .A(n_566), .B(n_648), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_566), .B(n_585), .Y(n_678) );
AOI322xp5_ASAP7_75t_L g632 ( .A1(n_567), .A2(n_601), .A3(n_608), .B1(n_633), .B2(n_636), .C1(n_637), .C2(n_639), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_567), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g698 ( .A(n_570), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g644 ( .A(n_571), .Y(n_644) );
INVx2_ASAP7_75t_L g575 ( .A(n_572), .Y(n_575) );
INVx1_ASAP7_75t_L g634 ( .A(n_572), .Y(n_634) );
CKINVDCx16_ASAP7_75t_R g581 ( .A(n_573), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
AND2x2_ASAP7_75t_L g670 ( .A(n_575), .B(n_583), .Y(n_670) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g582 ( .A(n_577), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g625 ( .A(n_577), .B(n_618), .Y(n_625) );
AND2x2_ASAP7_75t_L g629 ( .A(n_577), .B(n_589), .Y(n_629) );
OAI21xp33_ASAP7_75t_SL g639 ( .A1(n_578), .A2(n_640), .B(n_642), .Y(n_639) );
OAI22xp33_ASAP7_75t_L g709 ( .A1(n_578), .A2(n_710), .B1(n_711), .B2(n_713), .Y(n_709) );
INVx3_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g584 ( .A(n_579), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_579), .B(n_599), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_581), .B(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
INVx1_ASAP7_75t_L g721 ( .A(n_588), .Y(n_721) );
INVx4_ASAP7_75t_L g594 ( .A(n_589), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_589), .B(n_616), .Y(n_664) );
INVx1_ASAP7_75t_SL g676 ( .A(n_590), .Y(n_676) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NOR2xp67_ASAP7_75t_L g689 ( .A(n_594), .B(n_690), .Y(n_689) );
OAI211xp5_ASAP7_75t_SL g595 ( .A1(n_596), .A2(n_597), .B(n_602), .C(n_619), .Y(n_595) );
OAI221xp5_ASAP7_75t_SL g715 ( .A1(n_597), .A2(n_635), .B1(n_714), .B2(n_716), .C(n_718), .Y(n_715) );
INVx1_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_599), .B(n_712), .Y(n_711) );
OAI31xp33_ASAP7_75t_L g691 ( .A1(n_600), .A2(n_677), .A3(n_692), .B(n_693), .Y(n_691) );
INVx1_ASAP7_75t_L g631 ( .A(n_601), .Y(n_631) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_608), .Y(n_605) );
INVx1_ASAP7_75t_L g681 ( .A(n_606), .Y(n_681) );
AND2x2_ASAP7_75t_L g694 ( .A(n_608), .B(n_617), .Y(n_694) );
AOI21xp33_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_612), .B(n_614), .Y(n_610) );
INVx1_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
INVxp67_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_618), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_618), .B(n_721), .Y(n_720) );
OAI21xp33_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_621), .B(n_625), .Y(n_619) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OAI221xp5_ASAP7_75t_SL g626 ( .A1(n_627), .A2(n_628), .B1(n_630), .B2(n_631), .C(n_632), .Y(n_626) );
A2O1A1Ixp33_ASAP7_75t_L g695 ( .A1(n_627), .A2(n_696), .B(n_698), .C(n_701), .Y(n_695) );
CKINVDCx16_ASAP7_75t_R g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_SL g679 ( .A(n_630), .B(n_680), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
INVx1_ASAP7_75t_L g657 ( .A(n_638), .Y(n_657) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g643 ( .A(n_641), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g685 ( .A(n_641), .B(n_686), .Y(n_685) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OAI211xp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_649), .B(n_651), .C(n_660), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OAI221xp5_ASAP7_75t_L g722 ( .A1(n_649), .A2(n_659), .B1(n_723), .B2(n_724), .C(n_726), .Y(n_722) );
INVx1_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_654), .B1(n_655), .B2(n_658), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
OAI21xp5_ASAP7_75t_SL g660 ( .A1(n_661), .A2(n_662), .B(n_663), .Y(n_660) );
INVx1_ASAP7_75t_SL g723 ( .A(n_662), .Y(n_723) );
INVxp67_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NOR4xp25_ASAP7_75t_L g665 ( .A(n_666), .B(n_695), .C(n_715), .D(n_722), .Y(n_665) );
OAI211xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_671), .B(n_673), .C(n_691), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_668), .B(n_670), .Y(n_667) );
INVxp67_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
O2A1O1Ixp33_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_677), .B(n_679), .C(n_683), .Y(n_673) );
INVx1_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_SL g702 ( .A(n_680), .Y(n_702) );
OR2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
OR2x2_ASAP7_75t_L g713 ( .A(n_681), .B(n_714), .Y(n_713) );
OAI21xp33_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_687), .B(n_688), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AOI221xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_703), .B1(n_705), .B2(n_707), .C(n_709), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVxp67_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_712), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_741), .Y(n_745) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
endmodule