module real_aes_15582_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_849, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_849;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g839 ( .A(n_0), .B(n_840), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g145 ( .A1(n_1), .A2(n_32), .B1(n_123), .B2(n_146), .Y(n_145) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_2), .A2(n_9), .B1(n_165), .B2(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g840 ( .A(n_3), .Y(n_840) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_4), .Y(n_121) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_5), .A2(n_10), .B1(n_182), .B2(n_185), .Y(n_181) );
OR2x2_ASAP7_75t_L g797 ( .A(n_6), .B(n_29), .Y(n_797) );
BUFx2_ASAP7_75t_L g843 ( .A(n_6), .Y(n_843) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_7), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_8), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_11), .B(n_126), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g164 ( .A1(n_12), .A2(n_96), .B1(n_165), .B2(n_166), .Y(n_164) );
AOI22xp33_ASAP7_75t_L g197 ( .A1(n_13), .A2(n_28), .B1(n_131), .B2(n_198), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g125 ( .A(n_14), .B(n_126), .Y(n_125) );
OAI21x1_ASAP7_75t_L g117 ( .A1(n_15), .A2(n_44), .B(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g787 ( .A(n_16), .Y(n_787) );
CKINVDCx5p33_ASAP7_75t_R g799 ( .A(n_16), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_17), .B(n_489), .Y(n_488) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_18), .Y(n_175) );
AOI22xp33_ASAP7_75t_L g150 ( .A1(n_19), .A2(n_37), .B1(n_151), .B2(n_152), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g527 ( .A(n_20), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g260 ( .A1(n_21), .A2(n_42), .B1(n_152), .B2(n_165), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_22), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_23), .B(n_131), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_24), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_25), .B(n_183), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_26), .B(n_140), .Y(n_536) );
CKINVDCx5p33_ASAP7_75t_R g604 ( .A(n_27), .Y(n_604) );
HB1xp67_ASAP7_75t_L g845 ( .A(n_29), .Y(n_845) );
AOI22xp5_ASAP7_75t_L g220 ( .A1(n_30), .A2(n_80), .B1(n_123), .B2(n_221), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g186 ( .A1(n_31), .A2(n_35), .B1(n_122), .B2(n_123), .Y(n_186) );
AOI22xp33_ASAP7_75t_L g168 ( .A1(n_33), .A2(n_47), .B1(n_165), .B2(n_169), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g530 ( .A(n_34), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g100 ( .A1(n_36), .A2(n_101), .B1(n_834), .B2(n_846), .Y(n_100) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_38), .B(n_126), .Y(n_472) );
INVx2_ASAP7_75t_L g792 ( .A(n_39), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_40), .B(n_127), .Y(n_484) );
BUFx3_ASAP7_75t_L g795 ( .A(n_41), .Y(n_795) );
INVx1_ASAP7_75t_L g809 ( .A(n_41), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_43), .B(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g532 ( .A(n_45), .B(n_492), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_46), .B(n_199), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_48), .B(n_183), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_49), .B(n_151), .Y(n_608) );
INVx1_ASAP7_75t_L g810 ( .A(n_50), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_51), .A2(n_67), .B1(n_151), .B2(n_169), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g212 ( .A1(n_52), .A2(n_70), .B1(n_122), .B2(n_123), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_53), .B(n_517), .Y(n_516) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_54), .A2(n_224), .B(n_473), .C(n_526), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_55), .A2(n_92), .B1(n_165), .B2(n_185), .Y(n_211) );
INVx1_ASAP7_75t_L g118 ( .A(n_56), .Y(n_118) );
AND2x4_ASAP7_75t_L g137 ( .A(n_57), .B(n_138), .Y(n_137) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_58), .A2(n_59), .B1(n_152), .B2(n_202), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_60), .B(n_140), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_61), .B(n_492), .Y(n_558) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_62), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_63), .B(n_152), .Y(n_477) );
INVx1_ASAP7_75t_L g138 ( .A(n_64), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g499 ( .A(n_65), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_66), .B(n_140), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_68), .B(n_123), .Y(n_512) );
NAND3xp33_ASAP7_75t_L g485 ( .A(n_69), .B(n_127), .C(n_146), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_71), .B(n_123), .Y(n_539) );
INVx2_ASAP7_75t_L g128 ( .A(n_72), .Y(n_128) );
CKINVDCx14_ASAP7_75t_R g459 ( .A(n_73), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_74), .B(n_188), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g607 ( .A(n_75), .B(n_126), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_76), .B(n_543), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_77), .A2(n_93), .B1(n_152), .B2(n_224), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_78), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_79), .Y(n_155) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_81), .A2(n_87), .B1(n_183), .B2(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_82), .B(n_126), .Y(n_605) );
NAND2xp33_ASAP7_75t_SL g557 ( .A(n_83), .B(n_132), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_84), .B(n_167), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g139 ( .A(n_85), .B(n_140), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g820 ( .A(n_86), .Y(n_820) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_88), .Y(n_192) );
INVx1_ASAP7_75t_L g456 ( .A(n_89), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g807 ( .A(n_89), .B(n_808), .Y(n_807) );
NAND2xp33_ASAP7_75t_L g133 ( .A(n_90), .B(n_126), .Y(n_133) );
NAND2xp33_ASAP7_75t_L g540 ( .A(n_91), .B(n_132), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_94), .B(n_492), .Y(n_520) );
NAND3xp33_ASAP7_75t_L g554 ( .A(n_95), .B(n_132), .C(n_188), .Y(n_554) );
CKINVDCx5p33_ASAP7_75t_R g828 ( .A(n_97), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_98), .B(n_123), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_99), .B(n_183), .Y(n_515) );
AO21x2_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_788), .B(n_800), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
NOR2xp33_ASAP7_75t_L g103 ( .A(n_104), .B(n_787), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_104), .B(n_799), .Y(n_798) );
AND2x4_ASAP7_75t_L g104 ( .A(n_105), .B(n_457), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g105 ( .A(n_106), .B(n_452), .Y(n_105) );
NAND2x1p5_ASAP7_75t_L g106 ( .A(n_107), .B(n_396), .Y(n_106) );
NOR3x1_ASAP7_75t_L g107 ( .A(n_108), .B(n_314), .C(n_351), .Y(n_107) );
NAND4xp75_ASAP7_75t_L g108 ( .A(n_109), .B(n_234), .C(n_268), .D(n_298), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OAI32xp33_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_156), .A3(n_206), .B1(n_215), .B2(n_229), .Y(n_110) );
OR2x2_ASAP7_75t_L g215 ( .A(n_111), .B(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OAI21xp5_ASAP7_75t_L g425 ( .A1(n_112), .A2(n_426), .B(n_428), .Y(n_425) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_141), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_113), .B(n_267), .Y(n_266) );
AND2x4_ASAP7_75t_L g297 ( .A(n_113), .B(n_243), .Y(n_297) );
AND2x2_ASAP7_75t_L g392 ( .A(n_113), .B(n_208), .Y(n_392) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
BUFx2_ASAP7_75t_L g241 ( .A(n_114), .Y(n_241) );
OAI21x1_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_119), .B(n_139), .Y(n_114) );
OAI21x1_ASAP7_75t_L g274 ( .A1(n_115), .A2(n_119), .B(n_139), .Y(n_274) );
INVx2_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
INVx4_ASAP7_75t_L g140 ( .A(n_116), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_116), .B(n_155), .Y(n_154) );
BUFx3_ASAP7_75t_L g203 ( .A(n_116), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_116), .B(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_116), .B(n_214), .Y(n_213) );
INVx2_ASAP7_75t_L g468 ( .A(n_116), .Y(n_468) );
AND2x4_ASAP7_75t_SL g547 ( .A(n_116), .B(n_478), .Y(n_547) );
INVx1_ASAP7_75t_SL g550 ( .A(n_116), .Y(n_550) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g173 ( .A(n_117), .Y(n_173) );
OAI21x1_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_129), .B(n_135), .Y(n_119) );
O2A1O1Ixp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_122), .B(n_125), .C(n_127), .Y(n_120) );
INVx4_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g169 ( .A(n_123), .Y(n_169) );
INVx1_ASAP7_75t_L g185 ( .A(n_123), .Y(n_185) );
OAI22xp33_ASAP7_75t_L g529 ( .A1(n_123), .A2(n_152), .B1(n_530), .B2(n_531), .Y(n_529) );
INVx3_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_124), .Y(n_126) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_124), .Y(n_132) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_124), .Y(n_146) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_124), .Y(n_152) );
INVx1_ASAP7_75t_L g167 ( .A(n_124), .Y(n_167) );
INVx1_ASAP7_75t_L g184 ( .A(n_124), .Y(n_184) );
INVx1_ASAP7_75t_L g199 ( .A(n_124), .Y(n_199) );
INVx1_ASAP7_75t_L g202 ( .A(n_124), .Y(n_202) );
INVx2_ASAP7_75t_L g222 ( .A(n_124), .Y(n_222) );
INVx1_ASAP7_75t_L g224 ( .A(n_124), .Y(n_224) );
INVx3_ASAP7_75t_L g165 ( .A(n_126), .Y(n_165) );
INVx1_ASAP7_75t_L g489 ( .A(n_126), .Y(n_489) );
OAI21xp5_ASAP7_75t_L g552 ( .A1(n_126), .A2(n_553), .B(n_554), .Y(n_552) );
INVx6_ASAP7_75t_L g134 ( .A(n_127), .Y(n_134) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_127), .A2(n_476), .B(n_477), .Y(n_475) );
O2A1O1Ixp5_ASAP7_75t_L g603 ( .A1(n_127), .A2(n_166), .B(n_604), .C(n_605), .Y(n_603) );
BUFx8_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g149 ( .A(n_128), .Y(n_149) );
INVx1_ASAP7_75t_L g188 ( .A(n_128), .Y(n_188) );
INVx1_ASAP7_75t_L g474 ( .A(n_128), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_133), .B(n_134), .Y(n_129) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g151 ( .A(n_132), .Y(n_151) );
OAI22xp5_ASAP7_75t_L g144 ( .A1(n_134), .A2(n_145), .B1(n_147), .B2(n_150), .Y(n_144) );
OAI22xp5_ASAP7_75t_L g163 ( .A1(n_134), .A2(n_147), .B1(n_164), .B2(n_168), .Y(n_163) );
OAI22xp5_ASAP7_75t_L g180 ( .A1(n_134), .A2(n_181), .B1(n_186), .B2(n_187), .Y(n_180) );
OAI22xp5_ASAP7_75t_L g196 ( .A1(n_134), .A2(n_147), .B1(n_197), .B2(n_200), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g210 ( .A1(n_134), .A2(n_187), .B1(n_211), .B2(n_212), .Y(n_210) );
OAI22xp5_ASAP7_75t_L g219 ( .A1(n_134), .A2(n_220), .B1(n_223), .B2(n_225), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g258 ( .A1(n_134), .A2(n_147), .B1(n_259), .B2(n_260), .Y(n_258) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_134), .A2(n_147), .B1(n_495), .B2(n_497), .Y(n_494) );
INVx2_ASAP7_75t_SL g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_SL g226 ( .A(n_136), .Y(n_226) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
BUFx10_ASAP7_75t_L g143 ( .A(n_137), .Y(n_143) );
BUFx10_ASAP7_75t_L g478 ( .A(n_137), .Y(n_478) );
INVx2_ASAP7_75t_L g153 ( .A(n_140), .Y(n_153) );
INVx2_ASAP7_75t_L g265 ( .A(n_141), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_141), .B(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_142), .Y(n_252) );
INVx1_ASAP7_75t_L g296 ( .A(n_142), .Y(n_296) );
AND2x2_ASAP7_75t_L g340 ( .A(n_142), .B(n_274), .Y(n_340) );
OR2x2_ASAP7_75t_L g394 ( .A(n_142), .B(n_218), .Y(n_394) );
AO31x2_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_144), .A3(n_153), .B(n_154), .Y(n_142) );
INVx2_ASAP7_75t_L g162 ( .A(n_143), .Y(n_162) );
AO31x2_ASAP7_75t_L g179 ( .A1(n_143), .A2(n_180), .A3(n_189), .B(n_191), .Y(n_179) );
AO31x2_ASAP7_75t_L g195 ( .A1(n_143), .A2(n_196), .A3(n_203), .B(n_204), .Y(n_195) );
AO31x2_ASAP7_75t_L g493 ( .A1(n_143), .A2(n_172), .A3(n_494), .B(n_498), .Y(n_493) );
INVx2_ASAP7_75t_L g517 ( .A(n_146), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_147), .B(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g518 ( .A(n_148), .Y(n_518) );
BUFx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g544 ( .A(n_149), .Y(n_544) );
OAI21xp5_ASAP7_75t_L g483 ( .A1(n_152), .A2(n_484), .B(n_485), .Y(n_483) );
INVx2_ASAP7_75t_L g496 ( .A(n_152), .Y(n_496) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_157), .A2(n_320), .B1(n_412), .B2(n_414), .Y(n_411) );
AND2x2_ASAP7_75t_L g157 ( .A(n_158), .B(n_177), .Y(n_157) );
INVx4_ASAP7_75t_L g237 ( .A(n_158), .Y(n_237) );
AOI22xp5_ASAP7_75t_L g248 ( .A1(n_158), .A2(n_217), .B1(n_249), .B2(n_251), .Y(n_248) );
OR2x2_ASAP7_75t_L g254 ( .A(n_158), .B(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g373 ( .A(n_158), .B(n_272), .Y(n_373) );
INVx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g293 ( .A(n_159), .B(n_178), .Y(n_293) );
AND2x2_ASAP7_75t_L g384 ( .A(n_159), .B(n_256), .Y(n_384) );
AND2x2_ASAP7_75t_L g439 ( .A(n_159), .B(n_195), .Y(n_439) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g233 ( .A(n_160), .Y(n_233) );
AND2x4_ASAP7_75t_L g360 ( .A(n_160), .B(n_256), .Y(n_360) );
AO31x2_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_163), .A3(n_170), .B(n_174), .Y(n_160) );
AO31x2_ASAP7_75t_L g209 ( .A1(n_161), .A2(n_189), .A3(n_210), .B(n_213), .Y(n_209) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NOR2xp67_ASAP7_75t_SL g523 ( .A(n_162), .B(n_171), .Y(n_523) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AO31x2_ASAP7_75t_L g257 ( .A1(n_170), .A2(n_226), .A3(n_258), .B(n_261), .Y(n_257) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NOR2xp33_ASAP7_75t_SL g191 ( .A(n_172), .B(n_192), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_172), .B(n_228), .Y(n_227) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g176 ( .A(n_173), .Y(n_176) );
INVx2_ASAP7_75t_L g190 ( .A(n_173), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_175), .B(n_176), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_176), .B(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g492 ( .A(n_176), .Y(n_492) );
INVx2_ASAP7_75t_L g519 ( .A(n_176), .Y(n_519) );
NAND2x1_ASAP7_75t_L g236 ( .A(n_177), .B(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g343 ( .A(n_177), .B(n_344), .Y(n_343) );
AND2x4_ASAP7_75t_L g177 ( .A(n_178), .B(n_193), .Y(n_177) );
INVx2_ASAP7_75t_L g231 ( .A(n_178), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_178), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g279 ( .A(n_178), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_178), .B(n_281), .Y(n_306) );
AND2x2_ASAP7_75t_L g309 ( .A(n_178), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g369 ( .A(n_178), .Y(n_369) );
INVx4_ASAP7_75t_SL g178 ( .A(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_179), .B(n_194), .Y(n_247) );
BUFx2_ASAP7_75t_L g285 ( .A(n_179), .Y(n_285) );
AND2x2_ASAP7_75t_L g334 ( .A(n_179), .B(n_195), .Y(n_334) );
AND2x2_ASAP7_75t_L g376 ( .A(n_179), .B(n_257), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_179), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx1_ASAP7_75t_SL g187 ( .A(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g225 ( .A(n_188), .Y(n_225) );
INVx1_ASAP7_75t_L g490 ( .A(n_188), .Y(n_490) );
BUFx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_190), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_195), .B(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g287 ( .A(n_195), .B(n_257), .Y(n_287) );
INVx1_ASAP7_75t_L g310 ( .A(n_195), .Y(n_310) );
INVx2_ASAP7_75t_L g330 ( .A(n_195), .Y(n_330) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_195), .Y(n_375) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AO31x2_ASAP7_75t_L g218 ( .A1(n_203), .A2(n_219), .A3(n_226), .B(n_227), .Y(n_218) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g294 ( .A(n_207), .B(n_295), .Y(n_294) );
NOR2x1p5_ASAP7_75t_L g400 ( .A(n_207), .B(n_394), .Y(n_400) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x4_ASAP7_75t_L g217 ( .A(n_208), .B(n_218), .Y(n_217) );
INVx3_ASAP7_75t_L g250 ( .A(n_208), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_208), .B(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_208), .B(n_326), .Y(n_325) );
INVx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g242 ( .A(n_209), .B(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g300 ( .A(n_209), .B(n_218), .Y(n_300) );
BUFx2_ASAP7_75t_L g413 ( .A(n_209), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_215), .B(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g451 ( .A(n_215), .Y(n_451) );
INVx2_ASAP7_75t_SL g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g387 ( .A(n_217), .Y(n_387) );
AND2x4_ASAP7_75t_L g410 ( .A(n_217), .B(n_340), .Y(n_410) );
AND2x2_ASAP7_75t_L g434 ( .A(n_217), .B(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g243 ( .A(n_218), .Y(n_243) );
BUFx2_ASAP7_75t_L g267 ( .A(n_218), .Y(n_267) );
INVx1_ASAP7_75t_L g323 ( .A(n_218), .Y(n_323) );
OR2x2_ASAP7_75t_L g445 ( .A(n_218), .B(n_302), .Y(n_445) );
INVx2_ASAP7_75t_SL g221 ( .A(n_222), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_222), .B(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g545 ( .A(n_224), .Y(n_545) );
HB1xp67_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_232), .Y(n_230) );
INVx2_ASAP7_75t_L g291 ( .A(n_231), .Y(n_291) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_232), .Y(n_308) );
INVx1_ASAP7_75t_L g312 ( .A(n_232), .Y(n_312) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g253 ( .A(n_233), .Y(n_253) );
OR2x2_ASAP7_75t_L g290 ( .A(n_233), .B(n_282), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_238), .B(n_244), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_239), .A2(n_333), .B1(n_335), .B2(n_338), .Y(n_332) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
OR2x2_ASAP7_75t_L g378 ( .A(n_241), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g386 ( .A(n_241), .Y(n_386) );
AND2x2_ASAP7_75t_L g399 ( .A(n_241), .B(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g361 ( .A(n_242), .B(n_340), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_248), .B1(n_254), .B2(n_263), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g313 ( .A(n_247), .Y(n_313) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x4_ASAP7_75t_L g271 ( .A(n_250), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g339 ( .A(n_250), .B(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g348 ( .A(n_250), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_250), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_251), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
AND2x2_ASAP7_75t_L g336 ( .A(n_253), .B(n_337), .Y(n_336) );
INVx3_ASAP7_75t_L g350 ( .A(n_253), .Y(n_350) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g282 ( .A(n_257), .Y(n_282) );
AND2x4_ASAP7_75t_L g329 ( .A(n_257), .B(n_330), .Y(n_329) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_257), .Y(n_345) );
INVx1_ASAP7_75t_L g409 ( .A(n_257), .Y(n_409) );
OR2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
AND2x4_ASAP7_75t_L g301 ( .A(n_265), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g318 ( .A(n_265), .Y(n_318) );
INVx1_ASAP7_75t_L g276 ( .A(n_267), .Y(n_276) );
AOI22xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_277), .B1(n_288), .B2(n_294), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2x1p5_ASAP7_75t_L g270 ( .A(n_271), .B(n_275), .Y(n_270) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVxp67_ASAP7_75t_SL g326 ( .A(n_273), .Y(n_326) );
INVx1_ASAP7_75t_L g302 ( .A(n_274), .Y(n_302) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_278), .B(n_283), .Y(n_277) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_279), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g431 ( .A(n_280), .Y(n_431) );
INVx1_ASAP7_75t_L g450 ( .A(n_280), .Y(n_450) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2x1_ASAP7_75t_L g427 ( .A(n_284), .B(n_350), .Y(n_427) );
AND2x4_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVx1_ASAP7_75t_L g443 ( .A(n_285), .Y(n_443) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_292), .Y(n_288) );
INVx2_ASAP7_75t_L g381 ( .A(n_289), .Y(n_381) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx2_ASAP7_75t_L g370 ( .A(n_290), .Y(n_370) );
AND2x4_ASAP7_75t_L g372 ( .A(n_291), .B(n_329), .Y(n_372) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_295), .A2(n_441), .B1(n_444), .B2(n_446), .Y(n_440) );
AND2x4_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
INVx2_ASAP7_75t_L g365 ( .A(n_296), .Y(n_365) );
INVx1_ASAP7_75t_L g319 ( .A(n_297), .Y(n_319) );
AND2x4_ASAP7_75t_L g412 ( .A(n_297), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g420 ( .A(n_297), .B(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_303), .Y(n_298) );
AND2x4_ASAP7_75t_SL g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx1_ASAP7_75t_SL g363 ( .A(n_300), .Y(n_363) );
INVx2_ASAP7_75t_L g379 ( .A(n_300), .Y(n_379) );
INVx1_ASAP7_75t_L g406 ( .A(n_301), .Y(n_406) );
AND2x2_ASAP7_75t_L g437 ( .A(n_301), .B(n_348), .Y(n_437) );
NAND3xp33_ASAP7_75t_L g303 ( .A(n_304), .B(n_307), .C(n_311), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_308), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g349 ( .A(n_309), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_309), .B(n_384), .Y(n_417) );
INVx1_ASAP7_75t_L g337 ( .A(n_310), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_312), .B(n_376), .Y(n_402) );
INVx1_ASAP7_75t_L g357 ( .A(n_313), .Y(n_357) );
NAND3xp33_ASAP7_75t_L g314 ( .A(n_315), .B(n_331), .C(n_341), .Y(n_314) );
OAI21xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_320), .B(n_327), .Y(n_315) );
INVxp67_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx1_ASAP7_75t_L g435 ( .A(n_318), .Y(n_435) );
AND2x4_ASAP7_75t_L g320 ( .A(n_321), .B(n_324), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AOI32xp33_ASAP7_75t_L g371 ( .A1(n_322), .A2(n_372), .A3(n_373), .B1(n_374), .B2(n_377), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_322), .B(n_406), .Y(n_405) );
BUFx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g355 ( .A(n_329), .Y(n_355) );
NAND2x1p5_ASAP7_75t_L g390 ( .A(n_329), .B(n_350), .Y(n_390) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_334), .B(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g395 ( .A(n_334), .B(n_344), .Y(n_395) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g423 ( .A(n_337), .Y(n_423) );
INVx1_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
AOI22xp33_ASAP7_75t_SL g341 ( .A1(n_339), .A2(n_342), .B1(n_346), .B2(n_349), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_340), .B(n_348), .Y(n_347) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_342), .A2(n_400), .B1(n_437), .B2(n_438), .Y(n_436) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g438 ( .A(n_344), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_346), .A2(n_389), .B1(n_391), .B2(n_395), .Y(n_388) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g430 ( .A(n_350), .Y(n_430) );
NAND4xp25_ASAP7_75t_L g351 ( .A(n_352), .B(n_371), .C(n_380), .D(n_388), .Y(n_351) );
O2A1O1Ixp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_358), .B(n_361), .C(n_362), .Y(n_352) );
NOR2x1_ASAP7_75t_L g353 ( .A(n_354), .B(n_356), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx3_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x4_ASAP7_75t_L g416 ( .A(n_360), .B(n_375), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_360), .B(n_443), .Y(n_442) );
AOI21xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_364), .B(n_366), .Y(n_362) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_367), .A2(n_405), .B1(n_407), .B2(n_410), .Y(n_404) );
AND2x4_ASAP7_75t_L g367 ( .A(n_368), .B(n_370), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OAI21xp5_ASAP7_75t_L g433 ( .A1(n_372), .A2(n_377), .B(n_434), .Y(n_433) );
AND2x4_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OAI21xp33_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_382), .B(n_385), .Y(n_380) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NOR2xp33_ASAP7_75t_R g385 ( .A(n_386), .B(n_387), .Y(n_385) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_395), .A2(n_412), .B1(n_449), .B2(n_451), .Y(n_448) );
NOR3x1_ASAP7_75t_L g396 ( .A(n_397), .B(n_418), .C(n_432), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_411), .Y(n_397) );
AOI21xp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_401), .B(n_403), .Y(n_398) );
INVx1_ASAP7_75t_L g424 ( .A(n_399), .Y(n_424) );
INVx2_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
INVxp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g447 ( .A(n_409), .Y(n_447) );
INVx1_ASAP7_75t_L g421 ( .A(n_413), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_415), .B(n_417), .Y(n_414) );
OAI221xp5_ASAP7_75t_L g418 ( .A1(n_415), .A2(n_419), .B1(n_422), .B2(n_424), .C(n_425), .Y(n_418) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
NAND4xp25_ASAP7_75t_SL g432 ( .A(n_433), .B(n_436), .C(n_440), .D(n_448), .Y(n_432) );
AND2x2_ASAP7_75t_L g446 ( .A(n_439), .B(n_447), .Y(n_446) );
INVxp67_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
INVxp67_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx4_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx12f_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g825 ( .A(n_455), .B(n_826), .Y(n_825) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx2_ASAP7_75t_L g786 ( .A(n_456), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_458), .B(n_783), .Y(n_457) );
INVxp33_ASAP7_75t_L g811 ( .A(n_458), .Y(n_811) );
XNOR2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
NAND2x1p5_ASAP7_75t_SL g460 ( .A(n_461), .B(n_717), .Y(n_460) );
NOR2x1_ASAP7_75t_L g461 ( .A(n_462), .B(n_653), .Y(n_461) );
NAND4xp25_ASAP7_75t_L g462 ( .A(n_463), .B(n_575), .C(n_614), .D(n_643), .Y(n_462) );
O2A1O1Ixp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_500), .B(n_507), .C(n_559), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_480), .Y(n_464) );
INVx2_ASAP7_75t_L g503 ( .A(n_465), .Y(n_503) );
AND2x2_ASAP7_75t_L g641 ( .A(n_465), .B(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_465), .B(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_465), .B(n_561), .Y(n_736) );
OR2x2_ASAP7_75t_L g772 ( .A(n_465), .B(n_688), .Y(n_772) );
INVx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g669 ( .A(n_466), .B(n_481), .Y(n_669) );
NOR2xp67_ASAP7_75t_L g695 ( .A(n_466), .B(n_505), .Y(n_695) );
BUFx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g630 ( .A(n_467), .Y(n_630) );
OAI21x1_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_469), .B(n_479), .Y(n_467) );
OAI21x1_ASAP7_75t_L g481 ( .A1(n_468), .A2(n_482), .B(n_491), .Y(n_481) );
OAI21x1_ASAP7_75t_L g563 ( .A1(n_468), .A2(n_469), .B(n_479), .Y(n_563) );
OA21x2_ASAP7_75t_L g598 ( .A1(n_468), .A2(n_482), .B(n_491), .Y(n_598) );
OAI21x1_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_475), .B(n_478), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B(n_473), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_473), .A2(n_512), .B(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_473), .A2(n_539), .B(n_540), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_473), .A2(n_556), .B(n_557), .Y(n_555) );
BUFx4f_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
OAI21x1_ASAP7_75t_L g482 ( .A1(n_478), .A2(n_483), .B(n_486), .Y(n_482) );
OAI21x1_ASAP7_75t_L g510 ( .A1(n_478), .A2(n_511), .B(n_514), .Y(n_510) );
OAI21x1_ASAP7_75t_L g551 ( .A1(n_478), .A2(n_552), .B(n_555), .Y(n_551) );
OAI21x1_ASAP7_75t_L g602 ( .A1(n_478), .A2(n_603), .B(n_606), .Y(n_602) );
AND2x2_ASAP7_75t_L g569 ( .A(n_480), .B(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_480), .B(n_599), .Y(n_613) );
AND2x2_ASAP7_75t_L g621 ( .A(n_480), .B(n_622), .Y(n_621) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_480), .Y(n_644) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_493), .Y(n_480) );
INVx1_ASAP7_75t_L g505 ( .A(n_481), .Y(n_505) );
INVx1_ASAP7_75t_L g561 ( .A(n_481), .Y(n_561) );
AND2x2_ASAP7_75t_L g631 ( .A(n_481), .B(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g692 ( .A(n_481), .B(n_600), .Y(n_692) );
AOI21x1_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_488), .B(n_490), .Y(n_486) );
INVx1_ASAP7_75t_L g506 ( .A(n_493), .Y(n_506) );
AND2x2_ASAP7_75t_L g562 ( .A(n_493), .B(n_563), .Y(n_562) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_493), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_493), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g675 ( .A(n_493), .B(n_630), .Y(n_675) );
OR2x2_ASAP7_75t_L g688 ( .A(n_493), .B(n_598), .Y(n_688) );
OR2x2_ASAP7_75t_L g698 ( .A(n_493), .B(n_563), .Y(n_698) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_503), .B(n_504), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_503), .B(n_714), .Y(n_760) );
INVx1_ASAP7_75t_L g616 ( .A(n_504), .Y(n_616) );
AND2x4_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
AND2x2_ASAP7_75t_L g700 ( .A(n_506), .B(n_563), .Y(n_700) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_533), .Y(n_507) );
AND2x2_ASAP7_75t_L g573 ( .A(n_508), .B(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g635 ( .A(n_508), .Y(n_635) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_521), .Y(n_508) );
BUFx2_ASAP7_75t_L g742 ( .A(n_509), .Y(n_742) );
OAI21xp33_ASAP7_75t_SL g509 ( .A1(n_510), .A2(n_519), .B(n_520), .Y(n_509) );
OAI21x1_ASAP7_75t_L g583 ( .A1(n_510), .A2(n_519), .B(n_520), .Y(n_583) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B(n_518), .Y(n_514) );
OAI21x1_ASAP7_75t_L g601 ( .A1(n_519), .A2(n_602), .B(n_609), .Y(n_601) );
OAI21xp5_ASAP7_75t_L g632 ( .A1(n_519), .A2(n_602), .B(n_609), .Y(n_632) );
AND2x2_ASAP7_75t_L g581 ( .A(n_521), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g567 ( .A(n_522), .B(n_549), .Y(n_567) );
INVx2_ASAP7_75t_L g593 ( .A(n_522), .Y(n_593) );
AOI21x1_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_524), .B(n_532), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_525), .B(n_528), .Y(n_524) );
AND2x2_ASAP7_75t_L g739 ( .A(n_533), .B(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_548), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx4_ASAP7_75t_L g566 ( .A(n_535), .Y(n_566) );
BUFx2_ASAP7_75t_L g574 ( .A(n_535), .Y(n_574) );
OR2x2_ASAP7_75t_L g578 ( .A(n_535), .B(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g638 ( .A(n_535), .B(n_582), .Y(n_638) );
AND2x4_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
OAI21x1_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_541), .B(n_547), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_544), .B1(n_545), .B2(n_546), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g606 ( .A1(n_543), .A2(n_607), .B(n_608), .Y(n_606) );
INVx2_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g625 ( .A(n_548), .Y(n_625) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_548), .Y(n_639) );
INVx2_ASAP7_75t_L g664 ( .A(n_548), .Y(n_664) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g579 ( .A(n_549), .Y(n_579) );
OAI21x1_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_551), .B(n_558), .Y(n_549) );
OAI22xp33_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_564), .B1(n_568), .B2(n_572), .Y(n_559) );
INVx1_ASAP7_75t_L g649 ( .A(n_560), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
INVx2_ASAP7_75t_L g660 ( .A(n_561), .Y(n_660) );
AND2x2_ASAP7_75t_L g677 ( .A(n_562), .B(n_678), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_562), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g571 ( .A(n_563), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_564), .B(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_567), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_565), .B(n_581), .Y(n_672) );
AND2x2_ASAP7_75t_L g680 ( .A(n_565), .B(n_646), .Y(n_680) );
AND2x2_ASAP7_75t_L g756 ( .A(n_565), .B(n_703), .Y(n_756) );
BUFx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g591 ( .A(n_566), .B(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g612 ( .A(n_566), .B(n_582), .Y(n_612) );
OR2x2_ASAP7_75t_L g624 ( .A(n_566), .B(n_625), .Y(n_624) );
NAND2x1_ASAP7_75t_L g658 ( .A(n_566), .B(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g663 ( .A(n_566), .Y(n_663) );
INVx2_ASAP7_75t_L g657 ( .A(n_567), .Y(n_657) );
AND2x2_ASAP7_75t_L g683 ( .A(n_567), .B(n_647), .Y(n_683) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_570), .Y(n_619) );
INVx1_ASAP7_75t_L g686 ( .A(n_570), .Y(n_686) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g670 ( .A(n_571), .B(n_600), .Y(n_670) );
AOI21xp33_ASAP7_75t_L g681 ( .A1(n_572), .A2(n_682), .B(n_684), .Y(n_681) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x4_ASAP7_75t_L g743 ( .A(n_574), .B(n_683), .Y(n_743) );
INVx1_ASAP7_75t_L g779 ( .A(n_574), .Y(n_779) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_584), .B(n_588), .Y(n_575) );
AOI322xp5_ASAP7_75t_L g727 ( .A1(n_576), .A2(n_623), .A3(n_728), .B1(n_729), .B2(n_730), .C1(n_731), .C2(n_734), .Y(n_727) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_580), .Y(n_577) );
NOR3xp33_ASAP7_75t_L g715 ( .A(n_578), .B(n_580), .C(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g594 ( .A(n_579), .B(n_595), .Y(n_594) );
OR2x2_ASAP7_75t_L g723 ( .A(n_579), .B(n_724), .Y(n_723) );
HB1xp67_ASAP7_75t_L g775 ( .A(n_579), .Y(n_775) );
OR2x2_ASAP7_75t_L g671 ( .A(n_580), .B(n_624), .Y(n_671) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g659 ( .A(n_582), .Y(n_659) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g595 ( .A(n_583), .Y(n_595) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVxp67_ASAP7_75t_SL g720 ( .A(n_585), .Y(n_720) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g691 ( .A(n_586), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g754 ( .A(n_587), .B(n_714), .Y(n_754) );
OAI21xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_596), .B(n_610), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_590), .B(n_768), .Y(n_767) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_594), .Y(n_590) );
AND2x2_ASAP7_75t_L g646 ( .A(n_592), .B(n_647), .Y(n_646) );
AND3x2_ASAP7_75t_L g690 ( .A(n_592), .B(n_594), .C(n_663), .Y(n_690) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g652 ( .A(n_593), .Y(n_652) );
AND2x2_ASAP7_75t_L g703 ( .A(n_593), .B(n_664), .Y(n_703) );
INVx2_ASAP7_75t_L g726 ( .A(n_593), .Y(n_726) );
AND2x2_ASAP7_75t_L g730 ( .A(n_594), .B(n_726), .Y(n_730) );
INVx2_ASAP7_75t_L g647 ( .A(n_595), .Y(n_647) );
OR2x2_ASAP7_75t_L g781 ( .A(n_595), .B(n_664), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_596), .B(n_709), .Y(n_708) );
OR2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_599), .Y(n_596) );
INVx1_ASAP7_75t_L g733 ( .A(n_597), .Y(n_733) );
AND2x2_ASAP7_75t_L g642 ( .A(n_598), .B(n_632), .Y(n_642) );
AND2x2_ASAP7_75t_L g678 ( .A(n_598), .B(n_600), .Y(n_678) );
AND2x2_ASAP7_75t_L g674 ( .A(n_599), .B(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_599), .B(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g746 ( .A(n_599), .Y(n_746) );
BUFx3_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g617 ( .A(n_600), .Y(n_617) );
INVxp67_ASAP7_75t_SL g622 ( .A(n_600), .Y(n_622) );
INVxp67_ASAP7_75t_SL g668 ( .A(n_600), .Y(n_668) );
INVx1_ASAP7_75t_L g714 ( .A(n_600), .Y(n_714) );
INVx3_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
OR2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AOI21xp5_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_623), .B(n_626), .Y(n_614) );
OAI31xp33_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_617), .A3(n_618), .B(n_620), .Y(n_615) );
INVx1_ASAP7_75t_L g697 ( .A(n_617), .Y(n_697) );
OAI32xp33_ASAP7_75t_L g655 ( .A1(n_618), .A2(n_627), .A3(n_656), .B1(n_660), .B2(n_661), .Y(n_655) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g648 ( .A(n_624), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_633), .B1(n_636), .B2(n_640), .Y(n_626) );
OAI22xp33_ASAP7_75t_SL g711 ( .A1(n_627), .A2(n_672), .B1(n_712), .B2(n_713), .Y(n_711) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
INVx2_ASAP7_75t_L g769 ( .A(n_629), .Y(n_769) );
BUFx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g724 ( .A(n_632), .Y(n_724) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx3_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
AND2x2_ASAP7_75t_L g650 ( .A(n_638), .B(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g725 ( .A(n_638), .B(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g776 ( .A(n_638), .Y(n_776) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g716 ( .A(n_642), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_645), .B1(n_649), .B2(n_650), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_645), .B(n_758), .Y(n_757) );
AND2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_648), .Y(n_645) );
AND2x2_ASAP7_75t_L g702 ( .A(n_647), .B(n_663), .Y(n_702) );
AOI211xp5_ASAP7_75t_L g707 ( .A1(n_650), .A2(n_708), .B(n_711), .C(n_715), .Y(n_707) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_652), .Y(n_765) );
INVx1_ASAP7_75t_L g782 ( .A(n_652), .Y(n_782) );
NAND4xp25_ASAP7_75t_L g653 ( .A(n_654), .B(n_676), .C(n_689), .D(n_707), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_655), .B(n_665), .Y(n_654) );
OR2x6_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_659), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g764 ( .A(n_662), .B(n_765), .Y(n_764) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
OAI22xp33_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_671), .B1(n_672), .B2(n_673), .Y(n_665) );
NOR2xp33_ASAP7_75t_SL g666 ( .A(n_667), .B(n_670), .Y(n_666) );
BUFx2_ASAP7_75t_L g679 ( .A(n_667), .Y(n_679) );
AND2x4_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_673), .B(n_759), .Y(n_758) );
INVx3_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g728 ( .A(n_675), .B(n_714), .Y(n_728) );
O2A1O1Ixp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_679), .B(n_680), .C(n_681), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_678), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g738 ( .A(n_685), .B(n_739), .Y(n_738) );
AND2x4_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_691), .B1(n_693), .B2(n_701), .C(n_704), .Y(n_689) );
AND2x2_ASAP7_75t_L g768 ( .A(n_692), .B(n_769), .Y(n_768) );
NAND3xp33_ASAP7_75t_SL g693 ( .A(n_694), .B(n_696), .C(n_699), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
OR2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_697), .B(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_697), .B(n_733), .Y(n_763) );
INVx1_ASAP7_75t_L g706 ( .A(n_698), .Y(n_706) );
INVx1_ASAP7_75t_L g710 ( .A(n_698), .Y(n_710) );
AND2x2_ASAP7_75t_L g751 ( .A(n_700), .B(n_740), .Y(n_751) );
NAND2xp33_ASAP7_75t_SL g752 ( .A(n_700), .B(n_722), .Y(n_752) );
AND2x4_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
INVx1_ASAP7_75t_L g712 ( .A(n_703), .Y(n_712) );
NOR3x1_ASAP7_75t_L g717 ( .A(n_718), .B(n_747), .C(n_766), .Y(n_717) );
NAND3xp33_ASAP7_75t_L g718 ( .A(n_719), .B(n_727), .C(n_737), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .Y(n_719) );
AND2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_725), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g740 ( .A(n_724), .Y(n_740) );
INVx2_ASAP7_75t_L g729 ( .A(n_726), .Y(n_729) );
AOI22xp5_ASAP7_75t_L g777 ( .A1(n_728), .A2(n_771), .B1(n_778), .B2(n_849), .Y(n_777) );
O2A1O1Ixp5_ASAP7_75t_L g749 ( .A1(n_729), .A2(n_741), .B(n_750), .C(n_752), .Y(n_749) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AO21x1_ASAP7_75t_L g753 ( .A1(n_732), .A2(n_754), .B(n_755), .Y(n_753) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
OR2x2_ASAP7_75t_L g745 ( .A(n_736), .B(n_746), .Y(n_745) );
AOI22xp5_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_741), .B1(n_743), .B2(n_744), .Y(n_737) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
NAND4xp75_ASAP7_75t_L g747 ( .A(n_748), .B(n_753), .C(n_757), .D(n_761), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
HB1xp67_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_762), .B(n_764), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
NAND3xp33_ASAP7_75t_L g766 ( .A(n_767), .B(n_770), .C(n_777), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_771), .B(n_773), .Y(n_770) );
INVx2_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVxp67_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
OR2x2_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
AND2x4_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .Y(n_778) );
NOR2x1p5_ASAP7_75t_SL g780 ( .A(n_781), .B(n_782), .Y(n_780) );
CKINVDCx5p33_ASAP7_75t_R g783 ( .A(n_784), .Y(n_783) );
CKINVDCx5p33_ASAP7_75t_R g784 ( .A(n_785), .Y(n_784) );
BUFx6f_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
AND3x2_ASAP7_75t_L g832 ( .A(n_786), .B(n_796), .C(n_833), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_786), .B(n_839), .Y(n_838) );
AND2x2_ASAP7_75t_L g788 ( .A(n_789), .B(n_798), .Y(n_788) );
BUFx12f_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
AND2x6_ASAP7_75t_SL g790 ( .A(n_791), .B(n_793), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx3_ASAP7_75t_L g817 ( .A(n_792), .Y(n_817) );
NOR2xp33_ASAP7_75t_L g823 ( .A(n_792), .B(n_824), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_794), .B(n_796), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
NOR2x1_ASAP7_75t_L g826 ( .A(n_795), .B(n_797), .Y(n_826) );
AND2x6_ASAP7_75t_SL g806 ( .A(n_796), .B(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
A2O1A1Ixp33_ASAP7_75t_L g800 ( .A1(n_801), .A2(n_812), .B(n_814), .C(n_818), .Y(n_800) );
NAND2xp33_ASAP7_75t_SL g801 ( .A(n_802), .B(n_811), .Y(n_801) );
NOR2xp33_ASAP7_75t_SL g802 ( .A(n_803), .B(n_810), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_804), .B(n_810), .Y(n_813) );
BUFx2_ASAP7_75t_SL g804 ( .A(n_805), .Y(n_804) );
INVx3_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
HB1xp67_ASAP7_75t_L g833 ( .A(n_809), .Y(n_833) );
OR2x2_ASAP7_75t_L g812 ( .A(n_811), .B(n_813), .Y(n_812) );
INVxp67_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
BUFx2_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx2_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
NOR2xp33_ASAP7_75t_SL g818 ( .A(n_819), .B(n_827), .Y(n_818) );
NOR2xp33_ASAP7_75t_L g819 ( .A(n_820), .B(n_821), .Y(n_819) );
INVx6_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
BUFx10_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
NOR2xp33_ASAP7_75t_L g827 ( .A(n_828), .B(n_829), .Y(n_827) );
INVx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx3_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx4_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
NOR2x1p5_ASAP7_75t_L g837 ( .A(n_833), .B(n_838), .Y(n_837) );
INVx4_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx8_ASAP7_75t_L g847 ( .A(n_835), .Y(n_847) );
OR2x6_ASAP7_75t_L g835 ( .A(n_836), .B(n_841), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
NOR2xp33_ASAP7_75t_L g842 ( .A(n_843), .B(n_844), .Y(n_842) );
INVxp33_ASAP7_75t_SL g844 ( .A(n_845), .Y(n_844) );
INVx4_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
endmodule