module fake_jpeg_18034_n_165 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_165);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_10),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_10),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_22),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_48),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_13),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_47),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_12),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_12),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_74),
.Y(n_91)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_58),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_0),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_77),
.Y(n_92)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_0),
.Y(n_79)
);

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_79),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_67),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_80),
.A2(n_71),
.B1(n_70),
.B2(n_52),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_73),
.A2(n_66),
.B1(n_60),
.B2(n_65),
.Y(n_81)
);

AO22x1_ASAP7_75t_SL g107 ( 
.A1(n_81),
.A2(n_59),
.B1(n_50),
.B2(n_54),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_76),
.A2(n_66),
.B1(n_60),
.B2(n_63),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_82),
.A2(n_64),
.B1(n_54),
.B2(n_55),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_87),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_59),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

NAND2x1p5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_64),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_105),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_111),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_92),
.B(n_83),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_102),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_88),
.B(n_68),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_82),
.A2(n_69),
.B1(n_53),
.B2(n_61),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_103),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_91),
.B(n_54),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_106),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_107),
.A2(n_110),
.B1(n_57),
.B2(n_4),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_1),
.Y(n_109)
);

NAND3xp33_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_2),
.C(n_4),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_113),
.B(n_118),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_115),
.A2(n_117),
.B1(n_122),
.B2(n_124),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_108),
.A2(n_23),
.B1(n_46),
.B2(n_45),
.Y(n_117)
);

AND2x4_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_57),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_109),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_112),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_124)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_128),
.Y(n_136)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_121),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_127),
.B(n_131),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_125),
.Y(n_128)
);

OAI32xp33_ASAP7_75t_L g132 ( 
.A1(n_130),
.A2(n_118),
.A3(n_123),
.B1(n_116),
.B2(n_122),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_135),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_130),
.A2(n_118),
.B1(n_114),
.B2(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

AO21x1_ASAP7_75t_L g137 ( 
.A1(n_133),
.A2(n_131),
.B(n_129),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_137),
.A2(n_129),
.B(n_105),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_127),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_140),
.A2(n_139),
.B1(n_138),
.B2(n_96),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_135),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_141),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_145),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_143),
.B(n_144),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_104),
.C(n_106),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_104),
.C(n_32),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_120),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_107),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_150),
.A2(n_151),
.B(n_148),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_29),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_151),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_28),
.C(n_37),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_154),
.A2(n_126),
.B1(n_25),
.B2(n_31),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_24),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_20),
.C(n_35),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_19),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_33),
.B(n_34),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_18),
.C(n_40),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_17),
.C(n_44),
.Y(n_161)
);

O2A1O1Ixp33_ASAP7_75t_SL g162 ( 
.A1(n_161),
.A2(n_16),
.B(n_15),
.C(n_14),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_8),
.B(n_9),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_163),
.A2(n_9),
.B(n_11),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_11),
.Y(n_165)
);


endmodule