module real_jpeg_15733_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_16),
.B1(n_20),
.B2(n_21),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_1),
.B(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_1),
.B(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_1),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_1),
.B(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g131 ( 
.A(n_2),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_2),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g202 ( 
.A(n_2),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_3),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_3),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_3),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_3),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_3),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_3),
.B(n_271),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_3),
.B(n_301),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_4),
.Y(n_216)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_5),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_5),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g151 ( 
.A(n_5),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_5),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_6),
.B(n_127),
.Y(n_126)
);

AND2x4_ASAP7_75t_SL g166 ( 
.A(n_6),
.B(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_7),
.Y(n_125)
);

BUFx4f_ASAP7_75t_L g330 ( 
.A(n_7),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_8),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_8),
.B(n_102),
.Y(n_101)
);

AOI22x1_ASAP7_75t_SL g129 ( 
.A1(n_8),
.A2(n_17),
.B1(n_130),
.B2(n_132),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_8),
.B(n_161),
.Y(n_160)
);

AOI31xp33_ASAP7_75t_L g197 ( 
.A1(n_8),
.A2(n_129),
.A3(n_198),
.B(n_203),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_8),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_8),
.B(n_283),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_8),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_8),
.B(n_171),
.Y(n_311)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_9),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_9),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_9),
.B(n_183),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_9),
.B(n_201),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_10),
.B(n_171),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_11),
.B(n_65),
.Y(n_64)
);

AND2x4_ASAP7_75t_SL g93 ( 
.A(n_11),
.B(n_94),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_11),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_11),
.B(n_118),
.Y(n_117)
);

AND2x4_ASAP7_75t_L g143 ( 
.A(n_11),
.B(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_11),
.B(n_210),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_11),
.B(n_55),
.Y(n_272)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_12),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_13),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_13),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_13),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_13),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_13),
.B(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_13),
.B(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_13),
.B(n_328),
.Y(n_327)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_14),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_14),
.Y(n_99)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_14),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_14),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_15),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_15),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_17),
.B(n_123),
.Y(n_122)
);

NAND2x1_ASAP7_75t_L g148 ( 
.A(n_17),
.B(n_149),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_17),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_18),
.Y(n_92)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_18),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_223),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_188),
.B(n_221),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_24),
.B(n_189),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_111),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_73),
.C(n_96),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_26),
.B(n_191),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_47),
.C(n_58),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

XNOR2x1_ASAP7_75t_L g246 ( 
.A(n_28),
.B(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_35),
.Y(n_28)
);

MAJx2_ASAP7_75t_L g137 ( 
.A(n_29),
.B(n_40),
.C(n_46),
.Y(n_137)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_31),
.Y(n_281)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_34),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_40),
.B1(n_45),
.B2(n_46),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_36),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_39),
.Y(n_181)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_42),
.Y(n_299)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

XNOR2x1_ASAP7_75t_L g247 ( 
.A(n_47),
.B(n_58),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_53),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_48),
.B(n_53),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_51),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_57),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_64),
.C(n_69),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_59),
.A2(n_64),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_59),
.Y(n_233)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_64),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_64),
.A2(n_234),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_64),
.B(n_313),
.C(n_317),
.Y(n_337)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_69),
.B(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_73),
.B(n_96),
.Y(n_191)
);

XOR2x2_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_85),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_80),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_75),
.B(n_85),
.C(n_153),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_78),
.Y(n_206)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_80),
.Y(n_153)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_83),
.Y(n_285)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_90),
.C(n_93),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_86),
.A2(n_93),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_86),
.Y(n_196)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_90),
.B(n_194),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_93),
.Y(n_195)
);

XNOR2x1_ASAP7_75t_L g293 ( 
.A(n_93),
.B(n_294),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_95),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_100),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_97),
.B(n_101),
.C(n_109),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_104),
.B1(n_109),
.B2(n_110),
.Y(n_100)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_104),
.A2(n_109),
.B1(n_237),
.B2(n_289),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_105),
.Y(n_109)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_109),
.B(n_237),
.C(n_241),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_156),
.B1(n_186),
.B2(n_187),
.Y(n_111)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_112),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_138),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_128),
.C(n_137),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_114),
.B(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_121),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_122),
.C(n_126),
.Y(n_140)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_119),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.Y(n_121)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_125),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_125),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_127),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_128),
.A2(n_129),
.B1(n_137),
.B2(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g240 ( 
.A(n_136),
.Y(n_240)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_137),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_152),
.B1(n_154),
.B2(n_155),
.Y(n_138)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_147),
.B2(n_148),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_142),
.A2(n_143),
.B1(n_213),
.B2(n_214),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_143),
.B(n_208),
.C(n_213),
.Y(n_207)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVxp67_ASAP7_75t_SL g155 ( 
.A(n_152),
.Y(n_155)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_174),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

AOI22x1_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_170),
.B2(n_173),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx2_ASAP7_75t_SL g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_170),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XOR2x1_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_179),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.C(n_217),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_190),
.B(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_192),
.B(n_218),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_197),
.C(n_207),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_193),
.B(n_197),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_195),
.B(n_280),
.C(n_282),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_208),
.B(n_260),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_212),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_209),
.B(n_212),
.Y(n_263)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_209),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_209),
.A2(n_310),
.B1(n_311),
.B2(n_325),
.Y(n_324)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVxp33_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_250),
.B(n_346),
.Y(n_223)
);

INVxp33_ASAP7_75t_SL g224 ( 
.A(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_248),
.Y(n_225)
);

NOR2xp67_ASAP7_75t_L g347 ( 
.A(n_226),
.B(n_248),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.C(n_246),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_227),
.B(n_344),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_230),
.B(n_246),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_235),
.C(n_244),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_231),
.B(n_275),
.Y(n_274)
);

INVxp33_ASAP7_75t_SL g235 ( 
.A(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_236),
.B(n_245),
.Y(n_275)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_237),
.Y(n_289)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_240),
.Y(n_239)
);

XOR2x1_ASAP7_75t_L g287 ( 
.A(n_241),
.B(n_288),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_341),
.B(n_345),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_290),
.B(n_340),
.Y(n_253)
);

NAND2xp33_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_276),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_255),
.B(n_276),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_273),
.B2(n_274),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_261),
.B2(n_262),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_258),
.B(n_262),
.C(n_273),
.Y(n_342)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

MAJx2_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.C(n_268),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_264),
.Y(n_278)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g323 ( 
.A(n_267),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_272),
.Y(n_268)
);

AO22x1_ASAP7_75t_SL g302 ( 
.A1(n_269),
.A2(n_270),
.B1(n_272),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_272),
.Y(n_303)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_279),
.C(n_286),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_277),
.B(n_305),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_279),
.B(n_287),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_282),
.Y(n_294)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI21x1_ASAP7_75t_SL g290 ( 
.A1(n_291),
.A2(n_306),
.B(n_339),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_304),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g339 ( 
.A(n_292),
.B(n_304),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_295),
.C(n_302),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_293),
.B(n_335),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_295),
.A2(n_296),
.B1(n_302),
.B2(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_300),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_297),
.B(n_300),
.Y(n_314)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_302),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_303),
.B(n_327),
.Y(n_326)
);

AOI21x1_ASAP7_75t_SL g306 ( 
.A1(n_307),
.A2(n_333),
.B(n_338),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_308),
.A2(n_320),
.B(n_332),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_312),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_309),
.B(n_312),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_311),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_315),
.B2(n_316),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_326),
.B(n_331),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_324),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_324),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_334),
.B(n_337),
.Y(n_333)
);

NOR2x1_ASAP7_75t_SL g338 ( 
.A(n_334),
.B(n_337),
.Y(n_338)
);

NOR2xp67_ASAP7_75t_SL g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_342),
.B(n_343),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);


endmodule