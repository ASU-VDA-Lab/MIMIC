module fake_jpeg_13998_n_169 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_169);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx2_ASAP7_75t_SL g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_34),
.B(n_35),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_1),
.Y(n_35)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_27),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_36),
.B(n_42),
.Y(n_82)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_30),
.B(n_9),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_43),
.Y(n_62)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_16),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_16),
.B(n_25),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_45),
.B(n_58),
.Y(n_74)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_46),
.B(n_48),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_50),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_49),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_52),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

OA21x2_ASAP7_75t_L g53 ( 
.A1(n_16),
.A2(n_1),
.B(n_3),
.Y(n_53)
);

O2A1O1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_34),
.B(n_35),
.C(n_20),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_27),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_54),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_56),
.Y(n_73)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_59),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_18),
.B(n_22),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_10),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_22),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_80),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_23),
.C(n_31),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_76),
.C(n_87),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_68),
.A2(n_84),
.B1(n_85),
.B2(n_87),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_53),
.A2(n_23),
.B(n_31),
.C(n_28),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_72),
.B(n_89),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_39),
.B(n_48),
.C(n_52),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_32),
.B1(n_28),
.B2(n_24),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_32),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_24),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_75),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_57),
.A2(n_27),
.B1(n_4),
.B2(n_6),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_47),
.A2(n_3),
.B1(n_6),
.B2(n_8),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_86),
.B(n_88),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_47),
.A2(n_10),
.B1(n_50),
.B2(n_36),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_54),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_60),
.A2(n_26),
.B1(n_16),
.B2(n_12),
.Y(n_89)
);

AOI32xp33_ASAP7_75t_L g92 ( 
.A1(n_80),
.A2(n_61),
.A3(n_81),
.B1(n_68),
.B2(n_74),
.Y(n_92)
);

AND2x6_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_82),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_62),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_93),
.B(n_97),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_65),
.B(n_67),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_111),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_91),
.A2(n_72),
.B1(n_82),
.B2(n_64),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_102),
.A2(n_110),
.B1(n_82),
.B2(n_69),
.Y(n_112)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_108),
.B(n_109),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_67),
.B(n_63),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_76),
.A2(n_70),
.B1(n_73),
.B2(n_79),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_75),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_101),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_95),
.Y(n_127)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_123),
.Y(n_136)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_105),
.A2(n_91),
.B(n_63),
.C(n_66),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_124),
.A2(n_126),
.B(n_96),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_90),
.B(n_71),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_128),
.Y(n_141)
);

BUFx12f_ASAP7_75t_SL g128 ( 
.A(n_124),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_129),
.A2(n_130),
.B(n_131),
.Y(n_138)
);

AO22x1_ASAP7_75t_L g130 ( 
.A1(n_119),
.A2(n_107),
.B1(n_96),
.B2(n_108),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_110),
.B1(n_99),
.B2(n_95),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_132),
.A2(n_116),
.B1(n_114),
.B2(n_118),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_103),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_125),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_115),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_135),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_118),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_100),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_122),
.Y(n_143)
);

MAJx2_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_138),
.C(n_141),
.Y(n_150)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_142),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_143),
.A2(n_146),
.B(n_117),
.Y(n_147)
);

AOI22x1_ASAP7_75t_L g144 ( 
.A1(n_128),
.A2(n_131),
.B1(n_130),
.B2(n_137),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_144),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_120),
.C(n_77),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_117),
.B(n_94),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_147),
.B(n_149),
.Y(n_157)
);

A2O1A1O1Ixp25_ASAP7_75t_L g149 ( 
.A1(n_138),
.A2(n_133),
.B(n_129),
.C(n_101),
.D(n_106),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_150),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_120),
.C(n_104),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_153),
.Y(n_156)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_148),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_154),
.A2(n_155),
.B(n_149),
.Y(n_160)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_153),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_157),
.B(n_144),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_159),
.B(n_160),
.Y(n_163)
);

AOI22x1_ASAP7_75t_SL g161 ( 
.A1(n_158),
.A2(n_151),
.B1(n_150),
.B2(n_146),
.Y(n_161)
);

NOR2x1_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_156),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_158),
.A2(n_139),
.B(n_140),
.Y(n_162)
);

NOR2xp67_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_156),
.Y(n_164)
);

AOI21x1_ASAP7_75t_L g166 ( 
.A1(n_164),
.A2(n_165),
.B(n_77),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_166),
.B(n_167),
.Y(n_168)
);

INVxp33_ASAP7_75t_L g167 ( 
.A(n_163),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_165),
.Y(n_169)
);


endmodule