module real_aes_17366_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_502;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
AND2x4_ASAP7_75t_L g114 ( .A(n_0), .B(n_115), .Y(n_114) );
AOI22xp5_ASAP7_75t_L g280 ( .A1(n_1), .A2(n_4), .B1(n_281), .B2(n_282), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_2), .A2(n_43), .B1(n_138), .B2(n_208), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_3), .A2(n_23), .B1(n_208), .B2(n_217), .Y(n_225) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_5), .A2(n_15), .B1(n_514), .B2(n_560), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g165 ( .A1(n_6), .A2(n_62), .B1(n_166), .B2(n_167), .Y(n_165) );
AOI22xp5_ASAP7_75t_L g137 ( .A1(n_7), .A2(n_16), .B1(n_138), .B2(n_140), .Y(n_137) );
INVx1_ASAP7_75t_L g115 ( .A(n_8), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_9), .Y(n_216) );
CKINVDCx5p33_ASAP7_75t_R g527 ( .A(n_10), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_11), .A2(n_17), .B1(n_515), .B2(n_550), .Y(n_549) );
BUFx2_ASAP7_75t_L g118 ( .A(n_12), .Y(n_118) );
OR2x2_ASAP7_75t_L g817 ( .A(n_12), .B(n_38), .Y(n_817) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_13), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g562 ( .A(n_14), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_18), .A2(n_102), .B1(n_282), .B2(n_514), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_19), .A2(n_39), .B1(n_174), .B2(n_531), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_20), .B(n_173), .Y(n_528) );
OAI21x1_ASAP7_75t_L g150 ( .A1(n_21), .A2(n_59), .B(n_151), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_22), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g584 ( .A(n_24), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_25), .B(n_143), .Y(n_237) );
INVx4_ASAP7_75t_R g190 ( .A(n_26), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g830 ( .A1(n_27), .A2(n_55), .B1(n_831), .B2(n_832), .Y(n_830) );
CKINVDCx5p33_ASAP7_75t_R g831 ( .A(n_27), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_28), .A2(n_47), .B1(n_145), .B2(n_279), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_29), .A2(n_54), .B1(n_145), .B2(n_514), .Y(n_567) );
CKINVDCx5p33_ASAP7_75t_R g507 ( .A(n_30), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_31), .B(n_531), .Y(n_530) );
CKINVDCx5p33_ASAP7_75t_R g520 ( .A(n_32), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_33), .B(n_208), .Y(n_243) );
INVx1_ASAP7_75t_L g286 ( .A(n_34), .Y(n_286) );
A2O1A1Ixp33_ASAP7_75t_SL g214 ( .A1(n_35), .A2(n_138), .B(n_142), .C(n_215), .Y(n_214) );
AOI22xp33_ASAP7_75t_L g226 ( .A1(n_36), .A2(n_56), .B1(n_138), .B2(n_145), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_37), .A2(n_105), .B1(n_121), .B2(n_854), .Y(n_104) );
HB1xp67_ASAP7_75t_L g120 ( .A(n_38), .Y(n_120) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_40), .A2(n_87), .B1(n_138), .B2(n_504), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g801 ( .A1(n_41), .A2(n_80), .B1(n_802), .B2(n_803), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_41), .Y(n_802) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_42), .Y(n_211) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_44), .A2(n_46), .B1(n_138), .B2(n_140), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_45), .A2(n_60), .B1(n_514), .B2(n_566), .Y(n_582) );
INVx1_ASAP7_75t_L g240 ( .A(n_48), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_49), .B(n_138), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g843 ( .A1(n_50), .A2(n_844), .B(n_851), .Y(n_843) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_51), .Y(n_259) );
INVx2_ASAP7_75t_L g812 ( .A(n_52), .Y(n_812) );
INVx1_ASAP7_75t_L g110 ( .A(n_53), .Y(n_110) );
BUFx3_ASAP7_75t_L g815 ( .A(n_53), .Y(n_815) );
INVx1_ASAP7_75t_L g832 ( .A(n_55), .Y(n_832) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_57), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g144 ( .A1(n_58), .A2(n_88), .B1(n_138), .B2(n_145), .Y(n_144) );
OAI22xp5_ASAP7_75t_SL g799 ( .A1(n_61), .A2(n_800), .B1(n_801), .B2(n_804), .Y(n_799) );
CKINVDCx5p33_ASAP7_75t_R g804 ( .A(n_61), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_63), .A2(n_75), .B1(n_279), .B2(n_566), .Y(n_565) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_64), .Y(n_156) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_65), .A2(n_78), .B1(n_138), .B2(n_140), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_66), .A2(n_100), .B1(n_514), .B2(n_515), .Y(n_513) );
INVx1_ASAP7_75t_L g151 ( .A(n_67), .Y(n_151) );
AND2x4_ASAP7_75t_L g153 ( .A(n_68), .B(n_154), .Y(n_153) );
AOI22xp33_ASAP7_75t_L g278 ( .A1(n_69), .A2(n_90), .B1(n_145), .B2(n_279), .Y(n_278) );
AO22x1_ASAP7_75t_L g171 ( .A1(n_70), .A2(n_76), .B1(n_172), .B2(n_174), .Y(n_171) );
INVx1_ASAP7_75t_L g154 ( .A(n_71), .Y(n_154) );
AND2x2_ASAP7_75t_L g218 ( .A(n_72), .B(n_219), .Y(n_218) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_73), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_74), .B(n_166), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_77), .B(n_208), .Y(n_260) );
INVx2_ASAP7_75t_L g143 ( .A(n_79), .Y(n_143) );
INVx1_ASAP7_75t_L g803 ( .A(n_80), .Y(n_803) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_81), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_82), .B(n_219), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_83), .A2(n_99), .B1(n_145), .B2(n_166), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g569 ( .A(n_84), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_85), .B(n_149), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g542 ( .A(n_86), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_89), .B(n_219), .Y(n_534) );
CKINVDCx5p33_ASAP7_75t_R g553 ( .A(n_91), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_92), .B(n_219), .Y(n_256) );
HB1xp67_ASAP7_75t_L g835 ( .A(n_92), .Y(n_835) );
INVx1_ASAP7_75t_L g113 ( .A(n_93), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_93), .B(n_841), .Y(n_840) );
OAI22xp5_ASAP7_75t_L g797 ( .A1(n_94), .A2(n_798), .B1(n_805), .B2(n_806), .Y(n_797) );
CKINVDCx5p33_ASAP7_75t_R g805 ( .A(n_94), .Y(n_805) );
NAND2xp33_ASAP7_75t_L g532 ( .A(n_95), .B(n_173), .Y(n_532) );
A2O1A1Ixp33_ASAP7_75t_L g185 ( .A1(n_96), .A2(n_147), .B(n_166), .C(n_186), .Y(n_185) );
CKINVDCx16_ASAP7_75t_R g852 ( .A(n_97), .Y(n_852) );
AND2x2_ASAP7_75t_L g195 ( .A(n_98), .B(n_196), .Y(n_195) );
AOI22xp33_ASAP7_75t_SL g834 ( .A1(n_101), .A2(n_835), .B1(n_836), .B2(n_837), .Y(n_834) );
INVxp67_ASAP7_75t_SL g836 ( .A(n_101), .Y(n_836) );
NAND2xp33_ASAP7_75t_L g264 ( .A(n_103), .B(n_191), .Y(n_264) );
INVx3_ASAP7_75t_SL g854 ( .A(n_105), .Y(n_854) );
INVx4_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
OR2x6_ASAP7_75t_L g106 ( .A(n_107), .B(n_116), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
NOR2x1p5_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
AND3x2_ASAP7_75t_L g828 ( .A(n_109), .B(n_112), .C(n_816), .Y(n_828) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g841 ( .A(n_110), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_114), .Y(n_111) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g492 ( .A(n_113), .Y(n_492) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
INVxp33_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
OR2x6_ASAP7_75t_L g121 ( .A(n_122), .B(n_818), .Y(n_121) );
NOR2xp33_ASAP7_75t_L g122 ( .A(n_123), .B(n_808), .Y(n_122) );
AOI22xp33_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_796), .B1(n_797), .B2(n_807), .Y(n_123) );
INVx2_ASAP7_75t_L g807 ( .A(n_124), .Y(n_807) );
AO22x2_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_489), .B1(n_490), .B2(n_493), .Y(n_124) );
INVx1_ASAP7_75t_SL g125 ( .A(n_126), .Y(n_125) );
NOR2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_403), .Y(n_126) );
NAND4xp75_ASAP7_75t_L g127 ( .A(n_128), .B(n_308), .C(n_350), .D(n_374), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OAI211xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_197), .B(n_245), .C(n_287), .Y(n_129) );
INVxp67_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
BUFx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g394 ( .A(n_132), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g488 ( .A(n_132), .B(n_425), .Y(n_488) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_158), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g303 ( .A(n_134), .B(n_255), .Y(n_303) );
AND2x2_ASAP7_75t_L g344 ( .A(n_134), .B(n_305), .Y(n_344) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_L g251 ( .A(n_135), .B(n_180), .Y(n_251) );
OR2x2_ASAP7_75t_L g269 ( .A(n_135), .B(n_180), .Y(n_269) );
INVx2_ASAP7_75t_L g295 ( .A(n_135), .Y(n_295) );
AND2x2_ASAP7_75t_L g325 ( .A(n_135), .B(n_255), .Y(n_325) );
AND2x2_ASAP7_75t_L g354 ( .A(n_135), .B(n_179), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_135), .B(n_306), .Y(n_390) );
AO31x2_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_148), .A3(n_152), .B(n_155), .Y(n_135) );
OAI22x1_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_141), .B1(n_144), .B2(n_146), .Y(n_136) );
INVx4_ASAP7_75t_L g140 ( .A(n_138), .Y(n_140) );
INVx1_ASAP7_75t_L g515 ( .A(n_138), .Y(n_515) );
INVx1_ASAP7_75t_L g566 ( .A(n_138), .Y(n_566) );
INVx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_139), .Y(n_145) );
INVx1_ASAP7_75t_L g166 ( .A(n_139), .Y(n_166) );
INVx1_ASAP7_75t_L g168 ( .A(n_139), .Y(n_168) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_139), .Y(n_173) );
INVx1_ASAP7_75t_L g175 ( .A(n_139), .Y(n_175) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_139), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_139), .Y(n_192) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_139), .Y(n_208) );
INVx1_ASAP7_75t_L g210 ( .A(n_139), .Y(n_210) );
INVx2_ASAP7_75t_L g217 ( .A(n_139), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_L g258 ( .A1(n_140), .A2(n_259), .B(n_260), .C(n_261), .Y(n_258) );
O2A1O1Ixp5_ASAP7_75t_L g526 ( .A1(n_140), .A2(n_142), .B(n_527), .C(n_528), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g224 ( .A1(n_141), .A2(n_162), .B1(n_225), .B2(n_226), .Y(n_224) );
OAI22xp5_ASAP7_75t_L g277 ( .A1(n_141), .A2(n_146), .B1(n_278), .B2(n_280), .Y(n_277) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_141), .A2(n_146), .B1(n_503), .B2(n_505), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_141), .A2(n_513), .B1(n_516), .B2(n_517), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_141), .A2(n_530), .B(n_532), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_141), .A2(n_538), .B1(n_539), .B2(n_540), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_141), .A2(n_517), .B1(n_549), .B2(n_551), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_141), .A2(n_539), .B1(n_558), .B2(n_559), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_141), .A2(n_539), .B1(n_565), .B2(n_567), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_141), .A2(n_539), .B1(n_581), .B2(n_582), .Y(n_580) );
INVx6_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_142), .B(n_171), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_142), .A2(n_264), .B(n_265), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_L g307 ( .A1(n_142), .A2(n_161), .B(n_171), .C(n_177), .Y(n_307) );
BUFx8_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g147 ( .A(n_143), .Y(n_147) );
INVx2_ASAP7_75t_L g164 ( .A(n_143), .Y(n_164) );
INVx1_ASAP7_75t_L g213 ( .A(n_143), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_145), .B(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g281 ( .A(n_145), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_146), .B(n_189), .Y(n_188) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_SL g517 ( .A(n_147), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_148), .B(n_569), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_148), .B(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g157 ( .A(n_149), .Y(n_157) );
OAI21xp33_ASAP7_75t_L g177 ( .A1(n_149), .A2(n_169), .B(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g183 ( .A(n_149), .Y(n_183) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_150), .Y(n_220) );
INVx2_ASAP7_75t_L g194 ( .A(n_152), .Y(n_194) );
AO31x2_ASAP7_75t_L g536 ( .A1(n_152), .A2(n_227), .A3(n_537), .B(n_541), .Y(n_536) );
AO31x2_ASAP7_75t_L g547 ( .A1(n_152), .A2(n_203), .A3(n_548), .B(n_552), .Y(n_547) );
AO31x2_ASAP7_75t_L g556 ( .A1(n_152), .A2(n_501), .A3(n_557), .B(n_561), .Y(n_556) );
BUFx10_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g178 ( .A(n_153), .Y(n_178) );
BUFx10_ASAP7_75t_L g228 ( .A(n_153), .Y(n_228) );
INVx1_ASAP7_75t_L g284 ( .A(n_153), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
INVx2_ASAP7_75t_L g196 ( .A(n_157), .Y(n_196) );
BUFx2_ASAP7_75t_L g203 ( .A(n_157), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_157), .B(n_230), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_157), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g367 ( .A(n_158), .B(n_296), .Y(n_367) );
INVx2_ASAP7_75t_L g462 ( .A(n_158), .Y(n_462) );
AND2x2_ASAP7_75t_L g158 ( .A(n_159), .B(n_179), .Y(n_158) );
INVx2_ASAP7_75t_L g250 ( .A(n_159), .Y(n_250) );
AND2x4_ASAP7_75t_L g293 ( .A(n_159), .B(n_180), .Y(n_293) );
AOI21x1_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_170), .B(n_176), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
OAI21x1_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_165), .B(n_169), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_162), .A2(n_242), .B(n_243), .Y(n_241) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g539 ( .A(n_163), .Y(n_539) );
BUFx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g262 ( .A(n_164), .Y(n_262) );
INVx1_ASAP7_75t_L g550 ( .A(n_167), .Y(n_550) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_168), .B(n_187), .Y(n_186) );
INVxp67_ASAP7_75t_SL g172 ( .A(n_173), .Y(n_172) );
INVx3_ASAP7_75t_L g514 ( .A(n_173), .Y(n_514) );
OAI21xp33_ASAP7_75t_SL g236 ( .A1(n_174), .A2(n_237), .B(n_238), .Y(n_236) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_178), .A2(n_205), .B(n_214), .Y(n_204) );
AND2x2_ASAP7_75t_L g452 ( .A(n_179), .B(n_250), .Y(n_452) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g316 ( .A(n_180), .Y(n_316) );
AND2x2_ASAP7_75t_L g373 ( .A(n_180), .B(n_255), .Y(n_373) );
AND2x2_ASAP7_75t_L g388 ( .A(n_180), .B(n_296), .Y(n_388) );
AND2x2_ASAP7_75t_L g410 ( .A(n_180), .B(n_250), .Y(n_410) );
AO21x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_184), .B(n_195), .Y(n_180) );
AO31x2_ASAP7_75t_L g563 ( .A1(n_181), .A2(n_283), .A3(n_564), .B(n_568), .Y(n_563) );
AO31x2_ASAP7_75t_L g579 ( .A1(n_181), .A2(n_518), .A3(n_580), .B(n_583), .Y(n_579) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_183), .B(n_507), .Y(n_506) );
NOR2xp33_ASAP7_75t_SL g552 ( .A(n_183), .B(n_553), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_188), .B(n_194), .Y(n_184) );
OAI22xp33_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B1(n_192), .B2(n_193), .Y(n_189) );
INVx2_ASAP7_75t_L g279 ( .A(n_191), .Y(n_279) );
INVx1_ASAP7_75t_L g531 ( .A(n_191), .Y(n_531) );
INVx1_ASAP7_75t_L g560 ( .A(n_192), .Y(n_560) );
INVx1_ASAP7_75t_L g518 ( .A(n_194), .Y(n_518) );
OAI211xp5_ASAP7_75t_SL g457 ( .A1(n_197), .A2(n_458), .B(n_460), .C(n_467), .Y(n_457) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_231), .Y(n_198) );
INVxp67_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
OR2x2_ASAP7_75t_L g444 ( .A(n_200), .B(n_380), .Y(n_444) );
OR2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_221), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_201), .B(n_233), .Y(n_343) );
INVxp67_ASAP7_75t_L g357 ( .A(n_201), .Y(n_357) );
AND2x2_ASAP7_75t_L g377 ( .A(n_201), .B(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_201), .B(n_290), .Y(n_384) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g273 ( .A(n_202), .Y(n_273) );
AOI21x1_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B(n_218), .Y(n_202) );
AO31x2_ASAP7_75t_L g276 ( .A1(n_203), .A2(n_277), .A3(n_283), .B(n_285), .Y(n_276) );
AO31x2_ASAP7_75t_L g511 ( .A1(n_203), .A2(n_512), .A3(n_518), .B(n_519), .Y(n_511) );
OAI21xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_209), .B(n_212), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
INVx2_ASAP7_75t_L g282 ( .A(n_210), .Y(n_282) );
BUFx4f_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_213), .B(n_240), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_216), .B(n_217), .Y(n_215) );
INVx2_ASAP7_75t_SL g504 ( .A(n_217), .Y(n_504) );
INVx2_ASAP7_75t_L g227 ( .A(n_219), .Y(n_227) );
NOR2x1_ASAP7_75t_L g266 ( .A(n_219), .B(n_267), .Y(n_266) );
INVx4_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g244 ( .A(n_220), .B(n_228), .Y(n_244) );
BUFx3_ASAP7_75t_L g501 ( .A(n_220), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_220), .B(n_520), .Y(n_519) );
INVx2_ASAP7_75t_SL g524 ( .A(n_220), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_220), .B(n_542), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_220), .B(n_562), .Y(n_561) );
OR2x2_ASAP7_75t_L g318 ( .A(n_221), .B(n_300), .Y(n_318) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
OR2x2_ASAP7_75t_L g366 ( .A(n_222), .B(n_273), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_222), .B(n_276), .Y(n_372) );
INVx2_ASAP7_75t_SL g222 ( .A(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g272 ( .A(n_223), .B(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g341 ( .A(n_223), .B(n_276), .Y(n_341) );
BUFx2_ASAP7_75t_L g348 ( .A(n_223), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_223), .B(n_276), .Y(n_428) );
AO31x2_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_227), .A3(n_228), .B(n_229), .Y(n_223) );
INVx1_ASAP7_75t_L g267 ( .A(n_228), .Y(n_267) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x4_ASAP7_75t_L g358 ( .A(n_232), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g487 ( .A(n_232), .B(n_272), .Y(n_487) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx3_ASAP7_75t_L g290 ( .A(n_233), .Y(n_290) );
AND2x2_ASAP7_75t_L g301 ( .A(n_233), .B(n_276), .Y(n_301) );
AND2x2_ASAP7_75t_L g347 ( .A(n_233), .B(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g380 ( .A(n_233), .B(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_233), .B(n_291), .Y(n_397) );
AND2x2_ASAP7_75t_L g436 ( .A(n_233), .B(n_437), .Y(n_436) );
AND2x4_ASAP7_75t_L g233 ( .A(n_234), .B(n_235), .Y(n_233) );
OAI21xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_241), .B(n_244), .Y(n_235) );
OAI21xp5_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_252), .B(n_270), .Y(n_245) );
INVx2_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_247), .A2(n_415), .B1(n_416), .B2(n_418), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_248), .B(n_251), .Y(n_247) );
AND2x2_ASAP7_75t_L g412 ( .A(n_248), .B(n_303), .Y(n_412) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g327 ( .A(n_249), .Y(n_327) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g476 ( .A(n_250), .B(n_296), .Y(n_476) );
AND2x2_ASAP7_75t_L g440 ( .A(n_251), .B(n_335), .Y(n_440) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_268), .Y(n_252) );
OR2x2_ASAP7_75t_L g337 ( .A(n_253), .B(n_314), .Y(n_337) );
OR2x2_ASAP7_75t_L g449 ( .A(n_253), .B(n_269), .Y(n_449) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g312 ( .A(n_254), .Y(n_312) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g296 ( .A(n_255), .Y(n_296) );
BUFx3_ASAP7_75t_L g378 ( .A(n_255), .Y(n_378) );
NAND2x1p5_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
OAI21x1_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_263), .B(n_266), .Y(n_257) );
INVx2_ASAP7_75t_SL g261 ( .A(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g446 ( .A(n_269), .B(n_305), .Y(n_446) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
AND2x2_ASAP7_75t_L g288 ( .A(n_272), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g329 ( .A(n_272), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g466 ( .A(n_272), .Y(n_466) );
INVx1_ASAP7_75t_L g485 ( .A(n_272), .Y(n_485) );
INVx2_ASAP7_75t_L g300 ( .A(n_273), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_273), .B(n_276), .Y(n_349) );
INVx1_ASAP7_75t_L g413 ( .A(n_274), .Y(n_413) );
BUFx3_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g474 ( .A(n_275), .Y(n_474) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g291 ( .A(n_276), .Y(n_291) );
INVx1_ASAP7_75t_L g381 ( .A(n_276), .Y(n_381) );
AO31x2_ASAP7_75t_L g500 ( .A1(n_283), .A2(n_501), .A3(n_502), .B(n_506), .Y(n_500) );
INVx2_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
INVx2_ASAP7_75t_SL g533 ( .A(n_284), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_292), .B1(n_297), .B2(n_302), .Y(n_287) );
AND2x4_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx2_ASAP7_75t_L g330 ( .A(n_290), .Y(n_330) );
AND2x2_ASAP7_75t_L g332 ( .A(n_290), .B(n_317), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_290), .B(n_300), .Y(n_392) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx3_ASAP7_75t_L g323 ( .A(n_293), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_293), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g417 ( .A(n_293), .B(n_401), .Y(n_417) );
INVx1_ASAP7_75t_L g321 ( .A(n_294), .Y(n_321) );
AOI222xp33_ASAP7_75t_L g331 ( .A1(n_294), .A2(n_332), .B1(n_333), .B2(n_338), .C1(n_344), .C2(n_345), .Y(n_331) );
OAI21xp33_ASAP7_75t_SL g361 ( .A1(n_294), .A2(n_362), .B(n_363), .Y(n_361) );
AND2x2_ASAP7_75t_L g385 ( .A(n_294), .B(n_304), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_294), .B(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
OR2x2_ASAP7_75t_L g314 ( .A(n_295), .B(n_306), .Y(n_314) );
INVx1_ASAP7_75t_L g402 ( .A(n_295), .Y(n_402) );
BUFx2_ASAP7_75t_L g336 ( .A(n_296), .Y(n_336) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_301), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_299), .B(n_340), .Y(n_369) );
OR2x2_ASAP7_75t_L g481 ( .A(n_299), .B(n_341), .Y(n_481) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x4_ASAP7_75t_L g364 ( .A(n_301), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g479 ( .A(n_301), .Y(n_479) );
OAI31xp33_ASAP7_75t_L g460 ( .A1(n_302), .A2(n_461), .A3(n_463), .B(n_464), .Y(n_460) );
AND2x4_ASAP7_75t_SL g302 ( .A(n_303), .B(n_304), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_303), .B(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_331), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_317), .B(n_319), .Y(n_309) );
NOR2x1_ASAP7_75t_L g310 ( .A(n_311), .B(n_313), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OR2x6_ASAP7_75t_L g430 ( .A(n_312), .B(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx1_ASAP7_75t_L g362 ( .A(n_315), .Y(n_362) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g453 ( .A(n_316), .B(n_390), .Y(n_453) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_318), .A2(n_407), .B1(n_409), .B2(n_411), .Y(n_406) );
A2O1A1Ixp33_ASAP7_75t_L g467 ( .A1(n_318), .A2(n_379), .B(n_441), .C(n_468), .Y(n_467) );
AOI21xp33_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_324), .B(n_328), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND4xp25_ASAP7_75t_L g420 ( .A(n_323), .B(n_421), .C(n_422), .D(n_424), .Y(n_420) );
NAND2x1_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_325), .B(n_327), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_325), .B(n_410), .Y(n_433) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g399 ( .A(n_330), .B(n_359), .Y(n_399) );
NAND2xp33_ASAP7_75t_L g333 ( .A(n_334), .B(n_337), .Y(n_333) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OAI22xp5_ASAP7_75t_L g480 ( .A1(n_337), .A2(n_481), .B1(n_482), .B2(n_484), .Y(n_480) );
AOI221x1_ASAP7_75t_L g419 ( .A1(n_338), .A2(n_420), .B1(n_426), .B2(n_429), .C(n_432), .Y(n_419) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_342), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g359 ( .A(n_341), .Y(n_359) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g371 ( .A(n_343), .B(n_372), .Y(n_371) );
NAND2x1p5_ASAP7_75t_L g434 ( .A(n_344), .B(n_425), .Y(n_434) );
O2A1O1Ixp5_ASAP7_75t_L g447 ( .A1(n_345), .A2(n_429), .B(n_448), .C(n_450), .Y(n_447) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_349), .Y(n_346) );
INVx2_ASAP7_75t_L g396 ( .A(n_348), .Y(n_396) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_360), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_352), .B(n_355), .Y(n_351) );
AOI221xp5_ASAP7_75t_L g439 ( .A1(n_352), .A2(n_370), .B1(n_440), .B2(n_441), .C(n_443), .Y(n_439) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g376 ( .A(n_354), .B(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_354), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g475 ( .A(n_354), .B(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .Y(n_355) );
INVxp67_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
NAND2x1_ASAP7_75t_L g454 ( .A(n_357), .B(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_L g478 ( .A(n_357), .B(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g418 ( .A(n_358), .Y(n_418) );
AOI222xp33_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_364), .B1(n_367), .B2(n_368), .C1(n_370), .C2(n_373), .Y(n_360) );
INVx1_ASAP7_75t_L g445 ( .A(n_364), .Y(n_445) );
INVx1_ASAP7_75t_L g408 ( .A(n_365), .Y(n_408) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g442 ( .A(n_366), .Y(n_442) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
OR2x2_ASAP7_75t_L g383 ( .A(n_372), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g437 ( .A(n_372), .Y(n_437) );
AND2x2_ASAP7_75t_L g400 ( .A(n_373), .B(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_393), .Y(n_374) );
AOI222xp33_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_379), .B1(n_382), .B2(n_385), .C1(n_386), .C2(n_391), .Y(n_375) );
INVx3_ASAP7_75t_L g425 ( .A(n_378), .Y(n_425) );
BUFx2_ASAP7_75t_L g483 ( .A(n_378), .Y(n_483) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g455 ( .A(n_380), .Y(n_455) );
OR2x2_ASAP7_75t_L g465 ( .A(n_380), .B(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
INVx2_ASAP7_75t_SL g423 ( .A(n_388), .Y(n_423) );
AND2x2_ASAP7_75t_L g468 ( .A(n_389), .B(n_425), .Y(n_468) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_390), .Y(n_421) );
INVxp67_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
OR2x2_ASAP7_75t_L g427 ( .A(n_392), .B(n_428), .Y(n_427) );
NOR2x1_ASAP7_75t_L g393 ( .A(n_394), .B(n_398), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
OR2x2_ASAP7_75t_L g484 ( .A(n_397), .B(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
INVx1_ASAP7_75t_L g415 ( .A(n_399), .Y(n_415) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
OR2x2_ASAP7_75t_L g422 ( .A(n_402), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g472 ( .A(n_402), .Y(n_472) );
NAND4xp75_ASAP7_75t_L g403 ( .A(n_404), .B(n_438), .C(n_456), .D(n_469), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_419), .Y(n_404) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_413), .B(n_414), .Y(n_405) );
INVxp33_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_408), .B(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g431 ( .A(n_410), .Y(n_431) );
AND2x2_ASAP7_75t_L g471 ( .A(n_410), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g441 ( .A(n_413), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g459 ( .A(n_424), .Y(n_459) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OAI22xp33_ASAP7_75t_SL g450 ( .A1(n_427), .A2(n_451), .B1(n_453), .B2(n_454), .Y(n_450) );
INVx3_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AOI21xp33_ASAP7_75t_SL g432 ( .A1(n_433), .A2(n_434), .B(n_435), .Y(n_432) );
INVx1_ASAP7_75t_L g463 ( .A(n_434), .Y(n_463) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_447), .Y(n_438) );
AOI21xp5_ASAP7_75t_SL g443 ( .A1(n_444), .A2(n_445), .B(n_446), .Y(n_443) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx3_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_486), .Y(n_469) );
AOI221xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_473), .B1(n_475), .B2(n_477), .C(n_480), .Y(n_470) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx12f_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
CKINVDCx5p33_ASAP7_75t_R g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g849 ( .A(n_492), .B(n_850), .Y(n_849) );
NAND4xp75_ASAP7_75t_L g493 ( .A(n_494), .B(n_636), .C(n_712), .D(n_764), .Y(n_493) );
NAND4xp25_ASAP7_75t_L g833 ( .A(n_494), .B(n_636), .C(n_712), .D(n_764), .Y(n_833) );
AND3x1_ASAP7_75t_L g494 ( .A(n_495), .B(n_609), .C(n_622), .Y(n_494) );
AOI221x1_ASAP7_75t_SL g495 ( .A1(n_496), .A2(n_543), .B1(n_570), .B2(n_574), .C(n_586), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g609 ( .A1(n_496), .A2(n_610), .B(n_612), .C(n_613), .Y(n_609) );
AND2x4_ASAP7_75t_L g496 ( .A(n_497), .B(n_508), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g573 ( .A(n_500), .Y(n_573) );
BUFx2_ASAP7_75t_L g591 ( .A(n_500), .Y(n_591) );
OR2x2_ASAP7_75t_L g633 ( .A(n_500), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g640 ( .A(n_500), .B(n_511), .Y(n_640) );
AND2x4_ASAP7_75t_L g675 ( .A(n_500), .B(n_510), .Y(n_675) );
OR2x2_ASAP7_75t_L g718 ( .A(n_500), .B(n_536), .Y(n_718) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_521), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_510), .B(n_589), .Y(n_588) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_510), .Y(n_605) );
INVx2_ASAP7_75t_L g632 ( .A(n_510), .Y(n_632) );
INVx3_ASAP7_75t_L g645 ( .A(n_510), .Y(n_645) );
AND2x2_ASAP7_75t_L g763 ( .A(n_510), .B(n_592), .Y(n_763) );
INVx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g572 ( .A(n_511), .B(n_573), .Y(n_572) );
BUFx2_ASAP7_75t_L g628 ( .A(n_511), .Y(n_628) );
INVxp67_ASAP7_75t_SL g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g648 ( .A(n_522), .Y(n_648) );
INVx1_ASAP7_75t_L g775 ( .A(n_522), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_535), .Y(n_522) );
AND2x2_ASAP7_75t_L g571 ( .A(n_523), .B(n_536), .Y(n_571) );
INVx1_ASAP7_75t_L g634 ( .A(n_523), .Y(n_634) );
OAI21x1_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_525), .B(n_534), .Y(n_523) );
OAI21x1_ASAP7_75t_L g593 ( .A1(n_524), .A2(n_525), .B(n_534), .Y(n_593) );
OAI21x1_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_529), .B(n_533), .Y(n_525) );
INVx2_ASAP7_75t_L g589 ( .A(n_535), .Y(n_589) );
AND2x2_ASAP7_75t_L g641 ( .A(n_535), .B(n_592), .Y(n_641) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g603 ( .A(n_536), .Y(n_603) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_536), .Y(n_663) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_545), .A2(n_635), .B1(n_639), .B2(n_642), .Y(n_638) );
AND2x4_ASAP7_75t_L g545 ( .A(n_546), .B(n_554), .Y(n_545) );
INVx1_ASAP7_75t_L g656 ( .A(n_546), .Y(n_656) );
BUFx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g576 ( .A(n_547), .B(n_556), .Y(n_576) );
AND2x2_ASAP7_75t_L g607 ( .A(n_547), .B(n_563), .Y(n_607) );
INVx4_ASAP7_75t_SL g618 ( .A(n_547), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_547), .B(n_652), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_547), .B(n_791), .Y(n_790) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OR2x2_ASAP7_75t_L g689 ( .A(n_555), .B(n_667), .Y(n_689) );
OR2x2_ASAP7_75t_L g722 ( .A(n_555), .B(n_704), .Y(n_722) );
OR2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_563), .Y(n_555) );
INVx2_ASAP7_75t_L g596 ( .A(n_556), .Y(n_596) );
INVx1_ASAP7_75t_L g601 ( .A(n_556), .Y(n_601) );
AND2x2_ASAP7_75t_L g608 ( .A(n_556), .B(n_578), .Y(n_608) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_556), .Y(n_624) );
INVx1_ASAP7_75t_L g652 ( .A(n_556), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_556), .B(n_688), .Y(n_687) );
INVx2_ASAP7_75t_L g585 ( .A(n_563), .Y(n_585) );
AND2x4_ASAP7_75t_L g595 ( .A(n_563), .B(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g621 ( .A(n_563), .Y(n_621) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_563), .Y(n_698) );
INVx1_ASAP7_75t_L g791 ( .A(n_563), .Y(n_791) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_571), .B(n_644), .Y(n_711) );
AND2x2_ASAP7_75t_L g724 ( .A(n_571), .B(n_640), .Y(n_724) );
AND2x2_ASAP7_75t_L g794 ( .A(n_571), .B(n_645), .Y(n_794) );
AND2x4_ASAP7_75t_L g629 ( .A(n_573), .B(n_592), .Y(n_629) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
AND2x2_ASAP7_75t_L g696 ( .A(n_576), .B(n_697), .Y(n_696) );
INVx2_ASAP7_75t_L g710 ( .A(n_576), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_576), .B(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g612 ( .A(n_577), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_577), .B(n_650), .Y(n_649) );
AOI211xp5_ASAP7_75t_L g706 ( .A1(n_577), .A2(n_707), .B(n_710), .C(n_711), .Y(n_706) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_585), .Y(n_577) );
AND2x2_ASAP7_75t_L g677 ( .A(n_578), .B(n_618), .Y(n_677) );
INVx3_ASAP7_75t_L g704 ( .A(n_578), .Y(n_704) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g599 ( .A(n_579), .Y(n_599) );
AND2x4_ASAP7_75t_L g625 ( .A(n_579), .B(n_585), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_585), .B(n_618), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_594), .B1(n_602), .B2(n_606), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .Y(n_587) );
INVx1_ASAP7_75t_L g743 ( .A(n_588), .Y(n_743) );
AND2x4_ASAP7_75t_L g654 ( .A(n_589), .B(n_634), .Y(n_654) );
INVx1_ASAP7_75t_L g674 ( .A(n_589), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_591), .A2(n_647), .B1(n_657), .B2(n_659), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_591), .B(n_648), .Y(n_705) );
NAND2x1_ASAP7_75t_L g762 ( .A(n_591), .B(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g777 ( .A(n_591), .Y(n_777) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
BUFx2_ASAP7_75t_L g716 ( .A(n_593), .Y(n_716) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_595), .B(n_597), .Y(n_594) );
AND2x2_ASAP7_75t_L g635 ( .A(n_595), .B(n_617), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_595), .B(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g676 ( .A(n_595), .B(n_677), .Y(n_676) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_595), .Y(n_750) );
NAND2x1p5_ASAP7_75t_L g757 ( .A(n_595), .B(n_658), .Y(n_757) );
AND2x4_ASAP7_75t_L g780 ( .A(n_595), .B(n_708), .Y(n_780) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .Y(n_597) );
INVx3_ASAP7_75t_L g658 ( .A(n_598), .Y(n_658) );
AND2x2_ASAP7_75t_L g670 ( .A(n_598), .B(n_663), .Y(n_670) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g620 ( .A(n_599), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g668 ( .A(n_599), .Y(n_668) );
INVx1_ASAP7_75t_L g611 ( .A(n_600), .Y(n_611) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g768 ( .A(n_601), .B(n_618), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
AND2x2_ASAP7_75t_L g694 ( .A(n_603), .B(n_675), .Y(n_694) );
INVx2_ASAP7_75t_L g735 ( .A(n_603), .Y(n_735) );
AND2x4_ASAP7_75t_L g736 ( .A(n_603), .B(n_629), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_604), .B(n_654), .Y(n_784) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_607), .B(n_667), .Y(n_666) );
AND2x4_ASAP7_75t_L g679 ( .A(n_607), .B(n_624), .Y(n_679) );
INVx1_ASAP7_75t_L g771 ( .A(n_607), .Y(n_771) );
AND2x2_ASAP7_75t_L g770 ( .A(n_608), .B(n_697), .Y(n_770) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OAI22xp33_ASAP7_75t_L g741 ( .A1(n_612), .A2(n_742), .B1(n_744), .B2(n_746), .Y(n_741) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AND2x4_ASAP7_75t_L g615 ( .A(n_616), .B(n_619), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x4_ASAP7_75t_L g650 ( .A(n_618), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g686 ( .A(n_618), .Y(n_686) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_618), .Y(n_692) );
INVx2_ASAP7_75t_L g709 ( .A(n_618), .Y(n_709) );
OR2x2_ASAP7_75t_L g730 ( .A(n_618), .B(n_693), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_618), .B(n_688), .Y(n_740) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g707 ( .A(n_620), .B(n_708), .Y(n_707) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_620), .Y(n_761) );
INVx1_ASAP7_75t_L g688 ( .A(n_621), .Y(n_688) );
AOI21xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_626), .B(n_630), .Y(n_622) );
AND2x4_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_625), .B(n_656), .Y(n_655) );
INVx3_ASAP7_75t_L g693 ( .A(n_625), .Y(n_693) );
AND2x2_ASAP7_75t_L g767 ( .A(n_625), .B(n_768), .Y(n_767) );
AOI211x1_ASAP7_75t_SL g695 ( .A1(n_626), .A2(n_696), .B(n_699), .C(n_706), .Y(n_695) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x4_ASAP7_75t_L g752 ( .A(n_628), .B(n_629), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_629), .B(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g745 ( .A(n_629), .Y(n_745) );
AND2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_635), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
INVx1_ASAP7_75t_L g660 ( .A(n_632), .Y(n_660) );
NOR2x1p5_ASAP7_75t_L g717 ( .A(n_632), .B(n_718), .Y(n_717) );
NOR2x1_ASAP7_75t_L g661 ( .A(n_633), .B(n_662), .Y(n_661) );
NOR2xp67_ASAP7_75t_SL g734 ( .A(n_633), .B(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g795 ( .A(n_635), .B(n_703), .Y(n_795) );
NOR2x1_ASAP7_75t_L g636 ( .A(n_637), .B(n_680), .Y(n_636) );
NAND3xp33_ASAP7_75t_SL g637 ( .A(n_638), .B(n_646), .C(n_664), .Y(n_637) );
AND2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_640), .Y(n_671) );
AND2x2_ASAP7_75t_L g678 ( .A(n_640), .B(n_674), .Y(n_678) );
AND2x4_ASAP7_75t_SL g792 ( .A(n_640), .B(n_654), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_641), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_643), .A2(n_685), .B1(n_757), .B2(n_758), .Y(n_756) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AND2x4_ASAP7_75t_L g774 ( .A(n_645), .B(n_775), .Y(n_774) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_649), .B1(n_653), .B2(n_655), .Y(n_647) );
NAND2x1_ASAP7_75t_L g723 ( .A(n_650), .B(n_703), .Y(n_723) );
NAND2xp5_ASAP7_75t_SL g733 ( .A(n_650), .B(n_697), .Y(n_733) );
INVx1_ASAP7_75t_L g760 ( .A(n_650), .Y(n_760) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
OAI21xp5_ASAP7_75t_L g778 ( .A1(n_653), .A2(n_779), .B(n_782), .Y(n_778) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OAI21xp5_ASAP7_75t_L g665 ( .A1(n_654), .A2(n_666), .B(n_669), .Y(n_665) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx2_ASAP7_75t_L g739 ( .A(n_658), .Y(n_739) );
AND2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
INVx1_ASAP7_75t_L g683 ( .A(n_661), .Y(n_683) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AOI222xp33_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_671), .B1(n_672), .B2(n_676), .C1(n_678), .C2(n_679), .Y(n_664) );
AOI21xp33_ASAP7_75t_L g699 ( .A1(n_666), .A2(n_700), .B(n_705), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_667), .B(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g781 ( .A(n_667), .Y(n_781) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
HB1xp67_ASAP7_75t_L g787 ( .A(n_668), .Y(n_787) );
AND2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_675), .Y(n_672) );
AND2x2_ASAP7_75t_L g751 ( .A(n_673), .B(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OR2x2_ASAP7_75t_L g744 ( .A(n_674), .B(n_745), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_695), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_684), .B1(n_690), .B2(n_694), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND2xp33_ASAP7_75t_L g684 ( .A(n_685), .B(n_689), .Y(n_684) );
OR2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
INVx1_ASAP7_75t_L g701 ( .A(n_687), .Y(n_701) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
OR2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx4_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
OR2x2_ASAP7_75t_L g729 ( .A(n_704), .B(n_721), .Y(n_729) );
OR2x2_ASAP7_75t_L g789 ( .A(n_704), .B(n_790), .Y(n_789) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NAND5xp2_ASAP7_75t_L g765 ( .A(n_710), .B(n_757), .C(n_766), .D(n_769), .E(n_771), .Y(n_765) );
NOR2x1_ASAP7_75t_L g712 ( .A(n_713), .B(n_748), .Y(n_712) );
NAND2xp67_ASAP7_75t_SL g713 ( .A(n_714), .B(n_731), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_719), .B1(n_724), .B2(n_725), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
NAND3xp33_ASAP7_75t_SL g719 ( .A(n_720), .B(n_722), .C(n_723), .Y(n_719) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g754 ( .A(n_723), .Y(n_754) );
NAND3xp33_ASAP7_75t_SL g725 ( .A(n_726), .B(n_729), .C(n_730), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g747 ( .A(n_728), .Y(n_747) );
O2A1O1Ixp33_ASAP7_75t_SL g759 ( .A1(n_729), .A2(n_760), .B(n_761), .C(n_762), .Y(n_759) );
AOI221xp5_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_734), .B1(n_736), .B2(n_737), .C(n_741), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_738), .B(n_786), .Y(n_785) );
OR2x2_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
INVx1_ASAP7_75t_L g755 ( .A(n_742), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_749), .B(n_753), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g758 ( .A(n_752), .Y(n_758) );
AOI211xp5_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_755), .B(n_756), .C(n_759), .Y(n_753) );
AOI211x1_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_772), .B(n_778), .C(n_793), .Y(n_764) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
NAND2x1p5_ASAP7_75t_L g773 ( .A(n_774), .B(n_776), .Y(n_773) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
NAND2x1_ASAP7_75t_L g779 ( .A(n_780), .B(n_781), .Y(n_779) );
AOI22xp5_ASAP7_75t_L g782 ( .A1(n_783), .A2(n_785), .B1(n_788), .B2(n_792), .Y(n_782) );
INVxp67_ASAP7_75t_SL g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
AND2x2_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
CKINVDCx6p67_ASAP7_75t_R g806 ( .A(n_798), .Y(n_806) );
BUFx3_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
BUFx6f_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
AND2x6_ASAP7_75t_SL g810 ( .A(n_811), .B(n_813), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx3_ASAP7_75t_L g823 ( .A(n_812), .Y(n_823) );
NOR2xp33_ASAP7_75t_L g847 ( .A(n_812), .B(n_848), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_814), .B(n_816), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
NOR2x1_ASAP7_75t_L g850 ( .A(n_815), .B(n_817), .Y(n_850) );
AND2x6_ASAP7_75t_SL g839 ( .A(n_816), .B(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
OAI21x1_ASAP7_75t_SL g818 ( .A1(n_819), .A2(n_824), .B(n_843), .Y(n_818) );
INVx4_ASAP7_75t_SL g819 ( .A(n_820), .Y(n_819) );
BUFx6f_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
CKINVDCx11_ASAP7_75t_R g821 ( .A(n_822), .Y(n_821) );
BUFx6f_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
AOI22x1_ASAP7_75t_L g824 ( .A1(n_825), .A2(n_834), .B1(n_838), .B2(n_842), .Y(n_824) );
AND2x2_ASAP7_75t_L g825 ( .A(n_826), .B(n_829), .Y(n_825) );
BUFx2_ASAP7_75t_SL g826 ( .A(n_827), .Y(n_826) );
INVx4_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx2_ASAP7_75t_L g853 ( .A(n_828), .Y(n_853) );
INVxp67_ASAP7_75t_SL g842 ( .A(n_829), .Y(n_842) );
XNOR2xp5_ASAP7_75t_L g829 ( .A(n_830), .B(n_833), .Y(n_829) );
NOR2xp33_ASAP7_75t_R g838 ( .A(n_834), .B(n_839), .Y(n_838) );
CKINVDCx5p33_ASAP7_75t_R g837 ( .A(n_835), .Y(n_837) );
INVx3_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx6_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
BUFx10_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
NOR2xp33_ASAP7_75t_SL g851 ( .A(n_852), .B(n_853), .Y(n_851) );
endmodule