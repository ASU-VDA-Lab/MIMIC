module fake_jpeg_29434_n_538 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_538);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_538;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_480;
wire n_267;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_5),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_57),
.Y(n_143)
);

CKINVDCx9p33_ASAP7_75t_R g58 ( 
.A(n_46),
.Y(n_58)
);

INVx5_ASAP7_75t_SL g157 ( 
.A(n_58),
.Y(n_157)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_59),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_60),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_23),
.B(n_8),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_62),
.B(n_80),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_64),
.Y(n_134)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_67),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_68),
.Y(n_130)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_23),
.B(n_7),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_77),
.Y(n_111)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_71),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_73),
.Y(n_167)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_75),
.Y(n_141)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_76),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_26),
.B(n_7),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_78),
.Y(n_165)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_79),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_29),
.B(n_10),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_81),
.Y(n_122)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_82),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_83),
.Y(n_164)
);

AOI21xp33_ASAP7_75t_L g84 ( 
.A1(n_33),
.A2(n_17),
.B(n_6),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_84),
.B(n_12),
.Y(n_137)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_85),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_87),
.Y(n_144)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_88),
.Y(n_154)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_89),
.Y(n_159)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_90),
.Y(n_142)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_91),
.Y(n_152)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_92),
.Y(n_163)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_26),
.B(n_6),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_103),
.Y(n_124)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_95),
.Y(n_153)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_28),
.Y(n_96)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_96),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_38),
.B(n_6),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_102),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_98),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_99),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_100),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_101),
.Y(n_168)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_28),
.Y(n_102)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_31),
.Y(n_103)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_31),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_104),
.B(n_106),
.Y(n_172)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_108),
.Y(n_119)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_40),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_107),
.A2(n_29),
.B1(n_24),
.B2(n_54),
.Y(n_116)
);

BUFx12_ASAP7_75t_L g108 ( 
.A(n_46),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_42),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_43),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_80),
.A2(n_51),
.B1(n_53),
.B2(n_52),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_112),
.A2(n_133),
.B1(n_139),
.B2(n_170),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_116),
.A2(n_41),
.B1(n_27),
.B2(n_21),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_59),
.A2(n_78),
.B1(n_99),
.B2(n_98),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_123),
.A2(n_104),
.B1(n_101),
.B2(n_13),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_128),
.B(n_140),
.Y(n_174)
);

OAI21xp33_ASAP7_75t_L g129 ( 
.A1(n_106),
.A2(n_34),
.B(n_21),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_129),
.B(n_46),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_105),
.A2(n_29),
.B1(n_40),
.B2(n_45),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_137),
.B(n_147),
.Y(n_184)
);

AO22x1_ASAP7_75t_L g138 ( 
.A1(n_108),
.A2(n_46),
.B1(n_34),
.B2(n_35),
.Y(n_138)
);

AO22x1_ASAP7_75t_L g193 ( 
.A1(n_138),
.A2(n_157),
.B1(n_129),
.B2(n_133),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_93),
.A2(n_45),
.B1(n_54),
.B2(n_24),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_64),
.B(n_43),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_63),
.B(n_53),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_149),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_107),
.B(n_52),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_63),
.B(n_51),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_88),
.B(n_38),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_156),
.B(n_158),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_92),
.B(n_20),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_56),
.A2(n_45),
.B1(n_54),
.B2(n_36),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_103),
.B(n_20),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_171),
.Y(n_179)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_173),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_138),
.A2(n_42),
.B1(n_48),
.B2(n_49),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_175),
.Y(n_264)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_172),
.Y(n_178)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_178),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_163),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_180),
.B(n_187),
.Y(n_232)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_150),
.Y(n_181)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_181),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_122),
.Y(n_182)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_182),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_183),
.B(n_193),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_120),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_185),
.Y(n_262)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_186),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_163),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_124),
.B(n_35),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_188),
.B(n_190),
.Y(n_237)
);

BUFx12f_ASAP7_75t_L g189 ( 
.A(n_151),
.Y(n_189)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_189),
.Y(n_265)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_114),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_191),
.A2(n_196),
.B1(n_218),
.B2(n_220),
.Y(n_242)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_121),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_192),
.B(n_201),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_111),
.A2(n_61),
.B1(n_57),
.B2(n_60),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_194),
.A2(n_204),
.B1(n_210),
.B2(n_225),
.Y(n_266)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_120),
.Y(n_195)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_195),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_123),
.A2(n_49),
.B1(n_48),
.B2(n_21),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_115),
.A2(n_81),
.B1(n_66),
.B2(n_86),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_197),
.A2(n_226),
.B1(n_227),
.B2(n_3),
.Y(n_270)
);

INVx13_ASAP7_75t_L g198 ( 
.A(n_157),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g243 ( 
.A(n_198),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_142),
.A2(n_24),
.B1(n_54),
.B2(n_36),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_199),
.A2(n_216),
.B1(n_134),
.B2(n_155),
.Y(n_250)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_117),
.B(n_30),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_202),
.B(n_212),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_126),
.B(n_27),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_203),
.B(n_213),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_170),
.A2(n_73),
.B1(n_72),
.B2(n_83),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_166),
.Y(n_205)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_205),
.Y(n_257)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_132),
.Y(n_206)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_206),
.Y(n_261)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_135),
.Y(n_207)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_207),
.Y(n_238)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_168),
.Y(n_208)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_160),
.Y(n_209)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_209),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_139),
.A2(n_116),
.B1(n_100),
.B2(n_148),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_160),
.Y(n_211)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_211),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_119),
.B(n_30),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_118),
.B(n_41),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_110),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_214),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_159),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_215),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_144),
.A2(n_36),
.B1(n_54),
.B2(n_24),
.Y(n_216)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_113),
.Y(n_217)
);

INVx5_ASAP7_75t_L g247 ( 
.A(n_217),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_118),
.A2(n_41),
.B1(n_27),
.B2(n_36),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_131),
.B(n_36),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_219),
.B(n_221),
.C(n_4),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_153),
.A2(n_12),
.B1(n_16),
.B2(n_15),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_110),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_224),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_130),
.Y(n_223)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_223),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_145),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_148),
.A2(n_154),
.B1(n_164),
.B2(n_131),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_136),
.A2(n_12),
.B1(n_16),
.B2(n_15),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_136),
.A2(n_5),
.B1(n_16),
.B2(n_14),
.Y(n_227)
);

BUFx4f_ASAP7_75t_SL g228 ( 
.A(n_151),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_130),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_193),
.A2(n_165),
.B1(n_154),
.B2(n_167),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_230),
.A2(n_245),
.B1(n_225),
.B2(n_224),
.Y(n_272)
);

AND2x6_ASAP7_75t_L g233 ( 
.A(n_193),
.B(n_169),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_233),
.A2(n_248),
.B(n_254),
.Y(n_283)
);

OAI221xp5_ASAP7_75t_L g240 ( 
.A1(n_184),
.A2(n_127),
.B1(n_153),
.B2(n_159),
.C(n_155),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_240),
.B(n_189),
.Y(n_299)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_178),
.A2(n_165),
.B1(n_167),
.B2(n_122),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_246),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_183),
.A2(n_13),
.B(n_17),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_250),
.Y(n_295)
);

AO22x1_ASAP7_75t_SL g251 ( 
.A1(n_183),
.A2(n_125),
.B1(n_143),
.B2(n_161),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_220),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_177),
.A2(n_179),
.B1(n_210),
.B2(n_134),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_252),
.A2(n_253),
.B1(n_182),
.B2(n_189),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_179),
.A2(n_125),
.B1(n_161),
.B2(n_143),
.Y(n_253)
);

AND2x6_ASAP7_75t_L g255 ( 
.A(n_188),
.B(n_4),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_255),
.A2(n_3),
.B(n_4),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_204),
.A2(n_4),
.B1(n_13),
.B2(n_5),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_260),
.A2(n_228),
.B(n_215),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_270),
.A2(n_196),
.B1(n_221),
.B2(n_213),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_272),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_274),
.A2(n_277),
.B1(n_279),
.B2(n_286),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_275),
.A2(n_293),
.B1(n_280),
.B2(n_299),
.Y(n_311)
);

AOI32xp33_ASAP7_75t_L g276 ( 
.A1(n_233),
.A2(n_200),
.A3(n_176),
.B1(n_174),
.B2(n_180),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_276),
.B(n_299),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_242),
.A2(n_203),
.B1(n_192),
.B2(n_190),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_236),
.B(n_203),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_278),
.B(n_282),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_242),
.A2(n_191),
.B1(n_187),
.B2(n_207),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_232),
.Y(n_280)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_280),
.Y(n_312)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_261),
.Y(n_281)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_281),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_244),
.B(n_212),
.Y(n_282)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_229),
.Y(n_284)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_284),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_264),
.A2(n_206),
.B1(n_215),
.B2(n_186),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_285),
.A2(n_247),
.B(n_263),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_264),
.A2(n_201),
.B1(n_181),
.B2(n_173),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_236),
.B(n_202),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_287),
.B(n_300),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_288),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_268),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_289),
.B(n_291),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_256),
.B(n_219),
.C(n_222),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_290),
.B(n_294),
.C(n_304),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_241),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_268),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_292),
.B(n_302),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_266),
.A2(n_205),
.B1(n_195),
.B2(n_185),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_208),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_266),
.A2(n_211),
.B1(n_209),
.B2(n_214),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_296),
.A2(n_306),
.B1(n_243),
.B2(n_262),
.Y(n_334)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_261),
.Y(n_297)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_297),
.Y(n_321)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_238),
.Y(n_298)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_298),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_237),
.B(n_198),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_256),
.A2(n_217),
.B(n_228),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_301),
.A2(n_243),
.B(n_189),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_259),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_262),
.Y(n_303)
);

INVx3_ASAP7_75t_SL g338 ( 
.A(n_303),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_254),
.B(n_223),
.C(n_185),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_251),
.B(n_182),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_305),
.B(n_307),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_269),
.C(n_258),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_309),
.B(n_324),
.C(n_283),
.Y(n_362)
);

BUFx5_ASAP7_75t_L g310 ( 
.A(n_303),
.Y(n_310)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_310),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_311),
.B(n_317),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_287),
.B(n_248),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_314),
.B(n_319),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_315),
.A2(n_318),
.B(n_301),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_275),
.A2(n_251),
.B1(n_270),
.B2(n_255),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_288),
.A2(n_260),
.B(n_263),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_278),
.B(n_239),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_290),
.B(n_239),
.Y(n_324)
);

OAI32xp33_ASAP7_75t_L g327 ( 
.A1(n_305),
.A2(n_229),
.A3(n_257),
.B1(n_243),
.B2(n_249),
.Y(n_327)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_327),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_329),
.A2(n_285),
.B(n_286),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_302),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_330),
.B(n_337),
.Y(n_349)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_281),
.Y(n_333)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_333),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_334),
.A2(n_293),
.B1(n_279),
.B2(n_288),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_294),
.B(n_231),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_336),
.B(n_304),
.C(n_283),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_300),
.Y(n_337)
);

AO22x1_ASAP7_75t_SL g340 ( 
.A1(n_274),
.A2(n_257),
.B1(n_231),
.B2(n_234),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_340),
.B(n_296),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_342),
.B(n_298),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_343),
.A2(n_346),
.B(n_351),
.Y(n_393)
);

AOI32xp33_ASAP7_75t_L g344 ( 
.A1(n_335),
.A2(n_323),
.A3(n_329),
.B1(n_339),
.B2(n_295),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_344),
.B(n_359),
.Y(n_390)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_331),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_345),
.B(n_347),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_323),
.A2(n_301),
.B(n_306),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_308),
.B(n_294),
.C(n_304),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_348),
.B(n_324),
.C(n_336),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_312),
.B(n_282),
.Y(n_350)
);

CKINVDCx14_ASAP7_75t_R g398 ( 
.A(n_350),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_312),
.B(n_277),
.Y(n_352)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_352),
.Y(n_374)
);

A2O1A1Ixp33_ASAP7_75t_SL g386 ( 
.A1(n_353),
.A2(n_327),
.B(n_340),
.C(n_317),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_326),
.B(n_291),
.Y(n_355)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_355),
.B(n_357),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_313),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_356),
.B(n_363),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_313),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_321),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_311),
.B(n_273),
.Y(n_360)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_360),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_362),
.B(n_372),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_316),
.B(n_307),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_320),
.Y(n_364)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_364),
.Y(n_400)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_321),
.Y(n_365)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_365),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_333),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_366),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_325),
.B(n_276),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_367),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_318),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_368),
.B(n_340),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_316),
.B(n_285),
.Y(n_369)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_369),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_325),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_370),
.Y(n_396)
);

XNOR2x1_ASAP7_75t_L g372 ( 
.A(n_308),
.B(n_272),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_354),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_375),
.B(n_389),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_358),
.A2(n_322),
.B1(n_328),
.B2(n_334),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_377),
.A2(n_383),
.B1(n_353),
.B2(n_341),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_358),
.A2(n_322),
.B1(n_328),
.B2(n_315),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_384),
.B(n_404),
.C(n_348),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_386),
.A2(n_399),
.B(n_346),
.Y(n_416)
);

CKINVDCx14_ASAP7_75t_R g432 ( 
.A(n_387),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_364),
.Y(n_388)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_388),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_349),
.Y(n_389)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_349),
.Y(n_392)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_392),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_350),
.B(n_309),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_394),
.B(n_362),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_355),
.B(n_332),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_395),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_371),
.B(n_314),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_397),
.B(n_371),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_360),
.A2(n_332),
.B(n_292),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_345),
.B(n_319),
.Y(n_401)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_401),
.Y(n_425)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_361),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_402),
.B(n_403),
.Y(n_405)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_364),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_379),
.A2(n_367),
.B1(n_363),
.B2(n_351),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_406),
.A2(n_414),
.B1(n_424),
.B2(n_428),
.Y(n_440)
);

OAI32xp33_ASAP7_75t_L g407 ( 
.A1(n_379),
.A2(n_341),
.A3(n_369),
.B1(n_352),
.B2(n_347),
.Y(n_407)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_407),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_408),
.B(n_417),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_409),
.A2(n_386),
.B1(n_374),
.B2(n_381),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_411),
.B(n_415),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_392),
.B(n_357),
.Y(n_412)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_412),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_384),
.B(n_342),
.C(n_362),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_413),
.B(n_418),
.C(n_378),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_385),
.A2(n_372),
.B1(n_344),
.B2(n_343),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_416),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_382),
.B(n_366),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_404),
.B(n_372),
.C(n_356),
.Y(n_418)
);

OR2x2_ASAP7_75t_L g420 ( 
.A(n_391),
.B(n_370),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_420),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_382),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_421),
.B(n_430),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_391),
.B(n_356),
.Y(n_423)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_423),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_385),
.A2(n_365),
.B1(n_361),
.B2(n_359),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_398),
.B(n_297),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_426),
.B(n_429),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_374),
.A2(n_354),
.B1(n_338),
.B2(n_310),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_396),
.B(n_289),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_373),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_373),
.B(n_320),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_431),
.B(n_433),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_387),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_436),
.B(n_438),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_411),
.B(n_376),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_439),
.A2(n_448),
.B1(n_420),
.B2(n_430),
.Y(n_460)
);

A2O1A1Ixp33_ASAP7_75t_SL g442 ( 
.A1(n_416),
.A2(n_386),
.B(n_393),
.C(n_399),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_442),
.A2(n_433),
.B1(n_422),
.B2(n_407),
.Y(n_463)
);

XNOR2x1_ASAP7_75t_SL g445 ( 
.A(n_414),
.B(n_390),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_445),
.B(n_417),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_409),
.A2(n_393),
.B1(n_386),
.B2(n_377),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_422),
.Y(n_450)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_450),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_413),
.B(n_378),
.C(n_376),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_451),
.B(n_454),
.C(n_446),
.Y(n_458)
);

BUFx4f_ASAP7_75t_SL g452 ( 
.A(n_419),
.Y(n_452)
);

CKINVDCx14_ASAP7_75t_R g475 ( 
.A(n_452),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_406),
.A2(n_421),
.B1(n_410),
.B2(n_432),
.Y(n_453)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_453),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_418),
.B(n_397),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_410),
.A2(n_383),
.B1(n_401),
.B2(n_386),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_455),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_457),
.B(n_458),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_460),
.B(n_470),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_438),
.B(n_408),
.C(n_415),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_462),
.B(n_471),
.C(n_474),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_463),
.A2(n_472),
.B1(n_405),
.B2(n_403),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_434),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_464),
.B(n_465),
.Y(n_487)
);

BUFx24_ASAP7_75t_SL g465 ( 
.A(n_437),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_444),
.A2(n_427),
.B(n_429),
.Y(n_467)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_467),
.Y(n_484)
);

OAI21x1_ASAP7_75t_L g469 ( 
.A1(n_447),
.A2(n_412),
.B(n_427),
.Y(n_469)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_469),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_454),
.B(n_425),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_451),
.B(n_425),
.C(n_424),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_440),
.A2(n_426),
.B1(n_402),
.B2(n_380),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_436),
.B(n_446),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_473),
.B(n_456),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_440),
.B(n_423),
.C(n_431),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_459),
.A2(n_435),
.B1(n_449),
.B2(n_443),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_476),
.B(n_481),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_457),
.B(n_439),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_480),
.B(n_483),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_459),
.A2(n_456),
.B1(n_441),
.B2(n_445),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_482),
.B(n_486),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_463),
.Y(n_483)
);

CKINVDCx16_ASAP7_75t_R g485 ( 
.A(n_466),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_485),
.B(n_489),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_468),
.A2(n_475),
.B1(n_442),
.B2(n_474),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_472),
.A2(n_448),
.B1(n_420),
.B2(n_428),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_461),
.B(n_405),
.C(n_442),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_490),
.B(n_462),
.C(n_473),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_461),
.A2(n_442),
.B1(n_380),
.B2(n_471),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_491),
.B(n_492),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_493),
.B(n_502),
.Y(n_511)
);

XNOR2x1_ASAP7_75t_L g494 ( 
.A(n_479),
.B(n_470),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_494),
.B(n_481),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_488),
.A2(n_452),
.B1(n_419),
.B2(n_458),
.Y(n_495)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_495),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_477),
.A2(n_490),
.B(n_491),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_498),
.B(n_506),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_477),
.B(n_452),
.C(n_400),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_499),
.B(n_482),
.C(n_492),
.Y(n_510)
);

OR2x2_ASAP7_75t_L g502 ( 
.A(n_476),
.B(n_388),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_SL g503 ( 
.A(n_479),
.B(n_400),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_503),
.B(n_505),
.Y(n_512)
);

AOI21x1_ASAP7_75t_L g505 ( 
.A1(n_484),
.A2(n_338),
.B(n_303),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_478),
.B(n_284),
.C(n_265),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_478),
.B(n_265),
.C(n_249),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_507),
.B(n_499),
.Y(n_516)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_510),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_513),
.B(n_500),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_493),
.B(n_486),
.C(n_487),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_514),
.B(n_515),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_501),
.B(n_338),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_516),
.B(n_518),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_SL g517 ( 
.A(n_494),
.B(n_247),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_517),
.B(n_503),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_504),
.A2(n_234),
.B1(n_267),
.B2(n_235),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_510),
.B(n_497),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_519),
.B(n_520),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_509),
.A2(n_502),
.B1(n_496),
.B2(n_500),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_524),
.B(n_525),
.C(n_497),
.Y(n_528)
);

NOR3xp33_ASAP7_75t_SL g526 ( 
.A(n_522),
.B(n_511),
.C(n_508),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_526),
.A2(n_528),
.B(n_525),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_SL g529 ( 
.A1(n_521),
.A2(n_514),
.B(n_513),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_529),
.A2(n_523),
.B(n_519),
.Y(n_530)
);

OAI311xp33_ASAP7_75t_L g533 ( 
.A1(n_530),
.A2(n_531),
.A3(n_532),
.B1(n_512),
.C1(n_267),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_SL g532 ( 
.A1(n_527),
.A2(n_496),
.B(n_517),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_533),
.B(n_512),
.C(n_235),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_534),
.A2(n_17),
.B(n_1),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_535),
.A2(n_17),
.B(n_1),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_536),
.B(n_2),
.C(n_0),
.Y(n_537)
);

O2A1O1Ixp33_ASAP7_75t_SL g538 ( 
.A1(n_537),
.A2(n_1),
.B(n_2),
.C(n_522),
.Y(n_538)
);


endmodule