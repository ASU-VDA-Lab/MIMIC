module fake_jpeg_13341_n_181 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_181);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_181;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_24),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_43),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_27),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_49),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_13),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_33),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_7),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_4),
.Y(n_74)
);

INVx11_ASAP7_75t_SL g75 ( 
.A(n_6),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_48),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_12),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_73),
.B(n_0),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_86),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

BUFx8_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_68),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_79),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

BUFx12_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_1),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_2),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_88),
.B(n_78),
.Y(n_105)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_89),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_18),
.C(n_44),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_90),
.A2(n_52),
.B(n_77),
.Y(n_93)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_91),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_99),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_55),
.B1(n_74),
.B2(n_64),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_94),
.A2(n_97),
.B1(n_71),
.B2(n_65),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_66),
.B(n_59),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_104),
.B(n_91),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_55),
.B1(n_74),
.B2(n_67),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_84),
.B(n_90),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_105),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_82),
.A2(n_67),
.B1(n_62),
.B2(n_64),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_76),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_58),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_104),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_119),
.B1(n_3),
.B2(n_5),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_108),
.Y(n_111)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_100),
.B(n_84),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_112),
.B(n_117),
.Y(n_132)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_96),
.B(n_56),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_89),
.B(n_72),
.C(n_68),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_129),
.B(n_21),
.Y(n_140)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_126),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_123),
.Y(n_148)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_128),
.Y(n_144)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_92),
.B(n_60),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_127),
.B(n_130),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_63),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_101),
.A2(n_72),
.B1(n_68),
.B2(n_5),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_129),
.A2(n_120),
.B1(n_123),
.B2(n_122),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_100),
.B(n_2),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_3),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_131),
.B(n_6),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_116),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_149),
.Y(n_161)
);

MAJx2_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_72),
.C(n_20),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_139),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_17),
.C(n_42),
.Y(n_139)
);

NAND3xp33_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_29),
.C(n_32),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_142),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_146),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_25),
.C(n_41),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_127),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_127),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_11),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_151),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_162),
.Y(n_170)
);

AOI22x1_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_15),
.B1(n_39),
.B2(n_38),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_SL g171 ( 
.A1(n_156),
.A2(n_158),
.B(n_143),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_7),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_157),
.B(n_160),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_8),
.Y(n_160)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_163),
.B(n_164),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_9),
.B(n_10),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_144),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_169),
.C(n_154),
.Y(n_172)
);

XNOR2x1_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_138),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_SL g174 ( 
.A1(n_171),
.A2(n_158),
.B(n_140),
.C(n_156),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_173),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_159),
.C(n_153),
.Y(n_173)
);

INVxp33_ASAP7_75t_L g175 ( 
.A(n_174),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_135),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_141),
.Y(n_178)
);

AOI322xp5_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_167),
.A3(n_166),
.B1(n_159),
.B2(n_152),
.C1(n_175),
.C2(n_134),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_11),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_139),
.Y(n_181)
);


endmodule