module fake_jpeg_10855_n_356 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_356);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_356;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVxp67_ASAP7_75t_SL g88 ( 
.A(n_47),
.Y(n_88)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_16),
.C(n_15),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_33),
.Y(n_79)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

AOI21xp33_ASAP7_75t_L g55 ( 
.A1(n_32),
.A2(n_16),
.B(n_14),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_55),
.B(n_33),
.Y(n_95)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

BUFx4f_ASAP7_75t_SL g102 ( 
.A(n_58),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_23),
.A2(n_26),
.B1(n_35),
.B2(n_19),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_64),
.A2(n_23),
.B1(n_38),
.B2(n_37),
.Y(n_94)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_23),
.A2(n_19),
.B1(n_26),
.B2(n_35),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_66),
.A2(n_18),
.B1(n_40),
.B2(n_24),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_70),
.B(n_23),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_72),
.B(n_80),
.Y(n_131)
);

AOI21xp33_ASAP7_75t_L g73 ( 
.A1(n_51),
.A2(n_32),
.B(n_39),
.Y(n_73)
);

NAND3xp33_ASAP7_75t_L g144 ( 
.A(n_73),
.B(n_79),
.C(n_108),
.Y(n_144)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_47),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_75),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_39),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_81),
.B(n_84),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_28),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_82),
.B(n_107),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_28),
.Y(n_84)
);

INVx6_ASAP7_75t_SL g87 ( 
.A(n_46),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_87),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_64),
.A2(n_59),
.B1(n_68),
.B2(n_43),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_93),
.A2(n_44),
.B1(n_71),
.B2(n_69),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_94),
.A2(n_38),
.B1(n_50),
.B2(n_49),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_95),
.B(n_98),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_40),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_64),
.A2(n_19),
.B1(n_23),
.B2(n_37),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_99),
.A2(n_117),
.B1(n_38),
.B2(n_29),
.Y(n_125)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

INVx11_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_53),
.B(n_41),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_109),
.A2(n_21),
.B1(n_17),
.B2(n_31),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_67),
.B(n_18),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_111),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_65),
.B(n_20),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_3),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_45),
.A2(n_38),
.B1(n_41),
.B2(n_34),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_118),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_119),
.A2(n_125),
.B1(n_134),
.B2(n_149),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_80),
.A2(n_54),
.B(n_20),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_120),
.A2(n_78),
.B(n_9),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_121),
.A2(n_122),
.B1(n_124),
.B2(n_130),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_82),
.A2(n_31),
.B1(n_24),
.B2(n_34),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_123),
.A2(n_155),
.B1(n_9),
.B2(n_78),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_21),
.B1(n_17),
.B2(n_38),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_112),
.A2(n_29),
.B1(n_1),
.B2(n_2),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_129),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_105),
.A2(n_29),
.B1(n_16),
.B2(n_14),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_105),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_132),
.A2(n_152),
.B1(n_115),
.B2(n_77),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_88),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_90),
.Y(n_136)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_137),
.Y(n_176)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_138),
.Y(n_189)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_142),
.B(n_9),
.Y(n_186)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_143),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_97),
.B(n_113),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_154),
.Y(n_174)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_96),
.Y(n_147)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_103),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_149)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_77),
.Y(n_150)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_76),
.Y(n_151)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_100),
.A2(n_13),
.B1(n_11),
.B2(n_10),
.Y(n_152)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_104),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_102),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_92),
.B(n_4),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_100),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_103),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_156),
.A2(n_114),
.B1(n_115),
.B2(n_83),
.Y(n_177)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_76),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_96),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_159),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_116),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_161),
.B(n_164),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_144),
.C(n_146),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_163),
.B(n_183),
.C(n_124),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_86),
.Y(n_164)
);

O2A1O1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_131),
.A2(n_75),
.B(n_72),
.C(n_102),
.Y(n_166)
);

OA21x2_ASAP7_75t_L g226 ( 
.A1(n_166),
.A2(n_159),
.B(n_172),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_86),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_168),
.B(n_173),
.Y(n_201)
);

FAx1_ASAP7_75t_SL g171 ( 
.A(n_142),
.B(n_101),
.CI(n_106),
.CON(n_171),
.SN(n_171)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_178),
.Y(n_199)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_172),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_74),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_74),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_175),
.B(n_180),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_177),
.A2(n_185),
.B(n_157),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_141),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_102),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_184),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_121),
.A2(n_91),
.B1(n_85),
.B2(n_83),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_182),
.A2(n_192),
.B1(n_155),
.B2(n_150),
.Y(n_210)
);

AND2x2_ASAP7_75t_SL g183 ( 
.A(n_154),
.B(n_114),
.Y(n_183)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_145),
.A2(n_10),
.B(n_13),
.C(n_8),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_186),
.B(n_163),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_122),
.B(n_85),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_152),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_120),
.A2(n_131),
.B(n_127),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_190),
.A2(n_127),
.B(n_128),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_119),
.A2(n_91),
.B1(n_78),
.B2(n_9),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_193),
.A2(n_143),
.B1(n_153),
.B2(n_147),
.Y(n_218)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_169),
.Y(n_195)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_195),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_197),
.A2(n_207),
.B(n_226),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_198),
.B(n_224),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_208),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_166),
.A2(n_128),
.B1(n_140),
.B2(n_137),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_203),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_206),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_190),
.A2(n_118),
.B(n_130),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_205),
.A2(n_216),
.B(n_217),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_123),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_R g207 ( 
.A(n_168),
.B(n_141),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_132),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_136),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_219),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_210),
.A2(n_211),
.B1(n_193),
.B2(n_169),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_179),
.A2(n_150),
.B1(n_138),
.B2(n_135),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_164),
.B(n_126),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_212),
.B(n_214),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_173),
.B(n_126),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_175),
.B(n_151),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_222),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_185),
.A2(n_166),
.B(n_180),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_218),
.A2(n_178),
.B1(n_177),
.B2(n_176),
.Y(n_245)
);

NAND2x1p5_ASAP7_75t_L g219 ( 
.A(n_171),
.B(n_183),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_183),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_223),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_167),
.B(n_165),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_171),
.B(n_187),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_179),
.B(n_158),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_165),
.B(n_189),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_176),
.Y(n_234)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_225),
.Y(n_228)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_228),
.Y(n_260)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_195),
.Y(n_230)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_230),
.Y(n_264)
);

OA21x2_ASAP7_75t_L g232 ( 
.A1(n_199),
.A2(n_158),
.B(n_192),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_234),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_202),
.A2(n_223),
.B1(n_196),
.B2(n_208),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_235),
.A2(n_245),
.B1(n_252),
.B2(n_255),
.Y(n_257)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_211),
.Y(n_236)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_236),
.Y(n_266)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_237),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_167),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_240),
.Y(n_263)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_200),
.Y(n_242)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_242),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_210),
.A2(n_194),
.B1(n_181),
.B2(n_182),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_243),
.A2(n_253),
.B1(n_218),
.B2(n_220),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_213),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_247),
.Y(n_262)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_226),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_200),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_196),
.A2(n_194),
.B1(n_184),
.B2(n_189),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_205),
.A2(n_170),
.B1(n_162),
.B2(n_188),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_224),
.A2(n_170),
.B1(n_162),
.B2(n_188),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_197),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_258),
.A2(n_251),
.B(n_226),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_238),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_265),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_221),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_270),
.C(n_274),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_228),
.B(n_209),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_233),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_272),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_269),
.A2(n_255),
.B1(n_232),
.B2(n_226),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_239),
.B(n_198),
.C(n_204),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_234),
.B(n_201),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_201),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_229),
.B(n_242),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_277),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_219),
.C(n_227),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_227),
.C(n_235),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_229),
.B(n_206),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_246),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_274),
.Y(n_297)
);

XOR2x2_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_246),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_279),
.B(n_257),
.Y(n_307)
);

MAJx2_ASAP7_75t_L g306 ( 
.A(n_282),
.B(n_277),
.C(n_265),
.Y(n_306)
);

INVxp67_ASAP7_75t_SL g284 ( 
.A(n_262),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_284),
.B(n_288),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_231),
.C(n_250),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_296),
.C(n_281),
.Y(n_300)
);

AND2x6_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_248),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_286),
.A2(n_293),
.B1(n_257),
.B2(n_271),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_287),
.A2(n_292),
.B(n_294),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_275),
.Y(n_288)
);

NAND3xp33_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_231),
.C(n_250),
.Y(n_289)
);

NOR3xp33_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_291),
.C(n_260),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_271),
.A2(n_237),
.B1(n_236),
.B2(n_251),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_269),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_268),
.B(n_252),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_258),
.A2(n_248),
.B(n_219),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_258),
.A2(n_207),
.B(n_232),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_261),
.B(n_253),
.C(n_217),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_297),
.B(n_301),
.C(n_302),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_300),
.B(n_306),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_278),
.B(n_256),
.C(n_276),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_256),
.C(n_272),
.Y(n_302)
);

INVx11_ASAP7_75t_L g303 ( 
.A(n_294),
.Y(n_303)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_303),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_305),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_308),
.C(n_310),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_285),
.B(n_260),
.C(n_267),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_311),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_258),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_283),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_293),
.A2(n_266),
.B1(n_243),
.B2(n_259),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_290),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_303),
.A2(n_286),
.B(n_287),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_314),
.A2(n_321),
.B(n_298),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_322),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_298),
.A2(n_292),
.B(n_283),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_302),
.B(n_282),
.C(n_279),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_305),
.A2(n_295),
.B1(n_280),
.B2(n_266),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_323),
.A2(n_324),
.B1(n_273),
.B2(n_308),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_312),
.A2(n_295),
.B1(n_273),
.B2(n_216),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_325),
.B(n_332),
.Y(n_336)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_326),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_300),
.C(n_301),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_327),
.B(n_329),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_310),
.Y(n_328)
);

XNOR2x1_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_315),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_317),
.A2(n_299),
.B1(n_264),
.B2(n_307),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_313),
.A2(n_264),
.B1(n_241),
.B2(n_220),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_331),
.B(n_324),
.C(n_321),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_314),
.A2(n_297),
.B(n_306),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_323),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_334),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_315),
.B(n_241),
.C(n_191),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_335),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_330),
.B(n_327),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_340),
.B(n_328),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_334),
.B(n_319),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_341),
.A2(n_319),
.B(n_320),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_342),
.B(n_326),
.Y(n_346)
);

OAI21x1_ASAP7_75t_L g348 ( 
.A1(n_343),
.A2(n_344),
.B(n_347),
.Y(n_348)
);

NOR3xp33_ASAP7_75t_SL g344 ( 
.A(n_336),
.B(n_332),
.C(n_325),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_346),
.B(n_337),
.Y(n_349)
);

AO21x1_ASAP7_75t_L g351 ( 
.A1(n_349),
.A2(n_350),
.B(n_341),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_345),
.Y(n_350)
);

AOI321xp33_ASAP7_75t_L g353 ( 
.A1(n_351),
.A2(n_352),
.A3(n_339),
.B1(n_318),
.B2(n_322),
.C(n_191),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_348),
.A2(n_336),
.B(n_338),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_353),
.B(n_318),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_354),
.B(n_188),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_355),
.A2(n_160),
.B1(n_172),
.B2(n_263),
.Y(n_356)
);


endmodule