module real_jpeg_9111_n_7 (n_5, n_4, n_0, n_1, n_2, n_6, n_3, n_7);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_3;

output n_7;

wire n_17;
wire n_8;
wire n_43;
wire n_57;
wire n_37;
wire n_21;
wire n_54;
wire n_65;
wire n_33;
wire n_38;
wire n_35;
wire n_50;
wire n_29;
wire n_55;
wire n_69;
wire n_49;
wire n_52;
wire n_10;
wire n_9;
wire n_31;
wire n_67;
wire n_58;
wire n_63;
wire n_12;
wire n_68;
wire n_24;
wire n_66;
wire n_34;
wire n_28;
wire n_60;
wire n_44;
wire n_46;
wire n_62;
wire n_59;
wire n_64;
wire n_23;
wire n_11;
wire n_14;
wire n_47;
wire n_51;
wire n_45;
wire n_25;
wire n_61;
wire n_42;
wire n_53;
wire n_18;
wire n_22;
wire n_39;
wire n_40;
wire n_36;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_48;
wire n_30;
wire n_56;
wire n_16;
wire n_15;
wire n_13;

AOI22xp33_ASAP7_75t_SL g12 ( 
.A1(n_0),
.A2(n_13),
.B1(n_14),
.B2(n_17),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_0),
.A2(n_17),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_3),
.A2(n_13),
.B1(n_14),
.B2(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g37 ( 
.A1(n_3),
.A2(n_28),
.B(n_33),
.C(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_3),
.B(n_28),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_3),
.A2(n_6),
.B(n_14),
.Y(n_41)
);

BUFx6f_ASAP7_75t_SL g62 ( 
.A(n_4),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_6),
.A2(n_13),
.B1(n_14),
.B2(n_23),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_6),
.A2(n_23),
.B1(n_28),
.B2(n_29),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_6),
.B(n_60),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_53),
.Y(n_7)
);

AOI21xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_43),
.B(n_52),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_24),
.Y(n_9)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_10),
.B(n_24),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g10 ( 
.A1(n_11),
.A2(n_18),
.B(n_19),
.Y(n_10)
);

CKINVDCx16_ASAP7_75t_R g11 ( 
.A(n_12),
.Y(n_11)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_12),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_13),
.B(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_14),
.B(n_21),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

BUFx24_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_18),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_22),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_21),
.B(n_23),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_23),
.A2(n_29),
.B(n_34),
.C(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_23),
.B(n_33),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_25),
.B(n_40),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B(n_35),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_27),
.A2(n_33),
.B1(n_36),
.B2(n_37),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_28),
.A2(n_29),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_48),
.B(n_51),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_49),
.B(n_50),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_50),
.A2(n_56),
.B1(n_57),
.B2(n_66),
.Y(n_55)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_68),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_67),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_67),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_64),
.B2(n_65),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_62),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);


endmodule