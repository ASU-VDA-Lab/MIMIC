module fake_jpeg_18444_n_203 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_203);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_17),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_30),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_27),
.Y(n_54)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_46),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_16),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_32),
.A2(n_16),
.B1(n_17),
.B2(n_27),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_48),
.A2(n_19),
.B1(n_22),
.B2(n_18),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_15),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_40),
.C(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_54),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_57),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_54),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_41),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_65),
.Y(n_83)
);

FAx1_ASAP7_75t_SL g90 ( 
.A(n_60),
.B(n_66),
.CI(n_67),
.CON(n_90),
.SN(n_90)
);

AO22x1_ASAP7_75t_SL g61 ( 
.A1(n_46),
.A2(n_39),
.B1(n_34),
.B2(n_37),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_61),
.A2(n_64),
.B1(n_69),
.B2(n_76),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_62),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_23),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_68),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_36),
.Y(n_65)
);

AND2x4_ASAP7_75t_SL g66 ( 
.A(n_51),
.B(n_39),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_47),
.A2(n_29),
.B1(n_26),
.B2(n_24),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_74),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_42),
.B(n_23),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_72),
.B(n_73),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_52),
.A2(n_21),
.B(n_24),
.C(n_26),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_43),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_47),
.A2(n_29),
.B1(n_21),
.B2(n_22),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_52),
.A2(n_39),
.B(n_19),
.C(n_18),
.Y(n_78)
);

OAI32xp33_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_25),
.A3(n_20),
.B1(n_31),
.B2(n_15),
.Y(n_95)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_42),
.B(n_33),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_31),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_47),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_81),
.A2(n_61),
.B(n_78),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_14),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_86),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_50),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_95),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_75),
.A2(n_50),
.B1(n_52),
.B2(n_33),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_88),
.A2(n_91),
.B1(n_94),
.B2(n_102),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_64),
.A2(n_50),
.B1(n_40),
.B2(n_43),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_65),
.A2(n_43),
.B1(n_38),
.B2(n_36),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_71),
.Y(n_105)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_66),
.A2(n_25),
.B1(n_2),
.B2(n_3),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_76),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_103),
.B(n_1),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_60),
.C(n_66),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_84),
.C(n_85),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_107),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_82),
.A2(n_55),
.B(n_67),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_106),
.A2(n_110),
.B(n_122),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_69),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_103),
.A2(n_67),
.B1(n_95),
.B2(n_92),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_82),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_112),
.B(n_117),
.Y(n_141)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_115),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_61),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_125),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_73),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_119),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_77),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_93),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_99),
.Y(n_126)
);

OAI22x1_ASAP7_75t_SL g121 ( 
.A1(n_92),
.A2(n_79),
.B1(n_2),
.B2(n_3),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_121),
.A2(n_81),
.B1(n_98),
.B2(n_83),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_14),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_1),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_126),
.B(n_127),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_99),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_81),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_129),
.A2(n_118),
.B(n_113),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_133),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_90),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_100),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_134),
.B(n_144),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_94),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_135),
.B(n_138),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_102),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_108),
.A2(n_91),
.B1(n_85),
.B2(n_101),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_5),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_143),
.B(n_120),
.C(n_124),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_122),
.Y(n_144)
);

OA22x2_ASAP7_75t_L g146 ( 
.A1(n_137),
.A2(n_121),
.B1(n_117),
.B2(n_109),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_147),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_136),
.A2(n_110),
.B(n_108),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_150),
.Y(n_161)
);

AOI322xp5_ASAP7_75t_L g151 ( 
.A1(n_136),
.A2(n_124),
.A3(n_113),
.B1(n_84),
.B2(n_11),
.C1(n_12),
.C2(n_13),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_151),
.B(n_156),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_11),
.Y(n_153)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_157),
.A2(n_130),
.B1(n_145),
.B2(n_138),
.Y(n_166)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_158),
.A2(n_150),
.B1(n_156),
.B2(n_146),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_128),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_135),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_160),
.A2(n_140),
.B1(n_133),
.B2(n_143),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_162),
.A2(n_154),
.B1(n_129),
.B2(n_159),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_167),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_146),
.Y(n_167)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_169),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_157),
.A2(n_129),
.B1(n_131),
.B2(n_142),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_170),
.A2(n_171),
.B1(n_158),
.B2(n_149),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_163),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_176),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_178),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_148),
.C(n_159),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_170),
.B(n_147),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_179),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_167),
.A2(n_154),
.B1(n_146),
.B2(n_149),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_180),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_177),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_184),
.C(n_5),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_179),
.B(n_161),
.C(n_168),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_L g187 ( 
.A1(n_172),
.A2(n_164),
.B1(n_162),
.B2(n_155),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_187),
.A2(n_131),
.B(n_142),
.Y(n_190)
);

OAI21x1_ASAP7_75t_L g188 ( 
.A1(n_182),
.A2(n_174),
.B(n_155),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_188),
.B(n_190),
.Y(n_193)
);

OAI221xp5_ASAP7_75t_L g189 ( 
.A1(n_185),
.A2(n_175),
.B1(n_164),
.B2(n_178),
.C(n_145),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_189),
.B(n_191),
.Y(n_195)
);

FAx1_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_165),
.CI(n_6),
.CON(n_191),
.SN(n_191)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_192),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_188),
.A2(n_181),
.B(n_186),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_5),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_195),
.A2(n_187),
.B1(n_6),
.B2(n_7),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_197),
.B(n_198),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_196),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_200),
.Y(n_201)
);

AOI321xp33_ASAP7_75t_L g202 ( 
.A1(n_201),
.A2(n_193),
.A3(n_199),
.B1(n_10),
.B2(n_7),
.C(n_8),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_8),
.Y(n_203)
);


endmodule