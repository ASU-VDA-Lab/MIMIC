module real_aes_674_n_3 (n_0, n_2, n_1, n_3);
input n_0;
input n_2;
input n_1;
output n_3;
wire n_16;
wire n_13;
wire n_4;
wire n_5;
wire n_15;
wire n_7;
wire n_8;
wire n_9;
wire n_6;
wire n_12;
wire n_14;
wire n_10;
wire n_11;
INVx1_ASAP7_75t_L g16 ( .A(n_0), .Y(n_16) );
INVx1_ASAP7_75t_L g8 ( .A(n_1), .Y(n_8) );
INVx1_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
AND2x2_ASAP7_75t_L g12 ( .A(n_2), .B(n_8), .Y(n_12) );
A2O1A1Ixp33_ASAP7_75t_L g3 ( .A1(n_4), .A2(n_5), .B(n_9), .C(n_13), .Y(n_3) );
INVx1_ASAP7_75t_L g5 ( .A(n_6), .Y(n_5) );
INVx3_ASAP7_75t_L g6 ( .A(n_7), .Y(n_6) );
INVx2_ASAP7_75t_L g7 ( .A(n_8), .Y(n_7) );
INVxp67_ASAP7_75t_L g9 ( .A(n_10), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_11), .Y(n_10) );
BUFx3_ASAP7_75t_L g11 ( .A(n_12), .Y(n_11) );
CKINVDCx16_ASAP7_75t_R g13 ( .A(n_14), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_15), .Y(n_14) );
HB1xp67_ASAP7_75t_L g15 ( .A(n_16), .Y(n_15) );
endmodule