module fake_jpeg_12050_n_475 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_475);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_475;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_384;
wire n_296;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_10),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_8),
.Y(n_56)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_60),
.Y(n_140)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx11_ASAP7_75t_L g150 ( 
.A(n_62),
.Y(n_150)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_63),
.Y(n_152)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_64),
.Y(n_143)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_65),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_66),
.Y(n_146)
);

INVx4_ASAP7_75t_SL g67 ( 
.A(n_39),
.Y(n_67)
);

INVx13_ASAP7_75t_L g176 ( 
.A(n_67),
.Y(n_176)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_68),
.Y(n_177)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_70),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_42),
.B(n_16),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_72),
.B(n_98),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_19),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_75),
.Y(n_147)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_78),
.Y(n_185)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_79),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_80),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_82),
.Y(n_174)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_83),
.Y(n_158)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_84),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_26),
.B(n_14),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_85),
.B(n_102),
.Y(n_134)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_86),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g160 ( 
.A(n_87),
.Y(n_160)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_24),
.Y(n_90)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_90),
.Y(n_157)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_17),
.Y(n_91)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_91),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g171 ( 
.A(n_92),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

NAND2xp33_ASAP7_75t_SL g167 ( 
.A(n_93),
.B(n_100),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_94),
.Y(n_184)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_33),
.Y(n_95)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_95),
.Y(n_170)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_96),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_97),
.Y(n_173)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_23),
.Y(n_98)
);

BUFx12_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

BUFx16f_ASAP7_75t_L g138 ( 
.A(n_99),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_24),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_106),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_40),
.B(n_14),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_20),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_104),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_24),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_23),
.A2(n_12),
.B(n_3),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_105),
.A2(n_57),
.B(n_22),
.C(n_43),
.Y(n_165)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_41),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_41),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_108),
.Y(n_132)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_56),
.B(n_1),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_109),
.B(n_113),
.Y(n_118)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_110),
.B(n_111),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_45),
.B(n_3),
.Y(n_111)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_21),
.Y(n_112)
);

BUFx12_ASAP7_75t_L g183 ( 
.A(n_112),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_45),
.B(n_3),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_22),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_114),
.B(n_57),
.Y(n_180)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_28),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_115),
.B(n_47),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_25),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_120),
.B(n_135),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_61),
.A2(n_27),
.B1(n_54),
.B2(n_53),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_121),
.A2(n_145),
.B(n_164),
.Y(n_216)
);

CKINVDCx12_ASAP7_75t_R g130 ( 
.A(n_99),
.Y(n_130)
);

BUFx8_ASAP7_75t_L g212 ( 
.A(n_130),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_109),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_113),
.B(n_25),
.Y(n_136)
);

NAND3xp33_ASAP7_75t_L g238 ( 
.A(n_136),
.B(n_178),
.C(n_179),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_74),
.B(n_20),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_141),
.B(n_144),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_73),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_112),
.A2(n_29),
.B1(n_54),
.B2(n_53),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_74),
.B(n_38),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_149),
.B(n_151),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_80),
.B(n_38),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_80),
.B(n_48),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_155),
.B(n_162),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_90),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_161),
.B(n_166),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_101),
.B(n_48),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_76),
.A2(n_27),
.B1(n_54),
.B2(n_53),
.Y(n_164)
);

OAI21xp33_ASAP7_75t_L g237 ( 
.A1(n_165),
.A2(n_138),
.B(n_183),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_97),
.B(n_43),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_83),
.A2(n_27),
.B1(n_54),
.B2(n_53),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_172),
.A2(n_181),
.B1(n_182),
.B2(n_7),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_67),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_95),
.B(n_47),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_96),
.B(n_34),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_180),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_60),
.A2(n_34),
.B1(n_28),
.B2(n_29),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_100),
.A2(n_29),
.B1(n_27),
.B2(n_24),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_186),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_187),
.B(n_190),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_167),
.A2(n_29),
.B1(n_94),
.B2(n_75),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_189),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_3),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_118),
.B(n_4),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_191),
.B(n_235),
.Y(n_265)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_143),
.Y(n_192)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_192),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_165),
.A2(n_77),
.B1(n_89),
.B2(n_87),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_193),
.A2(n_194),
.B(n_208),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_122),
.A2(n_92),
.B1(n_82),
.B2(n_81),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_182),
.A2(n_66),
.B1(n_7),
.B2(n_8),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_195),
.A2(n_198),
.B1(n_199),
.B2(n_211),
.Y(n_268)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_140),
.Y(n_196)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_196),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_173),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_197),
.A2(n_206),
.B1(n_221),
.B2(n_231),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_164),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_167),
.A2(n_9),
.B1(n_10),
.B2(n_158),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_200),
.A2(n_218),
.B1(n_228),
.B2(n_236),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_180),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_201),
.B(n_205),
.Y(n_258)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_140),
.Y(n_203)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_203),
.Y(n_282)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_123),
.Y(n_204)
);

INVx6_ASAP7_75t_L g286 ( 
.A(n_204),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_117),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_129),
.A2(n_9),
.B1(n_153),
.B2(n_184),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_157),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_207),
.B(n_213),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_134),
.A2(n_132),
.B1(n_116),
.B2(n_170),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_125),
.B(n_163),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_209),
.B(n_187),
.C(n_202),
.Y(n_259)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_170),
.Y(n_210)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_210),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_172),
.A2(n_121),
.B1(n_145),
.B2(n_184),
.Y(n_211)
);

FAx1_ASAP7_75t_SL g213 ( 
.A(n_128),
.B(n_150),
.CI(n_154),
.CON(n_213),
.SN(n_213)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_183),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_215),
.B(n_240),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_123),
.A2(n_174),
.B1(n_139),
.B2(n_147),
.Y(n_218)
);

O2A1O1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_168),
.A2(n_176),
.B(n_150),
.C(n_128),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_219),
.A2(n_244),
.B(n_193),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_159),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_220),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_139),
.A2(n_174),
.B1(n_147),
.B2(n_146),
.Y(n_221)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_131),
.Y(n_223)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_223),
.Y(n_247)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_169),
.Y(n_224)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_224),
.Y(n_257)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_126),
.Y(n_225)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_131),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_126),
.Y(n_227)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_227),
.Y(n_283)
);

OA22x2_ASAP7_75t_L g228 ( 
.A1(n_146),
.A2(n_119),
.B1(n_152),
.B2(n_169),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_158),
.Y(n_229)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_229),
.Y(n_256)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_177),
.Y(n_230)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_230),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_160),
.A2(n_133),
.B1(n_127),
.B2(n_116),
.Y(n_231)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_131),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_232),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_160),
.A2(n_133),
.B1(n_127),
.B2(n_119),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_234),
.A2(n_246),
.B1(n_243),
.B2(n_194),
.Y(n_279)
);

AO22x1_ASAP7_75t_SL g235 ( 
.A1(n_142),
.A2(n_185),
.B1(n_124),
.B2(n_176),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_152),
.A2(n_171),
.B1(n_177),
.B2(n_185),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_237),
.A2(n_202),
.B1(n_201),
.B2(n_244),
.Y(n_260)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_142),
.Y(n_239)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_239),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_124),
.Y(n_240)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_240),
.Y(n_278)
);

NAND2x1_ASAP7_75t_SL g241 ( 
.A(n_138),
.B(n_183),
.Y(n_241)
);

BUFx8_ASAP7_75t_L g255 ( 
.A(n_241),
.Y(n_255)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_171),
.Y(n_242)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_242),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_171),
.A2(n_137),
.B1(n_148),
.B2(n_138),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_243),
.A2(n_216),
.B1(n_239),
.B2(n_229),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_137),
.A2(n_175),
.B1(n_156),
.B2(n_165),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_148),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_245),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_173),
.A2(n_76),
.B1(n_83),
.B2(n_95),
.Y(n_246)
);

AND2x2_ASAP7_75t_SL g250 ( 
.A(n_190),
.B(n_209),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_250),
.B(n_267),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_259),
.B(n_274),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_260),
.Y(n_303)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_210),
.Y(n_261)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_261),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_209),
.B(n_187),
.C(n_208),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_264),
.B(n_242),
.C(n_213),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_191),
.B(n_222),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_271),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_238),
.B(n_217),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_273),
.B(n_275),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_241),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_214),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_277),
.B(n_281),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_279),
.A2(n_294),
.B1(n_219),
.B2(n_228),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_233),
.B(n_188),
.Y(n_281)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_235),
.Y(n_285)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_285),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_288),
.A2(n_292),
.B1(n_232),
.B2(n_212),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_207),
.B(n_230),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_265),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_236),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_291),
.B(n_293),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_211),
.A2(n_216),
.B1(n_218),
.B2(n_228),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_225),
.B(n_224),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_228),
.A2(n_204),
.B1(n_203),
.B2(n_196),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_250),
.B(n_227),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_297),
.B(n_306),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_258),
.B(n_235),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_298),
.B(n_313),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_299),
.A2(n_311),
.B1(n_318),
.B2(n_287),
.Y(n_347)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_249),
.Y(n_300)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_300),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_290),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_301),
.B(n_312),
.Y(n_339)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_249),
.Y(n_302)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_302),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_304),
.B(n_317),
.C(n_319),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_262),
.A2(n_213),
.B(n_212),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_305),
.A2(n_321),
.B(n_248),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_250),
.B(n_223),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_267),
.A2(n_285),
.B(n_289),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_307),
.A2(n_325),
.B(n_257),
.Y(n_354)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_256),
.Y(n_308)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_308),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_309),
.B(n_310),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_265),
.B(n_226),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_272),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_270),
.B(n_212),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_252),
.B(n_264),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_314),
.B(n_331),
.Y(n_355)
);

INVx6_ASAP7_75t_L g315 ( 
.A(n_286),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_252),
.B(n_259),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_316),
.B(n_323),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_289),
.B(n_271),
.C(n_280),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_288),
.A2(n_294),
.B1(n_280),
.B2(n_269),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_255),
.A2(n_254),
.B(n_278),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_274),
.B(n_261),
.Y(n_323)
);

OR2x4_ASAP7_75t_L g325 ( 
.A(n_255),
.B(n_268),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_255),
.A2(n_268),
.B(n_278),
.Y(n_327)
);

OR2x2_ASAP7_75t_L g348 ( 
.A(n_327),
.B(n_251),
.Y(n_348)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_256),
.Y(n_328)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_328),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_266),
.B(n_284),
.C(n_253),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_330),
.B(n_287),
.C(n_283),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_284),
.B(n_251),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_323),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_332),
.B(n_333),
.Y(n_367)
);

AND2x6_ASAP7_75t_L g333 ( 
.A(n_317),
.B(n_248),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_295),
.A2(n_286),
.B1(n_282),
.B2(n_263),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_336),
.A2(n_308),
.B1(n_328),
.B2(n_312),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_319),
.B(n_266),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_341),
.B(n_358),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_318),
.A2(n_282),
.B1(n_263),
.B2(n_248),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_342),
.A2(n_344),
.B1(n_347),
.B2(n_329),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_307),
.A2(n_309),
.B1(n_299),
.B2(n_295),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_345),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_331),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_346),
.B(n_349),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_348),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_329),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_321),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_350),
.B(n_359),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_322),
.B(n_276),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_352),
.B(n_313),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_354),
.A2(n_327),
.B(n_298),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_314),
.B(n_283),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_356),
.B(n_360),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_316),
.B(n_257),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_320),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_361),
.A2(n_362),
.B1(n_384),
.B2(n_383),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_344),
.A2(n_329),
.B1(n_301),
.B2(n_310),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_364),
.A2(n_365),
.B(n_379),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_354),
.A2(n_324),
.B(n_305),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_334),
.Y(n_366)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_366),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_369),
.B(n_382),
.Y(n_386)
);

OAI22x1_ASAP7_75t_L g370 ( 
.A1(n_348),
.A2(n_325),
.B1(n_303),
.B2(n_304),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_370),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_373),
.B(n_380),
.Y(n_389)
);

CKINVDCx14_ASAP7_75t_R g375 ( 
.A(n_339),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_375),
.B(n_346),
.Y(n_403)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_334),
.Y(n_377)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_377),
.Y(n_396)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_335),
.Y(n_378)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_378),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_350),
.A2(n_306),
.B(n_297),
.Y(n_379)
);

OA21x2_ASAP7_75t_SL g380 ( 
.A1(n_359),
.A2(n_296),
.B(n_302),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_335),
.Y(n_381)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_381),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_348),
.A2(n_296),
.B1(n_330),
.B2(n_300),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_336),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_383),
.B(n_332),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_342),
.A2(n_315),
.B1(n_326),
.B2(n_247),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_353),
.Y(n_385)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_385),
.Y(n_406)
);

AOI21x1_ASAP7_75t_L g387 ( 
.A1(n_364),
.A2(n_345),
.B(n_351),
.Y(n_387)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_387),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_363),
.B(n_340),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_SL g410 ( 
.A(n_388),
.B(n_343),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_376),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_390),
.B(n_398),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_374),
.B(n_363),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_391),
.B(n_399),
.C(n_401),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_376),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_392),
.B(n_351),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_379),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_374),
.B(n_340),
.C(n_356),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_382),
.B(n_355),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_370),
.B(n_358),
.C(n_341),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_402),
.B(n_360),
.C(n_343),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_403),
.B(n_337),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_404),
.Y(n_419)
);

AOI21x1_ASAP7_75t_SL g414 ( 
.A1(n_405),
.A2(n_390),
.B(n_371),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_389),
.A2(n_367),
.B1(n_361),
.B2(n_372),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_408),
.A2(n_409),
.B1(n_412),
.B2(n_420),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_386),
.A2(n_367),
.B1(n_372),
.B2(n_365),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_410),
.B(n_415),
.Y(n_425)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_405),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_411),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_386),
.A2(n_362),
.B1(n_368),
.B2(n_371),
.Y(n_412)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_414),
.Y(n_429)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_416),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_399),
.B(n_368),
.C(n_349),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_418),
.B(n_388),
.C(n_394),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_394),
.Y(n_420)
);

OR2x2_ASAP7_75t_L g431 ( 
.A(n_421),
.B(n_401),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_391),
.B(n_333),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_422),
.B(n_423),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_402),
.B(n_337),
.Y(n_423)
);

MAJx2_ASAP7_75t_L g440 ( 
.A(n_424),
.B(n_434),
.C(n_436),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_417),
.A2(n_395),
.B(n_422),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_427),
.A2(n_432),
.B(n_407),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_431),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_417),
.A2(n_395),
.B(n_398),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_413),
.B(n_387),
.C(n_338),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_433),
.B(n_437),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_413),
.B(n_406),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_423),
.B(n_406),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_415),
.B(n_400),
.C(n_397),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_426),
.B(n_418),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_438),
.B(n_424),
.C(n_440),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_441),
.A2(n_433),
.B(n_436),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_437),
.B(n_412),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_443),
.B(n_444),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_434),
.B(n_419),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_429),
.A2(n_407),
.B1(n_414),
.B2(n_369),
.Y(n_445)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_445),
.Y(n_450)
);

AOI221xp5_ASAP7_75t_L g446 ( 
.A1(n_430),
.A2(n_410),
.B1(n_400),
.B2(n_397),
.C(n_396),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_446),
.B(n_447),
.Y(n_453)
);

AOI221xp5_ASAP7_75t_L g447 ( 
.A1(n_435),
.A2(n_396),
.B1(n_393),
.B2(n_366),
.C(n_378),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_439),
.B(n_428),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_448),
.B(n_449),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_442),
.B(n_431),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_452),
.B(n_440),
.Y(n_456)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_454),
.Y(n_458)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_445),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_455),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_456),
.B(n_457),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_452),
.B(n_438),
.C(n_425),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_451),
.B(n_425),
.C(n_426),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_459),
.B(n_460),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_454),
.B(n_441),
.C(n_393),
.Y(n_460)
);

INVxp33_ASAP7_75t_L g463 ( 
.A(n_461),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_463),
.A2(n_466),
.B(n_458),
.Y(n_469)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_462),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_465),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_458),
.A2(n_450),
.B1(n_453),
.B2(n_384),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_469),
.B(n_377),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_464),
.A2(n_385),
.B(n_381),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_470),
.A2(n_467),
.B(n_463),
.Y(n_471)
);

NOR3xp33_ASAP7_75t_L g473 ( 
.A(n_471),
.B(n_472),
.C(n_468),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_473),
.A2(n_357),
.B(n_353),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_474),
.B(n_357),
.Y(n_475)
);


endmodule