module fake_jpeg_25103_n_125 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_125);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVxp33_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_25),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_29),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx4f_ASAP7_75t_SL g71 ( 
.A(n_56),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_46),
.Y(n_68)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_50),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_65),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_55),
.A2(n_51),
.B1(n_49),
.B2(n_48),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_63),
.A2(n_67),
.B1(n_1),
.B2(n_2),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_44),
.C(n_46),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_54),
.A2(n_47),
.B1(n_42),
.B2(n_40),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_72),
.Y(n_85)
);

OR2x2_ASAP7_75t_SL g69 ( 
.A(n_57),
.B(n_1),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_69),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_84)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_83),
.Y(n_93)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_77),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_39),
.B1(n_45),
.B2(n_20),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_76),
.A2(n_79),
.B1(n_7),
.B2(n_8),
.Y(n_97)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_82),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_70),
.A2(n_36),
.B1(n_18),
.B2(n_21),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_81),
.A2(n_82),
.B1(n_87),
.B2(n_76),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_64),
.B(n_2),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_86),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_3),
.Y(n_86)
);

INVx3_ASAP7_75t_SL g87 ( 
.A(n_71),
.Y(n_87)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_6),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_7),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_23),
.C(n_35),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_84),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_6),
.Y(n_95)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_98),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_99),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_103),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_94),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_89),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_104),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_89),
.A2(n_79),
.B(n_12),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_105),
.A2(n_96),
.B(n_98),
.Y(n_108)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_108),
.A2(n_101),
.B(n_106),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_102),
.A2(n_90),
.B1(n_91),
.B2(n_93),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_105),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_113),
.A2(n_114),
.B1(n_111),
.B2(n_108),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_100),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_117),
.A2(n_110),
.B(n_116),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_9),
.C(n_13),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_119),
.A2(n_14),
.B(n_16),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_120),
.A2(n_17),
.B(n_22),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_121),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_24),
.B(n_28),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_31),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_34),
.Y(n_125)
);


endmodule