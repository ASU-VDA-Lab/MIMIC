module fake_aes_3283_n_778 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_93, n_51, n_96, n_39, n_778);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_93;
input n_51;
input n_96;
input n_39;
output n_778;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_529;
wire n_455;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_581;
wire n_458;
wire n_504;
wire n_493;
wire n_418;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_79), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_42), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_53), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_85), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_25), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_5), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_77), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_33), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_28), .Y(n_105) );
NOR2xp67_ASAP7_75t_L g106 ( .A(n_94), .B(n_15), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_83), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_29), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_32), .Y(n_109) );
INVx1_ASAP7_75t_SL g110 ( .A(n_82), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_89), .Y(n_111) );
BUFx6f_ASAP7_75t_L g112 ( .A(n_41), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_81), .Y(n_113) );
INVxp67_ASAP7_75t_L g114 ( .A(n_48), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_59), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_51), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_45), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_8), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_62), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_56), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_9), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_57), .Y(n_122) );
BUFx2_ASAP7_75t_L g123 ( .A(n_1), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_58), .Y(n_124) );
INVxp67_ASAP7_75t_SL g125 ( .A(n_1), .Y(n_125) );
CKINVDCx16_ASAP7_75t_R g126 ( .A(n_64), .Y(n_126) );
XOR2xp5_ASAP7_75t_L g127 ( .A(n_50), .B(n_86), .Y(n_127) );
INVx1_ASAP7_75t_SL g128 ( .A(n_54), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_78), .Y(n_129) );
INVxp33_ASAP7_75t_SL g130 ( .A(n_34), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_5), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_76), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_131), .B(n_0), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_131), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_98), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_112), .Y(n_136) );
INVx3_ASAP7_75t_L g137 ( .A(n_102), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_112), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_112), .Y(n_139) );
AND2x6_ASAP7_75t_L g140 ( .A(n_99), .B(n_17), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_100), .Y(n_141) );
OAI22xp5_ASAP7_75t_L g142 ( .A1(n_123), .A2(n_0), .B1(n_2), .B2(n_3), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_126), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_118), .B(n_2), .Y(n_144) );
AND2x4_ASAP7_75t_L g145 ( .A(n_103), .B(n_3), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_112), .B(n_4), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_104), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_105), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_107), .Y(n_149) );
INVx4_ASAP7_75t_L g150 ( .A(n_112), .Y(n_150) );
OAI21x1_ASAP7_75t_L g151 ( .A1(n_108), .A2(n_44), .B(n_95), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_118), .B(n_4), .Y(n_152) );
OAI22xp5_ASAP7_75t_L g153 ( .A1(n_121), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_153) );
AOI22xp5_ASAP7_75t_L g154 ( .A1(n_130), .A2(n_6), .B1(n_7), .B2(n_9), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_109), .Y(n_155) );
INVx4_ASAP7_75t_SL g156 ( .A(n_140), .Y(n_156) );
AOI22xp33_ASAP7_75t_L g157 ( .A1(n_133), .A2(n_130), .B1(n_121), .B2(n_125), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_133), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_150), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_133), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_145), .B(n_106), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_133), .Y(n_162) );
AOI22xp33_ASAP7_75t_L g163 ( .A1(n_145), .A2(n_111), .B1(n_113), .B2(n_116), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_150), .Y(n_164) );
BUFx3_ASAP7_75t_L g165 ( .A(n_140), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_150), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_135), .B(n_97), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_145), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_145), .Y(n_169) );
BUFx3_ASAP7_75t_L g170 ( .A(n_140), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_134), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_135), .B(n_114), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_134), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_147), .B(n_119), .Y(n_174) );
AOI22xp33_ASAP7_75t_L g175 ( .A1(n_140), .A2(n_120), .B1(n_124), .B2(n_97), .Y(n_175) );
INVx3_ASAP7_75t_L g176 ( .A(n_137), .Y(n_176) );
INVx2_ASAP7_75t_SL g177 ( .A(n_147), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_148), .B(n_132), .Y(n_178) );
INVx1_ASAP7_75t_SL g179 ( .A(n_143), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_137), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_148), .B(n_132), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_155), .B(n_117), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_137), .Y(n_183) );
BUFx3_ASAP7_75t_L g184 ( .A(n_140), .Y(n_184) );
AOI22xp33_ASAP7_75t_L g185 ( .A1(n_140), .A2(n_117), .B1(n_101), .B2(n_122), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_136), .Y(n_186) );
OR2x2_ASAP7_75t_L g187 ( .A(n_143), .B(n_129), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_141), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_141), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_149), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_149), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_155), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_144), .B(n_129), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_167), .B(n_152), .Y(n_194) );
A2O1A1Ixp33_ASAP7_75t_SL g195 ( .A1(n_174), .A2(n_154), .B(n_142), .C(n_153), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_176), .Y(n_196) );
INVx8_ASAP7_75t_L g197 ( .A(n_161), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_180), .Y(n_198) );
INVx3_ASAP7_75t_L g199 ( .A(n_176), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_182), .B(n_101), .Y(n_200) );
INVx3_ASAP7_75t_L g201 ( .A(n_176), .Y(n_201) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_157), .A2(n_115), .B1(n_127), .B2(n_122), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_179), .B(n_115), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_161), .B(n_151), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_177), .B(n_140), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_170), .B(n_151), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_180), .Y(n_207) );
INVx2_ASAP7_75t_SL g208 ( .A(n_187), .Y(n_208) );
O2A1O1Ixp5_ASAP7_75t_L g209 ( .A1(n_178), .A2(n_146), .B(n_128), .C(n_110), .Y(n_209) );
INVxp33_ASAP7_75t_L g210 ( .A(n_187), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_183), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_170), .B(n_139), .Y(n_212) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_170), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_177), .B(n_139), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_181), .B(n_139), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_165), .B(n_139), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_193), .B(n_52), .Y(n_217) );
NAND2x1p5_ASAP7_75t_L g218 ( .A(n_176), .B(n_139), .Y(n_218) );
CKINVDCx5p33_ASAP7_75t_R g219 ( .A(n_163), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_158), .A2(n_138), .B(n_136), .C(n_12), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_168), .A2(n_138), .B(n_136), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_183), .Y(n_222) );
BUFx12f_ASAP7_75t_L g223 ( .A(n_161), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_165), .B(n_138), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_188), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_188), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_161), .B(n_49), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_192), .B(n_138), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_189), .Y(n_229) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_184), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_171), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_192), .B(n_138), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_171), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_172), .B(n_47), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_184), .B(n_136), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g236 ( .A1(n_219), .A2(n_168), .B1(n_169), .B2(n_162), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_208), .B(n_156), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_231), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_230), .B(n_156), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g240 ( .A1(n_231), .A2(n_169), .B(n_160), .C(n_162), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_205), .A2(n_158), .B(n_160), .Y(n_241) );
OR2x6_ASAP7_75t_SL g242 ( .A(n_202), .B(n_191), .Y(n_242) );
OR2x6_ASAP7_75t_L g243 ( .A(n_197), .B(n_173), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_194), .B(n_185), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_210), .B(n_175), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_198), .Y(n_246) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_233), .A2(n_191), .B(n_190), .C(n_189), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_233), .A2(n_190), .B(n_173), .C(n_159), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_200), .B(n_197), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_206), .A2(n_164), .B(n_166), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_207), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_230), .B(n_156), .Y(n_252) );
AO32x1_ASAP7_75t_L g253 ( .A1(n_225), .A2(n_186), .A3(n_136), .B1(n_159), .B2(n_166), .Y(n_253) );
INVx5_ASAP7_75t_L g254 ( .A(n_213), .Y(n_254) );
NAND3xp33_ASAP7_75t_L g255 ( .A(n_227), .B(n_164), .C(n_186), .Y(n_255) );
INVx1_ASAP7_75t_SL g256 ( .A(n_203), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_197), .B(n_156), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_197), .B(n_156), .Y(n_258) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_223), .Y(n_259) );
BUFx12f_ASAP7_75t_L g260 ( .A(n_223), .Y(n_260) );
OAI22xp5_ASAP7_75t_SL g261 ( .A1(n_210), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_226), .B(n_164), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_L g263 ( .A1(n_195), .A2(n_164), .B(n_11), .C(n_13), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_229), .B(n_10), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_206), .A2(n_55), .B(n_93), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_199), .B(n_13), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g267 ( .A(n_217), .Y(n_267) );
NOR3xp33_ASAP7_75t_L g268 ( .A(n_195), .B(n_14), .C(n_15), .Y(n_268) );
AOI221xp5_ASAP7_75t_L g269 ( .A1(n_256), .A2(n_209), .B1(n_211), .B2(n_222), .C(n_204), .Y(n_269) );
OAI21xp5_ASAP7_75t_L g270 ( .A1(n_241), .A2(n_204), .B(n_221), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_256), .B(n_201), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_242), .B(n_199), .Y(n_272) );
OAI21xp33_ASAP7_75t_SL g273 ( .A1(n_243), .A2(n_234), .B(n_196), .Y(n_273) );
INVx1_ASAP7_75t_SL g274 ( .A(n_260), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_238), .B(n_204), .Y(n_275) );
INVx4_ASAP7_75t_L g276 ( .A(n_243), .Y(n_276) );
OAI22xp5_ASAP7_75t_L g277 ( .A1(n_243), .A2(n_196), .B1(n_201), .B2(n_215), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_264), .Y(n_278) );
BUFx8_ASAP7_75t_L g279 ( .A(n_246), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_251), .Y(n_280) );
AO31x2_ASAP7_75t_L g281 ( .A1(n_240), .A2(n_220), .A3(n_232), .B(n_228), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_259), .Y(n_282) );
A2O1A1Ixp33_ASAP7_75t_L g283 ( .A1(n_263), .A2(n_220), .B(n_214), .C(n_212), .Y(n_283) );
OA22x2_ASAP7_75t_L g284 ( .A1(n_261), .A2(n_235), .B1(n_224), .B2(n_216), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_267), .Y(n_285) );
OAI21x1_ASAP7_75t_SL g286 ( .A1(n_236), .A2(n_14), .B(n_16), .Y(n_286) );
AOI31xp67_ASAP7_75t_L g287 ( .A1(n_253), .A2(n_212), .A3(n_224), .B(n_216), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_262), .Y(n_288) );
INVxp67_ASAP7_75t_L g289 ( .A(n_249), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_250), .A2(n_235), .B(n_213), .Y(n_290) );
INVxp67_ASAP7_75t_SL g291 ( .A(n_266), .Y(n_291) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_279), .Y(n_292) );
INVx2_ASAP7_75t_SL g293 ( .A(n_279), .Y(n_293) );
BUFx3_ASAP7_75t_L g294 ( .A(n_276), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_280), .B(n_244), .Y(n_295) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_289), .Y(n_296) );
AO31x2_ASAP7_75t_L g297 ( .A1(n_283), .A2(n_247), .A3(n_248), .B(n_265), .Y(n_297) );
A2O1A1Ixp33_ASAP7_75t_L g298 ( .A1(n_278), .A2(n_245), .B(n_268), .C(n_255), .Y(n_298) );
BUFx2_ASAP7_75t_R g299 ( .A(n_285), .Y(n_299) );
OAI21x1_ASAP7_75t_L g300 ( .A1(n_270), .A2(n_253), .B(n_239), .Y(n_300) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_276), .Y(n_301) );
OAI21x1_ASAP7_75t_L g302 ( .A1(n_290), .A2(n_253), .B(n_252), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_272), .B(n_237), .Y(n_303) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_274), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_288), .B(n_254), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_275), .B(n_254), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_287), .Y(n_307) );
AND2x4_ASAP7_75t_L g308 ( .A(n_275), .B(n_254), .Y(n_308) );
NAND2x1p5_ASAP7_75t_L g309 ( .A(n_271), .B(n_254), .Y(n_309) );
CKINVDCx11_ASAP7_75t_R g310 ( .A(n_282), .Y(n_310) );
OAI21x1_ASAP7_75t_L g311 ( .A1(n_277), .A2(n_218), .B(n_257), .Y(n_311) );
OAI21x1_ASAP7_75t_L g312 ( .A1(n_291), .A2(n_218), .B(n_258), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_281), .Y(n_313) );
OAI21x1_ASAP7_75t_L g314 ( .A1(n_291), .A2(n_213), .B(n_230), .Y(n_314) );
A2O1A1Ixp33_ASAP7_75t_L g315 ( .A1(n_273), .A2(n_213), .B(n_230), .C(n_16), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_271), .B(n_18), .Y(n_316) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_284), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_317), .B(n_281), .Y(n_318) );
AO21x2_ASAP7_75t_L g319 ( .A1(n_307), .A2(n_283), .B(n_286), .Y(n_319) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_309), .Y(n_320) );
OA21x2_ASAP7_75t_L g321 ( .A1(n_307), .A2(n_269), .B(n_281), .Y(n_321) );
BUFx2_ASAP7_75t_R g322 ( .A(n_294), .Y(n_322) );
BUFx12f_ASAP7_75t_L g323 ( .A(n_310), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_307), .Y(n_324) );
AO21x2_ASAP7_75t_L g325 ( .A1(n_313), .A2(n_281), .B(n_284), .Y(n_325) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_309), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_313), .Y(n_327) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_309), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_300), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_300), .Y(n_330) );
AO21x2_ASAP7_75t_L g331 ( .A1(n_315), .A2(n_19), .B(n_20), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_305), .B(n_21), .Y(n_332) );
AO21x2_ASAP7_75t_L g333 ( .A1(n_302), .A2(n_22), .B(n_23), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_295), .Y(n_334) );
OA21x2_ASAP7_75t_L g335 ( .A1(n_302), .A2(n_24), .B(n_26), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_314), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_295), .B(n_27), .Y(n_337) );
OR2x2_ASAP7_75t_L g338 ( .A(n_303), .B(n_30), .Y(n_338) );
INVx3_ASAP7_75t_L g339 ( .A(n_301), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_314), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_312), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_299), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_303), .B(n_31), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_305), .B(n_35), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_312), .Y(n_345) );
AND2x4_ASAP7_75t_L g346 ( .A(n_306), .B(n_96), .Y(n_346) );
AO21x2_ASAP7_75t_L g347 ( .A1(n_298), .A2(n_36), .B(n_37), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_297), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_297), .Y(n_349) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_301), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_297), .Y(n_351) );
INVx3_ASAP7_75t_L g352 ( .A(n_301), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_301), .Y(n_353) );
AO21x2_ASAP7_75t_L g354 ( .A1(n_311), .A2(n_38), .B(n_39), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_297), .Y(n_355) );
AND2x2_ASAP7_75t_SL g356 ( .A(n_316), .B(n_40), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_297), .Y(n_357) );
OAI21x1_ASAP7_75t_L g358 ( .A1(n_311), .A2(n_43), .B(n_46), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_297), .B(n_60), .Y(n_359) );
OR2x2_ASAP7_75t_L g360 ( .A(n_318), .B(n_296), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_324), .Y(n_361) );
INVx2_ASAP7_75t_SL g362 ( .A(n_320), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_327), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_324), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_324), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_318), .B(n_308), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_318), .B(n_308), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_334), .B(n_304), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_324), .Y(n_369) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_336), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_327), .Y(n_371) );
INVxp67_ASAP7_75t_L g372 ( .A(n_320), .Y(n_372) );
INVx4_ASAP7_75t_L g373 ( .A(n_356), .Y(n_373) );
INVx4_ASAP7_75t_R g374 ( .A(n_332), .Y(n_374) );
INVx4_ASAP7_75t_L g375 ( .A(n_356), .Y(n_375) );
INVx2_ASAP7_75t_SL g376 ( .A(n_326), .Y(n_376) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_326), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_325), .B(n_308), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_325), .B(n_308), .Y(n_379) );
INVx1_ASAP7_75t_SL g380 ( .A(n_322), .Y(n_380) );
INVx2_ASAP7_75t_SL g381 ( .A(n_328), .Y(n_381) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_336), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_325), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_336), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_325), .Y(n_385) );
BUFx2_ASAP7_75t_L g386 ( .A(n_350), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_325), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_359), .B(n_306), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_359), .B(n_306), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_359), .B(n_306), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_334), .B(n_355), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_355), .B(n_301), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_348), .B(n_301), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_348), .B(n_294), .Y(n_394) );
INVx3_ASAP7_75t_L g395 ( .A(n_339), .Y(n_395) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_328), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_348), .B(n_294), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_348), .B(n_316), .Y(n_398) );
AND2x4_ASAP7_75t_L g399 ( .A(n_349), .B(n_293), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_349), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_336), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_349), .B(n_293), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_350), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_349), .B(n_292), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_351), .B(n_61), .Y(n_405) );
INVxp33_ASAP7_75t_L g406 ( .A(n_332), .Y(n_406) );
AND2x4_ASAP7_75t_L g407 ( .A(n_351), .B(n_63), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_351), .B(n_65), .Y(n_408) );
INVx4_ASAP7_75t_L g409 ( .A(n_356), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_351), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_357), .B(n_66), .Y(n_411) );
INVxp67_ASAP7_75t_SL g412 ( .A(n_353), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_357), .B(n_67), .Y(n_413) );
AND2x4_ASAP7_75t_L g414 ( .A(n_357), .B(n_68), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_329), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_353), .Y(n_416) );
BUFx2_ASAP7_75t_L g417 ( .A(n_339), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_357), .B(n_69), .Y(n_418) );
NOR2xp67_ASAP7_75t_L g419 ( .A(n_339), .B(n_70), .Y(n_419) );
BUFx3_ASAP7_75t_L g420 ( .A(n_339), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_329), .Y(n_421) );
INVx3_ASAP7_75t_L g422 ( .A(n_339), .Y(n_422) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_332), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_338), .B(n_71), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_329), .Y(n_425) );
NOR2x1_ASAP7_75t_SL g426 ( .A(n_338), .B(n_299), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_338), .B(n_72), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_341), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_341), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_342), .B(n_73), .Y(n_430) );
INVx1_ASAP7_75t_SL g431 ( .A(n_322), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_319), .B(n_74), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_344), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_360), .B(n_343), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_363), .B(n_319), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_363), .B(n_319), .Y(n_436) );
AND2x4_ASAP7_75t_L g437 ( .A(n_399), .B(n_352), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_391), .B(n_319), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_368), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_360), .B(n_343), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_386), .Y(n_441) );
INVx2_ASAP7_75t_SL g442 ( .A(n_386), .Y(n_442) );
AND2x4_ASAP7_75t_L g443 ( .A(n_399), .B(n_352), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_373), .A2(n_356), .B1(n_342), .B2(n_344), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_404), .B(n_344), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_404), .B(n_352), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_433), .B(n_343), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_366), .B(n_352), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_423), .B(n_352), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_361), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_362), .B(n_319), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_371), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_361), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_391), .B(n_321), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_371), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_366), .B(n_346), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_361), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_371), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_402), .Y(n_459) );
NAND2x1p5_ASAP7_75t_L g460 ( .A(n_373), .B(n_346), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_367), .B(n_402), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_364), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_367), .B(n_346), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_377), .B(n_346), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_396), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_403), .Y(n_466) );
INVx2_ASAP7_75t_SL g467 ( .A(n_416), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_399), .B(n_321), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_362), .B(n_346), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_364), .Y(n_470) );
BUFx2_ASAP7_75t_SL g471 ( .A(n_380), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_399), .B(n_321), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_376), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_426), .B(n_337), .Y(n_474) );
AND2x4_ASAP7_75t_L g475 ( .A(n_378), .B(n_345), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_376), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_381), .B(n_333), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_381), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_406), .B(n_333), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_372), .B(n_321), .Y(n_480) );
INVx2_ASAP7_75t_SL g481 ( .A(n_374), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_388), .B(n_333), .Y(n_482) );
INVx3_ASAP7_75t_L g483 ( .A(n_373), .Y(n_483) );
NOR2x1_ASAP7_75t_L g484 ( .A(n_380), .B(n_354), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_388), .B(n_389), .Y(n_485) );
AND2x4_ASAP7_75t_L g486 ( .A(n_378), .B(n_345), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_389), .B(n_333), .Y(n_487) );
BUFx2_ASAP7_75t_L g488 ( .A(n_412), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_390), .B(n_321), .Y(n_489) );
BUFx2_ASAP7_75t_L g490 ( .A(n_431), .Y(n_490) );
INVx3_ASAP7_75t_L g491 ( .A(n_373), .Y(n_491) );
INVxp67_ASAP7_75t_SL g492 ( .A(n_384), .Y(n_492) );
OR2x6_ASAP7_75t_L g493 ( .A(n_375), .B(n_323), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_390), .B(n_333), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_400), .B(n_321), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_379), .B(n_354), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_379), .B(n_354), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_428), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_428), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_400), .B(n_329), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_431), .B(n_354), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_394), .B(n_330), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_429), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_394), .B(n_354), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_364), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_410), .B(n_330), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_429), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_365), .Y(n_508) );
AND2x2_ASAP7_75t_SL g509 ( .A(n_375), .B(n_335), .Y(n_509) );
AND2x4_ASAP7_75t_L g510 ( .A(n_397), .B(n_330), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_365), .Y(n_511) );
NOR2xp67_ASAP7_75t_L g512 ( .A(n_375), .B(n_323), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_365), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_369), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_375), .B(n_409), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_369), .Y(n_516) );
AND2x4_ASAP7_75t_L g517 ( .A(n_397), .B(n_330), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_426), .B(n_347), .Y(n_518) );
AND2x4_ASAP7_75t_L g519 ( .A(n_393), .B(n_340), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_393), .B(n_409), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_409), .B(n_347), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_409), .B(n_347), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_369), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_417), .B(n_347), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_392), .B(n_337), .Y(n_525) );
INVx3_ASAP7_75t_L g526 ( .A(n_420), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_417), .B(n_347), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_432), .B(n_340), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_392), .Y(n_529) );
INVx5_ASAP7_75t_L g530 ( .A(n_407), .Y(n_530) );
INVx2_ASAP7_75t_SL g531 ( .A(n_374), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_410), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_432), .B(n_335), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_405), .B(n_335), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_461), .B(n_420), .Y(n_535) );
NOR2xp67_ASAP7_75t_SL g536 ( .A(n_530), .B(n_323), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_448), .B(n_420), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_490), .B(n_323), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_529), .B(n_383), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_471), .B(n_430), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_466), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_466), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_467), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_465), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_438), .B(n_383), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_498), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_438), .B(n_385), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_485), .B(n_395), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_499), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_503), .Y(n_550) );
AND2x4_ASAP7_75t_L g551 ( .A(n_493), .B(n_395), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_445), .B(n_395), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_507), .B(n_385), .Y(n_553) );
INVx1_ASAP7_75t_SL g554 ( .A(n_488), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_467), .B(n_398), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_435), .B(n_387), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_435), .B(n_387), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_520), .B(n_395), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_456), .B(n_422), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_463), .B(n_459), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_439), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_446), .B(n_422), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_532), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_436), .B(n_398), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_434), .B(n_401), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_475), .B(n_422), .Y(n_566) );
NOR2x1_ASAP7_75t_L g567 ( .A(n_493), .B(n_419), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_436), .B(n_415), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_452), .Y(n_569) );
AND2x4_ASAP7_75t_L g570 ( .A(n_493), .B(n_422), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_475), .B(n_414), .Y(n_571) );
AND2x4_ASAP7_75t_L g572 ( .A(n_512), .B(n_425), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_455), .Y(n_573) );
OAI21xp5_ASAP7_75t_L g574 ( .A1(n_444), .A2(n_427), .B(n_424), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_475), .B(n_414), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_454), .B(n_415), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_486), .B(n_414), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_458), .Y(n_578) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_441), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_486), .B(n_414), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_440), .B(n_384), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_474), .B(n_427), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_486), .B(n_407), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_473), .Y(n_584) );
NAND3xp33_ASAP7_75t_L g585 ( .A(n_484), .B(n_370), .C(n_382), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_464), .B(n_407), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_450), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_476), .Y(n_588) );
INVx2_ASAP7_75t_SL g589 ( .A(n_442), .Y(n_589) );
AND2x4_ASAP7_75t_L g590 ( .A(n_515), .B(n_425), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_478), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_454), .B(n_425), .Y(n_592) );
INVxp67_ASAP7_75t_L g593 ( .A(n_441), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_508), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_495), .B(n_421), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_495), .B(n_421), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_513), .Y(n_597) );
NOR2x1_ASAP7_75t_L g598 ( .A(n_515), .B(n_419), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_442), .B(n_401), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_469), .B(n_407), .Y(n_600) );
INVx1_ASAP7_75t_SL g601 ( .A(n_437), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_474), .B(n_424), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_437), .B(n_411), .Y(n_603) );
AND2x2_ASAP7_75t_SL g604 ( .A(n_518), .B(n_405), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_514), .B(n_421), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_437), .B(n_418), .Y(n_606) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_492), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_450), .Y(n_608) );
NAND2x1_ASAP7_75t_SL g609 ( .A(n_483), .B(n_418), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_453), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_453), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_443), .B(n_413), .Y(n_612) );
NOR2x1p5_ASAP7_75t_L g613 ( .A(n_483), .B(n_413), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_501), .B(n_415), .Y(n_614) );
NOR2xp67_ASAP7_75t_L g615 ( .A(n_481), .B(n_401), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_443), .B(n_411), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_457), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_443), .B(n_408), .Y(n_618) );
OR2x2_ASAP7_75t_L g619 ( .A(n_489), .B(n_384), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_457), .Y(n_620) );
INVx3_ASAP7_75t_L g621 ( .A(n_530), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_462), .Y(n_622) );
INVx3_ASAP7_75t_SL g623 ( .A(n_481), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_519), .B(n_408), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_531), .B(n_75), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_519), .B(n_382), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_519), .B(n_382), .Y(n_627) );
INVx2_ASAP7_75t_SL g628 ( .A(n_531), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_496), .B(n_382), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_462), .Y(n_630) );
INVx1_ASAP7_75t_SL g631 ( .A(n_554), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_535), .B(n_491), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_541), .Y(n_633) );
NOR2x1_ASAP7_75t_L g634 ( .A(n_538), .B(n_491), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_542), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_561), .Y(n_636) );
INVxp67_ASAP7_75t_L g637 ( .A(n_554), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_544), .B(n_480), .Y(n_638) );
OR2x2_ASAP7_75t_L g639 ( .A(n_619), .B(n_468), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_546), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_549), .Y(n_641) );
INVxp67_ASAP7_75t_L g642 ( .A(n_589), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_550), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_584), .B(n_528), .Y(n_644) );
NOR3xp33_ASAP7_75t_L g645 ( .A(n_540), .B(n_526), .C(n_522), .Y(n_645) );
INVx2_ASAP7_75t_SL g646 ( .A(n_623), .Y(n_646) );
NAND2x1_ASAP7_75t_L g647 ( .A(n_536), .B(n_526), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_607), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_563), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_588), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_591), .Y(n_651) );
NOR2x1_ASAP7_75t_L g652 ( .A(n_567), .B(n_331), .Y(n_652) );
INVxp67_ASAP7_75t_L g653 ( .A(n_543), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_555), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_545), .B(n_497), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_539), .Y(n_656) );
OR2x2_ASAP7_75t_L g657 ( .A(n_565), .B(n_472), .Y(n_657) );
INVx2_ASAP7_75t_SL g658 ( .A(n_628), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_548), .B(n_502), .Y(n_659) );
NOR3xp33_ASAP7_75t_L g660 ( .A(n_593), .B(n_521), .C(n_479), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_582), .A2(n_482), .B1(n_487), .B2(n_494), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_539), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_569), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_573), .Y(n_664) );
OR2x2_ASAP7_75t_L g665 ( .A(n_581), .B(n_472), .Y(n_665) );
AOI22xp33_ASAP7_75t_SL g666 ( .A1(n_604), .A2(n_460), .B1(n_530), .B2(n_509), .Y(n_666) );
AOI21xp5_ASAP7_75t_L g667 ( .A1(n_598), .A2(n_460), .B(n_509), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_578), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_553), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_553), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_560), .B(n_449), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_607), .Y(n_672) );
OAI21xp5_ASAP7_75t_L g673 ( .A1(n_615), .A2(n_533), .B(n_477), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_579), .Y(n_674) );
OAI22xp33_ASAP7_75t_L g675 ( .A1(n_621), .A2(n_530), .B1(n_447), .B2(n_468), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_602), .A2(n_504), .B1(n_502), .B2(n_517), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_558), .B(n_525), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_579), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_566), .B(n_502), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_537), .B(n_510), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_594), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_552), .B(n_510), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_545), .B(n_470), .Y(n_683) );
NAND2xp5_ASAP7_75t_SL g684 ( .A(n_551), .B(n_451), .Y(n_684) );
NAND2xp33_ASAP7_75t_SL g685 ( .A(n_609), .B(n_527), .Y(n_685) );
NAND2x1p5_ASAP7_75t_L g686 ( .A(n_613), .B(n_358), .Y(n_686) );
OR2x2_ASAP7_75t_L g687 ( .A(n_614), .B(n_576), .Y(n_687) );
OR2x2_ASAP7_75t_L g688 ( .A(n_614), .B(n_492), .Y(n_688) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_593), .Y(n_689) );
NAND2xp33_ASAP7_75t_R g690 ( .A(n_621), .B(n_510), .Y(n_690) );
OR2x2_ASAP7_75t_L g691 ( .A(n_576), .B(n_517), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_547), .B(n_511), .Y(n_692) );
AOI21xp33_ASAP7_75t_SL g693 ( .A1(n_551), .A2(n_331), .B(n_524), .Y(n_693) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_599), .Y(n_694) );
OAI21xp33_ASAP7_75t_L g695 ( .A1(n_631), .A2(n_547), .B(n_556), .Y(n_695) );
INVx1_ASAP7_75t_SL g696 ( .A(n_631), .Y(n_696) );
INVxp67_ASAP7_75t_L g697 ( .A(n_689), .Y(n_697) );
NAND2x1p5_ASAP7_75t_L g698 ( .A(n_647), .B(n_570), .Y(n_698) );
INVx2_ASAP7_75t_L g699 ( .A(n_688), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_680), .B(n_601), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_679), .B(n_601), .Y(n_701) );
NOR2x1p5_ASAP7_75t_L g702 ( .A(n_690), .B(n_655), .Y(n_702) );
OAI221xp5_ASAP7_75t_SL g703 ( .A1(n_645), .A2(n_575), .B1(n_577), .B2(n_583), .C(n_571), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_646), .B(n_570), .Y(n_704) );
INVxp67_ASAP7_75t_L g705 ( .A(n_658), .Y(n_705) );
NOR2x1_ASAP7_75t_L g706 ( .A(n_634), .B(n_585), .Y(n_706) );
OAI22xp33_ASAP7_75t_L g707 ( .A1(n_667), .A2(n_574), .B1(n_592), .B2(n_629), .Y(n_707) );
NAND2x1_ASAP7_75t_L g708 ( .A(n_648), .B(n_572), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_642), .B(n_559), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_669), .Y(n_710) );
OAI322xp33_ASAP7_75t_L g711 ( .A1(n_637), .A2(n_655), .A3(n_661), .B1(n_638), .B2(n_687), .C1(n_644), .C2(n_654), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_656), .B(n_557), .Y(n_712) );
INVx2_ASAP7_75t_SL g713 ( .A(n_632), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_682), .B(n_562), .Y(n_714) );
AOI32xp33_ASAP7_75t_L g715 ( .A1(n_685), .A2(n_580), .A3(n_624), .B1(n_625), .B2(n_590), .Y(n_715) );
AOI221xp5_ASAP7_75t_L g716 ( .A1(n_693), .A2(n_557), .B1(n_556), .B2(n_564), .C(n_574), .Y(n_716) );
INVx3_ASAP7_75t_L g717 ( .A(n_672), .Y(n_717) );
XNOR2x2_ASAP7_75t_L g718 ( .A(n_652), .B(n_592), .Y(n_718) );
AOI221xp5_ASAP7_75t_L g719 ( .A1(n_660), .A2(n_564), .B1(n_595), .B2(n_596), .C(n_568), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g720 ( .A1(n_666), .A2(n_572), .B1(n_590), .B2(n_596), .Y(n_720) );
OAI221xp5_ASAP7_75t_L g721 ( .A1(n_676), .A2(n_673), .B1(n_686), .B2(n_653), .C(n_684), .Y(n_721) );
NOR3xp33_ASAP7_75t_L g722 ( .A(n_674), .B(n_568), .C(n_595), .Y(n_722) );
OAI21xp5_ASAP7_75t_L g723 ( .A1(n_686), .A2(n_358), .B(n_597), .Y(n_723) );
AOI222xp33_ASAP7_75t_L g724 ( .A1(n_636), .A2(n_629), .B1(n_622), .B2(n_620), .C1(n_617), .C2(n_610), .Y(n_724) );
OAI221xp5_ASAP7_75t_L g725 ( .A1(n_673), .A2(n_627), .B1(n_626), .B2(n_605), .C(n_587), .Y(n_725) );
OAI221xp5_ASAP7_75t_L g726 ( .A1(n_662), .A2(n_605), .B1(n_630), .B2(n_608), .C(n_611), .Y(n_726) );
OAI22xp33_ASAP7_75t_L g727 ( .A1(n_675), .A2(n_618), .B1(n_616), .B2(n_612), .Y(n_727) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_694), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_659), .B(n_606), .Y(n_729) );
INVxp67_ASAP7_75t_L g730 ( .A(n_633), .Y(n_730) );
OAI22xp33_ASAP7_75t_L g731 ( .A1(n_721), .A2(n_639), .B1(n_665), .B2(n_657), .Y(n_731) );
AOI221xp5_ASAP7_75t_SL g732 ( .A1(n_711), .A2(n_678), .B1(n_650), .B2(n_651), .C(n_649), .Y(n_732) );
AO21x1_ASAP7_75t_L g733 ( .A1(n_707), .A2(n_640), .B(n_641), .Y(n_733) );
OAI22xp33_ASAP7_75t_L g734 ( .A1(n_720), .A2(n_691), .B1(n_671), .B2(n_683), .Y(n_734) );
AND2x4_ASAP7_75t_L g735 ( .A(n_702), .B(n_670), .Y(n_735) );
OAI21x1_ASAP7_75t_SL g736 ( .A1(n_718), .A2(n_643), .B(n_692), .Y(n_736) );
OAI322xp33_ASAP7_75t_L g737 ( .A1(n_697), .A2(n_677), .A3(n_635), .B1(n_681), .B2(n_663), .C1(n_668), .C2(n_664), .Y(n_737) );
OA21x2_ASAP7_75t_SL g738 ( .A1(n_696), .A2(n_692), .B(n_683), .Y(n_738) );
NOR4xp25_ASAP7_75t_L g739 ( .A(n_696), .B(n_500), .C(n_506), .D(n_523), .Y(n_739) );
INVx2_ASAP7_75t_L g740 ( .A(n_717), .Y(n_740) );
AOI222xp33_ASAP7_75t_L g741 ( .A1(n_719), .A2(n_534), .B1(n_603), .B2(n_517), .C1(n_586), .C2(n_506), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_728), .Y(n_742) );
BUFx3_ASAP7_75t_L g743 ( .A(n_704), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_710), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_724), .B(n_600), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_717), .Y(n_746) );
OAI221xp5_ASAP7_75t_L g747 ( .A1(n_715), .A2(n_500), .B1(n_516), .B2(n_511), .C(n_505), .Y(n_747) );
AOI211xp5_ASAP7_75t_L g748 ( .A1(n_716), .A2(n_523), .B(n_516), .C(n_505), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_712), .Y(n_749) );
NAND3xp33_ASAP7_75t_L g750 ( .A(n_724), .B(n_382), .C(n_370), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g751 ( .A1(n_727), .A2(n_331), .B1(n_470), .B2(n_370), .Y(n_751) );
NOR3xp33_ASAP7_75t_L g752 ( .A(n_703), .B(n_358), .C(n_331), .Y(n_752) );
AOI221xp5_ASAP7_75t_L g753 ( .A1(n_695), .A2(n_382), .B1(n_370), .B2(n_331), .C(n_335), .Y(n_753) );
AOI21xp33_ASAP7_75t_SL g754 ( .A1(n_698), .A2(n_335), .B(n_84), .Y(n_754) );
NOR4xp25_ASAP7_75t_L g755 ( .A(n_705), .B(n_335), .C(n_370), .D(n_88), .Y(n_755) );
AO21x1_ASAP7_75t_L g756 ( .A1(n_698), .A2(n_370), .B(n_87), .Y(n_756) );
OAI211xp5_ASAP7_75t_L g757 ( .A1(n_706), .A2(n_80), .B(n_90), .C(n_91), .Y(n_757) );
NAND4xp25_ASAP7_75t_SL g758 ( .A(n_725), .B(n_92), .C(n_722), .D(n_726), .Y(n_758) );
NAND2xp5_ASAP7_75t_SL g759 ( .A(n_723), .B(n_713), .Y(n_759) );
OAI211xp5_ASAP7_75t_SL g760 ( .A1(n_747), .A2(n_731), .B(n_759), .C(n_734), .Y(n_760) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_742), .Y(n_761) );
NOR2x1_ASAP7_75t_L g762 ( .A(n_758), .B(n_757), .Y(n_762) );
NOR4xp25_ASAP7_75t_L g763 ( .A(n_737), .B(n_750), .C(n_745), .D(n_738), .Y(n_763) );
OAI22xp5_ASAP7_75t_L g764 ( .A1(n_735), .A2(n_743), .B1(n_748), .B2(n_749), .Y(n_764) );
AOI211xp5_ASAP7_75t_L g765 ( .A1(n_763), .A2(n_733), .B(n_752), .C(n_732), .Y(n_765) );
NOR3x1_ASAP7_75t_L g766 ( .A(n_764), .B(n_736), .C(n_708), .Y(n_766) );
NOR2xp33_ASAP7_75t_R g767 ( .A(n_761), .B(n_735), .Y(n_767) );
NAND4xp75_ASAP7_75t_L g768 ( .A(n_766), .B(n_762), .C(n_732), .D(n_756), .Y(n_768) );
NAND3x1_ASAP7_75t_SL g769 ( .A(n_767), .B(n_760), .C(n_753), .Y(n_769) );
XNOR2xp5_ASAP7_75t_L g770 ( .A(n_769), .B(n_765), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_768), .B(n_744), .Y(n_771) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_770), .A2(n_751), .B1(n_746), .B2(n_740), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_771), .B(n_739), .Y(n_773) );
AO22x2_ASAP7_75t_L g774 ( .A1(n_773), .A2(n_730), .B1(n_699), .B2(n_723), .Y(n_774) );
OAI22xp33_ASAP7_75t_L g775 ( .A1(n_774), .A2(n_772), .B1(n_754), .B2(n_709), .Y(n_775) );
AOI21xp33_ASAP7_75t_L g776 ( .A1(n_775), .A2(n_741), .B(n_700), .Y(n_776) );
OAI22xp5_ASAP7_75t_L g777 ( .A1(n_776), .A2(n_701), .B1(n_729), .B2(n_714), .Y(n_777) );
AOI22xp5_ASAP7_75t_L g778 ( .A1(n_777), .A2(n_741), .B1(n_739), .B2(n_755), .Y(n_778) );
endmodule