module fake_netlist_6_108_n_1958 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1958);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1958;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_683;
wire n_811;
wire n_527;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1892;
wire n_1459;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1737;
wire n_236;
wire n_653;
wire n_1464;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_104),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_100),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_62),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_92),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_185),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_111),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_50),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_34),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_149),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_24),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_153),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_118),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_129),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_172),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_139),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_79),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_5),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_60),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_78),
.Y(n_209)
);

BUFx5_ASAP7_75t_L g210 ( 
.A(n_117),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_89),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_54),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_16),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_123),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_75),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_24),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_97),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_127),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_16),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_73),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_171),
.Y(n_221)
);

BUFx10_ASAP7_75t_L g222 ( 
.A(n_134),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_7),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_84),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_151),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_13),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_177),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_91),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_2),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_103),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_25),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_186),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_1),
.Y(n_233)
);

BUFx10_ASAP7_75t_L g234 ( 
.A(n_105),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_66),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_8),
.Y(n_236)
);

BUFx5_ASAP7_75t_L g237 ( 
.A(n_166),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_181),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_152),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_64),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_169),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_31),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_27),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_38),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_170),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_74),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_21),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_136),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_168),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_132),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_101),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_179),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_10),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_162),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_38),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_121),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_5),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_19),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_154),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_27),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_52),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_42),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_68),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_175),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_150),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_35),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_83),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_28),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_45),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_34),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_50),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_119),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_110),
.Y(n_273)
);

BUFx8_ASAP7_75t_SL g274 ( 
.A(n_64),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_190),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_109),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_20),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_93),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_183),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_10),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_14),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_143),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_88),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_39),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_87),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_19),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_81),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_128),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_145),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_141),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_58),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_106),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_90),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_140),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_189),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_57),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_21),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_126),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_114),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_60),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_77),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_54),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_57),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_130),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_11),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_94),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_8),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_14),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_35),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_70),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_36),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_116),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_56),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_86),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_3),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_98),
.Y(n_316)
);

BUFx5_ASAP7_75t_L g317 ( 
.A(n_51),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_44),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_187),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_11),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_49),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_47),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_48),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_17),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_20),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_156),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_28),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_137),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_107),
.Y(n_329)
);

BUFx10_ASAP7_75t_L g330 ( 
.A(n_182),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_9),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_30),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_115),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_71),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_184),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_164),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_147),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_85),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_133),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_142),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_158),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_138),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_96),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_176),
.Y(n_344)
);

BUFx10_ASAP7_75t_L g345 ( 
.A(n_161),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_0),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_45),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_157),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_46),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_58),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_135),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_40),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_49),
.Y(n_353)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_173),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_165),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_159),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_52),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_37),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_7),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_80),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_113),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_160),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_102),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_43),
.Y(n_364)
);

CKINVDCx14_ASAP7_75t_R g365 ( 
.A(n_23),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_67),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_48),
.Y(n_367)
);

INVx2_ASAP7_75t_SL g368 ( 
.A(n_40),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_26),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_59),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_31),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_6),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_23),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_22),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_112),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_120),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_39),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_33),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_99),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_32),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_155),
.Y(n_381)
);

INVx2_ASAP7_75t_SL g382 ( 
.A(n_62),
.Y(n_382)
);

BUFx10_ASAP7_75t_L g383 ( 
.A(n_53),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_4),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_42),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_174),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_66),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_12),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_317),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_317),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_317),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_317),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_224),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_224),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_317),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_225),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_317),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_317),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_225),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_240),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_245),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_274),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_258),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_258),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_240),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_274),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_240),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g408 ( 
.A(n_197),
.B(n_0),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_240),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_R g410 ( 
.A(n_365),
.B(n_188),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_318),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_245),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_318),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_318),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_318),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_347),
.Y(n_416)
);

NOR2xp67_ASAP7_75t_L g417 ( 
.A(n_368),
.B(n_1),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_285),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_347),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_347),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_347),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_372),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_285),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_309),
.Y(n_424)
);

INVxp67_ASAP7_75t_SL g425 ( 
.A(n_256),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_383),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_212),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_372),
.Y(n_428)
);

OR2x2_ASAP7_75t_L g429 ( 
.A(n_200),
.B(n_2),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_372),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_299),
.B(n_3),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_288),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_372),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_288),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_301),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_383),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_208),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_193),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_198),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_207),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_299),
.B(n_4),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_212),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_383),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_301),
.Y(n_444)
);

INVxp33_ASAP7_75t_SL g445 ( 
.A(n_216),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_213),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_223),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_219),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_328),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_328),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_226),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_222),
.Y(n_452)
);

INVxp67_ASAP7_75t_SL g453 ( 
.A(n_256),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_247),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_195),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_216),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_323),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_231),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_261),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_262),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_233),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_235),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_291),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_236),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_305),
.Y(n_465)
);

INVxp67_ASAP7_75t_SL g466 ( 
.A(n_306),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_242),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_311),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_204),
.B(n_6),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_320),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_196),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_321),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_327),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_300),
.Y(n_474)
);

CKINVDCx16_ASAP7_75t_R g475 ( 
.A(n_222),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_346),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_199),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_243),
.Y(n_478)
);

NOR2xp67_ASAP7_75t_L g479 ( 
.A(n_368),
.B(n_9),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_352),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_366),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_202),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_244),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_306),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_253),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_255),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_206),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_192),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_373),
.Y(n_489)
);

INVxp33_ASAP7_75t_L g490 ( 
.A(n_377),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_385),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_455),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_488),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_389),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_410),
.B(n_222),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_400),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_389),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_400),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_409),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_427),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_409),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_442),
.Y(n_502)
);

AND2x6_ASAP7_75t_L g503 ( 
.A(n_488),
.B(n_204),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_425),
.B(n_211),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_488),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_390),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_411),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_488),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_390),
.B(n_211),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_391),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_411),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_391),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_413),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_392),
.B(n_220),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_413),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_453),
.B(n_191),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_395),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_414),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_414),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_466),
.B(n_220),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_488),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_397),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_398),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_424),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_393),
.B(n_229),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_415),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_415),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_474),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_416),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_416),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_405),
.Y(n_531)
);

BUFx2_ASAP7_75t_L g532 ( 
.A(n_438),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_407),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_419),
.Y(n_534)
);

BUFx2_ASAP7_75t_L g535 ( 
.A(n_438),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_417),
.B(n_234),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_420),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_421),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_422),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_456),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_428),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_439),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_430),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_433),
.Y(n_544)
);

OAI21x1_ASAP7_75t_L g545 ( 
.A1(n_469),
.A2(n_294),
.B(n_273),
.Y(n_545)
);

CKINVDCx11_ASAP7_75t_R g546 ( 
.A(n_394),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_484),
.B(n_273),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_457),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_457),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_437),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_446),
.Y(n_551)
);

NAND2xp33_ASAP7_75t_SL g552 ( 
.A(n_431),
.B(n_229),
.Y(n_552)
);

CKINVDCx16_ASAP7_75t_R g553 ( 
.A(n_432),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_447),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_454),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_479),
.B(n_234),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_484),
.B(n_191),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_459),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_460),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_463),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_465),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_403),
.B(n_215),
.Y(n_562)
);

INVx1_ASAP7_75t_SL g563 ( 
.A(n_396),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_468),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_470),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_472),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_441),
.B(n_234),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_404),
.B(n_473),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_480),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_481),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_491),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_452),
.B(n_249),
.Y(n_572)
);

NAND2xp33_ASAP7_75t_SL g573 ( 
.A(n_408),
.B(n_270),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_568),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_568),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_500),
.B(n_439),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_516),
.B(n_445),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_568),
.Y(n_578)
);

AND2x6_ASAP7_75t_L g579 ( 
.A(n_504),
.B(n_294),
.Y(n_579)
);

BUFx2_ASAP7_75t_L g580 ( 
.A(n_532),
.Y(n_580)
);

NAND2xp33_ASAP7_75t_L g581 ( 
.A(n_516),
.B(n_440),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_500),
.B(n_440),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_557),
.B(n_445),
.Y(n_583)
);

NAND2xp33_ASAP7_75t_L g584 ( 
.A(n_567),
.B(n_448),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_SL g585 ( 
.A(n_492),
.B(n_402),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_505),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_502),
.B(n_448),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_505),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_547),
.B(n_476),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_567),
.A2(n_477),
.B1(n_482),
.B2(n_471),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_SL g591 ( 
.A(n_492),
.B(n_406),
.Y(n_591)
);

INVxp67_ASAP7_75t_L g592 ( 
.A(n_540),
.Y(n_592)
);

NAND2xp33_ASAP7_75t_L g593 ( 
.A(n_562),
.B(n_451),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_550),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_494),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_504),
.B(n_458),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_505),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_514),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_532),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_528),
.B(n_458),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_550),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_528),
.B(n_461),
.Y(n_602)
);

OAI22xp33_ASAP7_75t_SL g603 ( 
.A1(n_536),
.A2(n_475),
.B1(n_429),
.B2(n_408),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_505),
.Y(n_604)
);

AND2x6_ASAP7_75t_L g605 ( 
.A(n_504),
.B(n_520),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_540),
.B(n_435),
.Y(n_606)
);

INVx5_ASAP7_75t_L g607 ( 
.A(n_503),
.Y(n_607)
);

INVx8_ASAP7_75t_L g608 ( 
.A(n_520),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_554),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_562),
.B(n_461),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_554),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_520),
.B(n_462),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_547),
.B(n_462),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_559),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_495),
.B(n_464),
.Y(n_615)
);

OAI22xp33_ASAP7_75t_L g616 ( 
.A1(n_572),
.A2(n_429),
.B1(n_284),
.B2(n_332),
.Y(n_616)
);

INVx4_ASAP7_75t_L g617 ( 
.A(n_509),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_509),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_509),
.B(n_379),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_546),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_494),
.Y(n_621)
);

AND2x4_ASAP7_75t_L g622 ( 
.A(n_547),
.B(n_489),
.Y(n_622)
);

NAND3xp33_ASAP7_75t_L g623 ( 
.A(n_573),
.B(n_467),
.C(n_464),
.Y(n_623)
);

NAND2xp33_ASAP7_75t_L g624 ( 
.A(n_495),
.B(n_467),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_493),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_509),
.Y(n_626)
);

INVxp67_ASAP7_75t_SL g627 ( 
.A(n_506),
.Y(n_627)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_546),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_509),
.B(n_379),
.Y(n_629)
);

BUFx10_ASAP7_75t_L g630 ( 
.A(n_524),
.Y(n_630)
);

INVx4_ASAP7_75t_L g631 ( 
.A(n_514),
.Y(n_631)
);

INVx2_ASAP7_75t_SL g632 ( 
.A(n_524),
.Y(n_632)
);

INVxp67_ASAP7_75t_L g633 ( 
.A(n_573),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_493),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_536),
.B(n_478),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_553),
.Y(n_636)
);

NOR3xp33_ASAP7_75t_L g637 ( 
.A(n_552),
.B(n_456),
.C(n_436),
.Y(n_637)
);

INVx4_ASAP7_75t_L g638 ( 
.A(n_514),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_559),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_561),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_506),
.B(n_510),
.Y(n_641)
);

INVx5_ASAP7_75t_L g642 ( 
.A(n_503),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_561),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_506),
.B(n_478),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_570),
.Y(n_645)
);

AND2x4_ASAP7_75t_L g646 ( 
.A(n_570),
.B(n_382),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_517),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_517),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_530),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_494),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_514),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_532),
.B(n_483),
.Y(n_652)
);

INVx4_ASAP7_75t_L g653 ( 
.A(n_514),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_506),
.B(n_483),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_556),
.B(n_382),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_514),
.B(n_192),
.Y(n_656)
);

AND2x6_ASAP7_75t_L g657 ( 
.A(n_510),
.B(n_192),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_530),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_556),
.B(n_485),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_553),
.Y(n_660)
);

OAI22xp33_ASAP7_75t_L g661 ( 
.A1(n_572),
.A2(n_284),
.B1(n_332),
.B2(n_270),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_517),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_517),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_535),
.B(n_485),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_510),
.B(n_486),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_530),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_510),
.B(n_486),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_530),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_552),
.A2(n_370),
.B1(n_371),
.B2(n_323),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_512),
.B(n_354),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_522),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_512),
.B(n_522),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_522),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_530),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_493),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_522),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_563),
.Y(n_677)
);

BUFx4f_ASAP7_75t_L g678 ( 
.A(n_535),
.Y(n_678)
);

HB1xp67_ASAP7_75t_L g679 ( 
.A(n_564),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_564),
.B(n_487),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_523),
.Y(n_681)
);

CKINVDCx20_ASAP7_75t_R g682 ( 
.A(n_563),
.Y(n_682)
);

NAND2x1p5_ASAP7_75t_L g683 ( 
.A(n_545),
.B(n_194),
.Y(n_683)
);

AO22x2_ASAP7_75t_L g684 ( 
.A1(n_512),
.A2(n_371),
.B1(n_370),
.B2(n_363),
.Y(n_684)
);

BUFx4f_ASAP7_75t_L g685 ( 
.A(n_535),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_564),
.B(n_192),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_530),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_534),
.B(n_337),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_523),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_523),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_564),
.B(n_228),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_564),
.Y(n_692)
);

NAND2xp33_ASAP7_75t_L g693 ( 
.A(n_503),
.B(n_203),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_496),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_497),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_508),
.B(n_230),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_496),
.B(n_498),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_508),
.B(n_239),
.Y(n_698)
);

INVx4_ASAP7_75t_L g699 ( 
.A(n_538),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_498),
.Y(n_700)
);

OR2x6_ASAP7_75t_L g701 ( 
.A(n_542),
.B(n_426),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_508),
.B(n_241),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_551),
.B(n_203),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_525),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_499),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_508),
.B(n_246),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_542),
.B(n_443),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_545),
.A2(n_298),
.B1(n_267),
.B2(n_263),
.Y(n_708)
);

INVx4_ASAP7_75t_L g709 ( 
.A(n_538),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_521),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_521),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_499),
.Y(n_712)
);

NOR2x1p5_ASAP7_75t_L g713 ( 
.A(n_548),
.B(n_406),
.Y(n_713)
);

BUFx2_ASAP7_75t_L g714 ( 
.A(n_682),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_679),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_679),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_598),
.Y(n_717)
);

INVx2_ASAP7_75t_SL g718 ( 
.A(n_630),
.Y(n_718)
);

NAND2x1p5_ASAP7_75t_L g719 ( 
.A(n_678),
.B(n_542),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_594),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_601),
.Y(n_721)
);

OAI221xp5_ASAP7_75t_L g722 ( 
.A1(n_669),
.A2(n_254),
.B1(n_569),
.B2(n_566),
.C(n_565),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_609),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_611),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_630),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_605),
.B(n_497),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_605),
.B(n_497),
.Y(n_727)
);

NAND2x1p5_ASAP7_75t_L g728 ( 
.A(n_678),
.B(n_548),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_614),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_577),
.A2(n_583),
.B1(n_605),
.B2(n_610),
.Y(n_730)
);

OAI221xp5_ASAP7_75t_L g731 ( 
.A1(n_669),
.A2(n_577),
.B1(n_578),
.B2(n_575),
.C(n_574),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_639),
.Y(n_732)
);

CKINVDCx16_ASAP7_75t_R g733 ( 
.A(n_660),
.Y(n_733)
);

CKINVDCx20_ASAP7_75t_R g734 ( 
.A(n_628),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_640),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_583),
.B(n_399),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_643),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_610),
.B(n_401),
.Y(n_738)
);

AND2x4_ASAP7_75t_L g739 ( 
.A(n_645),
.B(n_589),
.Y(n_739)
);

AND2x4_ASAP7_75t_L g740 ( 
.A(n_589),
.B(n_551),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_598),
.Y(n_741)
);

AO22x2_ASAP7_75t_L g742 ( 
.A1(n_633),
.A2(n_205),
.B1(n_209),
.B2(n_201),
.Y(n_742)
);

AO22x2_ASAP7_75t_L g743 ( 
.A1(n_633),
.A2(n_221),
.B1(n_227),
.B2(n_214),
.Y(n_743)
);

BUFx6f_ASAP7_75t_SL g744 ( 
.A(n_632),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_652),
.B(n_664),
.Y(n_745)
);

AO22x2_ASAP7_75t_L g746 ( 
.A1(n_637),
.A2(n_238),
.B1(n_251),
.B2(n_232),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_600),
.B(n_615),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_622),
.B(n_571),
.Y(n_748)
);

NOR2xp67_ASAP7_75t_L g749 ( 
.A(n_615),
.B(n_534),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_622),
.B(n_551),
.Y(n_750)
);

BUFx8_ASAP7_75t_L g751 ( 
.A(n_580),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_651),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_694),
.Y(n_753)
);

OAI221xp5_ASAP7_75t_L g754 ( 
.A1(n_596),
.A2(n_571),
.B1(n_569),
.B2(n_566),
.C(n_565),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_605),
.A2(n_635),
.B1(n_659),
.B2(n_581),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_700),
.Y(n_756)
);

AND2x4_ASAP7_75t_L g757 ( 
.A(n_646),
.B(n_551),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_705),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_712),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_605),
.Y(n_760)
);

AO22x2_ASAP7_75t_L g761 ( 
.A1(n_637),
.A2(n_287),
.B1(n_290),
.B2(n_292),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_692),
.Y(n_762)
);

OAI221xp5_ASAP7_75t_L g763 ( 
.A1(n_612),
.A2(n_571),
.B1(n_569),
.B2(n_566),
.C(n_565),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_608),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_646),
.B(n_555),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_608),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_689),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_608),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_R g769 ( 
.A(n_636),
.B(n_412),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_697),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_697),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_713),
.B(n_571),
.Y(n_772)
);

INVx3_ASAP7_75t_L g773 ( 
.A(n_710),
.Y(n_773)
);

AO22x2_ASAP7_75t_L g774 ( 
.A1(n_590),
.A2(n_275),
.B1(n_276),
.B2(n_304),
.Y(n_774)
);

OAI221xp5_ASAP7_75t_L g775 ( 
.A1(n_613),
.A2(n_569),
.B1(n_566),
.B2(n_565),
.C(n_560),
.Y(n_775)
);

OAI221xp5_ASAP7_75t_L g776 ( 
.A1(n_644),
.A2(n_667),
.B1(n_665),
.B2(n_654),
.C(n_635),
.Y(n_776)
);

AO22x2_ASAP7_75t_L g777 ( 
.A1(n_616),
.A2(n_312),
.B1(n_259),
.B2(n_334),
.Y(n_777)
);

OAI22xp33_ASAP7_75t_SL g778 ( 
.A1(n_659),
.A2(n_655),
.B1(n_685),
.B2(n_680),
.Y(n_778)
);

A2O1A1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_655),
.A2(n_545),
.B(n_386),
.C(n_342),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_627),
.Y(n_780)
);

INVxp33_ASAP7_75t_SL g781 ( 
.A(n_585),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_627),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_677),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_680),
.B(n_215),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_618),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_618),
.Y(n_786)
);

AO22x2_ASAP7_75t_L g787 ( 
.A1(n_616),
.A2(n_339),
.B1(n_343),
.B2(n_360),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_576),
.B(n_490),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_710),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_592),
.Y(n_790)
);

AO22x2_ASAP7_75t_L g791 ( 
.A1(n_661),
.A2(n_381),
.B1(n_525),
.B2(n_374),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_688),
.B(n_555),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_579),
.B(n_497),
.Y(n_793)
);

INVxp67_ASAP7_75t_L g794 ( 
.A(n_707),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_688),
.B(n_560),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_618),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_579),
.B(n_526),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_618),
.Y(n_798)
);

AO22x2_ASAP7_75t_L g799 ( 
.A1(n_661),
.A2(n_525),
.B1(n_374),
.B2(n_384),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_595),
.Y(n_800)
);

NAND2x1p5_ASAP7_75t_L g801 ( 
.A(n_685),
.B(n_555),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_626),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_626),
.Y(n_803)
);

INVx8_ASAP7_75t_L g804 ( 
.A(n_701),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_592),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_626),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_626),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_579),
.B(n_526),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_711),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_711),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_603),
.B(n_217),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_684),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_579),
.A2(n_210),
.B1(n_237),
.B2(n_362),
.Y(n_813)
);

INVxp33_ASAP7_75t_SL g814 ( 
.A(n_591),
.Y(n_814)
);

OAI221xp5_ASAP7_75t_L g815 ( 
.A1(n_593),
.A2(n_560),
.B1(n_558),
.B2(n_555),
.C(n_544),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_684),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_621),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_620),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_650),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_597),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_579),
.A2(n_584),
.B1(n_624),
.B2(n_587),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_670),
.B(n_526),
.Y(n_822)
);

AND2x4_ASAP7_75t_L g823 ( 
.A(n_631),
.B(n_558),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_684),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_625),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_625),
.Y(n_826)
);

OAI221xp5_ASAP7_75t_L g827 ( 
.A1(n_708),
.A2(n_558),
.B1(n_544),
.B2(n_543),
.C(n_541),
.Y(n_827)
);

AO22x2_ASAP7_75t_L g828 ( 
.A1(n_623),
.A2(n_582),
.B1(n_602),
.B2(n_606),
.Y(n_828)
);

OR2x6_ASAP7_75t_L g829 ( 
.A(n_701),
.B(n_418),
.Y(n_829)
);

AO22x2_ASAP7_75t_L g830 ( 
.A1(n_619),
.A2(n_384),
.B1(n_423),
.B2(n_434),
.Y(n_830)
);

AO22x2_ASAP7_75t_L g831 ( 
.A1(n_619),
.A2(n_444),
.B1(n_449),
.B2(n_450),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_634),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_675),
.Y(n_833)
);

AO22x2_ASAP7_75t_L g834 ( 
.A1(n_629),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_834)
);

INVxp67_ASAP7_75t_L g835 ( 
.A(n_599),
.Y(n_835)
);

NAND2x1p5_ASAP7_75t_L g836 ( 
.A(n_617),
.B(n_537),
.Y(n_836)
);

BUFx3_ASAP7_75t_L g837 ( 
.A(n_701),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_631),
.B(n_537),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_638),
.B(n_539),
.Y(n_839)
);

BUFx8_ASAP7_75t_L g840 ( 
.A(n_704),
.Y(n_840)
);

HB1xp67_ASAP7_75t_L g841 ( 
.A(n_683),
.Y(n_841)
);

NOR2xp67_ASAP7_75t_L g842 ( 
.A(n_691),
.B(n_539),
.Y(n_842)
);

AO22x2_ASAP7_75t_L g843 ( 
.A1(n_629),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_843)
);

AO22x2_ASAP7_75t_L g844 ( 
.A1(n_656),
.A2(n_18),
.B1(n_22),
.B2(n_25),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_696),
.Y(n_845)
);

BUFx2_ASAP7_75t_L g846 ( 
.A(n_683),
.Y(n_846)
);

OAI221xp5_ASAP7_75t_L g847 ( 
.A1(n_708),
.A2(n_541),
.B1(n_543),
.B2(n_286),
.C(n_313),
.Y(n_847)
);

AOI22xp5_ASAP7_75t_SL g848 ( 
.A1(n_657),
.A2(n_300),
.B1(n_315),
.B2(n_387),
.Y(n_848)
);

AO22x2_ASAP7_75t_L g849 ( 
.A1(n_656),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_L g850 ( 
.A1(n_617),
.A2(n_653),
.B1(n_638),
.B2(n_702),
.Y(n_850)
);

AO22x2_ASAP7_75t_L g851 ( 
.A1(n_686),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_851)
);

AO22x2_ASAP7_75t_L g852 ( 
.A1(n_686),
.A2(n_36),
.B1(n_37),
.B2(n_41),
.Y(n_852)
);

INVx4_ASAP7_75t_L g853 ( 
.A(n_653),
.Y(n_853)
);

AO22x2_ASAP7_75t_L g854 ( 
.A1(n_703),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_854)
);

INVxp67_ASAP7_75t_L g855 ( 
.A(n_698),
.Y(n_855)
);

OAI221xp5_ASAP7_75t_L g856 ( 
.A1(n_672),
.A2(n_296),
.B1(n_325),
.B2(n_257),
.C(n_260),
.Y(n_856)
);

AO22x2_ASAP7_75t_L g857 ( 
.A1(n_703),
.A2(n_46),
.B1(n_47),
.B2(n_51),
.Y(n_857)
);

INVxp67_ASAP7_75t_L g858 ( 
.A(n_706),
.Y(n_858)
);

AO22x2_ASAP7_75t_L g859 ( 
.A1(n_586),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_747),
.B(n_588),
.Y(n_860)
);

NAND2xp33_ASAP7_75t_SL g861 ( 
.A(n_760),
.B(n_203),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_730),
.B(n_778),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_788),
.B(n_315),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_770),
.B(n_588),
.Y(n_864)
);

NAND2xp33_ASAP7_75t_SL g865 ( 
.A(n_745),
.B(n_217),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_755),
.B(n_597),
.Y(n_866)
);

NAND2xp33_ASAP7_75t_SL g867 ( 
.A(n_845),
.B(n_771),
.Y(n_867)
);

NAND2xp33_ASAP7_75t_SL g868 ( 
.A(n_841),
.B(n_218),
.Y(n_868)
);

NAND2xp33_ASAP7_75t_SL g869 ( 
.A(n_846),
.B(n_218),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_780),
.B(n_604),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_749),
.B(n_316),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_782),
.B(n_641),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_736),
.B(n_738),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_717),
.B(n_316),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_717),
.B(n_248),
.Y(n_875)
);

NAND2xp33_ASAP7_75t_SL g876 ( 
.A(n_744),
.B(n_387),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_717),
.B(n_250),
.Y(n_877)
);

NAND2xp33_ASAP7_75t_SL g878 ( 
.A(n_744),
.B(n_388),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_794),
.B(n_388),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_855),
.B(n_647),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_858),
.B(n_648),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_740),
.B(n_252),
.Y(n_882)
);

NAND2xp33_ASAP7_75t_SL g883 ( 
.A(n_769),
.B(n_264),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_740),
.B(n_272),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_748),
.B(n_750),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_748),
.B(n_750),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_739),
.B(n_278),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_739),
.B(n_279),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_821),
.B(n_282),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_776),
.B(n_266),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_792),
.B(n_289),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_792),
.B(n_293),
.Y(n_892)
);

NAND2xp33_ASAP7_75t_SL g893 ( 
.A(n_783),
.B(n_295),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_795),
.B(n_310),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_715),
.B(n_662),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_795),
.B(n_314),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_715),
.B(n_663),
.Y(n_897)
);

NAND2xp33_ASAP7_75t_SL g898 ( 
.A(n_784),
.B(n_319),
.Y(n_898)
);

NAND2xp33_ASAP7_75t_SL g899 ( 
.A(n_764),
.B(n_766),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_757),
.B(n_765),
.Y(n_900)
);

NAND2xp33_ASAP7_75t_SL g901 ( 
.A(n_812),
.B(n_326),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_757),
.B(n_329),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_765),
.B(n_333),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_716),
.B(n_335),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_716),
.B(n_336),
.Y(n_905)
);

NAND2xp33_ASAP7_75t_SL g906 ( 
.A(n_768),
.B(n_338),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_781),
.B(n_340),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_814),
.B(n_341),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_823),
.B(n_344),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_753),
.B(n_671),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_756),
.B(n_673),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_790),
.B(n_805),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_758),
.B(n_759),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_728),
.B(n_348),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_719),
.B(n_351),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_822),
.B(n_676),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_720),
.B(n_681),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_772),
.B(n_355),
.Y(n_918)
);

NAND2xp33_ASAP7_75t_SL g919 ( 
.A(n_718),
.B(n_356),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_772),
.B(n_361),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_721),
.B(n_723),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_724),
.B(n_690),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_853),
.B(n_838),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_729),
.B(n_695),
.Y(n_924)
);

NAND2xp33_ASAP7_75t_SL g925 ( 
.A(n_816),
.B(n_375),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_732),
.B(n_695),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_853),
.B(n_376),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_838),
.B(n_839),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_839),
.B(n_607),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_801),
.B(n_607),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_735),
.B(n_607),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_737),
.B(n_642),
.Y(n_932)
);

NAND2xp33_ASAP7_75t_SL g933 ( 
.A(n_824),
.B(n_649),
.Y(n_933)
);

NAND2xp33_ASAP7_75t_SL g934 ( 
.A(n_725),
.B(n_649),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_835),
.B(n_642),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_741),
.B(n_642),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_752),
.B(n_249),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_785),
.B(n_249),
.Y(n_938)
);

NAND2xp33_ASAP7_75t_SL g939 ( 
.A(n_797),
.B(n_808),
.Y(n_939)
);

NAND2xp33_ASAP7_75t_SL g940 ( 
.A(n_811),
.B(n_268),
.Y(n_940)
);

NAND2xp33_ASAP7_75t_R g941 ( 
.A(n_714),
.B(n_269),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_731),
.B(n_271),
.Y(n_942)
);

NAND2xp33_ASAP7_75t_SL g943 ( 
.A(n_726),
.B(n_649),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_786),
.B(n_265),
.Y(n_944)
);

AND2x4_ASAP7_75t_L g945 ( 
.A(n_809),
.B(n_531),
.Y(n_945)
);

NAND2xp33_ASAP7_75t_SL g946 ( 
.A(n_727),
.B(n_658),
.Y(n_946)
);

NAND2xp33_ASAP7_75t_SL g947 ( 
.A(n_813),
.B(n_658),
.Y(n_947)
);

NAND2xp33_ASAP7_75t_SL g948 ( 
.A(n_793),
.B(n_658),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_796),
.B(n_265),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_798),
.B(n_265),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_802),
.B(n_283),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_803),
.B(n_283),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_806),
.B(n_283),
.Y(n_953)
);

NAND2xp33_ASAP7_75t_SL g954 ( 
.A(n_762),
.B(n_658),
.Y(n_954)
);

OR2x2_ASAP7_75t_L g955 ( 
.A(n_733),
.B(n_829),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_807),
.B(n_330),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_842),
.B(n_330),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_820),
.B(n_330),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_820),
.B(n_345),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_810),
.B(n_531),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_767),
.B(n_666),
.Y(n_961)
);

NAND2xp33_ASAP7_75t_SL g962 ( 
.A(n_825),
.B(n_666),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_820),
.B(n_345),
.Y(n_963)
);

NAND2xp33_ASAP7_75t_SL g964 ( 
.A(n_826),
.B(n_666),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_773),
.B(n_345),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_828),
.B(n_277),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_773),
.B(n_789),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_850),
.B(n_668),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_848),
.B(n_668),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_836),
.B(n_674),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_837),
.B(n_674),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_832),
.B(n_833),
.Y(n_972)
);

NAND2xp33_ASAP7_75t_SL g973 ( 
.A(n_818),
.B(n_280),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_817),
.B(n_687),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_779),
.B(n_531),
.Y(n_975)
);

NAND2xp33_ASAP7_75t_SL g976 ( 
.A(n_734),
.B(n_281),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_819),
.B(n_501),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_804),
.B(n_210),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_804),
.B(n_210),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_751),
.B(n_210),
.Y(n_980)
);

NAND2xp33_ASAP7_75t_SL g981 ( 
.A(n_777),
.B(n_297),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_751),
.B(n_210),
.Y(n_982)
);

NAND2xp33_ASAP7_75t_SL g983 ( 
.A(n_777),
.B(n_302),
.Y(n_983)
);

NAND2xp33_ASAP7_75t_SL g984 ( 
.A(n_787),
.B(n_303),
.Y(n_984)
);

NAND2xp33_ASAP7_75t_SL g985 ( 
.A(n_787),
.B(n_307),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_800),
.B(n_237),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_828),
.B(n_308),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_742),
.B(n_743),
.Y(n_988)
);

NAND2xp33_ASAP7_75t_SL g989 ( 
.A(n_774),
.B(n_322),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_742),
.B(n_743),
.Y(n_990)
);

NAND2xp33_ASAP7_75t_SL g991 ( 
.A(n_774),
.B(n_324),
.Y(n_991)
);

NAND2xp33_ASAP7_75t_SL g992 ( 
.A(n_831),
.B(n_331),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_840),
.B(n_237),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_840),
.B(n_237),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_831),
.B(n_511),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_830),
.B(n_501),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_830),
.B(n_513),
.Y(n_997)
);

NAND2xp33_ASAP7_75t_SL g998 ( 
.A(n_791),
.B(n_349),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_856),
.B(n_513),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_746),
.B(n_709),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_746),
.B(n_709),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_761),
.B(n_699),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_761),
.B(n_511),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_754),
.B(n_699),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_847),
.B(n_529),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_791),
.B(n_507),
.Y(n_1006)
);

NAND2xp33_ASAP7_75t_SL g1007 ( 
.A(n_834),
.B(n_350),
.Y(n_1007)
);

NAND2xp33_ASAP7_75t_SL g1008 ( 
.A(n_834),
.B(n_353),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_843),
.B(n_527),
.Y(n_1009)
);

NAND2xp33_ASAP7_75t_SL g1010 ( 
.A(n_843),
.B(n_357),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_859),
.B(n_507),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_859),
.B(n_527),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_844),
.B(n_519),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_844),
.B(n_519),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_849),
.B(n_518),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_849),
.B(n_518),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_851),
.B(n_515),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_851),
.B(n_515),
.Y(n_1018)
);

NAND2xp33_ASAP7_75t_SL g1019 ( 
.A(n_852),
.B(n_358),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_799),
.B(n_829),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_852),
.B(n_529),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_L g1022 ( 
.A1(n_974),
.A2(n_533),
.B(n_521),
.Y(n_1022)
);

INVx3_ASAP7_75t_L g1023 ( 
.A(n_977),
.Y(n_1023)
);

OAI21xp33_ASAP7_75t_L g1024 ( 
.A1(n_873),
.A2(n_799),
.B(n_364),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_977),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_945),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_924),
.Y(n_1027)
);

HB1xp67_ASAP7_75t_L g1028 ( 
.A(n_912),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_945),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_863),
.B(n_879),
.Y(n_1030)
);

NOR4xp25_ASAP7_75t_L g1031 ( 
.A(n_890),
.B(n_763),
.C(n_775),
.D(n_815),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_860),
.B(n_857),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_867),
.B(n_722),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_866),
.A2(n_827),
.B(n_693),
.Y(n_1034)
);

AO21x2_ASAP7_75t_L g1035 ( 
.A1(n_862),
.A2(n_857),
.B(n_854),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_880),
.B(n_854),
.Y(n_1036)
);

AOI21xp33_ASAP7_75t_L g1037 ( 
.A1(n_942),
.A2(n_359),
.B(n_367),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_867),
.B(n_928),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_926),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_966),
.B(n_369),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_910),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_945),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_1007),
.A2(n_378),
.B(n_380),
.C(n_533),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_913),
.B(n_549),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_960),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_885),
.B(n_886),
.Y(n_1046)
);

CKINVDCx11_ASAP7_75t_R g1047 ( 
.A(n_976),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_921),
.B(n_549),
.Y(n_1048)
);

INVxp67_ASAP7_75t_L g1049 ( 
.A(n_1003),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_911),
.Y(n_1050)
);

AO21x2_ASAP7_75t_L g1051 ( 
.A1(n_968),
.A2(n_657),
.B(n_503),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_939),
.A2(n_549),
.B(n_538),
.Y(n_1052)
);

OAI21xp33_ASAP7_75t_SL g1053 ( 
.A1(n_923),
.A2(n_55),
.B(n_59),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_960),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_881),
.B(n_549),
.Y(n_1055)
);

AO32x2_ASAP7_75t_L g1056 ( 
.A1(n_1007),
.A2(n_61),
.A3(n_63),
.B1(n_65),
.B2(n_67),
.Y(n_1056)
);

NOR2x1_ASAP7_75t_SL g1057 ( 
.A(n_967),
.B(n_549),
.Y(n_1057)
);

NOR2xp67_ASAP7_75t_SL g1058 ( 
.A(n_900),
.B(n_549),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_864),
.B(n_549),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_916),
.B(n_872),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_1006),
.B(n_61),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_917),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_895),
.B(n_549),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_922),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_SL g1065 ( 
.A1(n_1011),
.A2(n_63),
.B(n_65),
.C(n_69),
.Y(n_1065)
);

NAND3x1_ASAP7_75t_L g1066 ( 
.A(n_1020),
.B(n_72),
.C(n_76),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_897),
.B(n_538),
.Y(n_1067)
);

AO21x2_ASAP7_75t_L g1068 ( 
.A1(n_889),
.A2(n_503),
.B(n_538),
.Y(n_1068)
);

AND2x4_ASAP7_75t_L g1069 ( 
.A(n_960),
.B(n_82),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_947),
.A2(n_95),
.B(n_108),
.Y(n_1070)
);

OA21x2_ASAP7_75t_L g1071 ( 
.A1(n_1004),
.A2(n_1012),
.B(n_1001),
.Y(n_1071)
);

AOI221x1_ASAP7_75t_L g1072 ( 
.A1(n_1008),
.A2(n_122),
.B1(n_124),
.B2(n_125),
.C(n_131),
.Y(n_1072)
);

OA21x2_ASAP7_75t_L g1073 ( 
.A1(n_1000),
.A2(n_144),
.B(n_146),
.Y(n_1073)
);

INVxp67_ASAP7_75t_SL g1074 ( 
.A(n_870),
.Y(n_1074)
);

HB1xp67_ASAP7_75t_L g1075 ( 
.A(n_988),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_1002),
.B(n_148),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_972),
.Y(n_1077)
);

INVxp67_ASAP7_75t_L g1078 ( 
.A(n_1009),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_961),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_975),
.Y(n_1080)
);

NAND2xp33_ASAP7_75t_L g1081 ( 
.A(n_934),
.B(n_163),
.Y(n_1081)
);

BUFx2_ASAP7_75t_L g1082 ( 
.A(n_955),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_943),
.B(n_167),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_975),
.Y(n_1084)
);

NOR3xp33_ASAP7_75t_L g1085 ( 
.A(n_992),
.B(n_178),
.C(n_180),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_943),
.B(n_946),
.Y(n_1086)
);

OAI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_1005),
.A2(n_946),
.B(n_948),
.Y(n_1087)
);

OAI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_948),
.A2(n_929),
.B(n_1013),
.Y(n_1088)
);

NOR2xp67_ASAP7_75t_L g1089 ( 
.A(n_957),
.B(n_915),
.Y(n_1089)
);

NAND2xp33_ASAP7_75t_SL g1090 ( 
.A(n_990),
.B(n_1017),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_933),
.B(n_1008),
.Y(n_1091)
);

BUFx3_ASAP7_75t_L g1092 ( 
.A(n_987),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_996),
.B(n_997),
.Y(n_1093)
);

NAND2x1p5_ASAP7_75t_L g1094 ( 
.A(n_970),
.B(n_930),
.Y(n_1094)
);

AND2x4_ASAP7_75t_L g1095 ( 
.A(n_971),
.B(n_887),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1018),
.B(n_1021),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1014),
.B(n_1015),
.Y(n_1097)
);

NAND3x1_ASAP7_75t_L g1098 ( 
.A(n_1019),
.B(n_1010),
.C(n_998),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1016),
.B(n_871),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_899),
.Y(n_1100)
);

AO31x2_ASAP7_75t_L g1101 ( 
.A1(n_1010),
.A2(n_1019),
.A3(n_933),
.B(n_995),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_907),
.B(n_908),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_986),
.Y(n_1103)
);

OAI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_969),
.A2(n_999),
.B(n_936),
.Y(n_1104)
);

INVx5_ASAP7_75t_L g1105 ( 
.A(n_954),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_904),
.B(n_905),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_874),
.B(n_958),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_931),
.A2(n_932),
.B(n_935),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_875),
.A2(n_877),
.B(n_978),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_SL g1110 ( 
.A1(n_914),
.A2(n_927),
.B(n_909),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_901),
.A2(n_925),
.B(n_981),
.C(n_984),
.Y(n_1111)
);

NOR2xp67_ASAP7_75t_L g1112 ( 
.A(n_959),
.B(n_963),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_L g1113 ( 
.A1(n_979),
.A2(n_896),
.B(n_894),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_918),
.B(n_920),
.Y(n_1114)
);

OA22x2_ASAP7_75t_L g1115 ( 
.A1(n_993),
.A2(n_994),
.B1(n_937),
.B2(n_980),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_901),
.B(n_925),
.Y(n_1116)
);

AO31x2_ASAP7_75t_L g1117 ( 
.A1(n_962),
.A2(n_964),
.A3(n_861),
.B(n_985),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_983),
.A2(n_991),
.B(n_989),
.C(n_868),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_891),
.A2(n_892),
.B(n_903),
.Y(n_1119)
);

OAI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_882),
.A2(n_884),
.B(n_902),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_868),
.A2(n_865),
.B(n_940),
.C(n_869),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_888),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_965),
.Y(n_1123)
);

AOI211x1_ASAP7_75t_L g1124 ( 
.A1(n_938),
.A2(n_952),
.B(n_949),
.C(n_950),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_944),
.A2(n_956),
.B(n_953),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_865),
.B(n_951),
.Y(n_1126)
);

AO31x2_ASAP7_75t_L g1127 ( 
.A1(n_962),
.A2(n_861),
.A3(n_934),
.B(n_898),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_982),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_869),
.B(n_893),
.Y(n_1129)
);

AOI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_883),
.A2(n_906),
.B1(n_941),
.B2(n_973),
.Y(n_1130)
);

O2A1O1Ixp5_ASAP7_75t_L g1131 ( 
.A1(n_919),
.A2(n_747),
.B(n_862),
.C(n_890),
.Y(n_1131)
);

AO21x2_ASAP7_75t_L g1132 ( 
.A1(n_876),
.A2(n_862),
.B(n_866),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_876),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_878),
.A2(n_747),
.B(n_730),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_878),
.Y(n_1135)
);

AO31x2_ASAP7_75t_L g1136 ( 
.A1(n_942),
.A2(n_779),
.A3(n_890),
.B(n_988),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_939),
.A2(n_947),
.B(n_928),
.Y(n_1137)
);

NAND2x1p5_ASAP7_75t_L g1138 ( 
.A(n_928),
.B(n_923),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_873),
.A2(n_730),
.B1(n_747),
.B2(n_755),
.Y(n_1139)
);

AOI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_873),
.A2(n_747),
.B1(n_730),
.B2(n_738),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_873),
.B(n_747),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_939),
.A2(n_947),
.B(n_928),
.Y(n_1142)
);

BUFx4f_ASAP7_75t_SL g1143 ( 
.A(n_955),
.Y(n_1143)
);

AOI211x1_ASAP7_75t_L g1144 ( 
.A1(n_988),
.A2(n_990),
.B(n_731),
.C(n_1018),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_866),
.A2(n_747),
.B(n_730),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_885),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_867),
.B(n_730),
.Y(n_1147)
);

OAI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_866),
.A2(n_747),
.B(n_730),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_873),
.B(n_747),
.Y(n_1149)
);

AOI221xp5_ASAP7_75t_L g1150 ( 
.A1(n_873),
.A2(n_661),
.B1(n_616),
.B2(n_747),
.C(n_791),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_873),
.B(n_747),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_873),
.B(n_747),
.Y(n_1152)
);

BUFx2_ASAP7_75t_L g1153 ( 
.A(n_912),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_939),
.A2(n_947),
.B(n_928),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_939),
.A2(n_947),
.B(n_928),
.Y(n_1155)
);

AO31x2_ASAP7_75t_L g1156 ( 
.A1(n_942),
.A2(n_779),
.A3(n_890),
.B(n_988),
.Y(n_1156)
);

AOI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_873),
.A2(n_747),
.B1(n_730),
.B2(n_738),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_873),
.B(n_747),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_885),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_863),
.B(n_788),
.Y(n_1160)
);

INVxp67_ASAP7_75t_L g1161 ( 
.A(n_1153),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_1028),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1160),
.B(n_1030),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_SL g1164 ( 
.A(n_1152),
.B(n_1028),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_L g1165 ( 
.A1(n_1152),
.A2(n_1150),
.B1(n_1149),
.B2(n_1151),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1141),
.B(n_1158),
.Y(n_1166)
);

A2O1A1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_1140),
.A2(n_1157),
.B(n_1139),
.C(n_1145),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1154),
.A2(n_1155),
.B(n_1052),
.Y(n_1168)
);

AOI21x1_ASAP7_75t_L g1169 ( 
.A1(n_1086),
.A2(n_1147),
.B(n_1059),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1084),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_SL g1171 ( 
.A(n_1134),
.B(n_1143),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1075),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1060),
.A2(n_1062),
.B1(n_1041),
.B2(n_1064),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_1131),
.B(n_1148),
.Y(n_1174)
);

OA21x2_ASAP7_75t_L g1175 ( 
.A1(n_1147),
.A2(n_1131),
.B(n_1034),
.Y(n_1175)
);

HB1xp67_ASAP7_75t_L g1176 ( 
.A(n_1075),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1049),
.Y(n_1177)
);

INVx4_ASAP7_75t_SL g1178 ( 
.A(n_1101),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1059),
.A2(n_1088),
.B(n_1070),
.Y(n_1179)
);

OAI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1033),
.A2(n_1099),
.B(n_1032),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_1078),
.B(n_1049),
.Y(n_1181)
);

A2O1A1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1033),
.A2(n_1061),
.B(n_1093),
.C(n_1024),
.Y(n_1182)
);

AOI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1107),
.A2(n_1046),
.B1(n_1102),
.B2(n_1126),
.Y(n_1183)
);

OAI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1050),
.A2(n_1074),
.B(n_1043),
.Y(n_1184)
);

HB1xp67_ASAP7_75t_L g1185 ( 
.A(n_1082),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1108),
.A2(n_1083),
.B(n_1048),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_1047),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1074),
.A2(n_1110),
.B(n_1081),
.Y(n_1188)
);

OAI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1043),
.A2(n_1104),
.B(n_1111),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_1143),
.Y(n_1190)
);

BUFx2_ASAP7_75t_L g1191 ( 
.A(n_1092),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_1078),
.Y(n_1192)
);

BUFx3_ASAP7_75t_L g1193 ( 
.A(n_1128),
.Y(n_1193)
);

NOR2x1_ASAP7_75t_R g1194 ( 
.A(n_1047),
.B(n_1133),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1083),
.A2(n_1048),
.B(n_1044),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1096),
.Y(n_1196)
);

CKINVDCx20_ASAP7_75t_R g1197 ( 
.A(n_1092),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1061),
.A2(n_1037),
.B1(n_1035),
.B2(n_1116),
.Y(n_1198)
);

INVx2_ASAP7_75t_SL g1199 ( 
.A(n_1128),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1054),
.Y(n_1200)
);

AOI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1107),
.A2(n_1046),
.B1(n_1126),
.B2(n_1095),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1097),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1113),
.A2(n_1091),
.B(n_1109),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1040),
.B(n_1026),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1077),
.Y(n_1205)
);

INVxp67_ASAP7_75t_L g1206 ( 
.A(n_1093),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1023),
.A2(n_1036),
.B1(n_1029),
.B2(n_1144),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1111),
.A2(n_1098),
.B(n_1116),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1054),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1091),
.A2(n_1119),
.B(n_1038),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1038),
.A2(n_1063),
.B(n_1067),
.Y(n_1211)
);

INVxp67_ASAP7_75t_L g1212 ( 
.A(n_1135),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1076),
.A2(n_1094),
.B(n_1055),
.Y(n_1213)
);

BUFx2_ASAP7_75t_L g1214 ( 
.A(n_1122),
.Y(n_1214)
);

BUFx8_ASAP7_75t_L g1215 ( 
.A(n_1133),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1079),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1042),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1045),
.Y(n_1218)
);

OA21x2_ASAP7_75t_L g1219 ( 
.A1(n_1072),
.A2(n_1076),
.B(n_1118),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1025),
.Y(n_1220)
);

INVx2_ASAP7_75t_SL g1221 ( 
.A(n_1128),
.Y(n_1221)
);

AND2x4_ASAP7_75t_L g1222 ( 
.A(n_1146),
.B(n_1159),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_1122),
.Y(n_1223)
);

AOI221xp5_ASAP7_75t_L g1224 ( 
.A1(n_1090),
.A2(n_1121),
.B1(n_1118),
.B2(n_1065),
.C(n_1031),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1035),
.A2(n_1090),
.B1(n_1085),
.B2(n_1039),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_1133),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1094),
.A2(n_1071),
.B(n_1138),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1071),
.A2(n_1138),
.B(n_1120),
.Y(n_1228)
);

INVxp67_ASAP7_75t_SL g1229 ( 
.A(n_1080),
.Y(n_1229)
);

NOR2xp67_ASAP7_75t_L g1230 ( 
.A(n_1130),
.B(n_1123),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1128),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1105),
.A2(n_1080),
.B1(n_1027),
.B2(n_1114),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1125),
.A2(n_1073),
.B(n_1103),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1095),
.B(n_1159),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1073),
.A2(n_1115),
.B(n_1066),
.Y(n_1235)
);

BUFx12f_ASAP7_75t_L g1236 ( 
.A(n_1133),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_1146),
.B(n_1159),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1069),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1121),
.A2(n_1053),
.B(n_1069),
.C(n_1106),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1146),
.B(n_1159),
.Y(n_1240)
);

INVxp67_ASAP7_75t_SL g1241 ( 
.A(n_1058),
.Y(n_1241)
);

INVxp67_ASAP7_75t_SL g1242 ( 
.A(n_1146),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1073),
.A2(n_1115),
.B(n_1129),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1132),
.Y(n_1244)
);

INVx6_ASAP7_75t_L g1245 ( 
.A(n_1100),
.Y(n_1245)
);

INVx5_ASAP7_75t_L g1246 ( 
.A(n_1105),
.Y(n_1246)
);

HB1xp67_ASAP7_75t_L g1247 ( 
.A(n_1101),
.Y(n_1247)
);

OR2x2_ASAP7_75t_L g1248 ( 
.A(n_1132),
.B(n_1101),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1089),
.A2(n_1112),
.B(n_1068),
.Y(n_1249)
);

BUFx10_ASAP7_75t_L g1250 ( 
.A(n_1124),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_R g1251 ( 
.A(n_1100),
.B(n_1105),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1065),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1068),
.A2(n_1057),
.B(n_1117),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1051),
.A2(n_1085),
.B(n_1136),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1117),
.A2(n_1136),
.B(n_1156),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1101),
.B(n_1136),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1117),
.A2(n_1136),
.B(n_1156),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1117),
.A2(n_1156),
.B(n_1127),
.Y(n_1258)
);

AO21x1_ASAP7_75t_L g1259 ( 
.A1(n_1056),
.A2(n_1156),
.B(n_1127),
.Y(n_1259)
);

O2A1O1Ixp33_ASAP7_75t_SL g1260 ( 
.A1(n_1056),
.A2(n_1091),
.B(n_1111),
.C(n_1116),
.Y(n_1260)
);

INVx2_ASAP7_75t_SL g1261 ( 
.A(n_1127),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1127),
.A2(n_1022),
.B(n_1137),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_1056),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1056),
.B(n_1152),
.Y(n_1264)
);

NOR2x1_ASAP7_75t_L g1265 ( 
.A(n_1110),
.B(n_682),
.Y(n_1265)
);

BUFx8_ASAP7_75t_L g1266 ( 
.A(n_1082),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_1152),
.B(n_1141),
.Y(n_1267)
);

CKINVDCx14_ASAP7_75t_R g1268 ( 
.A(n_1047),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1075),
.Y(n_1269)
);

INVx2_ASAP7_75t_SL g1270 ( 
.A(n_1028),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1075),
.Y(n_1271)
);

OAI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1141),
.A2(n_1151),
.B1(n_1158),
.B2(n_1149),
.Y(n_1272)
);

O2A1O1Ixp33_ASAP7_75t_SL g1273 ( 
.A1(n_1091),
.A2(n_1111),
.B(n_1116),
.C(n_1043),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1152),
.A2(n_1150),
.B1(n_747),
.B2(n_1149),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1152),
.B(n_1141),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1152),
.A2(n_747),
.B(n_730),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1060),
.A2(n_1148),
.B(n_1145),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1160),
.B(n_745),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1046),
.B(n_1029),
.Y(n_1279)
);

OA21x2_ASAP7_75t_L g1280 ( 
.A1(n_1145),
.A2(n_1148),
.B(n_1087),
.Y(n_1280)
);

AO21x2_ASAP7_75t_L g1281 ( 
.A1(n_1087),
.A2(n_1086),
.B(n_1147),
.Y(n_1281)
);

OAI21xp5_ASAP7_75t_SL g1282 ( 
.A1(n_1152),
.A2(n_873),
.B(n_738),
.Y(n_1282)
);

AOI21xp33_ASAP7_75t_L g1283 ( 
.A1(n_1152),
.A2(n_747),
.B(n_873),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1152),
.B(n_1141),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1075),
.Y(n_1285)
);

INVx4_ASAP7_75t_L g1286 ( 
.A(n_1080),
.Y(n_1286)
);

AOI21xp33_ASAP7_75t_L g1287 ( 
.A1(n_1152),
.A2(n_747),
.B(n_873),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1022),
.A2(n_1142),
.B(n_1137),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1084),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1028),
.Y(n_1290)
);

INVx2_ASAP7_75t_SL g1291 ( 
.A(n_1028),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1022),
.A2(n_1142),
.B(n_1137),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1160),
.B(n_745),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1022),
.A2(n_1142),
.B(n_1137),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1152),
.A2(n_1141),
.B1(n_1151),
.B2(n_1149),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1075),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1075),
.Y(n_1297)
);

AND2x4_ASAP7_75t_L g1298 ( 
.A(n_1046),
.B(n_1029),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1160),
.B(n_745),
.Y(n_1299)
);

OR2x2_ASAP7_75t_L g1300 ( 
.A(n_1028),
.B(n_1153),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_1046),
.B(n_1029),
.Y(n_1301)
);

AND2x4_ASAP7_75t_L g1302 ( 
.A(n_1046),
.B(n_1029),
.Y(n_1302)
);

AO31x2_ASAP7_75t_L g1303 ( 
.A1(n_1139),
.A2(n_1043),
.A3(n_779),
.B(n_1137),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1022),
.A2(n_1142),
.B(n_1137),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1084),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1075),
.Y(n_1306)
);

AO21x2_ASAP7_75t_L g1307 ( 
.A1(n_1087),
.A2(n_1086),
.B(n_1147),
.Y(n_1307)
);

AO31x2_ASAP7_75t_L g1308 ( 
.A1(n_1139),
.A2(n_1043),
.A3(n_779),
.B(n_1137),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1282),
.B(n_1267),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1180),
.B(n_1165),
.Y(n_1310)
);

AO22x1_ASAP7_75t_L g1311 ( 
.A1(n_1246),
.A2(n_1215),
.B1(n_1265),
.B2(n_1276),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_1300),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1176),
.Y(n_1313)
);

INVx8_ASAP7_75t_L g1314 ( 
.A(n_1246),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1267),
.B(n_1272),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1247),
.Y(n_1316)
);

HB1xp67_ASAP7_75t_L g1317 ( 
.A(n_1185),
.Y(n_1317)
);

INVx2_ASAP7_75t_SL g1318 ( 
.A(n_1245),
.Y(n_1318)
);

BUFx3_ASAP7_75t_L g1319 ( 
.A(n_1190),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1244),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1165),
.B(n_1274),
.Y(n_1321)
);

AOI222xp33_ASAP7_75t_L g1322 ( 
.A1(n_1274),
.A2(n_1295),
.B1(n_1275),
.B2(n_1284),
.C1(n_1167),
.C2(n_1166),
.Y(n_1322)
);

HB1xp67_ASAP7_75t_L g1323 ( 
.A(n_1162),
.Y(n_1323)
);

OR2x2_ASAP7_75t_L g1324 ( 
.A(n_1167),
.B(n_1264),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1200),
.B(n_1170),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1227),
.Y(n_1326)
);

OAI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1283),
.A2(n_1287),
.B1(n_1164),
.B2(n_1171),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1227),
.Y(n_1328)
);

INVx3_ASAP7_75t_L g1329 ( 
.A(n_1246),
.Y(n_1329)
);

OR2x6_ASAP7_75t_L g1330 ( 
.A(n_1188),
.B(n_1210),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1260),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1260),
.Y(n_1332)
);

INVx2_ASAP7_75t_SL g1333 ( 
.A(n_1245),
.Y(n_1333)
);

OAI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1183),
.A2(n_1201),
.B1(n_1230),
.B2(n_1206),
.Y(n_1334)
);

HB1xp67_ASAP7_75t_L g1335 ( 
.A(n_1290),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1270),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1279),
.B(n_1298),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1228),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1279),
.B(n_1298),
.Y(n_1339)
);

BUFx2_ASAP7_75t_L g1340 ( 
.A(n_1172),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1228),
.Y(n_1341)
);

OA21x2_ASAP7_75t_L g1342 ( 
.A1(n_1258),
.A2(n_1257),
.B(n_1255),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1291),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1259),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1261),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1210),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1289),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1258),
.Y(n_1348)
);

HB1xp67_ASAP7_75t_L g1349 ( 
.A(n_1161),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1178),
.Y(n_1350)
);

AO21x1_ASAP7_75t_SL g1351 ( 
.A1(n_1208),
.A2(n_1252),
.B(n_1189),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1178),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1305),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1255),
.Y(n_1354)
);

INVx1_ASAP7_75t_SL g1355 ( 
.A(n_1163),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1257),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1203),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1182),
.B(n_1256),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1203),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1216),
.Y(n_1360)
);

INVx3_ASAP7_75t_L g1361 ( 
.A(n_1246),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1233),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_1187),
.Y(n_1363)
);

AOI21xp33_ASAP7_75t_SL g1364 ( 
.A1(n_1173),
.A2(n_1182),
.B(n_1232),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1233),
.Y(n_1365)
);

INVx2_ASAP7_75t_SL g1366 ( 
.A(n_1245),
.Y(n_1366)
);

INVx3_ASAP7_75t_L g1367 ( 
.A(n_1168),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1248),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1279),
.B(n_1298),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1205),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1226),
.A2(n_1198),
.B1(n_1238),
.B2(n_1225),
.Y(n_1371)
);

INVx3_ASAP7_75t_L g1372 ( 
.A(n_1286),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1243),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1209),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1196),
.B(n_1202),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1217),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_SL g1377 ( 
.A(n_1266),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1281),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1281),
.Y(n_1379)
);

BUFx2_ASAP7_75t_L g1380 ( 
.A(n_1269),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1307),
.Y(n_1381)
);

BUFx3_ASAP7_75t_L g1382 ( 
.A(n_1190),
.Y(n_1382)
);

INVx3_ASAP7_75t_L g1383 ( 
.A(n_1286),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1218),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1220),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1307),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1263),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1263),
.Y(n_1388)
);

HB1xp67_ASAP7_75t_L g1389 ( 
.A(n_1192),
.Y(n_1389)
);

INVx3_ASAP7_75t_L g1390 ( 
.A(n_1286),
.Y(n_1390)
);

OAI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1226),
.A2(n_1234),
.B1(n_1191),
.B2(n_1197),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1278),
.B(n_1293),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1169),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1175),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1175),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1301),
.B(n_1302),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1299),
.B(n_1204),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1175),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1174),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1174),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1280),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1271),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1280),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_1214),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1235),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1285),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1198),
.A2(n_1224),
.B1(n_1250),
.B2(n_1302),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1223),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_1187),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1301),
.B(n_1302),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1301),
.B(n_1239),
.Y(n_1411)
);

INVx3_ASAP7_75t_L g1412 ( 
.A(n_1236),
.Y(n_1412)
);

AO21x2_ASAP7_75t_L g1413 ( 
.A1(n_1254),
.A2(n_1184),
.B(n_1168),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1296),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1297),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1306),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1273),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1273),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1207),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1250),
.A2(n_1197),
.B1(n_1277),
.B2(n_1219),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1250),
.A2(n_1219),
.B1(n_1225),
.B2(n_1181),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1177),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1239),
.B(n_1240),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1262),
.Y(n_1424)
);

INVx2_ASAP7_75t_SL g1425 ( 
.A(n_1215),
.Y(n_1425)
);

INVx2_ASAP7_75t_SL g1426 ( 
.A(n_1215),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1186),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1303),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1186),
.Y(n_1429)
);

AND2x4_ASAP7_75t_L g1430 ( 
.A(n_1222),
.B(n_1237),
.Y(n_1430)
);

BUFx6f_ASAP7_75t_L g1431 ( 
.A(n_1236),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1303),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1222),
.A2(n_1237),
.B1(n_1266),
.B2(n_1242),
.Y(n_1433)
);

BUFx2_ASAP7_75t_L g1434 ( 
.A(n_1251),
.Y(n_1434)
);

BUFx3_ASAP7_75t_L g1435 ( 
.A(n_1266),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1303),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1303),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_SL g1438 ( 
.A1(n_1251),
.A2(n_1268),
.B1(n_1222),
.B2(n_1237),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1308),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1229),
.B(n_1231),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1308),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1193),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1308),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1253),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1213),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1213),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_R g1447 ( 
.A(n_1363),
.B(n_1268),
.Y(n_1447)
);

BUFx3_ASAP7_75t_L g1448 ( 
.A(n_1319),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1360),
.Y(n_1449)
);

BUFx3_ASAP7_75t_L g1450 ( 
.A(n_1319),
.Y(n_1450)
);

NAND2xp33_ASAP7_75t_R g1451 ( 
.A(n_1363),
.B(n_1194),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1430),
.B(n_1231),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1310),
.B(n_1212),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_R g1454 ( 
.A(n_1409),
.B(n_1193),
.Y(n_1454)
);

INVxp67_ASAP7_75t_L g1455 ( 
.A(n_1317),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1370),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1430),
.B(n_1199),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_R g1458 ( 
.A(n_1409),
.B(n_1221),
.Y(n_1458)
);

BUFx10_ASAP7_75t_L g1459 ( 
.A(n_1431),
.Y(n_1459)
);

XNOR2xp5_ASAP7_75t_L g1460 ( 
.A(n_1377),
.B(n_1249),
.Y(n_1460)
);

BUFx3_ASAP7_75t_L g1461 ( 
.A(n_1382),
.Y(n_1461)
);

NAND2xp33_ASAP7_75t_R g1462 ( 
.A(n_1434),
.B(n_1249),
.Y(n_1462)
);

INVxp67_ASAP7_75t_L g1463 ( 
.A(n_1389),
.Y(n_1463)
);

NOR2xp33_ASAP7_75t_R g1464 ( 
.A(n_1412),
.B(n_1241),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1397),
.B(n_1195),
.Y(n_1465)
);

INVx5_ASAP7_75t_L g1466 ( 
.A(n_1314),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1355),
.B(n_1195),
.Y(n_1467)
);

INVxp67_ASAP7_75t_L g1468 ( 
.A(n_1312),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1309),
.B(n_1179),
.Y(n_1469)
);

INVxp67_ASAP7_75t_L g1470 ( 
.A(n_1349),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_1382),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1402),
.Y(n_1472)
);

AND2x4_ASAP7_75t_L g1473 ( 
.A(n_1430),
.B(n_1288),
.Y(n_1473)
);

NAND2xp33_ASAP7_75t_R g1474 ( 
.A(n_1434),
.B(n_1288),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1430),
.B(n_1211),
.Y(n_1475)
);

NAND2xp33_ASAP7_75t_SL g1476 ( 
.A(n_1431),
.B(n_1315),
.Y(n_1476)
);

INVxp67_ASAP7_75t_L g1477 ( 
.A(n_1323),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1402),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1396),
.B(n_1304),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1337),
.B(n_1292),
.Y(n_1480)
);

NAND2xp33_ASAP7_75t_R g1481 ( 
.A(n_1337),
.B(n_1292),
.Y(n_1481)
);

AND2x4_ASAP7_75t_L g1482 ( 
.A(n_1337),
.B(n_1294),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_R g1483 ( 
.A(n_1431),
.B(n_1425),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1310),
.B(n_1322),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1435),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_R g1486 ( 
.A(n_1425),
.B(n_1426),
.Y(n_1486)
);

AND2x4_ASAP7_75t_L g1487 ( 
.A(n_1337),
.B(n_1339),
.Y(n_1487)
);

OR2x6_ASAP7_75t_L g1488 ( 
.A(n_1311),
.B(n_1314),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1396),
.B(n_1410),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1423),
.B(n_1440),
.Y(n_1490)
);

NAND2xp33_ASAP7_75t_SL g1491 ( 
.A(n_1318),
.B(n_1333),
.Y(n_1491)
);

INVxp67_ASAP7_75t_L g1492 ( 
.A(n_1335),
.Y(n_1492)
);

BUFx10_ASAP7_75t_L g1493 ( 
.A(n_1318),
.Y(n_1493)
);

INVxp67_ASAP7_75t_L g1494 ( 
.A(n_1404),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_SL g1495 ( 
.A(n_1327),
.B(n_1334),
.Y(n_1495)
);

NAND2xp33_ASAP7_75t_R g1496 ( 
.A(n_1339),
.B(n_1369),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_R g1497 ( 
.A(n_1426),
.B(n_1333),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1370),
.Y(n_1498)
);

NAND2xp33_ASAP7_75t_R g1499 ( 
.A(n_1339),
.B(n_1369),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_SL g1500 ( 
.A(n_1391),
.B(n_1369),
.Y(n_1500)
);

NAND2xp33_ASAP7_75t_R g1501 ( 
.A(n_1440),
.B(n_1392),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_R g1502 ( 
.A(n_1366),
.B(n_1435),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_1336),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1376),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1406),
.Y(n_1505)
);

XOR2xp5_ASAP7_75t_L g1506 ( 
.A(n_1438),
.B(n_1311),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1406),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1376),
.Y(n_1508)
);

CKINVDCx8_ASAP7_75t_R g1509 ( 
.A(n_1313),
.Y(n_1509)
);

NAND2xp33_ASAP7_75t_R g1510 ( 
.A(n_1313),
.B(n_1375),
.Y(n_1510)
);

AND2x4_ASAP7_75t_L g1511 ( 
.A(n_1411),
.B(n_1442),
.Y(n_1511)
);

XNOR2xp5_ASAP7_75t_L g1512 ( 
.A(n_1433),
.B(n_1408),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1414),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_SL g1514 ( 
.A(n_1364),
.B(n_1321),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_R g1515 ( 
.A(n_1366),
.B(n_1329),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_R g1516 ( 
.A(n_1329),
.B(n_1361),
.Y(n_1516)
);

INVxp67_ASAP7_75t_L g1517 ( 
.A(n_1343),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1324),
.B(n_1419),
.Y(n_1518)
);

NAND2xp33_ASAP7_75t_R g1519 ( 
.A(n_1364),
.B(n_1340),
.Y(n_1519)
);

BUFx12f_ASAP7_75t_L g1520 ( 
.A(n_1340),
.Y(n_1520)
);

XNOR2xp5_ASAP7_75t_L g1521 ( 
.A(n_1371),
.B(n_1422),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1325),
.B(n_1414),
.Y(n_1522)
);

NAND2xp33_ASAP7_75t_R g1523 ( 
.A(n_1380),
.B(n_1361),
.Y(n_1523)
);

XOR2xp5_ASAP7_75t_L g1524 ( 
.A(n_1420),
.B(n_1358),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1415),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1384),
.Y(n_1526)
);

XNOR2xp5_ASAP7_75t_L g1527 ( 
.A(n_1407),
.B(n_1380),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1399),
.B(n_1400),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1400),
.B(n_1417),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1417),
.B(n_1418),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1384),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1415),
.Y(n_1532)
);

NAND2xp33_ASAP7_75t_R g1533 ( 
.A(n_1325),
.B(n_1372),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_SL g1534 ( 
.A(n_1416),
.B(n_1421),
.Y(n_1534)
);

XNOR2xp5_ASAP7_75t_L g1535 ( 
.A(n_1385),
.B(n_1358),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1387),
.Y(n_1536)
);

NAND2xp33_ASAP7_75t_R g1537 ( 
.A(n_1383),
.B(n_1390),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1374),
.B(n_1351),
.Y(n_1538)
);

NAND2xp33_ASAP7_75t_R g1539 ( 
.A(n_1390),
.B(n_1350),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1368),
.B(n_1331),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1390),
.B(n_1374),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1331),
.B(n_1332),
.Y(n_1542)
);

CKINVDCx8_ASAP7_75t_R g1543 ( 
.A(n_1330),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1387),
.Y(n_1544)
);

XNOR2xp5_ASAP7_75t_L g1545 ( 
.A(n_1347),
.B(n_1353),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_R g1546 ( 
.A(n_1352),
.B(n_1393),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1388),
.Y(n_1547)
);

AND2x4_ASAP7_75t_L g1548 ( 
.A(n_1388),
.B(n_1316),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1320),
.Y(n_1549)
);

BUFx3_ASAP7_75t_L g1550 ( 
.A(n_1345),
.Y(n_1550)
);

CKINVDCx16_ASAP7_75t_R g1551 ( 
.A(n_1330),
.Y(n_1551)
);

NAND2xp33_ASAP7_75t_R g1552 ( 
.A(n_1393),
.B(n_1330),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1428),
.B(n_1432),
.Y(n_1553)
);

XNOR2xp5_ASAP7_75t_L g1554 ( 
.A(n_1436),
.B(n_1437),
.Y(n_1554)
);

BUFx3_ASAP7_75t_L g1555 ( 
.A(n_1345),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_R g1556 ( 
.A(n_1436),
.B(n_1437),
.Y(n_1556)
);

OR2x6_ASAP7_75t_L g1557 ( 
.A(n_1330),
.B(n_1441),
.Y(n_1557)
);

CKINVDCx11_ASAP7_75t_R g1558 ( 
.A(n_1330),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_1445),
.B(n_1446),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1344),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1378),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_R g1562 ( 
.A(n_1439),
.B(n_1443),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1561),
.Y(n_1563)
);

AND2x4_ASAP7_75t_L g1564 ( 
.A(n_1473),
.B(n_1446),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1468),
.B(n_1378),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1495),
.A2(n_1441),
.B1(n_1413),
.B2(n_1405),
.Y(n_1566)
);

NOR2x1_ASAP7_75t_L g1567 ( 
.A(n_1469),
.B(n_1381),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1536),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1490),
.B(n_1405),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1544),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1547),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1560),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1473),
.B(n_1445),
.Y(n_1573)
);

INVx1_ASAP7_75t_SL g1574 ( 
.A(n_1503),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_L g1575 ( 
.A(n_1489),
.B(n_1381),
.Y(n_1575)
);

AOI21xp33_ASAP7_75t_L g1576 ( 
.A1(n_1484),
.A2(n_1413),
.B(n_1379),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1540),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1484),
.B(n_1386),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1524),
.A2(n_1413),
.B1(n_1386),
.B2(n_1367),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1538),
.B(n_1401),
.Y(n_1580)
);

INVx2_ASAP7_75t_SL g1581 ( 
.A(n_1546),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1465),
.B(n_1401),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1467),
.B(n_1403),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1528),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1475),
.B(n_1403),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1463),
.B(n_1398),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1477),
.B(n_1398),
.Y(n_1587)
);

OAI221xp5_ASAP7_75t_L g1588 ( 
.A1(n_1476),
.A2(n_1514),
.B1(n_1470),
.B2(n_1453),
.C(n_1512),
.Y(n_1588)
);

BUFx6f_ASAP7_75t_L g1589 ( 
.A(n_1488),
.Y(n_1589)
);

INVxp67_ASAP7_75t_L g1590 ( 
.A(n_1510),
.Y(n_1590)
);

INVxp67_ASAP7_75t_L g1591 ( 
.A(n_1517),
.Y(n_1591)
);

INVxp67_ASAP7_75t_SL g1592 ( 
.A(n_1533),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1528),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1549),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1551),
.B(n_1373),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1500),
.A2(n_1367),
.B1(n_1341),
.B2(n_1338),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1553),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1492),
.B(n_1394),
.Y(n_1598)
);

INVx2_ASAP7_75t_SL g1599 ( 
.A(n_1520),
.Y(n_1599)
);

BUFx2_ASAP7_75t_L g1600 ( 
.A(n_1556),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1559),
.Y(n_1601)
);

NOR2xp33_ASAP7_75t_L g1602 ( 
.A(n_1509),
.B(n_1395),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1453),
.B(n_1535),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1559),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1523),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_L g1606 ( 
.A(n_1548),
.Y(n_1606)
);

NOR2xp67_ASAP7_75t_L g1607 ( 
.A(n_1460),
.B(n_1429),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1548),
.B(n_1395),
.Y(n_1608)
);

BUFx2_ASAP7_75t_L g1609 ( 
.A(n_1562),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1506),
.A2(n_1367),
.B1(n_1338),
.B2(n_1341),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1511),
.A2(n_1367),
.B1(n_1346),
.B2(n_1328),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_SL g1612 ( 
.A1(n_1501),
.A2(n_1346),
.B1(n_1326),
.B2(n_1328),
.Y(n_1612)
);

NOR2x1_ASAP7_75t_L g1613 ( 
.A(n_1488),
.B(n_1326),
.Y(n_1613)
);

OAI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1527),
.A2(n_1424),
.B1(n_1348),
.B2(n_1354),
.Y(n_1614)
);

BUFx2_ASAP7_75t_L g1615 ( 
.A(n_1557),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1537),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1479),
.B(n_1348),
.Y(n_1617)
);

INVx1_ASAP7_75t_SL g1618 ( 
.A(n_1545),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1511),
.B(n_1354),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1521),
.A2(n_1427),
.B1(n_1429),
.B2(n_1424),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1480),
.B(n_1427),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1480),
.B(n_1359),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1518),
.B(n_1554),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1518),
.B(n_1356),
.Y(n_1624)
);

AND2x2_ASAP7_75t_SL g1625 ( 
.A(n_1496),
.B(n_1499),
.Y(n_1625)
);

INVxp67_ASAP7_75t_SL g1626 ( 
.A(n_1529),
.Y(n_1626)
);

OAI222xp33_ASAP7_75t_L g1627 ( 
.A1(n_1534),
.A2(n_1359),
.B1(n_1357),
.B2(n_1365),
.C1(n_1362),
.C2(n_1444),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1472),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1478),
.B(n_1342),
.Y(n_1629)
);

INVx1_ASAP7_75t_SL g1630 ( 
.A(n_1491),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1629),
.Y(n_1631)
);

BUFx2_ASAP7_75t_L g1632 ( 
.A(n_1615),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1597),
.B(n_1557),
.Y(n_1633)
);

BUFx3_ASAP7_75t_L g1634 ( 
.A(n_1589),
.Y(n_1634)
);

NAND3xp33_ASAP7_75t_L g1635 ( 
.A(n_1588),
.B(n_1519),
.C(n_1455),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1572),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1629),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1626),
.B(n_1505),
.Y(n_1638)
);

BUFx2_ASAP7_75t_L g1639 ( 
.A(n_1615),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1572),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1563),
.Y(n_1641)
);

AOI221xp5_ASAP7_75t_L g1642 ( 
.A1(n_1614),
.A2(n_1494),
.B1(n_1507),
.B2(n_1532),
.C(n_1513),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1563),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1585),
.B(n_1617),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1568),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1623),
.A2(n_1558),
.B1(n_1485),
.B2(n_1488),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1594),
.Y(n_1647)
);

OAI31xp33_ASAP7_75t_L g1648 ( 
.A1(n_1618),
.A2(n_1461),
.A3(n_1450),
.B(n_1448),
.Y(n_1648)
);

BUFx2_ASAP7_75t_L g1649 ( 
.A(n_1564),
.Y(n_1649)
);

OAI31xp33_ASAP7_75t_L g1650 ( 
.A1(n_1618),
.A2(n_1550),
.A3(n_1555),
.B(n_1457),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1582),
.B(n_1580),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1580),
.B(n_1564),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1578),
.B(n_1525),
.Y(n_1653)
);

INVx3_ASAP7_75t_L g1654 ( 
.A(n_1564),
.Y(n_1654)
);

INVxp67_ASAP7_75t_SL g1655 ( 
.A(n_1567),
.Y(n_1655)
);

AOI22xp5_ASAP7_75t_L g1656 ( 
.A1(n_1603),
.A2(n_1539),
.B1(n_1451),
.B2(n_1487),
.Y(n_1656)
);

INVx5_ASAP7_75t_L g1657 ( 
.A(n_1589),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1594),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1570),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1571),
.Y(n_1660)
);

BUFx3_ASAP7_75t_L g1661 ( 
.A(n_1589),
.Y(n_1661)
);

INVx3_ASAP7_75t_L g1662 ( 
.A(n_1573),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1571),
.Y(n_1663)
);

AOI33xp33_ASAP7_75t_L g1664 ( 
.A1(n_1620),
.A2(n_1456),
.A3(n_1449),
.B1(n_1498),
.B2(n_1531),
.B3(n_1526),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1577),
.Y(n_1665)
);

NAND3xp33_ASAP7_75t_L g1666 ( 
.A(n_1576),
.B(n_1462),
.C(n_1474),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1584),
.B(n_1522),
.Y(n_1667)
);

INVxp67_ASAP7_75t_SL g1668 ( 
.A(n_1567),
.Y(n_1668)
);

INVxp67_ASAP7_75t_SL g1669 ( 
.A(n_1577),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1573),
.B(n_1482),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1628),
.Y(n_1671)
);

AND2x2_ASAP7_75t_SL g1672 ( 
.A(n_1625),
.B(n_1543),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1583),
.B(n_1586),
.Y(n_1673)
);

INVx5_ASAP7_75t_SL g1674 ( 
.A(n_1625),
.Y(n_1674)
);

OAI31xp33_ASAP7_75t_L g1675 ( 
.A1(n_1630),
.A2(n_1457),
.A3(n_1452),
.B(n_1541),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1593),
.B(n_1624),
.Y(n_1676)
);

OAI221xp5_ASAP7_75t_SL g1677 ( 
.A1(n_1579),
.A2(n_1508),
.B1(n_1504),
.B2(n_1542),
.C(n_1530),
.Y(n_1677)
);

INVx1_ASAP7_75t_SL g1678 ( 
.A(n_1616),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1649),
.B(n_1601),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1631),
.B(n_1601),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1649),
.B(n_1622),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1649),
.B(n_1622),
.Y(n_1682)
);

OR2x6_ASAP7_75t_L g1683 ( 
.A(n_1666),
.B(n_1589),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1652),
.B(n_1622),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1631),
.B(n_1637),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1631),
.B(n_1583),
.Y(n_1686)
);

NAND2xp33_ASAP7_75t_SL g1687 ( 
.A(n_1646),
.B(n_1581),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1665),
.B(n_1624),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1640),
.Y(n_1689)
);

AND2x2_ASAP7_75t_SL g1690 ( 
.A(n_1672),
.B(n_1625),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1631),
.B(n_1604),
.Y(n_1691)
);

INVx3_ASAP7_75t_L g1692 ( 
.A(n_1654),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1637),
.B(n_1604),
.Y(n_1693)
);

INVx2_ASAP7_75t_SL g1694 ( 
.A(n_1654),
.Y(n_1694)
);

INVx3_ASAP7_75t_SL g1695 ( 
.A(n_1672),
.Y(n_1695)
);

INVx3_ASAP7_75t_L g1696 ( 
.A(n_1654),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1652),
.B(n_1619),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1644),
.B(n_1619),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1644),
.B(n_1608),
.Y(n_1699)
);

NOR2xp67_ASAP7_75t_L g1700 ( 
.A(n_1666),
.B(n_1605),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1644),
.B(n_1608),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1678),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1637),
.B(n_1595),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1651),
.B(n_1621),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1637),
.B(n_1595),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1660),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1651),
.B(n_1621),
.Y(n_1707)
);

NOR2xp33_ASAP7_75t_L g1708 ( 
.A(n_1678),
.B(n_1599),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1635),
.B(n_1599),
.Y(n_1709)
);

AND2x4_ASAP7_75t_L g1710 ( 
.A(n_1657),
.B(n_1613),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1654),
.B(n_1662),
.Y(n_1711)
);

AND2x4_ASAP7_75t_L g1712 ( 
.A(n_1657),
.B(n_1613),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1673),
.B(n_1587),
.Y(n_1713)
);

NAND2x1p5_ASAP7_75t_L g1714 ( 
.A(n_1657),
.B(n_1600),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1673),
.B(n_1598),
.Y(n_1715)
);

NAND2x1p5_ASAP7_75t_L g1716 ( 
.A(n_1657),
.B(n_1600),
.Y(n_1716)
);

NOR2xp67_ASAP7_75t_L g1717 ( 
.A(n_1657),
.B(n_1581),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1662),
.B(n_1670),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1662),
.B(n_1569),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1691),
.Y(n_1720)
);

AOI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1687),
.A2(n_1672),
.B1(n_1656),
.B2(n_1635),
.Y(n_1721)
);

NOR2xp33_ASAP7_75t_R g1722 ( 
.A(n_1695),
.B(n_1471),
.Y(n_1722)
);

CKINVDCx14_ASAP7_75t_R g1723 ( 
.A(n_1708),
.Y(n_1723)
);

AO221x2_ASAP7_75t_L g1724 ( 
.A1(n_1700),
.A2(n_1627),
.B1(n_1648),
.B2(n_1656),
.C(n_1676),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1713),
.B(n_1673),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1702),
.B(n_1623),
.Y(n_1726)
);

OAI22xp33_ASAP7_75t_L g1727 ( 
.A1(n_1695),
.A2(n_1607),
.B1(n_1609),
.B2(n_1590),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1700),
.B(n_1676),
.Y(n_1728)
);

OAI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1695),
.A2(n_1646),
.B1(n_1674),
.B2(n_1672),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1691),
.Y(n_1730)
);

NAND2xp33_ASAP7_75t_SL g1731 ( 
.A(n_1690),
.B(n_1454),
.Y(n_1731)
);

AOI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1690),
.A2(n_1674),
.B1(n_1607),
.B2(n_1670),
.Y(n_1732)
);

NAND2xp33_ASAP7_75t_SL g1733 ( 
.A(n_1690),
.B(n_1502),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_SL g1734 ( 
.A(n_1709),
.B(n_1648),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1713),
.B(n_1574),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1715),
.B(n_1591),
.Y(n_1736)
);

INVx3_ASAP7_75t_L g1737 ( 
.A(n_1693),
.Y(n_1737)
);

NOR2xp33_ASAP7_75t_L g1738 ( 
.A(n_1715),
.B(n_1653),
.Y(n_1738)
);

AND2x4_ASAP7_75t_L g1739 ( 
.A(n_1717),
.B(n_1657),
.Y(n_1739)
);

NOR4xp25_ASAP7_75t_SL g1740 ( 
.A(n_1714),
.B(n_1609),
.C(n_1668),
.D(n_1655),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1719),
.Y(n_1741)
);

AO221x2_ASAP7_75t_L g1742 ( 
.A1(n_1683),
.A2(n_1653),
.B1(n_1674),
.B2(n_1667),
.C(n_1645),
.Y(n_1742)
);

OAI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1683),
.A2(n_1674),
.B1(n_1612),
.B2(n_1610),
.Y(n_1743)
);

OAI221xp5_ASAP7_75t_L g1744 ( 
.A1(n_1683),
.A2(n_1650),
.B1(n_1675),
.B2(n_1630),
.C(n_1642),
.Y(n_1744)
);

INVx4_ASAP7_75t_L g1745 ( 
.A(n_1714),
.Y(n_1745)
);

AO221x2_ASAP7_75t_L g1746 ( 
.A1(n_1683),
.A2(n_1674),
.B1(n_1667),
.B2(n_1636),
.C(n_1645),
.Y(n_1746)
);

NAND2xp33_ASAP7_75t_SL g1747 ( 
.A(n_1710),
.B(n_1458),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1699),
.B(n_1647),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_L g1749 ( 
.A(n_1697),
.B(n_1684),
.Y(n_1749)
);

AOI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1683),
.A2(n_1674),
.B1(n_1670),
.B2(n_1592),
.Y(n_1750)
);

INVxp67_ASAP7_75t_L g1751 ( 
.A(n_1688),
.Y(n_1751)
);

AO221x2_ASAP7_75t_L g1752 ( 
.A1(n_1688),
.A2(n_1636),
.B1(n_1641),
.B2(n_1643),
.C(n_1659),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1699),
.B(n_1647),
.Y(n_1753)
);

AO221x2_ASAP7_75t_L g1754 ( 
.A1(n_1689),
.A2(n_1663),
.B1(n_1643),
.B2(n_1641),
.C(n_1659),
.Y(n_1754)
);

AO221x2_ASAP7_75t_L g1755 ( 
.A1(n_1689),
.A2(n_1663),
.B1(n_1650),
.B2(n_1671),
.C(n_1638),
.Y(n_1755)
);

INVxp67_ASAP7_75t_L g1756 ( 
.A(n_1679),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1703),
.B(n_1632),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1693),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1701),
.B(n_1658),
.Y(n_1759)
);

BUFx2_ASAP7_75t_L g1760 ( 
.A(n_1714),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_L g1761 ( 
.A(n_1697),
.B(n_1670),
.Y(n_1761)
);

AOI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1717),
.A2(n_1670),
.B1(n_1642),
.B2(n_1661),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_1710),
.Y(n_1763)
);

CKINVDCx8_ASAP7_75t_R g1764 ( 
.A(n_1710),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1742),
.B(n_1718),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1754),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1754),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1752),
.Y(n_1768)
);

INVx1_ASAP7_75t_SL g1769 ( 
.A(n_1722),
.Y(n_1769)
);

INVxp67_ASAP7_75t_L g1770 ( 
.A(n_1734),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1742),
.B(n_1718),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1752),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1746),
.B(n_1711),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1755),
.B(n_1703),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1720),
.Y(n_1775)
);

AND2x4_ASAP7_75t_L g1776 ( 
.A(n_1739),
.B(n_1710),
.Y(n_1776)
);

INVxp33_ASAP7_75t_L g1777 ( 
.A(n_1736),
.Y(n_1777)
);

INVx1_ASAP7_75t_SL g1778 ( 
.A(n_1726),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1755),
.B(n_1705),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1746),
.B(n_1711),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1738),
.B(n_1701),
.Y(n_1781)
);

NAND2x1p5_ASAP7_75t_L g1782 ( 
.A(n_1745),
.B(n_1657),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_L g1783 ( 
.A(n_1723),
.B(n_1684),
.Y(n_1783)
);

AOI222xp33_ASAP7_75t_L g1784 ( 
.A1(n_1743),
.A2(n_1729),
.B1(n_1744),
.B2(n_1731),
.C1(n_1733),
.C2(n_1728),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1737),
.Y(n_1785)
);

OA22x2_ASAP7_75t_L g1786 ( 
.A1(n_1721),
.A2(n_1762),
.B1(n_1750),
.B2(n_1732),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1741),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1760),
.B(n_1681),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1730),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1725),
.B(n_1705),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1758),
.Y(n_1791)
);

INVx1_ASAP7_75t_SL g1792 ( 
.A(n_1747),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1748),
.Y(n_1793)
);

AOI22xp33_ASAP7_75t_SL g1794 ( 
.A1(n_1724),
.A2(n_1716),
.B1(n_1657),
.B2(n_1655),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1764),
.B(n_1681),
.Y(n_1795)
);

INVx1_ASAP7_75t_SL g1796 ( 
.A(n_1763),
.Y(n_1796)
);

OR2x2_ASAP7_75t_L g1797 ( 
.A(n_1751),
.B(n_1686),
.Y(n_1797)
);

INVx2_ASAP7_75t_SL g1798 ( 
.A(n_1739),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1724),
.B(n_1698),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1753),
.Y(n_1800)
);

INVx1_ASAP7_75t_SL g1801 ( 
.A(n_1735),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1759),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1757),
.Y(n_1803)
);

HB1xp67_ASAP7_75t_L g1804 ( 
.A(n_1756),
.Y(n_1804)
);

HB1xp67_ASAP7_75t_L g1805 ( 
.A(n_1749),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1761),
.B(n_1682),
.Y(n_1806)
);

INVx1_ASAP7_75t_SL g1807 ( 
.A(n_1727),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1740),
.B(n_1698),
.Y(n_1808)
);

INVxp67_ASAP7_75t_L g1809 ( 
.A(n_1734),
.Y(n_1809)
);

AND2x4_ASAP7_75t_L g1810 ( 
.A(n_1739),
.B(n_1712),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1798),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1775),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1775),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1789),
.Y(n_1814)
);

AOI221xp5_ASAP7_75t_L g1815 ( 
.A1(n_1770),
.A2(n_1677),
.B1(n_1668),
.B2(n_1638),
.C(n_1658),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1809),
.B(n_1704),
.Y(n_1816)
);

OR2x2_ASAP7_75t_L g1817 ( 
.A(n_1778),
.B(n_1680),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1789),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1791),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1791),
.Y(n_1820)
);

NAND2xp33_ASAP7_75t_SL g1821 ( 
.A(n_1774),
.B(n_1447),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1805),
.B(n_1704),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1801),
.B(n_1707),
.Y(n_1823)
);

OR2x2_ASAP7_75t_L g1824 ( 
.A(n_1781),
.B(n_1680),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1804),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1803),
.Y(n_1826)
);

AOI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1794),
.A2(n_1712),
.B1(n_1716),
.B2(n_1602),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1803),
.Y(n_1828)
);

OAI211xp5_ASAP7_75t_L g1829 ( 
.A1(n_1784),
.A2(n_1675),
.B(n_1596),
.C(n_1566),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1787),
.Y(n_1830)
);

O2A1O1Ixp5_ASAP7_75t_L g1831 ( 
.A1(n_1799),
.A2(n_1677),
.B(n_1712),
.C(n_1692),
.Y(n_1831)
);

OAI322xp33_ASAP7_75t_L g1832 ( 
.A1(n_1768),
.A2(n_1716),
.A3(n_1685),
.B1(n_1686),
.B2(n_1565),
.C1(n_1669),
.C2(n_1706),
.Y(n_1832)
);

AOI21xp5_ASAP7_75t_L g1833 ( 
.A1(n_1786),
.A2(n_1712),
.B(n_1669),
.Y(n_1833)
);

INVxp67_ASAP7_75t_L g1834 ( 
.A(n_1768),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1787),
.Y(n_1835)
);

INVx1_ASAP7_75t_SL g1836 ( 
.A(n_1769),
.Y(n_1836)
);

INVx1_ASAP7_75t_SL g1837 ( 
.A(n_1792),
.Y(n_1837)
);

INVx1_ASAP7_75t_SL g1838 ( 
.A(n_1796),
.Y(n_1838)
);

AOI22xp5_ASAP7_75t_L g1839 ( 
.A1(n_1786),
.A2(n_1634),
.B1(n_1661),
.B2(n_1657),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1798),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1766),
.Y(n_1841)
);

HB1xp67_ASAP7_75t_L g1842 ( 
.A(n_1767),
.Y(n_1842)
);

OAI211xp5_ASAP7_75t_SL g1843 ( 
.A1(n_1807),
.A2(n_1664),
.B(n_1611),
.C(n_1633),
.Y(n_1843)
);

AOI21xp33_ASAP7_75t_SL g1844 ( 
.A1(n_1786),
.A2(n_1694),
.B(n_1692),
.Y(n_1844)
);

INVxp67_ASAP7_75t_L g1845 ( 
.A(n_1767),
.Y(n_1845)
);

XNOR2xp5_ASAP7_75t_L g1846 ( 
.A(n_1777),
.B(n_1487),
.Y(n_1846)
);

OAI221xp5_ASAP7_75t_L g1847 ( 
.A1(n_1774),
.A2(n_1661),
.B1(n_1634),
.B2(n_1639),
.C(n_1632),
.Y(n_1847)
);

AOI22xp5_ASAP7_75t_L g1848 ( 
.A1(n_1783),
.A2(n_1661),
.B1(n_1634),
.B2(n_1575),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1837),
.B(n_1772),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1836),
.B(n_1772),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1812),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1813),
.Y(n_1852)
);

INVx1_ASAP7_75t_SL g1853 ( 
.A(n_1821),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_SL g1854 ( 
.A(n_1838),
.B(n_1779),
.Y(n_1854)
);

NOR3xp33_ASAP7_75t_SL g1855 ( 
.A(n_1821),
.B(n_1808),
.C(n_1800),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1814),
.Y(n_1856)
);

NOR2xp33_ASAP7_75t_L g1857 ( 
.A(n_1825),
.B(n_1779),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_L g1858 ( 
.A(n_1846),
.B(n_1793),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1841),
.B(n_1793),
.Y(n_1859)
);

NOR2xp33_ASAP7_75t_L g1860 ( 
.A(n_1834),
.B(n_1800),
.Y(n_1860)
);

NAND2x1_ASAP7_75t_L g1861 ( 
.A(n_1839),
.B(n_1795),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1822),
.B(n_1802),
.Y(n_1862)
);

AND2x4_ASAP7_75t_L g1863 ( 
.A(n_1811),
.B(n_1795),
.Y(n_1863)
);

AOI22xp33_ASAP7_75t_L g1864 ( 
.A1(n_1834),
.A2(n_1802),
.B1(n_1765),
.B2(n_1771),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1840),
.B(n_1785),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1844),
.B(n_1765),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1848),
.B(n_1806),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1818),
.Y(n_1868)
);

BUFx2_ASAP7_75t_L g1869 ( 
.A(n_1842),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1819),
.Y(n_1870)
);

OAI21xp5_ASAP7_75t_SL g1871 ( 
.A1(n_1827),
.A2(n_1771),
.B(n_1773),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1820),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1830),
.Y(n_1873)
);

OR2x2_ASAP7_75t_L g1874 ( 
.A(n_1816),
.B(n_1797),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1835),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1826),
.B(n_1785),
.Y(n_1876)
);

CKINVDCx20_ASAP7_75t_R g1877 ( 
.A(n_1853),
.Y(n_1877)
);

INVxp33_ASAP7_75t_SL g1878 ( 
.A(n_1854),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1869),
.Y(n_1879)
);

BUFx4f_ASAP7_75t_SL g1880 ( 
.A(n_1863),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1857),
.B(n_1845),
.Y(n_1881)
);

INVx1_ASAP7_75t_SL g1882 ( 
.A(n_1863),
.Y(n_1882)
);

CKINVDCx6p67_ASAP7_75t_R g1883 ( 
.A(n_1850),
.Y(n_1883)
);

BUFx2_ASAP7_75t_L g1884 ( 
.A(n_1849),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1851),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1852),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1874),
.Y(n_1887)
);

BUFx6f_ASAP7_75t_L g1888 ( 
.A(n_1861),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1856),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1867),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1868),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1870),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1872),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1873),
.Y(n_1894)
);

CKINVDCx20_ASAP7_75t_R g1895 ( 
.A(n_1855),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1875),
.Y(n_1896)
);

INVxp33_ASAP7_75t_SL g1897 ( 
.A(n_1860),
.Y(n_1897)
);

NAND4xp25_ASAP7_75t_L g1898 ( 
.A(n_1878),
.B(n_1864),
.C(n_1866),
.D(n_1871),
.Y(n_1898)
);

AOI21xp5_ASAP7_75t_L g1899 ( 
.A1(n_1878),
.A2(n_1866),
.B(n_1864),
.Y(n_1899)
);

O2A1O1Ixp33_ASAP7_75t_L g1900 ( 
.A1(n_1895),
.A2(n_1855),
.B(n_1860),
.C(n_1845),
.Y(n_1900)
);

NAND4xp75_ASAP7_75t_L g1901 ( 
.A(n_1879),
.B(n_1881),
.C(n_1887),
.D(n_1890),
.Y(n_1901)
);

NOR2x1_ASAP7_75t_L g1902 ( 
.A(n_1877),
.B(n_1865),
.Y(n_1902)
);

NOR3xp33_ASAP7_75t_L g1903 ( 
.A(n_1884),
.B(n_1859),
.C(n_1876),
.Y(n_1903)
);

NOR2x1_ASAP7_75t_L g1904 ( 
.A(n_1879),
.B(n_1828),
.Y(n_1904)
);

NAND4xp75_ASAP7_75t_L g1905 ( 
.A(n_1887),
.B(n_1831),
.C(n_1833),
.D(n_1815),
.Y(n_1905)
);

NOR3x1_ASAP7_75t_L g1906 ( 
.A(n_1884),
.B(n_1847),
.C(n_1829),
.Y(n_1906)
);

NAND4xp25_ASAP7_75t_L g1907 ( 
.A(n_1890),
.B(n_1882),
.C(n_1897),
.D(n_1886),
.Y(n_1907)
);

NAND5xp2_ASAP7_75t_L g1908 ( 
.A(n_1897),
.B(n_1858),
.C(n_1782),
.D(n_1773),
.E(n_1780),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1883),
.B(n_1842),
.Y(n_1909)
);

OR2x2_ASAP7_75t_L g1910 ( 
.A(n_1883),
.B(n_1862),
.Y(n_1910)
);

AOI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1900),
.A2(n_1888),
.B(n_1892),
.Y(n_1911)
);

AOI22xp5_ASAP7_75t_L g1912 ( 
.A1(n_1905),
.A2(n_1880),
.B1(n_1888),
.B2(n_1889),
.Y(n_1912)
);

AOI21xp5_ASAP7_75t_L g1913 ( 
.A1(n_1899),
.A2(n_1888),
.B(n_1892),
.Y(n_1913)
);

OAI22xp5_ASAP7_75t_L g1914 ( 
.A1(n_1902),
.A2(n_1888),
.B1(n_1823),
.B2(n_1782),
.Y(n_1914)
);

OAI211xp5_ASAP7_75t_SL g1915 ( 
.A1(n_1910),
.A2(n_1896),
.B(n_1893),
.C(n_1891),
.Y(n_1915)
);

XOR2xp5_ASAP7_75t_L g1916 ( 
.A(n_1898),
.B(n_1888),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1904),
.Y(n_1917)
);

INVx1_ASAP7_75t_SL g1918 ( 
.A(n_1909),
.Y(n_1918)
);

OAI221xp5_ASAP7_75t_SL g1919 ( 
.A1(n_1907),
.A2(n_1893),
.B1(n_1891),
.B2(n_1885),
.C(n_1894),
.Y(n_1919)
);

OAI311xp33_ASAP7_75t_L g1920 ( 
.A1(n_1906),
.A2(n_1894),
.A3(n_1885),
.B1(n_1817),
.C1(n_1780),
.Y(n_1920)
);

NAND4xp75_ASAP7_75t_L g1921 ( 
.A(n_1901),
.B(n_1831),
.C(n_1788),
.D(n_1832),
.Y(n_1921)
);

AOI221xp5_ASAP7_75t_L g1922 ( 
.A1(n_1908),
.A2(n_1843),
.B1(n_1782),
.B2(n_1810),
.C(n_1776),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1917),
.Y(n_1923)
);

AOI21xp5_ASAP7_75t_L g1924 ( 
.A1(n_1913),
.A2(n_1903),
.B(n_1843),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1911),
.B(n_1788),
.Y(n_1925)
);

NOR2x1_ASAP7_75t_L g1926 ( 
.A(n_1916),
.B(n_1776),
.Y(n_1926)
);

OR2x2_ASAP7_75t_L g1927 ( 
.A(n_1918),
.B(n_1919),
.Y(n_1927)
);

NOR2x1_ASAP7_75t_L g1928 ( 
.A(n_1915),
.B(n_1776),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1914),
.Y(n_1929)
);

NAND2x1p5_ASAP7_75t_L g1930 ( 
.A(n_1912),
.B(n_1810),
.Y(n_1930)
);

NAND3xp33_ASAP7_75t_SL g1931 ( 
.A(n_1924),
.B(n_1922),
.C(n_1920),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1925),
.B(n_1921),
.Y(n_1932)
);

NAND2xp33_ASAP7_75t_SL g1933 ( 
.A(n_1927),
.B(n_1486),
.Y(n_1933)
);

NOR2xp33_ASAP7_75t_R g1934 ( 
.A(n_1929),
.B(n_1493),
.Y(n_1934)
);

OAI21x1_ASAP7_75t_L g1935 ( 
.A1(n_1928),
.A2(n_1824),
.B(n_1797),
.Y(n_1935)
);

NAND3xp33_ASAP7_75t_SL g1936 ( 
.A(n_1930),
.B(n_1497),
.C(n_1483),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1923),
.B(n_1810),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_R g1938 ( 
.A(n_1926),
.B(n_1493),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1935),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1937),
.Y(n_1940)
);

AOI221xp5_ASAP7_75t_L g1941 ( 
.A1(n_1931),
.A2(n_1806),
.B1(n_1790),
.B2(n_1639),
.C(n_1632),
.Y(n_1941)
);

OAI22xp5_ASAP7_75t_SL g1942 ( 
.A1(n_1932),
.A2(n_1790),
.B1(n_1466),
.B2(n_1634),
.Y(n_1942)
);

AND2x4_ASAP7_75t_L g1943 ( 
.A(n_1938),
.B(n_1692),
.Y(n_1943)
);

AOI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1933),
.A2(n_1936),
.B1(n_1934),
.B2(n_1694),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1939),
.B(n_1692),
.Y(n_1945)
);

OAI21xp5_ASAP7_75t_SL g1946 ( 
.A1(n_1941),
.A2(n_1639),
.B(n_1696),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1943),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1940),
.Y(n_1948)
);

OAI22xp5_ASAP7_75t_SL g1949 ( 
.A1(n_1948),
.A2(n_1942),
.B1(n_1944),
.B2(n_1466),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_SL g1950 ( 
.A(n_1947),
.B(n_1696),
.Y(n_1950)
);

AOI31xp33_ASAP7_75t_L g1951 ( 
.A1(n_1950),
.A2(n_1945),
.A3(n_1946),
.B(n_1606),
.Y(n_1951)
);

XNOR2xp5_ASAP7_75t_L g1952 ( 
.A(n_1951),
.B(n_1949),
.Y(n_1952)
);

NAND4xp25_ASAP7_75t_SL g1953 ( 
.A(n_1951),
.B(n_1664),
.C(n_1682),
.D(n_1719),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1952),
.Y(n_1954)
);

HB1xp67_ASAP7_75t_L g1955 ( 
.A(n_1953),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1954),
.B(n_1696),
.Y(n_1956)
);

OAI221xp5_ASAP7_75t_R g1957 ( 
.A1(n_1956),
.A2(n_1955),
.B1(n_1552),
.B2(n_1481),
.C(n_1459),
.Y(n_1957)
);

AOI211xp5_ASAP7_75t_L g1958 ( 
.A1(n_1957),
.A2(n_1464),
.B(n_1515),
.C(n_1516),
.Y(n_1958)
);


endmodule