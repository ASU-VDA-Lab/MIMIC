module fake_aes_2941_n_44 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_44);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_44;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_30;
wire n_13;
wire n_26;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_3), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_5), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_3), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_8), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_6), .Y(n_15) );
INVx1_ASAP7_75t_SL g16 ( .A(n_6), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_9), .Y(n_17) );
OR2x2_ASAP7_75t_SL g18 ( .A(n_15), .B(n_0), .Y(n_18) );
AND3x2_ASAP7_75t_SL g19 ( .A(n_12), .B(n_0), .C(n_1), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_11), .B(n_1), .Y(n_20) );
AND2x4_ASAP7_75t_L g21 ( .A(n_12), .B(n_2), .Y(n_21) );
HB1xp67_ASAP7_75t_L g22 ( .A(n_12), .Y(n_22) );
INVx5_ASAP7_75t_L g23 ( .A(n_15), .Y(n_23) );
AOI22xp5_ASAP7_75t_L g24 ( .A1(n_21), .A2(n_14), .B1(n_13), .B2(n_16), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_22), .B(n_14), .Y(n_25) );
AOI22xp33_ASAP7_75t_L g26 ( .A1(n_21), .A2(n_13), .B1(n_17), .B2(n_5), .Y(n_26) );
AOI22xp33_ASAP7_75t_L g27 ( .A1(n_21), .A2(n_2), .B1(n_4), .B2(n_7), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
BUFx3_ASAP7_75t_L g29 ( .A(n_25), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_27), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_29), .Y(n_31) );
INVx1_ASAP7_75t_SL g32 ( .A(n_29), .Y(n_32) );
A2O1A1Ixp33_ASAP7_75t_L g33 ( .A1(n_31), .A2(n_30), .B(n_28), .C(n_26), .Y(n_33) );
NOR2xp33_ASAP7_75t_R g34 ( .A(n_31), .B(n_29), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_32), .Y(n_35) );
INVx1_ASAP7_75t_SL g36 ( .A(n_34), .Y(n_36) );
OAI322xp33_ASAP7_75t_L g37 ( .A1(n_35), .A2(n_24), .A3(n_28), .B1(n_30), .B2(n_20), .C1(n_22), .C2(n_19), .Y(n_37) );
INVx1_ASAP7_75t_L g38 ( .A(n_33), .Y(n_38) );
INVx1_ASAP7_75t_L g39 ( .A(n_37), .Y(n_39) );
AOI221xp5_ASAP7_75t_L g40 ( .A1(n_38), .A2(n_35), .B1(n_23), .B2(n_19), .C(n_18), .Y(n_40) );
OAI211xp5_ASAP7_75t_L g41 ( .A1(n_36), .A2(n_23), .B(n_7), .C(n_8), .Y(n_41) );
OAI22xp5_ASAP7_75t_L g42 ( .A1(n_39), .A2(n_38), .B1(n_23), .B2(n_4), .Y(n_42) );
AND2x4_ASAP7_75t_L g43 ( .A(n_41), .B(n_23), .Y(n_43) );
AOI22xp33_ASAP7_75t_L g44 ( .A1(n_43), .A2(n_10), .B1(n_40), .B2(n_42), .Y(n_44) );
endmodule