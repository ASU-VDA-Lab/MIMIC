module fake_jpeg_6698_n_300 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_118;
wire n_128;
wire n_82;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_17),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_33),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_36),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_35),
.Y(n_57)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_38),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_22),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_20),
.B(n_25),
.Y(n_39)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_40),
.A2(n_27),
.B1(n_21),
.B2(n_30),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_41),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_36),
.A2(n_27),
.B1(n_21),
.B2(n_26),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_42),
.A2(n_52),
.B(n_18),
.Y(n_73)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_47),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_27),
.B1(n_20),
.B2(n_25),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_51),
.B1(n_62),
.B2(n_34),
.Y(n_69)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_54),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_23),
.B1(n_15),
.B2(n_26),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_36),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_32),
.Y(n_79)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_36),
.A2(n_24),
.B1(n_28),
.B2(n_15),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_60),
.A2(n_40),
.B1(n_34),
.B2(n_31),
.Y(n_68)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_36),
.A2(n_40),
.B1(n_37),
.B2(n_39),
.Y(n_62)
);

AO22x1_ASAP7_75t_SL g64 ( 
.A1(n_62),
.A2(n_33),
.B1(n_36),
.B2(n_37),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_64),
.A2(n_56),
.B1(n_49),
.B2(n_44),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_37),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_75),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_68),
.A2(n_80),
.B1(n_81),
.B2(n_38),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_69),
.A2(n_40),
.B1(n_38),
.B2(n_57),
.Y(n_96)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_74),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_33),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_72),
.B(n_33),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_73),
.A2(n_78),
.B(n_18),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_31),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_33),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_45),
.A2(n_33),
.B(n_32),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_79),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_40),
.B1(n_34),
.B2(n_31),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_61),
.A2(n_40),
.B1(n_34),
.B2(n_31),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_33),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_57),
.Y(n_93)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_85),
.Y(n_101)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_86),
.A2(n_104),
.B(n_107),
.Y(n_116)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_92),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_58),
.B(n_46),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_105),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_58),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_64),
.C(n_69),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_77),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_106),
.Y(n_112)
);

AO22x1_ASAP7_75t_SL g94 ( 
.A1(n_64),
.A2(n_40),
.B1(n_28),
.B2(n_15),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_94),
.A2(n_76),
.B1(n_70),
.B2(n_66),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_72),
.B(n_47),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_98),
.Y(n_119)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_102),
.Y(n_120)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_72),
.B(n_74),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_74),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_32),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_32),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g107 ( 
.A1(n_83),
.A2(n_38),
.B(n_14),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_108),
.B(n_70),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_101),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_111),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_101),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_71),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_128),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_95),
.C(n_103),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_115),
.B(n_122),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_104),
.A2(n_64),
.B(n_73),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_121),
.A2(n_124),
.B(n_106),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_92),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_123),
.A2(n_96),
.B1(n_94),
.B2(n_99),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_125),
.B(n_100),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_126),
.B(n_97),
.Y(n_149)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_129),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_79),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_88),
.Y(n_129)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_63),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_93),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_132),
.Y(n_151)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_133),
.Y(n_146)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_136),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_135),
.A2(n_154),
.B(n_110),
.Y(n_177)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_137),
.A2(n_150),
.B1(n_153),
.B2(n_146),
.Y(n_179)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_139),
.Y(n_164)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

AOI32xp33_ASAP7_75t_L g140 ( 
.A1(n_121),
.A2(n_90),
.A3(n_130),
.B1(n_116),
.B2(n_86),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_140),
.A2(n_149),
.B(n_131),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_94),
.B1(n_87),
.B2(n_98),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_156),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_91),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_132),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_155),
.Y(n_160)
);

OA22x2_ASAP7_75t_L g150 ( 
.A1(n_133),
.A2(n_100),
.B1(n_76),
.B2(n_105),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_152),
.B(n_125),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_118),
.A2(n_85),
.B1(n_66),
.B2(n_82),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_116),
.A2(n_77),
.B(n_57),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_114),
.C(n_112),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_135),
.A2(n_133),
.B1(n_117),
.B2(n_123),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_184),
.B1(n_146),
.B2(n_137),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_158),
.B(n_129),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_163),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_140),
.A2(n_112),
.B(n_119),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_170),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_167),
.B(n_172),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_158),
.B(n_122),
.Y(n_169)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_130),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_147),
.B(n_119),
.Y(n_171)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_139),
.B(n_111),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_157),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_175),
.A2(n_177),
.B1(n_178),
.B2(n_182),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_147),
.B(n_117),
.Y(n_176)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_176),
.Y(n_208)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_179),
.A2(n_183),
.B1(n_154),
.B2(n_150),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_134),
.B(n_124),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_180),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_143),
.B(n_82),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_181),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_151),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_146),
.A2(n_66),
.B1(n_82),
.B2(n_115),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_181),
.Y(n_186)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_148),
.C(n_145),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_198),
.C(n_204),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_189),
.B(n_195),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_190),
.A2(n_203),
.B1(n_173),
.B2(n_172),
.Y(n_223)
);

NAND3xp33_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_150),
.C(n_151),
.Y(n_193)
);

NAND3xp33_ASAP7_75t_SL g228 ( 
.A(n_193),
.B(n_0),
.C(n_1),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_179),
.A2(n_149),
.B1(n_150),
.B2(n_156),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_194),
.A2(n_168),
.B1(n_162),
.B2(n_171),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_166),
.B(n_144),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_184),
.Y(n_196)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_196),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_150),
.C(n_152),
.Y(n_198)
);

AO22x1_ASAP7_75t_SL g200 ( 
.A1(n_161),
.A2(n_153),
.B1(n_136),
.B2(n_138),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_200),
.A2(n_176),
.B(n_163),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_183),
.A2(n_138),
.B1(n_49),
.B2(n_56),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_175),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_165),
.A2(n_63),
.B1(n_54),
.B2(n_50),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_44),
.C(n_54),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_167),
.B(n_44),
.C(n_50),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_164),
.Y(n_221)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_209),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_177),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_219),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_200),
.A2(n_178),
.B1(n_173),
.B2(n_180),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_212),
.A2(n_216),
.B1(n_225),
.B2(n_205),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_213),
.A2(n_188),
.B(n_198),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_192),
.B(n_159),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_217),
.B(n_218),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_191),
.B(n_159),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_169),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_204),
.C(n_199),
.Y(n_229)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_224),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_223),
.A2(n_22),
.B1(n_29),
.B2(n_19),
.Y(n_245)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_194),
.A2(n_84),
.B1(n_1),
.B2(n_2),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_200),
.Y(n_226)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_226),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_84),
.Y(n_227)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

NAND2xp33_ASAP7_75t_SL g232 ( 
.A(n_228),
.B(n_13),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_237),
.C(n_239),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_215),
.A2(n_196),
.B1(n_190),
.B2(n_208),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_230),
.A2(n_243),
.B1(n_236),
.B2(n_235),
.Y(n_249)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_216),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_220),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_212),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_234),
.A2(n_244),
.B1(n_245),
.B2(n_225),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_219),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_187),
.C(n_207),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_186),
.C(n_185),
.Y(n_239)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_226),
.Y(n_243)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_243),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_213),
.A2(n_185),
.B(n_203),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_22),
.C(n_16),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_29),
.C(n_19),
.Y(n_260)
);

AOI221xp5_ASAP7_75t_L g273 ( 
.A1(n_247),
.A2(n_9),
.B1(n_13),
.B2(n_12),
.C(n_6),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_249),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_251),
.B(n_252),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_231),
.A2(n_220),
.B1(n_214),
.B2(n_210),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_244),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_256),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_241),
.B(n_11),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_255),
.A2(n_259),
.B(n_9),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_11),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_29),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_260),
.C(n_261),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_234),
.A2(n_10),
.B1(n_14),
.B2(n_13),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_258),
.A2(n_245),
.B1(n_242),
.B2(n_246),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_2),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_16),
.C(n_29),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_262),
.A2(n_271),
.B(n_274),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_242),
.Y(n_264)
);

FAx1_ASAP7_75t_SL g283 ( 
.A(n_264),
.B(n_267),
.CI(n_6),
.CON(n_283),
.SN(n_283)
);

NOR3xp33_ASAP7_75t_SL g267 ( 
.A(n_253),
.B(n_238),
.C(n_229),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_270),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_250),
.A2(n_237),
.B1(n_10),
.B2(n_12),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_19),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_6),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_273),
.A2(n_8),
.B(n_9),
.Y(n_284)
);

MAJx2_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_8),
.C(n_10),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_262),
.A2(n_266),
.B1(n_264),
.B2(n_267),
.Y(n_275)
);

A2O1A1Ixp33_ASAP7_75t_SL g289 ( 
.A1(n_275),
.A2(n_274),
.B(n_8),
.C(n_4),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_248),
.C(n_261),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_277),
.C(n_279),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_260),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_281),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_269),
.A2(n_2),
.B(n_3),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_3),
.C(n_4),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_284),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_280),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_285),
.B(n_283),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_266),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_288),
.A2(n_289),
.B(n_286),
.Y(n_293)
);

INVxp33_ASAP7_75t_L g291 ( 
.A(n_282),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_3),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_292),
.A2(n_294),
.B(n_296),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_293),
.B(n_295),
.Y(n_298)
);

AOI332xp33_ASAP7_75t_L g294 ( 
.A1(n_289),
.A2(n_3),
.A3(n_4),
.B1(n_16),
.B2(n_275),
.B3(n_276),
.C1(n_277),
.C2(n_290),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_287),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_297),
.B(n_298),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_16),
.Y(n_300)
);


endmodule