module fake_netlist_6_4589_n_2505 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2505);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2505;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2382;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_2447;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_2495;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2394;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_2364;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_2496;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_2397;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_2455;
wire n_558;
wire n_2469;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_2459;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_2434;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2453;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1886;
wire n_1801;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_2467;
wire n_2468;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_2476;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_437;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_295;
wire n_701;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2411;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_1052;
wire n_462;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_2391;
wire n_304;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_673;
wire n_382;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_2436;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2407;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2501;
wire n_2238;
wire n_293;
wire n_2368;
wire n_458;
wire n_1070;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_1395;
wire n_2199;
wire n_2110;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_474;
wire n_683;
wire n_1207;
wire n_811;
wire n_2442;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_2432;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_2475;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_2416;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2357;
wire n_2025;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_2410;
wire n_1053;
wire n_2374;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_2502;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_2289;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_2420;
wire n_575;
wire n_368;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2381;
wire n_2052;
wire n_1847;
wire n_248;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_2423;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_2499;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_2486;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_239;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_2376;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_2479;
wire n_1974;
wire n_2456;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_2406;
wire n_533;
wire n_2390;
wire n_806;
wire n_959;
wire n_879;
wire n_2310;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_2383;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_306;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_346;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1962;
wire n_1236;
wire n_1794;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_2400;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_400;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_1147;
wire n_763;
wire n_1785;
wire n_360;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1702;
wire n_1570;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2081;
wire n_2168;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_653;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_839;
wire n_2437;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_265;
wire n_1184;
wire n_2483;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1362;
wire n_1156;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_2334;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_240;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_2471;
wire n_467;
wire n_269;
wire n_973;
wire n_359;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2461;
wire n_2215;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_2477;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2185;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2415;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_336;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_62),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_150),
.Y(n_238)
);

BUFx2_ASAP7_75t_SL g239 ( 
.A(n_16),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_7),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_65),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_117),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_236),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_142),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_141),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_31),
.Y(n_246)
);

BUFx2_ASAP7_75t_SL g247 ( 
.A(n_57),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_192),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_182),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_220),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_41),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_41),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_73),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_37),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_108),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_110),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_171),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_101),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_71),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_79),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_47),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_178),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_1),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_85),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_147),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_40),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_8),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_43),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_34),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_122),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_126),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_217),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_157),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_47),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_46),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_204),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_209),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_196),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_16),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_189),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_136),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_133),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_106),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_9),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_167),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_218),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_159),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_69),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_172),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_115),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_123),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_82),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_166),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_168),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_54),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_154),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_174),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_131),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_1),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_72),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_203),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_29),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_190),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_195),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_137),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_222),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_183),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_78),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_42),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_191),
.Y(n_310)
);

BUFx5_ASAP7_75t_L g311 ( 
.A(n_33),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_66),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_129),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_148),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_109),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_179),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_12),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_88),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_98),
.Y(n_319)
);

INVx2_ASAP7_75t_SL g320 ( 
.A(n_146),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_69),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_37),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_45),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_215),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_185),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_71),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_31),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_160),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_156),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_73),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_9),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_180),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_26),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_100),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_33),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_199),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_197),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_2),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_130),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_226),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_124),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_173),
.Y(n_342)
);

BUFx10_ASAP7_75t_L g343 ( 
.A(n_223),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_144),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_92),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_87),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_20),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_132),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_20),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_110),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_61),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_193),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_26),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_90),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_120),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_85),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_231),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_91),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_118),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_233),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_59),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_98),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_177),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_44),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_162),
.Y(n_365)
);

INVx2_ASAP7_75t_SL g366 ( 
.A(n_187),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_158),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_46),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_139),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_97),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_155),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_164),
.Y(n_372)
);

BUFx10_ASAP7_75t_L g373 ( 
.A(n_60),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_184),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_87),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_224),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_21),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_0),
.Y(n_378)
);

CKINVDCx14_ASAP7_75t_R g379 ( 
.A(n_5),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_225),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_107),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_39),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_127),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_52),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_109),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_119),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_4),
.Y(n_387)
);

INVx2_ASAP7_75t_SL g388 ( 
.A(n_205),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_94),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_43),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_163),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_210),
.Y(n_392)
);

CKINVDCx14_ASAP7_75t_R g393 ( 
.A(n_93),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_104),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_175),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_63),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_219),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_213),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_106),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_57),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_104),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_113),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_111),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_116),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_22),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_181),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_55),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_93),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_128),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_149),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_54),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_27),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_114),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_78),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_208),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_29),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_95),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_151),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_114),
.Y(n_419)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_198),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_214),
.Y(n_421)
);

BUFx5_ASAP7_75t_L g422 ( 
.A(n_200),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_81),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_140),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_13),
.Y(n_425)
);

INVx2_ASAP7_75t_SL g426 ( 
.A(n_169),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_30),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_227),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_119),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_118),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_81),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_88),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_60),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_15),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_202),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_112),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_59),
.Y(n_437)
);

CKINVDCx14_ASAP7_75t_R g438 ( 
.A(n_176),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_125),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_25),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_65),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_188),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_212),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_115),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_5),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_72),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_111),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_19),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_22),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_145),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_152),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_63),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_194),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_103),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_23),
.Y(n_455)
);

INVxp33_ASAP7_75t_SL g456 ( 
.A(n_116),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_77),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_40),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_11),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_64),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_4),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_108),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_67),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_113),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_311),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_243),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_432),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_432),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_311),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_311),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_374),
.B(n_0),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_257),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_423),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_262),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_423),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_311),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_265),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_280),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_270),
.Y(n_479)
);

INVxp67_ASAP7_75t_SL g480 ( 
.A(n_374),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_311),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_239),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_311),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_311),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_272),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_311),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_311),
.Y(n_487)
);

INVxp67_ASAP7_75t_SL g488 ( 
.A(n_282),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_311),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_287),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_463),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_463),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_276),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_414),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_463),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_263),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_463),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_277),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_282),
.B(n_2),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_239),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_310),
.Y(n_501)
);

BUFx5_ASAP7_75t_L g502 ( 
.A(n_244),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_463),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_289),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_291),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_463),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_297),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_409),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_414),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_414),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_338),
.B(n_3),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_298),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_303),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_304),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_428),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_451),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_285),
.B(n_3),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_281),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_314),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_281),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_414),
.Y(n_521)
);

INVxp67_ASAP7_75t_SL g522 ( 
.A(n_285),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_247),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_249),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_252),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_249),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_251),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_251),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_324),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_251),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_336),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_339),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_318),
.Y(n_533)
);

INVxp33_ASAP7_75t_SL g534 ( 
.A(n_237),
.Y(n_534)
);

INVxp67_ASAP7_75t_SL g535 ( 
.A(n_325),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_341),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_318),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_273),
.Y(n_538)
);

CKINVDCx16_ASAP7_75t_R g539 ( 
.A(n_252),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_318),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_344),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_407),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_348),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_352),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_273),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_407),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_438),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_407),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_325),
.B(n_6),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_379),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_357),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_379),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_434),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_360),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_250),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g556 ( 
.A(n_247),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_369),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_434),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_371),
.Y(n_559)
);

INVxp67_ASAP7_75t_L g560 ( 
.A(n_246),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_393),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_393),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_372),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_434),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_263),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_376),
.Y(n_566)
);

INVxp67_ASAP7_75t_SL g567 ( 
.A(n_250),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_380),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_406),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_435),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_263),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_284),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_284),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_284),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_442),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_453),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_350),
.Y(n_577)
);

NOR2xp67_ASAP7_75t_L g578 ( 
.A(n_242),
.B(n_6),
.Y(n_578)
);

INVxp67_ASAP7_75t_L g579 ( 
.A(n_246),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_350),
.Y(n_580)
);

CKINVDCx16_ASAP7_75t_R g581 ( 
.A(n_322),
.Y(n_581)
);

BUFx6f_ASAP7_75t_SL g582 ( 
.A(n_343),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_240),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_267),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_241),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_350),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_425),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_425),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_250),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_253),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_425),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_320),
.B(n_7),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_491),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_527),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_491),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_492),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_492),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_466),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_495),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_465),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_567),
.B(n_320),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_495),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_497),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_497),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_472),
.Y(n_605)
);

INVx1_ASAP7_75t_SL g606 ( 
.A(n_550),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_474),
.Y(n_607)
);

OR2x2_ASAP7_75t_L g608 ( 
.A(n_496),
.B(n_322),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_477),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_479),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_SL g611 ( 
.A(n_552),
.B(n_353),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_503),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_527),
.Y(n_613)
);

INVxp67_ASAP7_75t_L g614 ( 
.A(n_525),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_503),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_518),
.B(n_343),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_506),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_478),
.Y(n_618)
);

AND3x2_ASAP7_75t_L g619 ( 
.A(n_499),
.B(n_242),
.C(n_286),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_506),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_465),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_555),
.B(n_320),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_555),
.B(n_366),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_469),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_565),
.B(n_366),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_490),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_555),
.B(n_366),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_530),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_530),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_485),
.Y(n_630)
);

INVxp67_ASAP7_75t_L g631 ( 
.A(n_496),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_493),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_565),
.B(n_388),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_494),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_469),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_498),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_494),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_509),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_509),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_510),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_470),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_504),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_505),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_510),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_470),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_476),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_555),
.B(n_388),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_476),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_521),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_507),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_555),
.B(n_388),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_501),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_512),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_513),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_521),
.Y(n_655)
);

BUFx2_ASAP7_75t_L g656 ( 
.A(n_561),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_481),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_520),
.B(n_343),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_514),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_519),
.Y(n_660)
);

BUFx2_ASAP7_75t_L g661 ( 
.A(n_562),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_481),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_511),
.B(n_343),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_571),
.B(n_426),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_483),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_589),
.B(n_426),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_529),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_483),
.Y(n_668)
);

CKINVDCx20_ASAP7_75t_R g669 ( 
.A(n_508),
.Y(n_669)
);

INVx4_ASAP7_75t_L g670 ( 
.A(n_589),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_515),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_531),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_484),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_532),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_536),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_484),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_541),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_486),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_589),
.B(n_426),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_486),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_543),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_487),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_544),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_551),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_487),
.Y(n_685)
);

NAND2xp33_ASAP7_75t_SL g686 ( 
.A(n_592),
.B(n_295),
.Y(n_686)
);

CKINVDCx20_ASAP7_75t_R g687 ( 
.A(n_516),
.Y(n_687)
);

CKINVDCx20_ASAP7_75t_R g688 ( 
.A(n_547),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_489),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_489),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_657),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_606),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_601),
.B(n_554),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_657),
.Y(n_694)
);

INVx1_ASAP7_75t_SL g695 ( 
.A(n_606),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_665),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_593),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_631),
.B(n_557),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_600),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_601),
.B(n_591),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_601),
.B(n_559),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_665),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_668),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_688),
.Y(n_704)
);

AND2x6_ASAP7_75t_L g705 ( 
.A(n_625),
.B(n_286),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_609),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_668),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_625),
.B(n_589),
.Y(n_708)
);

INVxp67_ASAP7_75t_L g709 ( 
.A(n_611),
.Y(n_709)
);

OR2x2_ASAP7_75t_SL g710 ( 
.A(n_608),
.B(n_539),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_625),
.B(n_591),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_673),
.Y(n_712)
);

OR2x2_ASAP7_75t_L g713 ( 
.A(n_608),
.B(n_581),
.Y(n_713)
);

INVx4_ASAP7_75t_L g714 ( 
.A(n_670),
.Y(n_714)
);

OR2x2_ASAP7_75t_L g715 ( 
.A(n_608),
.B(n_475),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_673),
.B(n_566),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_631),
.B(n_475),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_678),
.B(n_568),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_663),
.A2(n_480),
.B1(n_522),
.B2(n_488),
.Y(n_719)
);

INVxp67_ASAP7_75t_L g720 ( 
.A(n_611),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_593),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_593),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_618),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_SL g724 ( 
.A(n_598),
.B(n_524),
.Y(n_724)
);

AND2x4_ASAP7_75t_L g725 ( 
.A(n_633),
.B(n_589),
.Y(n_725)
);

INVx4_ASAP7_75t_L g726 ( 
.A(n_670),
.Y(n_726)
);

BUFx4f_ASAP7_75t_L g727 ( 
.A(n_600),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_678),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_682),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_682),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_600),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_600),
.Y(n_732)
);

AND2x2_ASAP7_75t_SL g733 ( 
.A(n_670),
.B(n_286),
.Y(n_733)
);

BUFx10_ASAP7_75t_L g734 ( 
.A(n_605),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_633),
.B(n_664),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_690),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_690),
.B(n_569),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_624),
.Y(n_738)
);

INVxp67_ASAP7_75t_L g739 ( 
.A(n_656),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_595),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_635),
.B(n_570),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_600),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_595),
.Y(n_743)
);

INVx4_ASAP7_75t_L g744 ( 
.A(n_670),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_663),
.B(n_534),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_633),
.B(n_244),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_595),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_612),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_619),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_624),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_607),
.B(n_575),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_610),
.B(n_576),
.Y(n_752)
);

OR2x2_ASAP7_75t_L g753 ( 
.A(n_614),
.B(n_473),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_624),
.Y(n_754)
);

HB1xp67_ASAP7_75t_L g755 ( 
.A(n_614),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_612),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_646),
.Y(n_757)
);

NAND3xp33_ASAP7_75t_L g758 ( 
.A(n_686),
.B(n_549),
.C(n_517),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_646),
.Y(n_759)
);

AND2x2_ASAP7_75t_SL g760 ( 
.A(n_622),
.B(n_363),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_600),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_646),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_676),
.Y(n_763)
);

NAND2xp33_ASAP7_75t_L g764 ( 
.A(n_664),
.B(n_583),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_612),
.Y(n_765)
);

OAI22xp33_ASAP7_75t_SL g766 ( 
.A1(n_616),
.A2(n_535),
.B1(n_471),
.B2(n_467),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_630),
.B(n_585),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_635),
.B(n_590),
.Y(n_768)
);

INVx1_ASAP7_75t_SL g769 ( 
.A(n_626),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_632),
.B(n_563),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_676),
.Y(n_771)
);

BUFx3_ASAP7_75t_L g772 ( 
.A(n_635),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_635),
.B(n_502),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_664),
.B(n_245),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_636),
.B(n_482),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_638),
.B(n_245),
.Y(n_776)
);

BUFx2_ASAP7_75t_L g777 ( 
.A(n_656),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_638),
.B(n_571),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_642),
.B(n_582),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_652),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_676),
.B(n_502),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_619),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_600),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_680),
.B(n_685),
.Y(n_784)
);

AND2x6_ASAP7_75t_L g785 ( 
.A(n_680),
.B(n_363),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_643),
.B(n_500),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_615),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_621),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_680),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_621),
.Y(n_790)
);

AND2x6_ASAP7_75t_L g791 ( 
.A(n_685),
.B(n_363),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_685),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_615),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_596),
.Y(n_794)
);

AND2x2_ASAP7_75t_SL g795 ( 
.A(n_622),
.B(n_418),
.Y(n_795)
);

INVx5_ASAP7_75t_L g796 ( 
.A(n_621),
.Y(n_796)
);

BUFx8_ASAP7_75t_SL g797 ( 
.A(n_669),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_SL g798 ( 
.A(n_650),
.B(n_526),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_596),
.Y(n_799)
);

XOR2xp5_ASAP7_75t_L g800 ( 
.A(n_671),
.B(n_584),
.Y(n_800)
);

INVxp67_ASAP7_75t_SL g801 ( 
.A(n_623),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_653),
.B(n_654),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_621),
.B(n_502),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_597),
.Y(n_804)
);

OAI21xp33_ASAP7_75t_L g805 ( 
.A1(n_658),
.A2(n_556),
.B(n_523),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_597),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_599),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_R g808 ( 
.A(n_659),
.B(n_538),
.Y(n_808)
);

AO22x2_ASAP7_75t_L g809 ( 
.A1(n_623),
.A2(n_418),
.B1(n_450),
.B2(n_433),
.Y(n_809)
);

INVx4_ASAP7_75t_L g810 ( 
.A(n_621),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_615),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_639),
.B(n_572),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_599),
.Y(n_813)
);

INVx2_ASAP7_75t_SL g814 ( 
.A(n_627),
.Y(n_814)
);

BUFx6f_ASAP7_75t_L g815 ( 
.A(n_621),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_602),
.Y(n_816)
);

INVx3_ASAP7_75t_L g817 ( 
.A(n_621),
.Y(n_817)
);

AND2x4_ASAP7_75t_L g818 ( 
.A(n_639),
.B(n_640),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_641),
.Y(n_819)
);

CKINVDCx16_ASAP7_75t_R g820 ( 
.A(n_687),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_641),
.B(n_645),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_640),
.B(n_572),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_660),
.B(n_582),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_602),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_667),
.B(n_582),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_603),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_672),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_641),
.Y(n_828)
);

CKINVDCx16_ASAP7_75t_R g829 ( 
.A(n_661),
.Y(n_829)
);

INVx1_ASAP7_75t_SL g830 ( 
.A(n_661),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_641),
.B(n_502),
.Y(n_831)
);

BUFx4f_ASAP7_75t_L g832 ( 
.A(n_641),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_674),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_603),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_604),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_604),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_675),
.B(n_545),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_641),
.B(n_502),
.Y(n_838)
);

AND2x6_ASAP7_75t_L g839 ( 
.A(n_641),
.B(n_418),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_617),
.Y(n_840)
);

HB1xp67_ASAP7_75t_L g841 ( 
.A(n_644),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_617),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_620),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_644),
.A2(n_468),
.B1(n_502),
.B2(n_274),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_645),
.B(n_502),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_645),
.B(n_648),
.Y(n_846)
);

NAND2xp33_ASAP7_75t_SL g847 ( 
.A(n_677),
.B(n_355),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_649),
.B(n_573),
.Y(n_848)
);

HB1xp67_ASAP7_75t_L g849 ( 
.A(n_649),
.Y(n_849)
);

BUFx3_ASAP7_75t_L g850 ( 
.A(n_645),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_645),
.B(n_502),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_655),
.B(n_573),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_L g853 ( 
.A1(n_733),
.A2(n_814),
.B1(n_693),
.B2(n_701),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_691),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_691),
.Y(n_855)
);

OR2x2_ASAP7_75t_L g856 ( 
.A(n_717),
.B(n_681),
.Y(n_856)
);

NOR3x1_ASAP7_75t_L g857 ( 
.A(n_758),
.B(n_274),
.C(n_261),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_694),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_826),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_814),
.B(n_645),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_826),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_694),
.Y(n_862)
);

OR2x6_ASAP7_75t_L g863 ( 
.A(n_749),
.B(n_450),
.Y(n_863)
);

HB1xp67_ASAP7_75t_L g864 ( 
.A(n_749),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_801),
.B(n_645),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_772),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_745),
.B(n_683),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_809),
.A2(n_456),
.B1(n_578),
.B2(n_627),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_716),
.B(n_684),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_733),
.B(n_648),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_696),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_718),
.B(n_737),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_733),
.B(n_648),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_735),
.B(n_648),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_834),
.Y(n_875)
);

INVxp67_ASAP7_75t_L g876 ( 
.A(n_755),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_752),
.B(n_238),
.Y(n_877)
);

AND2x6_ASAP7_75t_SL g878 ( 
.A(n_837),
.B(n_261),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_696),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_767),
.B(n_238),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_735),
.B(n_648),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_729),
.B(n_648),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_834),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_729),
.B(n_648),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_782),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_730),
.B(n_662),
.Y(n_886)
);

OAI22xp5_ASAP7_75t_L g887 ( 
.A1(n_760),
.A2(n_398),
.B1(n_415),
.B2(n_278),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_702),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_708),
.B(n_248),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_760),
.A2(n_502),
.B1(n_450),
.B2(n_271),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_SL g891 ( 
.A1(n_766),
.A2(n_384),
.B1(n_436),
.B2(n_377),
.Y(n_891)
);

BUFx8_ASAP7_75t_L g892 ( 
.A(n_777),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_842),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_730),
.B(n_662),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_842),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_702),
.B(n_662),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_703),
.B(n_662),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_703),
.B(n_662),
.Y(n_898)
);

INVxp67_ASAP7_75t_L g899 ( 
.A(n_753),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_719),
.B(n_278),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_707),
.B(n_662),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_SL g902 ( 
.A(n_827),
.B(n_461),
.Y(n_902)
);

AOI22xp33_ASAP7_75t_L g903 ( 
.A1(n_760),
.A2(n_271),
.B1(n_293),
.B2(n_248),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_707),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_712),
.B(n_728),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_712),
.B(n_662),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_728),
.B(n_689),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_700),
.B(n_655),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_768),
.B(n_398),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_736),
.Y(n_910)
);

INVx5_ASAP7_75t_L g911 ( 
.A(n_839),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_700),
.B(n_574),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_736),
.B(n_689),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_794),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_809),
.A2(n_651),
.B1(n_666),
.B2(n_647),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_708),
.B(n_689),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_772),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_782),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_818),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_794),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_711),
.B(n_574),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_741),
.B(n_415),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_698),
.B(n_420),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_708),
.B(n_689),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_708),
.B(n_689),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_711),
.B(n_577),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_725),
.B(n_420),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_818),
.Y(n_928)
);

BUFx2_ASAP7_75t_L g929 ( 
.A(n_777),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_818),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_725),
.B(n_293),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_746),
.B(n_577),
.Y(n_932)
);

AND2x4_ASAP7_75t_SL g933 ( 
.A(n_734),
.B(n_373),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_805),
.B(n_353),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_799),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_818),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_821),
.A2(n_651),
.B(n_647),
.Y(n_937)
);

BUFx3_ASAP7_75t_L g938 ( 
.A(n_725),
.Y(n_938)
);

INVxp67_ASAP7_75t_SL g939 ( 
.A(n_699),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_753),
.B(n_433),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_779),
.B(n_294),
.Y(n_941)
);

INVx5_ASAP7_75t_L g942 ( 
.A(n_839),
.Y(n_942)
);

AND2x6_ASAP7_75t_SL g943 ( 
.A(n_770),
.B(n_279),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_799),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_804),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_797),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_804),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_746),
.B(n_580),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_795),
.B(n_689),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_808),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_795),
.B(n_666),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_795),
.B(n_679),
.Y(n_952)
);

NOR2xp67_ASAP7_75t_L g953 ( 
.A(n_714),
.B(n_679),
.Y(n_953)
);

INVx4_ASAP7_75t_L g954 ( 
.A(n_714),
.Y(n_954)
);

AOI22xp33_ASAP7_75t_L g955 ( 
.A1(n_705),
.A2(n_296),
.B1(n_301),
.B2(n_294),
.Y(n_955)
);

AOI22xp33_ASAP7_75t_L g956 ( 
.A1(n_705),
.A2(n_746),
.B1(n_774),
.B2(n_809),
.Y(n_956)
);

BUFx3_ASAP7_75t_L g957 ( 
.A(n_734),
.Y(n_957)
);

AND2x6_ASAP7_75t_SL g958 ( 
.A(n_802),
.B(n_279),
.Y(n_958)
);

INVxp67_ASAP7_75t_L g959 ( 
.A(n_717),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_R g960 ( 
.A(n_827),
.B(n_254),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_746),
.A2(n_301),
.B(n_305),
.C(n_296),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_774),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_823),
.B(n_305),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_806),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_774),
.B(n_620),
.Y(n_965)
);

NAND2x1_ASAP7_75t_L g966 ( 
.A(n_714),
.B(n_634),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_774),
.B(n_634),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_806),
.B(n_637),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_807),
.B(n_637),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_807),
.B(n_813),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_709),
.B(n_457),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_809),
.A2(n_307),
.B1(n_313),
.B2(n_306),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_778),
.B(n_580),
.Y(n_973)
);

INVx8_ASAP7_75t_L g974 ( 
.A(n_705),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_720),
.B(n_457),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_825),
.B(n_306),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_813),
.B(n_628),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_816),
.B(n_628),
.Y(n_978)
);

AOI22xp33_ASAP7_75t_L g979 ( 
.A1(n_705),
.A2(n_313),
.B1(n_316),
.B2(n_307),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_846),
.A2(n_629),
.B(n_613),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_816),
.B(n_629),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_824),
.B(n_835),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_824),
.Y(n_983)
);

INVxp67_ASAP7_75t_L g984 ( 
.A(n_715),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_835),
.B(n_316),
.Y(n_985)
);

AOI22x1_ASAP7_75t_L g986 ( 
.A1(n_776),
.A2(n_329),
.B1(n_332),
.B2(n_328),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_699),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_836),
.B(n_328),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_836),
.B(n_329),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_840),
.B(n_332),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_840),
.Y(n_991)
);

AOI22xp33_ASAP7_75t_L g992 ( 
.A1(n_705),
.A2(n_340),
.B1(n_342),
.B2(n_337),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_843),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_843),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_738),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_775),
.B(n_255),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_705),
.B(n_337),
.Y(n_997)
);

INVx8_ASAP7_75t_L g998 ( 
.A(n_839),
.Y(n_998)
);

INVx4_ASAP7_75t_L g999 ( 
.A(n_726),
.Y(n_999)
);

INVx4_ASAP7_75t_L g1000 ( 
.A(n_726),
.Y(n_1000)
);

NOR3xp33_ASAP7_75t_SL g1001 ( 
.A(n_829),
.B(n_258),
.C(n_256),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_841),
.B(n_340),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_849),
.B(n_342),
.Y(n_1003)
);

INVxp67_ASAP7_75t_L g1004 ( 
.A(n_715),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_697),
.Y(n_1005)
);

NOR3xp33_ASAP7_75t_L g1006 ( 
.A(n_847),
.B(n_579),
.C(n_560),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_734),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_713),
.B(n_365),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_778),
.B(n_586),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_738),
.Y(n_1010)
);

OAI22xp33_ASAP7_75t_L g1011 ( 
.A1(n_713),
.A2(n_798),
.B1(n_724),
.B2(n_367),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_844),
.B(n_786),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_751),
.B(n_259),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_750),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_776),
.B(n_365),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_833),
.B(n_367),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_697),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_750),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_SL g1019 ( 
.A(n_833),
.B(n_373),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_812),
.B(n_586),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_776),
.B(n_383),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_721),
.Y(n_1022)
);

AND2x6_ASAP7_75t_SL g1023 ( 
.A(n_800),
.B(n_283),
.Y(n_1023)
);

INVxp67_ASAP7_75t_L g1024 ( 
.A(n_800),
.Y(n_1024)
);

INVx1_ASAP7_75t_SL g1025 ( 
.A(n_929),
.Y(n_1025)
);

INVx1_ASAP7_75t_SL g1026 ( 
.A(n_929),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_872),
.B(n_764),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_877),
.B(n_692),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_880),
.B(n_695),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_904),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_869),
.B(n_706),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_870),
.A2(n_710),
.B1(n_739),
.B2(n_727),
.Y(n_1032)
);

AO22x1_ASAP7_75t_L g1033 ( 
.A1(n_857),
.A2(n_776),
.B1(n_391),
.B2(n_392),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_904),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_995),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_914),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_R g1037 ( 
.A(n_950),
.B(n_723),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_914),
.Y(n_1038)
);

NAND2x1p5_ASAP7_75t_L g1039 ( 
.A(n_911),
.B(n_726),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_892),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_899),
.B(n_769),
.Y(n_1041)
);

INVx3_ASAP7_75t_L g1042 ( 
.A(n_866),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_995),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_912),
.B(n_812),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_853),
.B(n_822),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_923),
.A2(n_744),
.B1(n_848),
.B2(n_822),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_920),
.Y(n_1047)
);

NOR3xp33_ASAP7_75t_SL g1048 ( 
.A(n_1011),
.B(n_829),
.C(n_780),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1010),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_854),
.B(n_848),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_912),
.B(n_852),
.Y(n_1051)
);

INVx3_ASAP7_75t_L g1052 ( 
.A(n_866),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1010),
.Y(n_1053)
);

O2A1O1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_887),
.A2(n_852),
.B(n_784),
.C(n_757),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_856),
.B(n_830),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_932),
.B(n_587),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1014),
.Y(n_1057)
);

INVx4_ASAP7_75t_L g1058 ( 
.A(n_974),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_920),
.Y(n_1059)
);

OAI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_919),
.A2(n_391),
.B1(n_392),
.B2(n_383),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_971),
.B(n_723),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1014),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_946),
.Y(n_1063)
);

AOI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_962),
.A2(n_791),
.B1(n_785),
.B2(n_757),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_946),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_935),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_975),
.B(n_780),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1018),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1018),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_935),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_854),
.B(n_744),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_R g1072 ( 
.A(n_950),
.B(n_704),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_866),
.Y(n_1073)
);

INVx3_ASAP7_75t_L g1074 ( 
.A(n_938),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_876),
.B(n_820),
.Y(n_1075)
);

BUFx2_ASAP7_75t_L g1076 ( 
.A(n_892),
.Y(n_1076)
);

BUFx4f_ASAP7_75t_L g1077 ( 
.A(n_917),
.Y(n_1077)
);

INVx5_ASAP7_75t_L g1078 ( 
.A(n_974),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_R g1079 ( 
.A(n_957),
.B(n_704),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_945),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_855),
.B(n_744),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_957),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_938),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_859),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_859),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_861),
.Y(n_1086)
);

BUFx10_ASAP7_75t_L g1087 ( 
.A(n_940),
.Y(n_1087)
);

INVx2_ASAP7_75t_SL g1088 ( 
.A(n_908),
.Y(n_1088)
);

NOR3xp33_ASAP7_75t_SL g1089 ( 
.A(n_1016),
.B(n_264),
.C(n_260),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_919),
.B(n_783),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_974),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_861),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_SL g1093 ( 
.A1(n_891),
.A2(n_820),
.B1(n_710),
.B2(n_268),
.Y(n_1093)
);

NOR3xp33_ASAP7_75t_SL g1094 ( 
.A(n_1008),
.B(n_269),
.C(n_266),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_875),
.Y(n_1095)
);

AOI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_962),
.A2(n_783),
.B1(n_850),
.B2(n_788),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_945),
.Y(n_1097)
);

BUFx2_ASAP7_75t_L g1098 ( 
.A(n_892),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_947),
.Y(n_1099)
);

AND3x1_ASAP7_75t_SL g1100 ( 
.A(n_958),
.B(n_288),
.C(n_283),
.Y(n_1100)
);

AOI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_928),
.A2(n_791),
.B1(n_785),
.B2(n_759),
.Y(n_1101)
);

BUFx2_ASAP7_75t_L g1102 ( 
.A(n_892),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_917),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_875),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_883),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_855),
.B(n_754),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_974),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_858),
.B(n_754),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_947),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_867),
.B(n_810),
.Y(n_1110)
);

INVxp67_ASAP7_75t_SL g1111 ( 
.A(n_917),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_974),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_883),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_893),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_893),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_928),
.B(n_788),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_856),
.B(n_727),
.Y(n_1117)
);

AOI22xp33_ASAP7_75t_L g1118 ( 
.A1(n_903),
.A2(n_762),
.B1(n_763),
.B2(n_759),
.Y(n_1118)
);

O2A1O1Ixp33_ASAP7_75t_SL g1119 ( 
.A1(n_961),
.A2(n_773),
.B(n_397),
.C(n_410),
.Y(n_1119)
);

BUFx3_ASAP7_75t_L g1120 ( 
.A(n_1007),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_895),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_984),
.B(n_810),
.Y(n_1122)
);

AO221x1_ASAP7_75t_L g1123 ( 
.A1(n_1004),
.A2(n_351),
.B1(n_290),
.B2(n_315),
.C(n_321),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_994),
.Y(n_1124)
);

AOI22xp5_ASAP7_75t_SL g1125 ( 
.A1(n_1024),
.A2(n_292),
.B1(n_299),
.B2(n_275),
.Y(n_1125)
);

INVx8_ASAP7_75t_L g1126 ( 
.A(n_998),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_858),
.B(n_762),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_917),
.Y(n_1128)
);

INVxp67_ASAP7_75t_L g1129 ( 
.A(n_864),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_987),
.Y(n_1130)
);

INVx4_ASAP7_75t_L g1131 ( 
.A(n_987),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_930),
.B(n_850),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_895),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_930),
.B(n_727),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_994),
.Y(n_1135)
);

NAND2xp33_ASAP7_75t_L g1136 ( 
.A(n_873),
.B(n_839),
.Y(n_1136)
);

BUFx3_ASAP7_75t_L g1137 ( 
.A(n_1007),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_862),
.B(n_763),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_959),
.B(n_810),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_862),
.B(n_771),
.Y(n_1140)
);

NOR3xp33_ASAP7_75t_SL g1141 ( 
.A(n_934),
.B(n_302),
.C(n_300),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_871),
.B(n_879),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_932),
.B(n_587),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_871),
.B(n_771),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_R g1145 ( 
.A(n_902),
.B(n_732),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1005),
.Y(n_1146)
);

BUFx3_ASAP7_75t_L g1147 ( 
.A(n_917),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1005),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_936),
.B(n_832),
.Y(n_1149)
);

NOR3xp33_ASAP7_75t_SL g1150 ( 
.A(n_1003),
.B(n_309),
.C(n_308),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_879),
.B(n_789),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_987),
.Y(n_1152)
);

BUFx4_ASAP7_75t_SL g1153 ( 
.A(n_1023),
.Y(n_1153)
);

INVx4_ASAP7_75t_L g1154 ( 
.A(n_987),
.Y(n_1154)
);

CKINVDCx20_ASAP7_75t_R g1155 ( 
.A(n_960),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_885),
.B(n_732),
.Y(n_1156)
);

INVx4_ASAP7_75t_L g1157 ( 
.A(n_987),
.Y(n_1157)
);

HB1xp67_ASAP7_75t_L g1158 ( 
.A(n_918),
.Y(n_1158)
);

INVxp67_ASAP7_75t_L g1159 ( 
.A(n_996),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1017),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_1023),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_954),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1017),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_888),
.B(n_789),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1022),
.Y(n_1165)
);

AOI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_1012),
.A2(n_817),
.B1(n_819),
.B2(n_732),
.Y(n_1166)
);

OR2x6_ASAP7_75t_L g1167 ( 
.A(n_998),
.B(n_395),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1022),
.Y(n_1168)
);

OR2x2_ASAP7_75t_L g1169 ( 
.A(n_863),
.B(n_588),
.Y(n_1169)
);

AND2x4_ASAP7_75t_L g1170 ( 
.A(n_936),
.B(n_395),
.Y(n_1170)
);

NOR2xp67_ASAP7_75t_L g1171 ( 
.A(n_954),
.B(n_817),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_888),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_1013),
.B(n_832),
.Y(n_1173)
);

INVxp67_ASAP7_75t_SL g1174 ( 
.A(n_939),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_909),
.B(n_817),
.Y(n_1175)
);

INVx5_ASAP7_75t_L g1176 ( 
.A(n_998),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_R g1177 ( 
.A(n_1019),
.B(n_910),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_908),
.Y(n_1178)
);

INVx2_ASAP7_75t_SL g1179 ( 
.A(n_973),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_948),
.B(n_397),
.Y(n_1180)
);

BUFx4f_ASAP7_75t_L g1181 ( 
.A(n_863),
.Y(n_1181)
);

INVx4_ASAP7_75t_L g1182 ( 
.A(n_954),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_878),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_910),
.B(n_792),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_944),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_944),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_948),
.Y(n_1187)
);

INVx3_ASAP7_75t_L g1188 ( 
.A(n_999),
.Y(n_1188)
);

INVxp67_ASAP7_75t_SL g1189 ( 
.A(n_860),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_964),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_964),
.B(n_792),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_983),
.B(n_819),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_983),
.Y(n_1193)
);

BUFx4f_ASAP7_75t_L g1194 ( 
.A(n_863),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_921),
.B(n_588),
.Y(n_1195)
);

NOR3xp33_ASAP7_75t_SL g1196 ( 
.A(n_941),
.B(n_317),
.C(n_312),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_878),
.Y(n_1197)
);

NOR3xp33_ASAP7_75t_SL g1198 ( 
.A(n_963),
.B(n_323),
.C(n_319),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_922),
.B(n_819),
.Y(n_1199)
);

AND2x4_ASAP7_75t_L g1200 ( 
.A(n_921),
.B(n_926),
.Y(n_1200)
);

NOR2x1_ASAP7_75t_L g1201 ( 
.A(n_999),
.B(n_781),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_SL g1202 ( 
.A(n_999),
.B(n_832),
.Y(n_1202)
);

INVx3_ASAP7_75t_L g1203 ( 
.A(n_1000),
.Y(n_1203)
);

A2O1A1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_874),
.A2(n_421),
.B(n_424),
.C(n_410),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_1000),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_926),
.B(n_421),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_991),
.B(n_699),
.Y(n_1207)
);

INVx4_ASAP7_75t_L g1208 ( 
.A(n_1000),
.Y(n_1208)
);

NOR2xp67_ASAP7_75t_L g1209 ( 
.A(n_915),
.B(n_803),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_973),
.B(n_699),
.Y(n_1210)
);

AND2x4_ASAP7_75t_L g1211 ( 
.A(n_1009),
.B(n_424),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1009),
.B(n_721),
.Y(n_1212)
);

INVx3_ASAP7_75t_L g1213 ( 
.A(n_966),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_998),
.Y(n_1214)
);

INVx4_ASAP7_75t_L g1215 ( 
.A(n_998),
.Y(n_1215)
);

NOR3xp33_ASAP7_75t_SL g1216 ( 
.A(n_976),
.B(n_327),
.C(n_326),
.Y(n_1216)
);

BUFx2_ASAP7_75t_L g1217 ( 
.A(n_863),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_991),
.B(n_699),
.Y(n_1218)
);

BUFx2_ASAP7_75t_L g1219 ( 
.A(n_889),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_993),
.B(n_731),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_1028),
.B(n_900),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_SL g1222 ( 
.A(n_1027),
.B(n_881),
.Y(n_1222)
);

AO21x1_ASAP7_75t_L g1223 ( 
.A1(n_1045),
.A2(n_972),
.B(n_868),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_1082),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_1130),
.Y(n_1225)
);

AOI21x1_ASAP7_75t_SL g1226 ( 
.A1(n_1211),
.A2(n_997),
.B(n_1015),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1200),
.A2(n_949),
.B1(n_952),
.B2(n_951),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1200),
.B(n_1020),
.Y(n_1228)
);

AND2x2_ASAP7_75t_SL g1229 ( 
.A(n_1181),
.B(n_972),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1200),
.B(n_1020),
.Y(n_1230)
);

AO31x2_ASAP7_75t_L g1231 ( 
.A1(n_1204),
.A2(n_1021),
.A3(n_993),
.B(n_937),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1213),
.A2(n_897),
.B(n_896),
.Y(n_1232)
);

NOR2x1_ASAP7_75t_L g1233 ( 
.A(n_1082),
.B(n_1120),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1044),
.B(n_905),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1044),
.B(n_970),
.Y(n_1235)
);

NAND2x1p5_ASAP7_75t_L g1236 ( 
.A(n_1078),
.B(n_1176),
.Y(n_1236)
);

OAI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1209),
.A2(n_956),
.B(n_865),
.Y(n_1237)
);

AO31x2_ASAP7_75t_L g1238 ( 
.A1(n_1172),
.A2(n_985),
.A3(n_989),
.B(n_988),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1051),
.B(n_982),
.Y(n_1239)
);

OAI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1209),
.A2(n_924),
.B(n_916),
.Y(n_1240)
);

OAI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1088),
.A2(n_868),
.B1(n_1002),
.B2(n_915),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1035),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1192),
.A2(n_901),
.B(n_898),
.Y(n_1243)
);

AO31x2_ASAP7_75t_L g1244 ( 
.A1(n_1172),
.A2(n_990),
.A3(n_907),
.B(n_913),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1207),
.A2(n_906),
.B(n_925),
.Y(n_1245)
);

OA22x2_ASAP7_75t_L g1246 ( 
.A1(n_1093),
.A2(n_933),
.B1(n_943),
.B2(n_958),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1218),
.A2(n_884),
.B(n_882),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_SL g1248 ( 
.A(n_1078),
.B(n_953),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1051),
.B(n_857),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1179),
.B(n_890),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1220),
.A2(n_894),
.B(n_886),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_1187),
.B(n_889),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1136),
.A2(n_965),
.B(n_967),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1213),
.A2(n_966),
.B(n_980),
.Y(n_1254)
);

BUFx3_ASAP7_75t_L g1255 ( 
.A(n_1120),
.Y(n_1255)
);

AOI221x1_ASAP7_75t_L g1256 ( 
.A1(n_1032),
.A2(n_1006),
.B1(n_977),
.B2(n_978),
.C(n_981),
.Y(n_1256)
);

CKINVDCx11_ASAP7_75t_R g1257 ( 
.A(n_1155),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1035),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1213),
.A2(n_969),
.B(n_968),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1039),
.A2(n_942),
.B(n_911),
.Y(n_1260)
);

AO31x2_ASAP7_75t_L g1261 ( 
.A1(n_1190),
.A2(n_443),
.A3(n_439),
.B(n_722),
.Y(n_1261)
);

O2A1O1Ixp5_ASAP7_75t_L g1262 ( 
.A1(n_1173),
.A2(n_931),
.B(n_889),
.C(n_927),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1039),
.A2(n_942),
.B(n_911),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1176),
.A2(n_942),
.B(n_911),
.Y(n_1264)
);

OR2x2_ASAP7_75t_L g1265 ( 
.A(n_1025),
.B(n_889),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1176),
.A2(n_942),
.B(n_911),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1179),
.B(n_931),
.Y(n_1267)
);

AO31x2_ASAP7_75t_L g1268 ( 
.A1(n_1190),
.A2(n_443),
.A3(n_439),
.B(n_722),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1088),
.B(n_931),
.Y(n_1269)
);

NAND3x1_ASAP7_75t_L g1270 ( 
.A(n_1061),
.B(n_290),
.C(n_288),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1201),
.A2(n_986),
.B(n_838),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1201),
.A2(n_986),
.B(n_845),
.Y(n_1272)
);

AOI221xp5_ASAP7_75t_L g1273 ( 
.A1(n_1067),
.A2(n_933),
.B1(n_349),
.B2(n_464),
.C(n_330),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1043),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1042),
.A2(n_851),
.B(n_831),
.Y(n_1275)
);

OAI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1142),
.A2(n_1046),
.B1(n_1186),
.B2(n_1185),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1176),
.A2(n_942),
.B(n_911),
.Y(n_1277)
);

OAI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1185),
.A2(n_979),
.B1(n_992),
.B2(n_955),
.Y(n_1278)
);

OA22x2_ASAP7_75t_L g1279 ( 
.A1(n_1159),
.A2(n_943),
.B1(n_333),
.B2(n_462),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_SL g1280 ( 
.A1(n_1193),
.A2(n_321),
.B(n_315),
.Y(n_1280)
);

AOI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1031),
.A2(n_1001),
.B1(n_839),
.B2(n_828),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1043),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1178),
.B(n_740),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1187),
.B(n_1219),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1042),
.A2(n_743),
.B(n_740),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1178),
.B(n_743),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_SL g1287 ( 
.A1(n_1193),
.A2(n_334),
.B(n_333),
.Y(n_1287)
);

OR2x2_ASAP7_75t_L g1288 ( 
.A(n_1026),
.B(n_528),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1195),
.B(n_747),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1186),
.A2(n_731),
.B1(n_828),
.B2(n_815),
.Y(n_1290)
);

INVxp67_ASAP7_75t_L g1291 ( 
.A(n_1158),
.Y(n_1291)
);

INVx6_ASAP7_75t_SL g1292 ( 
.A(n_1167),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1049),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1049),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1195),
.B(n_747),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1134),
.A2(n_756),
.B(n_748),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1056),
.B(n_748),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1149),
.A2(n_765),
.B(n_756),
.Y(n_1298)
);

BUFx2_ASAP7_75t_L g1299 ( 
.A(n_1079),
.Y(n_1299)
);

OA21x2_ASAP7_75t_L g1300 ( 
.A1(n_1053),
.A2(n_787),
.B(n_765),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1078),
.A2(n_742),
.B(n_731),
.Y(n_1301)
);

A2O1A1Ixp33_ASAP7_75t_L g1302 ( 
.A1(n_1050),
.A2(n_386),
.B(n_347),
.C(n_462),
.Y(n_1302)
);

NOR2xp67_ASAP7_75t_L g1303 ( 
.A(n_1063),
.B(n_121),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1056),
.B(n_787),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1219),
.A2(n_731),
.B1(n_828),
.B2(n_815),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1143),
.B(n_793),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1053),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1078),
.A2(n_742),
.B(n_731),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_1130),
.Y(n_1309)
);

AND2x4_ASAP7_75t_L g1310 ( 
.A(n_1074),
.B(n_742),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1143),
.B(n_793),
.Y(n_1311)
);

INVx3_ASAP7_75t_L g1312 ( 
.A(n_1182),
.Y(n_1312)
);

AO32x2_ASAP7_75t_L g1313 ( 
.A1(n_1131),
.A2(n_785),
.A3(n_791),
.B1(n_419),
.B2(n_460),
.Y(n_1313)
);

AO31x2_ASAP7_75t_L g1314 ( 
.A1(n_1057),
.A2(n_811),
.A3(n_455),
.B(n_454),
.Y(n_1314)
);

CKINVDCx11_ASAP7_75t_R g1315 ( 
.A(n_1155),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1042),
.A2(n_811),
.B(n_533),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1057),
.Y(n_1317)
);

AOI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1029),
.A2(n_839),
.B1(n_828),
.B2(n_815),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1212),
.A2(n_839),
.B(n_791),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1212),
.A2(n_1054),
.B(n_1189),
.Y(n_1320)
);

OAI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1166),
.A2(n_791),
.B(n_785),
.Y(n_1321)
);

AO31x2_ASAP7_75t_L g1322 ( 
.A1(n_1062),
.A2(n_358),
.A3(n_368),
.B(n_351),
.Y(n_1322)
);

NAND2x1p5_ASAP7_75t_L g1323 ( 
.A(n_1091),
.B(n_742),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1211),
.B(n_742),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1162),
.A2(n_828),
.B(n_790),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1211),
.B(n_761),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1162),
.A2(n_790),
.B(n_761),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_L g1328 ( 
.A(n_1087),
.B(n_1041),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1106),
.A2(n_1127),
.B(n_1108),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1062),
.Y(n_1330)
);

AND2x4_ASAP7_75t_L g1331 ( 
.A(n_1074),
.B(n_761),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1181),
.A2(n_1194),
.B1(n_1069),
.B2(n_1068),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1030),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1068),
.Y(n_1334)
);

CKINVDCx20_ASAP7_75t_R g1335 ( 
.A(n_1037),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1188),
.A2(n_790),
.B(n_761),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1206),
.B(n_761),
.Y(n_1337)
);

INVx1_ASAP7_75t_SL g1338 ( 
.A(n_1072),
.Y(n_1338)
);

OA22x2_ASAP7_75t_L g1339 ( 
.A1(n_1183),
.A2(n_446),
.B1(n_458),
.B2(n_455),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1087),
.B(n_1055),
.Y(n_1340)
);

OAI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1210),
.A2(n_791),
.B(n_785),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_1145),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1052),
.A2(n_1073),
.B(n_1138),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_1063),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_SL g1345 ( 
.A1(n_1131),
.A2(n_347),
.B(n_334),
.Y(n_1345)
);

AO31x2_ASAP7_75t_L g1346 ( 
.A1(n_1069),
.A2(n_358),
.A3(n_368),
.B(n_386),
.Y(n_1346)
);

BUFx2_ASAP7_75t_L g1347 ( 
.A(n_1177),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1188),
.A2(n_815),
.B(n_790),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1181),
.A2(n_1194),
.B1(n_1205),
.B2(n_1203),
.Y(n_1349)
);

AO31x2_ASAP7_75t_L g1350 ( 
.A1(n_1140),
.A2(n_400),
.A3(n_412),
.B(n_413),
.Y(n_1350)
);

AO21x1_ASAP7_75t_L g1351 ( 
.A1(n_1110),
.A2(n_412),
.B(n_400),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1030),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1034),
.Y(n_1353)
);

CKINVDCx20_ASAP7_75t_R g1354 ( 
.A(n_1065),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1071),
.A2(n_791),
.B(n_785),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1206),
.B(n_790),
.Y(n_1356)
);

INVx5_ASAP7_75t_L g1357 ( 
.A(n_1130),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1052),
.A2(n_533),
.B(n_528),
.Y(n_1358)
);

INVx3_ASAP7_75t_L g1359 ( 
.A(n_1182),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1034),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1206),
.B(n_815),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1087),
.B(n_373),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1180),
.B(n_785),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1180),
.B(n_331),
.Y(n_1364)
);

OAI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1081),
.A2(n_796),
.B(n_613),
.Y(n_1365)
);

OAI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1144),
.A2(n_796),
.B(n_613),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1052),
.A2(n_1073),
.B(n_1151),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1073),
.A2(n_540),
.B(n_537),
.Y(n_1368)
);

NAND3xp33_ASAP7_75t_SL g1369 ( 
.A(n_1141),
.B(n_345),
.C(n_335),
.Y(n_1369)
);

OAI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1164),
.A2(n_796),
.B(n_613),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1184),
.A2(n_1191),
.B(n_1148),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1203),
.A2(n_796),
.B(n_594),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1203),
.A2(n_796),
.B(n_594),
.Y(n_1373)
);

OAI22x1_ASAP7_75t_L g1374 ( 
.A1(n_1183),
.A2(n_431),
.B1(n_430),
.B2(n_429),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1125),
.B(n_373),
.Y(n_1375)
);

NOR2x1_ASAP7_75t_SL g1376 ( 
.A(n_1091),
.B(n_796),
.Y(n_1376)
);

O2A1O1Ixp5_ASAP7_75t_L g1377 ( 
.A1(n_1175),
.A2(n_537),
.B(n_564),
.C(n_558),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1205),
.A2(n_594),
.B(n_542),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1205),
.A2(n_1077),
.B(n_1202),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1129),
.B(n_346),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1036),
.Y(n_1381)
);

BUFx2_ASAP7_75t_L g1382 ( 
.A(n_1137),
.Y(n_1382)
);

NAND2x1_ASAP7_75t_L g1383 ( 
.A(n_1058),
.B(n_594),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1036),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1077),
.A2(n_542),
.B(n_540),
.Y(n_1385)
);

INVx3_ASAP7_75t_L g1386 ( 
.A(n_1236),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_SL g1387 ( 
.A1(n_1332),
.A2(n_1047),
.B(n_1038),
.Y(n_1387)
);

INVx3_ASAP7_75t_L g1388 ( 
.A(n_1236),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1226),
.A2(n_1047),
.B(n_1038),
.Y(n_1389)
);

OA21x2_ASAP7_75t_L g1390 ( 
.A1(n_1232),
.A2(n_1123),
.B(n_1066),
.Y(n_1390)
);

NOR2xp33_ASAP7_75t_L g1391 ( 
.A(n_1328),
.B(n_1075),
.Y(n_1391)
);

CKINVDCx6p67_ASAP7_75t_R g1392 ( 
.A(n_1354),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1221),
.A2(n_1180),
.B1(n_1217),
.B2(n_1194),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1328),
.B(n_1065),
.Y(n_1394)
);

OAI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1221),
.A2(n_1174),
.B1(n_1074),
.B2(n_1083),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1226),
.A2(n_1066),
.B(n_1059),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_R g1397 ( 
.A1(n_1349),
.A2(n_1153),
.B(n_1170),
.Y(n_1397)
);

OAI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1246),
.A2(n_1197),
.B1(n_1161),
.B2(n_1076),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1343),
.A2(n_1367),
.B(n_1232),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1234),
.B(n_1169),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1247),
.A2(n_1070),
.B(n_1059),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1242),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1229),
.A2(n_1217),
.B1(n_1170),
.B2(n_1083),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1258),
.Y(n_1404)
);

NAND3xp33_ASAP7_75t_L g1405 ( 
.A(n_1273),
.B(n_1048),
.C(n_1094),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1251),
.A2(n_1080),
.B(n_1070),
.Y(n_1406)
);

AO21x2_ASAP7_75t_L g1407 ( 
.A1(n_1320),
.A2(n_1101),
.B(n_1064),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1274),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1275),
.A2(n_1097),
.B(n_1080),
.Y(n_1409)
);

OAI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1222),
.A2(n_1101),
.B(n_1064),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1235),
.B(n_1239),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1259),
.A2(n_1245),
.B(n_1271),
.Y(n_1412)
);

AOI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1222),
.A2(n_1117),
.B(n_1085),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1284),
.Y(n_1414)
);

AO21x2_ASAP7_75t_L g1415 ( 
.A1(n_1366),
.A2(n_1096),
.B(n_1119),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1229),
.A2(n_1170),
.B1(n_1083),
.B2(n_1116),
.Y(n_1416)
);

OAI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1253),
.A2(n_1099),
.B(n_1097),
.Y(n_1417)
);

AOI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1276),
.A2(n_1085),
.B(n_1084),
.Y(n_1418)
);

CKINVDCx20_ASAP7_75t_R g1419 ( 
.A(n_1335),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1246),
.A2(n_1090),
.B1(n_1132),
.B2(n_1116),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1333),
.Y(n_1421)
);

AO21x2_ASAP7_75t_L g1422 ( 
.A1(n_1370),
.A2(n_1060),
.B(n_1199),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1272),
.A2(n_1109),
.B(n_1099),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1228),
.A2(n_1077),
.B1(n_1058),
.B2(n_1182),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1333),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1254),
.A2(n_1124),
.B(n_1109),
.Y(n_1426)
);

OA21x2_ASAP7_75t_L g1427 ( 
.A1(n_1377),
.A2(n_1123),
.B(n_1124),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1282),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1293),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1294),
.Y(n_1430)
);

AO31x2_ASAP7_75t_L g1431 ( 
.A1(n_1223),
.A2(n_1135),
.A3(n_1086),
.B(n_1092),
.Y(n_1431)
);

OAI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1227),
.A2(n_1135),
.B(n_1118),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1230),
.A2(n_1058),
.B1(n_1208),
.B2(n_1107),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1254),
.A2(n_1086),
.B(n_1084),
.Y(n_1434)
);

CKINVDCx16_ASAP7_75t_R g1435 ( 
.A(n_1354),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1316),
.A2(n_1095),
.B(n_1092),
.Y(n_1436)
);

BUFx12f_ASAP7_75t_L g1437 ( 
.A(n_1257),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1249),
.B(n_1284),
.Y(n_1438)
);

INVx4_ASAP7_75t_L g1439 ( 
.A(n_1357),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1252),
.B(n_1284),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_1288),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1307),
.Y(n_1442)
);

INVxp67_ASAP7_75t_SL g1443 ( 
.A(n_1291),
.Y(n_1443)
);

CKINVDCx8_ASAP7_75t_R g1444 ( 
.A(n_1344),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1317),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1248),
.A2(n_1208),
.B(n_1126),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1285),
.A2(n_1104),
.B(n_1095),
.Y(n_1447)
);

BUFx3_ASAP7_75t_L g1448 ( 
.A(n_1224),
.Y(n_1448)
);

OAI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1252),
.A2(n_1208),
.B1(n_1107),
.B2(n_1112),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1252),
.B(n_1241),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1330),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1241),
.B(n_1169),
.Y(n_1452)
);

O2A1O1Ixp33_ASAP7_75t_SL g1453 ( 
.A1(n_1363),
.A2(n_1113),
.B(n_1104),
.C(n_1105),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1334),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1296),
.A2(n_1113),
.B(n_1105),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1312),
.B(n_1090),
.Y(n_1456)
);

OA21x2_ASAP7_75t_L g1457 ( 
.A1(n_1377),
.A2(n_1115),
.B(n_1114),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1340),
.A2(n_1132),
.B1(n_1116),
.B2(n_1090),
.Y(n_1458)
);

OAI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1347),
.A2(n_1197),
.B1(n_1161),
.B2(n_1076),
.Y(n_1459)
);

INVx1_ASAP7_75t_SL g1460 ( 
.A(n_1265),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_SL g1461 ( 
.A1(n_1345),
.A2(n_1215),
.B(n_1154),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1360),
.Y(n_1462)
);

OAI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1296),
.A2(n_1115),
.B(n_1114),
.Y(n_1463)
);

AO21x2_ASAP7_75t_L g1464 ( 
.A1(n_1365),
.A2(n_1351),
.B(n_1237),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1360),
.Y(n_1465)
);

BUFx10_ASAP7_75t_L g1466 ( 
.A(n_1344),
.Y(n_1466)
);

OAI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1298),
.A2(n_1133),
.B(n_1121),
.Y(n_1467)
);

INVxp67_ASAP7_75t_SL g1468 ( 
.A(n_1291),
.Y(n_1468)
);

INVx3_ASAP7_75t_L g1469 ( 
.A(n_1312),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1384),
.Y(n_1470)
);

INVx3_ASAP7_75t_L g1471 ( 
.A(n_1359),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1384),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1352),
.Y(n_1473)
);

OAI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1342),
.A2(n_1040),
.B1(n_1098),
.B2(n_1102),
.Y(n_1474)
);

OAI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1299),
.A2(n_1364),
.B1(n_1338),
.B2(n_1279),
.Y(n_1475)
);

INVx2_ASAP7_75t_SL g1476 ( 
.A(n_1224),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1353),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1298),
.A2(n_1368),
.B(n_1358),
.Y(n_1478)
);

INVxp67_ASAP7_75t_SL g1479 ( 
.A(n_1225),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1381),
.Y(n_1480)
);

AOI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1379),
.A2(n_1126),
.B(n_1131),
.Y(n_1481)
);

AOI22x1_ASAP7_75t_L g1482 ( 
.A1(n_1240),
.A2(n_1319),
.B1(n_1355),
.B2(n_1321),
.Y(n_1482)
);

O2A1O1Ixp33_ASAP7_75t_L g1483 ( 
.A1(n_1369),
.A2(n_1089),
.B(n_1150),
.C(n_1196),
.Y(n_1483)
);

INVxp67_ASAP7_75t_L g1484 ( 
.A(n_1380),
.Y(n_1484)
);

INVx4_ASAP7_75t_SL g1485 ( 
.A(n_1225),
.Y(n_1485)
);

OAI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1243),
.A2(n_1133),
.B(n_1121),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1382),
.Y(n_1487)
);

NOR2xp33_ASAP7_75t_L g1488 ( 
.A(n_1362),
.B(n_1137),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_L g1489 ( 
.A1(n_1371),
.A2(n_1148),
.B(n_1146),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1369),
.A2(n_1375),
.B1(n_1267),
.B2(n_1269),
.Y(n_1490)
);

BUFx6f_ASAP7_75t_L g1491 ( 
.A(n_1357),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1335),
.B(n_1122),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1289),
.B(n_1139),
.Y(n_1493)
);

OR2x6_ASAP7_75t_L g1494 ( 
.A(n_1359),
.B(n_1091),
.Y(n_1494)
);

AOI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1260),
.A2(n_1157),
.B(n_1154),
.Y(n_1495)
);

NOR2xp67_ASAP7_75t_L g1496 ( 
.A(n_1281),
.B(n_1103),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_SL g1497 ( 
.A(n_1255),
.B(n_1040),
.Y(n_1497)
);

OA21x2_ASAP7_75t_L g1498 ( 
.A1(n_1256),
.A2(n_1160),
.B(n_1146),
.Y(n_1498)
);

INVx1_ASAP7_75t_SL g1499 ( 
.A(n_1255),
.Y(n_1499)
);

BUFx6f_ASAP7_75t_L g1500 ( 
.A(n_1357),
.Y(n_1500)
);

OA21x2_ASAP7_75t_L g1501 ( 
.A1(n_1329),
.A2(n_1262),
.B(n_1302),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1250),
.A2(n_1112),
.B1(n_1091),
.B2(n_1107),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_L g1503 ( 
.A1(n_1279),
.A2(n_1132),
.B1(n_1156),
.B2(n_1098),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1292),
.A2(n_1102),
.B1(n_1147),
.B2(n_1167),
.Y(n_1504)
);

INVx3_ASAP7_75t_L g1505 ( 
.A(n_1225),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1225),
.Y(n_1506)
);

NOR2xp67_ASAP7_75t_L g1507 ( 
.A(n_1357),
.B(n_1103),
.Y(n_1507)
);

OA21x2_ASAP7_75t_L g1508 ( 
.A1(n_1329),
.A2(n_1163),
.B(n_1160),
.Y(n_1508)
);

OAI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1262),
.A2(n_1165),
.B(n_1163),
.Y(n_1509)
);

OAI22xp33_ASAP7_75t_SL g1510 ( 
.A1(n_1270),
.A2(n_413),
.B1(n_419),
.B2(n_446),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1295),
.B(n_1033),
.Y(n_1511)
);

OAI21x1_ASAP7_75t_L g1512 ( 
.A1(n_1300),
.A2(n_1168),
.B(n_1165),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1302),
.B(n_1168),
.Y(n_1513)
);

OAI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1300),
.A2(n_1327),
.B(n_1325),
.Y(n_1514)
);

OAI21x1_ASAP7_75t_L g1515 ( 
.A1(n_1300),
.A2(n_1128),
.B(n_1103),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1261),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1292),
.A2(n_1278),
.B1(n_1326),
.B2(n_1324),
.Y(n_1517)
);

BUFx6f_ASAP7_75t_L g1518 ( 
.A(n_1309),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1297),
.Y(n_1519)
);

NOR3xp33_ASAP7_75t_SL g1520 ( 
.A(n_1270),
.B(n_356),
.C(n_354),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1304),
.Y(n_1521)
);

A2O1A1Ixp33_ASAP7_75t_L g1522 ( 
.A1(n_1337),
.A2(n_1216),
.B(n_1198),
.C(n_1111),
.Y(n_1522)
);

BUFx2_ASAP7_75t_R g1523 ( 
.A(n_1356),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1306),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1311),
.Y(n_1525)
);

OAI21x1_ASAP7_75t_L g1526 ( 
.A1(n_1336),
.A2(n_1128),
.B(n_1171),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1292),
.A2(n_1147),
.B1(n_1167),
.B2(n_1128),
.Y(n_1527)
);

BUFx8_ASAP7_75t_SL g1528 ( 
.A(n_1257),
.Y(n_1528)
);

O2A1O1Ixp33_ASAP7_75t_L g1529 ( 
.A1(n_1280),
.A2(n_447),
.B(n_452),
.C(n_454),
.Y(n_1529)
);

AOI222xp33_ASAP7_75t_L g1530 ( 
.A1(n_1374),
.A2(n_460),
.B1(n_458),
.B2(n_452),
.C1(n_447),
.C2(n_437),
.Y(n_1530)
);

NAND3xp33_ASAP7_75t_SL g1531 ( 
.A(n_1385),
.B(n_361),
.C(n_359),
.Y(n_1531)
);

AO21x2_ASAP7_75t_L g1532 ( 
.A1(n_1290),
.A2(n_1341),
.B(n_1287),
.Y(n_1532)
);

OAI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1378),
.A2(n_1171),
.B(n_1167),
.Y(n_1533)
);

O2A1O1Ixp33_ASAP7_75t_SL g1534 ( 
.A1(n_1361),
.A2(n_1033),
.B(n_558),
.C(n_564),
.Y(n_1534)
);

AOI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1263),
.A2(n_1157),
.B(n_1154),
.Y(n_1535)
);

AOI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1264),
.A2(n_1157),
.B(n_1107),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1261),
.Y(n_1537)
);

NOR2x1_ASAP7_75t_SL g1538 ( 
.A(n_1309),
.B(n_1091),
.Y(n_1538)
);

INVx1_ASAP7_75t_SL g1539 ( 
.A(n_1315),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1310),
.B(n_1107),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1261),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1268),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1283),
.Y(n_1543)
);

NAND2x1p5_ASAP7_75t_L g1544 ( 
.A(n_1309),
.B(n_1112),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1286),
.B(n_1322),
.Y(n_1545)
);

OAI21x1_ASAP7_75t_L g1546 ( 
.A1(n_1348),
.A2(n_548),
.B(n_546),
.Y(n_1546)
);

AO31x2_ASAP7_75t_L g1547 ( 
.A1(n_1305),
.A2(n_553),
.A3(n_548),
.B(n_546),
.Y(n_1547)
);

OAI21xp5_ASAP7_75t_L g1548 ( 
.A1(n_1318),
.A2(n_553),
.B(n_364),
.Y(n_1548)
);

BUFx2_ASAP7_75t_L g1549 ( 
.A(n_1309),
.Y(n_1549)
);

OAI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1301),
.A2(n_1112),
.B(n_1214),
.Y(n_1550)
);

OAI21x1_ASAP7_75t_L g1551 ( 
.A1(n_1308),
.A2(n_1112),
.B(n_1214),
.Y(n_1551)
);

BUFx2_ASAP7_75t_SL g1552 ( 
.A(n_1303),
.Y(n_1552)
);

OAI21x1_ASAP7_75t_L g1553 ( 
.A1(n_1372),
.A2(n_1214),
.B(n_1152),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1268),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1233),
.B(n_1130),
.Y(n_1555)
);

NAND3xp33_ASAP7_75t_SL g1556 ( 
.A(n_1383),
.B(n_403),
.C(n_459),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1268),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1268),
.Y(n_1558)
);

OAI21x1_ASAP7_75t_L g1559 ( 
.A1(n_1373),
.A2(n_1214),
.B(n_1152),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_1315),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1322),
.B(n_1130),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1310),
.Y(n_1562)
);

INVxp67_ASAP7_75t_L g1563 ( 
.A(n_1339),
.Y(n_1563)
);

AO31x2_ASAP7_75t_L g1564 ( 
.A1(n_1376),
.A2(n_1100),
.A3(n_1152),
.B(n_422),
.Y(n_1564)
);

OAI21x1_ASAP7_75t_L g1565 ( 
.A1(n_1266),
.A2(n_1214),
.B(n_1152),
.Y(n_1565)
);

INVx3_ASAP7_75t_L g1566 ( 
.A(n_1310),
.Y(n_1566)
);

OAI21x1_ASAP7_75t_L g1567 ( 
.A1(n_1277),
.A2(n_1152),
.B(n_422),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1421),
.Y(n_1568)
);

OAI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1391),
.A2(n_1331),
.B(n_1339),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1394),
.A2(n_1331),
.B1(n_1323),
.B2(n_362),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1402),
.Y(n_1571)
);

CKINVDCx20_ASAP7_75t_R g1572 ( 
.A(n_1528),
.Y(n_1572)
);

AO31x2_ASAP7_75t_L g1573 ( 
.A1(n_1516),
.A2(n_1313),
.A3(n_1314),
.B(n_1238),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_SL g1574 ( 
.A1(n_1405),
.A2(n_408),
.B1(n_375),
.B2(n_378),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1421),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1441),
.A2(n_416),
.B1(n_381),
.B2(n_382),
.Y(n_1576)
);

CKINVDCx11_ASAP7_75t_R g1577 ( 
.A(n_1444),
.Y(n_1577)
);

BUFx2_ASAP7_75t_R g1578 ( 
.A(n_1444),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1411),
.B(n_1350),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1400),
.B(n_1350),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1414),
.B(n_1322),
.Y(n_1581)
);

AND2x4_ASAP7_75t_L g1582 ( 
.A(n_1440),
.B(n_1314),
.Y(n_1582)
);

OAI22xp5_ASAP7_75t_SL g1583 ( 
.A1(n_1435),
.A2(n_449),
.B1(n_448),
.B2(n_445),
.Y(n_1583)
);

OAI211xp5_ASAP7_75t_L g1584 ( 
.A1(n_1530),
.A2(n_404),
.B(n_385),
.C(n_387),
.Y(n_1584)
);

OAI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1493),
.A2(n_370),
.B(n_389),
.Y(n_1585)
);

OAI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1441),
.A2(n_440),
.B1(n_394),
.B2(n_396),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1460),
.B(n_1350),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1425),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1425),
.Y(n_1589)
);

AOI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1481),
.A2(n_1238),
.B(n_1231),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1460),
.B(n_1350),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_1437),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1402),
.Y(n_1593)
);

OAI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1405),
.A2(n_427),
.B1(n_399),
.B2(n_401),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1404),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1404),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1408),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1414),
.B(n_1322),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1408),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_SL g1600 ( 
.A1(n_1510),
.A2(n_390),
.B1(n_402),
.B2(n_405),
.Y(n_1600)
);

BUFx6f_ASAP7_75t_L g1601 ( 
.A(n_1491),
.Y(n_1601)
);

OR2x6_ASAP7_75t_L g1602 ( 
.A(n_1450),
.B(n_1314),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1428),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1562),
.B(n_1346),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1492),
.B(n_411),
.Y(n_1605)
);

OAI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1420),
.A2(n_1393),
.B1(n_1490),
.B2(n_1484),
.Y(n_1606)
);

INVx4_ASAP7_75t_L g1607 ( 
.A(n_1491),
.Y(n_1607)
);

AND2x4_ASAP7_75t_L g1608 ( 
.A(n_1440),
.B(n_1314),
.Y(n_1608)
);

OAI21x1_ASAP7_75t_SL g1609 ( 
.A1(n_1387),
.A2(n_1346),
.B(n_1313),
.Y(n_1609)
);

AO31x2_ASAP7_75t_L g1610 ( 
.A1(n_1516),
.A2(n_1313),
.A3(n_1238),
.B(n_1244),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_SL g1611 ( 
.A1(n_1510),
.A2(n_444),
.B1(n_441),
.B2(n_417),
.Y(n_1611)
);

OAI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1435),
.A2(n_1346),
.B1(n_1231),
.B2(n_1238),
.Y(n_1612)
);

AOI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1495),
.A2(n_1231),
.B(n_1244),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1530),
.A2(n_422),
.B1(n_1346),
.B2(n_1231),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_L g1615 ( 
.A(n_1438),
.B(n_134),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1428),
.Y(n_1616)
);

OAI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1503),
.A2(n_1244),
.B1(n_1313),
.B2(n_11),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1429),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1562),
.B(n_1244),
.Y(n_1619)
);

CKINVDCx16_ASAP7_75t_R g1620 ( 
.A(n_1437),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1452),
.A2(n_422),
.B1(n_10),
.B2(n_12),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1566),
.B(n_135),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1400),
.B(n_1487),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1429),
.Y(n_1624)
);

OAI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1488),
.A2(n_8),
.B1(n_10),
.B2(n_13),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1462),
.Y(n_1626)
);

INVx1_ASAP7_75t_SL g1627 ( 
.A(n_1499),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1475),
.A2(n_422),
.B1(n_15),
.B2(n_17),
.Y(n_1628)
);

BUFx6f_ASAP7_75t_L g1629 ( 
.A(n_1491),
.Y(n_1629)
);

AOI22xp33_ASAP7_75t_L g1630 ( 
.A1(n_1531),
.A2(n_422),
.B1(n_17),
.B2(n_18),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1462),
.Y(n_1631)
);

AO21x2_ASAP7_75t_L g1632 ( 
.A1(n_1418),
.A2(n_422),
.B(n_235),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1403),
.A2(n_422),
.B1(n_18),
.B2(n_19),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1545),
.B(n_422),
.Y(n_1634)
);

AND2x4_ASAP7_75t_L g1635 ( 
.A(n_1566),
.B(n_138),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1465),
.Y(n_1636)
);

AOI22xp33_ASAP7_75t_L g1637 ( 
.A1(n_1517),
.A2(n_14),
.B1(n_21),
.B2(n_23),
.Y(n_1637)
);

CKINVDCx16_ASAP7_75t_R g1638 ( 
.A(n_1419),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1430),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1545),
.B(n_143),
.Y(n_1640)
);

INVx4_ASAP7_75t_L g1641 ( 
.A(n_1491),
.Y(n_1641)
);

O2A1O1Ixp33_ASAP7_75t_SL g1642 ( 
.A1(n_1522),
.A2(n_14),
.B(n_24),
.C(n_25),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1430),
.Y(n_1643)
);

INVxp67_ASAP7_75t_L g1644 ( 
.A(n_1443),
.Y(n_1644)
);

NAND2xp33_ASAP7_75t_R g1645 ( 
.A(n_1520),
.B(n_153),
.Y(n_1645)
);

BUFx2_ASAP7_75t_L g1646 ( 
.A(n_1448),
.Y(n_1646)
);

OAI21x1_ASAP7_75t_L g1647 ( 
.A1(n_1399),
.A2(n_234),
.B(n_232),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1480),
.B(n_161),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1563),
.B(n_24),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1442),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1543),
.B(n_27),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1543),
.B(n_28),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1499),
.Y(n_1653)
);

NAND3x1_ASAP7_75t_L g1654 ( 
.A(n_1397),
.B(n_28),
.C(n_30),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1465),
.Y(n_1655)
);

OAI211xp5_ASAP7_75t_SL g1656 ( 
.A1(n_1483),
.A2(n_32),
.B(n_34),
.C(n_35),
.Y(n_1656)
);

OAI211xp5_ASAP7_75t_L g1657 ( 
.A1(n_1529),
.A2(n_32),
.B(n_35),
.C(n_36),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1398),
.B(n_230),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_R g1659 ( 
.A(n_1392),
.B(n_229),
.Y(n_1659)
);

NAND2xp33_ASAP7_75t_SL g1660 ( 
.A(n_1491),
.B(n_36),
.Y(n_1660)
);

AOI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1474),
.A2(n_38),
.B1(n_39),
.B2(n_42),
.Y(n_1661)
);

INVx2_ASAP7_75t_SL g1662 ( 
.A(n_1448),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1480),
.B(n_228),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1442),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_1392),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1470),
.Y(n_1666)
);

AOI22xp33_ASAP7_75t_L g1667 ( 
.A1(n_1416),
.A2(n_38),
.B1(n_44),
.B2(n_45),
.Y(n_1667)
);

AOI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1552),
.A2(n_1511),
.B1(n_1556),
.B2(n_1482),
.Y(n_1668)
);

INVx4_ASAP7_75t_L g1669 ( 
.A(n_1500),
.Y(n_1669)
);

OR2x6_ASAP7_75t_L g1670 ( 
.A(n_1446),
.B(n_221),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1445),
.Y(n_1671)
);

AND2x4_ASAP7_75t_L g1672 ( 
.A(n_1566),
.B(n_216),
.Y(n_1672)
);

INVx6_ASAP7_75t_L g1673 ( 
.A(n_1466),
.Y(n_1673)
);

OAI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1458),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_1674)
);

A2O1A1Ixp33_ASAP7_75t_L g1675 ( 
.A1(n_1432),
.A2(n_48),
.B(n_49),
.C(n_50),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1470),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1519),
.B(n_211),
.Y(n_1677)
);

BUFx3_ASAP7_75t_L g1678 ( 
.A(n_1448),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1519),
.B(n_51),
.Y(n_1679)
);

INVx3_ASAP7_75t_L g1680 ( 
.A(n_1439),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1445),
.Y(n_1681)
);

OAI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1539),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1552),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_1683)
);

INVx2_ASAP7_75t_SL g1684 ( 
.A(n_1466),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1472),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1482),
.A2(n_56),
.B1(n_58),
.B2(n_61),
.Y(n_1686)
);

AOI22xp33_ASAP7_75t_SL g1687 ( 
.A1(n_1466),
.A2(n_1539),
.B1(n_1560),
.B2(n_1468),
.Y(n_1687)
);

BUFx2_ASAP7_75t_L g1688 ( 
.A(n_1476),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1560),
.A2(n_58),
.B1(n_62),
.B2(n_64),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1451),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1521),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_1691)
);

A2O1A1Ixp33_ASAP7_75t_L g1692 ( 
.A1(n_1432),
.A2(n_68),
.B(n_70),
.C(n_74),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1521),
.A2(n_70),
.B1(n_74),
.B2(n_75),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1524),
.B(n_207),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1451),
.Y(n_1695)
);

AO221x2_ASAP7_75t_L g1696 ( 
.A1(n_1459),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.C(n_79),
.Y(n_1696)
);

INVx3_ASAP7_75t_L g1697 ( 
.A(n_1439),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1454),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1524),
.B(n_1525),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_1466),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1497),
.B(n_76),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1525),
.B(n_206),
.Y(n_1702)
);

OAI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1476),
.A2(n_80),
.B1(n_82),
.B2(n_83),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1454),
.Y(n_1704)
);

NAND2xp33_ASAP7_75t_SL g1705 ( 
.A(n_1500),
.B(n_80),
.Y(n_1705)
);

NOR3xp33_ASAP7_75t_SL g1706 ( 
.A(n_1555),
.B(n_83),
.C(n_84),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_1523),
.Y(n_1707)
);

AOI21xp5_ASAP7_75t_L g1708 ( 
.A1(n_1535),
.A2(n_201),
.B(n_186),
.Y(n_1708)
);

NAND2x1p5_ASAP7_75t_L g1709 ( 
.A(n_1439),
.B(n_1500),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1472),
.Y(n_1710)
);

AND2x4_ASAP7_75t_L g1711 ( 
.A(n_1566),
.B(n_170),
.Y(n_1711)
);

AND2x4_ASAP7_75t_L g1712 ( 
.A(n_1456),
.B(n_165),
.Y(n_1712)
);

INVx3_ASAP7_75t_L g1713 ( 
.A(n_1439),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1512),
.Y(n_1714)
);

CKINVDCx11_ASAP7_75t_R g1715 ( 
.A(n_1500),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1512),
.Y(n_1716)
);

AND2x2_ASAP7_75t_SL g1717 ( 
.A(n_1501),
.B(n_1504),
.Y(n_1717)
);

OAI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1395),
.A2(n_84),
.B(n_86),
.Y(n_1718)
);

NOR2xp67_ASAP7_75t_SL g1719 ( 
.A(n_1500),
.B(n_86),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1508),
.Y(n_1720)
);

CKINVDCx8_ASAP7_75t_R g1721 ( 
.A(n_1485),
.Y(n_1721)
);

AND2x4_ASAP7_75t_L g1722 ( 
.A(n_1456),
.B(n_89),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1508),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1508),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1473),
.Y(n_1725)
);

NAND2xp33_ASAP7_75t_R g1726 ( 
.A(n_1456),
.B(n_89),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1473),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_1549),
.Y(n_1728)
);

AOI22xp33_ASAP7_75t_L g1729 ( 
.A1(n_1407),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1477),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1508),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1477),
.B(n_94),
.Y(n_1732)
);

NAND2xp33_ASAP7_75t_L g1733 ( 
.A(n_1449),
.B(n_95),
.Y(n_1733)
);

BUFx6f_ASAP7_75t_L g1734 ( 
.A(n_1518),
.Y(n_1734)
);

NAND3xp33_ASAP7_75t_SL g1735 ( 
.A(n_1527),
.B(n_96),
.C(n_97),
.Y(n_1735)
);

OAI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1496),
.A2(n_96),
.B1(n_99),
.B2(n_100),
.Y(n_1736)
);

AOI22xp33_ASAP7_75t_L g1737 ( 
.A1(n_1407),
.A2(n_99),
.B1(n_101),
.B2(n_102),
.Y(n_1737)
);

OAI21x1_ASAP7_75t_L g1738 ( 
.A1(n_1399),
.A2(n_102),
.B(n_103),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1513),
.B(n_1561),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_1549),
.Y(n_1740)
);

AOI22xp33_ASAP7_75t_L g1741 ( 
.A1(n_1407),
.A2(n_105),
.B1(n_107),
.B2(n_112),
.Y(n_1741)
);

NAND3xp33_ASAP7_75t_L g1742 ( 
.A(n_1548),
.B(n_105),
.C(n_117),
.Y(n_1742)
);

NAND2xp33_ASAP7_75t_SL g1743 ( 
.A(n_1540),
.B(n_120),
.Y(n_1743)
);

OAI21xp33_ASAP7_75t_L g1744 ( 
.A1(n_1513),
.A2(n_1410),
.B(n_1561),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1422),
.A2(n_1464),
.B1(n_1456),
.B2(n_1496),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1479),
.B(n_1431),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1431),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_SL g1748 ( 
.A1(n_1422),
.A2(n_1464),
.B1(n_1538),
.B2(n_1410),
.Y(n_1748)
);

INVx3_ASAP7_75t_L g1749 ( 
.A(n_1540),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_1518),
.Y(n_1750)
);

NOR2x1_ASAP7_75t_SL g1751 ( 
.A(n_1494),
.B(n_1502),
.Y(n_1751)
);

NAND2xp33_ASAP7_75t_SL g1752 ( 
.A(n_1540),
.B(n_1433),
.Y(n_1752)
);

AO21x2_ASAP7_75t_L g1753 ( 
.A1(n_1418),
.A2(n_1412),
.B(n_1542),
.Y(n_1753)
);

AOI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1422),
.A2(n_1464),
.B1(n_1387),
.B2(n_1532),
.Y(n_1754)
);

AND2x2_ASAP7_75t_SL g1755 ( 
.A(n_1501),
.B(n_1540),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1431),
.B(n_1564),
.Y(n_1756)
);

AOI21xp33_ASAP7_75t_L g1757 ( 
.A1(n_1532),
.A2(n_1501),
.B(n_1415),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1431),
.Y(n_1758)
);

AOI22xp33_ASAP7_75t_L g1759 ( 
.A1(n_1532),
.A2(n_1501),
.B1(n_1415),
.B2(n_1417),
.Y(n_1759)
);

AOI22xp33_ASAP7_75t_L g1760 ( 
.A1(n_1415),
.A2(n_1417),
.B1(n_1461),
.B2(n_1533),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_L g1761 ( 
.A(n_1505),
.B(n_1506),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1461),
.A2(n_1533),
.B1(n_1469),
.B2(n_1471),
.Y(n_1762)
);

BUFx3_ASAP7_75t_L g1763 ( 
.A(n_1518),
.Y(n_1763)
);

OR2x6_ASAP7_75t_L g1764 ( 
.A(n_1494),
.B(n_1509),
.Y(n_1764)
);

CKINVDCx5p33_ASAP7_75t_R g1765 ( 
.A(n_1518),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1431),
.B(n_1564),
.Y(n_1766)
);

AO21x1_ASAP7_75t_L g1767 ( 
.A1(n_1509),
.A2(n_1554),
.B(n_1558),
.Y(n_1767)
);

AOI22xp33_ASAP7_75t_L g1768 ( 
.A1(n_1469),
.A2(n_1471),
.B1(n_1390),
.B2(n_1424),
.Y(n_1768)
);

BUFx12f_ASAP7_75t_L g1769 ( 
.A(n_1518),
.Y(n_1769)
);

BUFx3_ASAP7_75t_L g1770 ( 
.A(n_1505),
.Y(n_1770)
);

AND2x4_ASAP7_75t_L g1771 ( 
.A(n_1485),
.B(n_1386),
.Y(n_1771)
);

AOI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1696),
.A2(n_1471),
.B1(n_1469),
.B2(n_1388),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1696),
.A2(n_1471),
.B1(n_1469),
.B2(n_1388),
.Y(n_1773)
);

OAI211xp5_ASAP7_75t_L g1774 ( 
.A1(n_1584),
.A2(n_1534),
.B(n_1413),
.C(n_1453),
.Y(n_1774)
);

AOI22xp33_ASAP7_75t_L g1775 ( 
.A1(n_1696),
.A2(n_1386),
.B1(n_1388),
.B2(n_1390),
.Y(n_1775)
);

OAI21xp33_ASAP7_75t_SL g1776 ( 
.A1(n_1658),
.A2(n_1494),
.B(n_1507),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1571),
.Y(n_1777)
);

INVx5_ASAP7_75t_SL g1778 ( 
.A(n_1670),
.Y(n_1778)
);

BUFx3_ASAP7_75t_L g1779 ( 
.A(n_1678),
.Y(n_1779)
);

OAI22xp5_ASAP7_75t_L g1780 ( 
.A1(n_1605),
.A2(n_1494),
.B1(n_1507),
.B2(n_1386),
.Y(n_1780)
);

INVx1_ASAP7_75t_SL g1781 ( 
.A(n_1627),
.Y(n_1781)
);

AOI22xp33_ASAP7_75t_L g1782 ( 
.A1(n_1656),
.A2(n_1386),
.B1(n_1388),
.B2(n_1390),
.Y(n_1782)
);

AOI22xp33_ASAP7_75t_L g1783 ( 
.A1(n_1733),
.A2(n_1427),
.B1(n_1494),
.B2(n_1505),
.Y(n_1783)
);

AOI22xp33_ASAP7_75t_L g1784 ( 
.A1(n_1733),
.A2(n_1427),
.B1(n_1505),
.B2(n_1506),
.Y(n_1784)
);

OAI22xp33_ASAP7_75t_L g1785 ( 
.A1(n_1726),
.A2(n_1506),
.B1(n_1413),
.B2(n_1544),
.Y(n_1785)
);

AOI22xp33_ASAP7_75t_L g1786 ( 
.A1(n_1735),
.A2(n_1427),
.B1(n_1506),
.B2(n_1557),
.Y(n_1786)
);

AOI22xp33_ASAP7_75t_L g1787 ( 
.A1(n_1743),
.A2(n_1542),
.B1(n_1558),
.B2(n_1557),
.Y(n_1787)
);

OAI221xp5_ASAP7_75t_L g1788 ( 
.A1(n_1574),
.A2(n_1554),
.B1(n_1537),
.B2(n_1541),
.C(n_1536),
.Y(n_1788)
);

OAI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1687),
.A2(n_1544),
.B1(n_1541),
.B2(n_1498),
.Y(n_1789)
);

BUFx4f_ASAP7_75t_SL g1790 ( 
.A(n_1572),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1739),
.B(n_1634),
.Y(n_1791)
);

OAI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1661),
.A2(n_1544),
.B1(n_1498),
.B2(n_1457),
.Y(n_1792)
);

AOI221xp5_ASAP7_75t_L g1793 ( 
.A1(n_1594),
.A2(n_1564),
.B1(n_1547),
.B2(n_1546),
.C(n_1389),
.Y(n_1793)
);

OAI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1628),
.A2(n_1498),
.B1(n_1457),
.B2(n_1564),
.Y(n_1794)
);

AOI22xp33_ASAP7_75t_L g1795 ( 
.A1(n_1743),
.A2(n_1498),
.B1(n_1396),
.B2(n_1389),
.Y(n_1795)
);

INVx2_ASAP7_75t_SL g1796 ( 
.A(n_1673),
.Y(n_1796)
);

INVx2_ASAP7_75t_SL g1797 ( 
.A(n_1673),
.Y(n_1797)
);

OAI22xp5_ASAP7_75t_SL g1798 ( 
.A1(n_1707),
.A2(n_1457),
.B1(n_1564),
.B2(n_1485),
.Y(n_1798)
);

AOI22xp33_ASAP7_75t_L g1799 ( 
.A1(n_1606),
.A2(n_1396),
.B1(n_1457),
.B2(n_1567),
.Y(n_1799)
);

BUFx3_ASAP7_75t_L g1800 ( 
.A(n_1678),
.Y(n_1800)
);

AOI221xp5_ASAP7_75t_L g1801 ( 
.A1(n_1682),
.A2(n_1547),
.B1(n_1546),
.B2(n_1486),
.C(n_1401),
.Y(n_1801)
);

AOI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1645),
.A2(n_1485),
.B1(n_1559),
.B2(n_1553),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1593),
.Y(n_1803)
);

OAI22xp5_ASAP7_75t_L g1804 ( 
.A1(n_1637),
.A2(n_1700),
.B1(n_1611),
.B2(n_1600),
.Y(n_1804)
);

NAND2x1_ASAP7_75t_L g1805 ( 
.A(n_1673),
.B(n_1538),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1595),
.Y(n_1806)
);

BUFx6f_ASAP7_75t_L g1807 ( 
.A(n_1715),
.Y(n_1807)
);

A2O1A1Ixp33_ASAP7_75t_L g1808 ( 
.A1(n_1675),
.A2(n_1550),
.B(n_1551),
.C(n_1486),
.Y(n_1808)
);

HB1xp67_ASAP7_75t_L g1809 ( 
.A(n_1653),
.Y(n_1809)
);

AOI221xp5_ASAP7_75t_L g1810 ( 
.A1(n_1675),
.A2(n_1692),
.B1(n_1625),
.B2(n_1736),
.C(n_1674),
.Y(n_1810)
);

AOI22xp33_ASAP7_75t_L g1811 ( 
.A1(n_1660),
.A2(n_1567),
.B1(n_1436),
.B2(n_1401),
.Y(n_1811)
);

INVx3_ASAP7_75t_L g1812 ( 
.A(n_1582),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1739),
.B(n_1547),
.Y(n_1813)
);

OAI22xp33_ASAP7_75t_L g1814 ( 
.A1(n_1707),
.A2(n_1526),
.B1(n_1547),
.B2(n_1551),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1596),
.Y(n_1815)
);

CKINVDCx11_ASAP7_75t_R g1816 ( 
.A(n_1572),
.Y(n_1816)
);

AOI221xp5_ASAP7_75t_L g1817 ( 
.A1(n_1692),
.A2(n_1547),
.B1(n_1406),
.B2(n_1423),
.C(n_1489),
.Y(n_1817)
);

AOI22xp33_ASAP7_75t_L g1818 ( 
.A1(n_1660),
.A2(n_1436),
.B1(n_1406),
.B2(n_1526),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1597),
.Y(n_1819)
);

AOI22xp33_ASAP7_75t_SL g1820 ( 
.A1(n_1718),
.A2(n_1550),
.B1(n_1559),
.B2(n_1553),
.Y(n_1820)
);

INVx3_ASAP7_75t_L g1821 ( 
.A(n_1582),
.Y(n_1821)
);

AOI22xp33_ASAP7_75t_L g1822 ( 
.A1(n_1705),
.A2(n_1412),
.B1(n_1423),
.B2(n_1434),
.Y(n_1822)
);

OR2x2_ASAP7_75t_L g1823 ( 
.A(n_1580),
.B(n_1434),
.Y(n_1823)
);

A2O1A1Ixp33_ASAP7_75t_L g1824 ( 
.A1(n_1705),
.A2(n_1426),
.B(n_1489),
.C(n_1514),
.Y(n_1824)
);

NOR2x1_ASAP7_75t_SL g1825 ( 
.A(n_1670),
.B(n_1426),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1636),
.Y(n_1826)
);

OAI22xp33_ASAP7_75t_L g1827 ( 
.A1(n_1701),
.A2(n_1447),
.B1(n_1565),
.B2(n_1455),
.Y(n_1827)
);

OAI221xp5_ASAP7_75t_L g1828 ( 
.A1(n_1630),
.A2(n_1409),
.B1(n_1514),
.B2(n_1455),
.C(n_1463),
.Y(n_1828)
);

AOI22xp33_ASAP7_75t_L g1829 ( 
.A1(n_1621),
.A2(n_1463),
.B1(n_1467),
.B2(n_1409),
.Y(n_1829)
);

INVx3_ASAP7_75t_L g1830 ( 
.A(n_1582),
.Y(n_1830)
);

AOI22xp33_ASAP7_75t_SL g1831 ( 
.A1(n_1657),
.A2(n_1659),
.B1(n_1569),
.B2(n_1722),
.Y(n_1831)
);

AOI221xp5_ASAP7_75t_L g1832 ( 
.A1(n_1703),
.A2(n_1467),
.B1(n_1447),
.B2(n_1515),
.C(n_1478),
.Y(n_1832)
);

INVxp67_ASAP7_75t_L g1833 ( 
.A(n_1623),
.Y(n_1833)
);

AOI33xp33_ASAP7_75t_L g1834 ( 
.A1(n_1689),
.A2(n_1478),
.A3(n_1515),
.B1(n_1565),
.B2(n_1737),
.B3(n_1729),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1633),
.A2(n_1741),
.B1(n_1667),
.B2(n_1722),
.Y(n_1835)
);

HB1xp67_ASAP7_75t_L g1836 ( 
.A(n_1646),
.Y(n_1836)
);

AOI22xp33_ASAP7_75t_L g1837 ( 
.A1(n_1722),
.A2(n_1615),
.B1(n_1683),
.B2(n_1686),
.Y(n_1837)
);

AOI22xp33_ASAP7_75t_L g1838 ( 
.A1(n_1608),
.A2(n_1693),
.B1(n_1691),
.B2(n_1583),
.Y(n_1838)
);

INVx4_ASAP7_75t_L g1839 ( 
.A(n_1715),
.Y(n_1839)
);

NAND3xp33_ASAP7_75t_SL g1840 ( 
.A(n_1585),
.B(n_1706),
.C(n_1668),
.Y(n_1840)
);

CKINVDCx5p33_ASAP7_75t_R g1841 ( 
.A(n_1577),
.Y(n_1841)
);

BUFx6f_ASAP7_75t_L g1842 ( 
.A(n_1721),
.Y(n_1842)
);

AOI221xp5_ASAP7_75t_L g1843 ( 
.A1(n_1642),
.A2(n_1586),
.B1(n_1576),
.B2(n_1614),
.C(n_1617),
.Y(n_1843)
);

AOI22xp33_ASAP7_75t_SL g1844 ( 
.A1(n_1700),
.A2(n_1751),
.B1(n_1717),
.B2(n_1670),
.Y(n_1844)
);

AOI21xp5_ASAP7_75t_L g1845 ( 
.A1(n_1613),
.A2(n_1590),
.B(n_1752),
.Y(n_1845)
);

AOI22xp33_ASAP7_75t_L g1846 ( 
.A1(n_1608),
.A2(n_1719),
.B1(n_1712),
.B2(n_1752),
.Y(n_1846)
);

BUFx4f_ASAP7_75t_L g1847 ( 
.A(n_1709),
.Y(n_1847)
);

AOI22xp33_ASAP7_75t_L g1848 ( 
.A1(n_1608),
.A2(n_1712),
.B1(n_1744),
.B2(n_1640),
.Y(n_1848)
);

INVx4_ASAP7_75t_L g1849 ( 
.A(n_1769),
.Y(n_1849)
);

AOI22xp33_ASAP7_75t_L g1850 ( 
.A1(n_1712),
.A2(n_1640),
.B1(n_1677),
.B2(n_1694),
.Y(n_1850)
);

AOI22xp33_ASAP7_75t_L g1851 ( 
.A1(n_1677),
.A2(n_1694),
.B1(n_1702),
.B2(n_1749),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1599),
.Y(n_1852)
);

AOI221xp5_ASAP7_75t_L g1853 ( 
.A1(n_1642),
.A2(n_1612),
.B1(n_1679),
.B2(n_1651),
.C(n_1652),
.Y(n_1853)
);

OAI22xp33_ASAP7_75t_L g1854 ( 
.A1(n_1620),
.A2(n_1670),
.B1(n_1665),
.B2(n_1638),
.Y(n_1854)
);

AOI22xp33_ASAP7_75t_L g1855 ( 
.A1(n_1702),
.A2(n_1749),
.B1(n_1634),
.B2(n_1602),
.Y(n_1855)
);

AOI22xp33_ASAP7_75t_L g1856 ( 
.A1(n_1749),
.A2(n_1602),
.B1(n_1711),
.B2(n_1622),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1587),
.B(n_1591),
.Y(n_1857)
);

OAI22xp33_ASAP7_75t_L g1858 ( 
.A1(n_1665),
.A2(n_1649),
.B1(n_1592),
.B2(n_1644),
.Y(n_1858)
);

OAI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1654),
.A2(n_1721),
.B1(n_1740),
.B2(n_1728),
.Y(n_1859)
);

AOI21xp5_ASAP7_75t_L g1860 ( 
.A1(n_1699),
.A2(n_1764),
.B(n_1708),
.Y(n_1860)
);

OAI211xp5_ASAP7_75t_SL g1861 ( 
.A1(n_1732),
.A2(n_1577),
.B(n_1579),
.C(n_1745),
.Y(n_1861)
);

AOI22xp33_ASAP7_75t_L g1862 ( 
.A1(n_1602),
.A2(n_1622),
.B1(n_1635),
.B2(n_1672),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1581),
.B(n_1598),
.Y(n_1863)
);

AOI22xp33_ASAP7_75t_SL g1864 ( 
.A1(n_1717),
.A2(n_1622),
.B1(n_1672),
.B2(n_1711),
.Y(n_1864)
);

AND2x4_ASAP7_75t_L g1865 ( 
.A(n_1684),
.B(n_1604),
.Y(n_1865)
);

AOI21xp5_ASAP7_75t_L g1866 ( 
.A1(n_1764),
.A2(n_1748),
.B(n_1757),
.Y(n_1866)
);

OAI22xp5_ASAP7_75t_L g1867 ( 
.A1(n_1654),
.A2(n_1728),
.B1(n_1740),
.B2(n_1578),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1688),
.B(n_1581),
.Y(n_1868)
);

INVx11_ASAP7_75t_L g1869 ( 
.A(n_1769),
.Y(n_1869)
);

OAI221xp5_ASAP7_75t_L g1870 ( 
.A1(n_1570),
.A2(n_1592),
.B1(n_1762),
.B2(n_1760),
.C(n_1602),
.Y(n_1870)
);

OAI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1684),
.A2(n_1764),
.B1(n_1662),
.B2(n_1765),
.Y(n_1871)
);

INVx3_ASAP7_75t_L g1872 ( 
.A(n_1755),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1598),
.B(n_1603),
.Y(n_1873)
);

NOR2xp33_ASAP7_75t_L g1874 ( 
.A(n_1648),
.B(n_1663),
.Y(n_1874)
);

OAI22xp5_ASAP7_75t_L g1875 ( 
.A1(n_1750),
.A2(n_1765),
.B1(n_1764),
.B2(n_1768),
.Y(n_1875)
);

OAI22x1_ASAP7_75t_L g1876 ( 
.A1(n_1747),
.A2(n_1758),
.B1(n_1756),
.B2(n_1766),
.Y(n_1876)
);

OAI21xp5_ASAP7_75t_L g1877 ( 
.A1(n_1648),
.A2(n_1663),
.B(n_1738),
.Y(n_1877)
);

OAI33xp33_ASAP7_75t_L g1878 ( 
.A1(n_1616),
.A2(n_1690),
.A3(n_1643),
.B1(n_1639),
.B2(n_1664),
.B3(n_1671),
.Y(n_1878)
);

OR2x6_ASAP7_75t_L g1879 ( 
.A(n_1619),
.B(n_1604),
.Y(n_1879)
);

AO21x2_ASAP7_75t_L g1880 ( 
.A1(n_1609),
.A2(n_1632),
.B(n_1767),
.Y(n_1880)
);

BUFx6f_ASAP7_75t_L g1881 ( 
.A(n_1601),
.Y(n_1881)
);

AOI22xp33_ASAP7_75t_L g1882 ( 
.A1(n_1635),
.A2(n_1672),
.B1(n_1711),
.B2(n_1755),
.Y(n_1882)
);

OAI22xp33_ASAP7_75t_L g1883 ( 
.A1(n_1662),
.A2(n_1750),
.B1(n_1698),
.B2(n_1695),
.Y(n_1883)
);

AOI22xp33_ASAP7_75t_L g1884 ( 
.A1(n_1635),
.A2(n_1619),
.B1(n_1766),
.B2(n_1756),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1618),
.Y(n_1885)
);

OAI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1754),
.A2(n_1650),
.B1(n_1681),
.B2(n_1624),
.Y(n_1886)
);

AOI322xp5_ASAP7_75t_L g1887 ( 
.A1(n_1704),
.A2(n_1727),
.A3(n_1725),
.B1(n_1730),
.B2(n_1746),
.C1(n_1759),
.C2(n_1676),
.Y(n_1887)
);

AOI22xp33_ASAP7_75t_SL g1888 ( 
.A1(n_1738),
.A2(n_1632),
.B1(n_1647),
.B2(n_1669),
.Y(n_1888)
);

NOR2x1_ASAP7_75t_SL g1889 ( 
.A(n_1632),
.B(n_1753),
.Y(n_1889)
);

AOI21xp5_ASAP7_75t_L g1890 ( 
.A1(n_1767),
.A2(n_1753),
.B(n_1720),
.Y(n_1890)
);

BUFx2_ASAP7_75t_L g1891 ( 
.A(n_1763),
.Y(n_1891)
);

OAI211xp5_ASAP7_75t_SL g1892 ( 
.A1(n_1761),
.A2(n_1676),
.B(n_1710),
.C(n_1685),
.Y(n_1892)
);

OAI211xp5_ASAP7_75t_SL g1893 ( 
.A1(n_1636),
.A2(n_1685),
.B(n_1710),
.C(n_1655),
.Y(n_1893)
);

INVx3_ASAP7_75t_L g1894 ( 
.A(n_1655),
.Y(n_1894)
);

AOI22xp33_ASAP7_75t_L g1895 ( 
.A1(n_1770),
.A2(n_1771),
.B1(n_1666),
.B2(n_1669),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1666),
.B(n_1568),
.Y(n_1896)
);

OAI22xp5_ASAP7_75t_L g1897 ( 
.A1(n_1709),
.A2(n_1669),
.B1(n_1641),
.B2(n_1607),
.Y(n_1897)
);

OAI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1607),
.A2(n_1641),
.B1(n_1771),
.B2(n_1697),
.Y(n_1898)
);

BUFx4f_ASAP7_75t_SL g1899 ( 
.A(n_1763),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1568),
.Y(n_1900)
);

AOI22xp33_ASAP7_75t_L g1901 ( 
.A1(n_1770),
.A2(n_1771),
.B1(n_1641),
.B2(n_1607),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1575),
.Y(n_1902)
);

AOI221xp5_ASAP7_75t_L g1903 ( 
.A1(n_1588),
.A2(n_1589),
.B1(n_1631),
.B2(n_1626),
.C(n_1716),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1589),
.B(n_1631),
.Y(n_1904)
);

AOI22xp33_ASAP7_75t_SL g1905 ( 
.A1(n_1647),
.A2(n_1629),
.B1(n_1601),
.B2(n_1713),
.Y(n_1905)
);

OAI22xp33_ASAP7_75t_L g1906 ( 
.A1(n_1601),
.A2(n_1629),
.B1(n_1713),
.B2(n_1680),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1626),
.B(n_1573),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1573),
.B(n_1610),
.Y(n_1908)
);

OAI22xp5_ASAP7_75t_L g1909 ( 
.A1(n_1680),
.A2(n_1713),
.B1(n_1697),
.B2(n_1629),
.Y(n_1909)
);

AOI22xp33_ASAP7_75t_L g1910 ( 
.A1(n_1680),
.A2(n_1697),
.B1(n_1601),
.B2(n_1629),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_SL g1911 ( 
.A(n_1734),
.B(n_1714),
.Y(n_1911)
);

AOI211xp5_ASAP7_75t_L g1912 ( 
.A1(n_1734),
.A2(n_1714),
.B(n_1716),
.C(n_1720),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1734),
.B(n_1573),
.Y(n_1913)
);

OAI22xp33_ASAP7_75t_L g1914 ( 
.A1(n_1734),
.A2(n_1723),
.B1(n_1724),
.B2(n_1731),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1723),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1573),
.B(n_1610),
.Y(n_1916)
);

OAI33xp33_ASAP7_75t_L g1917 ( 
.A1(n_1724),
.A2(n_1682),
.A3(n_1594),
.B1(n_1475),
.B2(n_1011),
.B3(n_1656),
.Y(n_1917)
);

AOI21x1_ASAP7_75t_L g1918 ( 
.A1(n_1731),
.A2(n_1753),
.B(n_1610),
.Y(n_1918)
);

INVx4_ASAP7_75t_L g1919 ( 
.A(n_1610),
.Y(n_1919)
);

BUFx3_ASAP7_75t_L g1920 ( 
.A(n_1678),
.Y(n_1920)
);

AOI22xp33_ASAP7_75t_L g1921 ( 
.A1(n_1696),
.A2(n_877),
.B1(n_880),
.B2(n_1658),
.Y(n_1921)
);

OAI221xp5_ASAP7_75t_L g1922 ( 
.A1(n_1584),
.A2(n_745),
.B1(n_1159),
.B2(n_891),
.C(n_1028),
.Y(n_1922)
);

AOI22xp33_ASAP7_75t_L g1923 ( 
.A1(n_1696),
.A2(n_877),
.B1(n_880),
.B2(n_1658),
.Y(n_1923)
);

AOI22xp33_ASAP7_75t_L g1924 ( 
.A1(n_1696),
.A2(n_877),
.B1(n_880),
.B2(n_1658),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1623),
.B(n_1699),
.Y(n_1925)
);

INVx1_ASAP7_75t_SL g1926 ( 
.A(n_1627),
.Y(n_1926)
);

OAI21x1_ASAP7_75t_L g1927 ( 
.A1(n_1590),
.A2(n_1412),
.B(n_1399),
.Y(n_1927)
);

INVx4_ASAP7_75t_L g1928 ( 
.A(n_1715),
.Y(n_1928)
);

AOI22xp5_ASAP7_75t_L g1929 ( 
.A1(n_1584),
.A2(n_880),
.B1(n_877),
.B2(n_1028),
.Y(n_1929)
);

AOI22xp33_ASAP7_75t_L g1930 ( 
.A1(n_1696),
.A2(n_877),
.B1(n_880),
.B2(n_1658),
.Y(n_1930)
);

AND2x4_ASAP7_75t_L g1931 ( 
.A(n_1582),
.B(n_1608),
.Y(n_1931)
);

AOI22xp33_ASAP7_75t_L g1932 ( 
.A1(n_1696),
.A2(n_877),
.B1(n_880),
.B2(n_1658),
.Y(n_1932)
);

AOI221xp5_ASAP7_75t_L g1933 ( 
.A1(n_1584),
.A2(n_1028),
.B1(n_758),
.B2(n_766),
.C(n_745),
.Y(n_1933)
);

AOI22xp5_ASAP7_75t_L g1934 ( 
.A1(n_1584),
.A2(n_880),
.B1(n_877),
.B2(n_1028),
.Y(n_1934)
);

AOI22xp33_ASAP7_75t_SL g1935 ( 
.A1(n_1696),
.A2(n_1584),
.B1(n_1733),
.B2(n_1658),
.Y(n_1935)
);

NAND3xp33_ASAP7_75t_L g1936 ( 
.A(n_1742),
.B(n_880),
.C(n_877),
.Y(n_1936)
);

AOI22xp5_ASAP7_75t_L g1937 ( 
.A1(n_1584),
.A2(n_880),
.B1(n_877),
.B2(n_1028),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1571),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_SL g1939 ( 
.A(n_1742),
.B(n_1027),
.Y(n_1939)
);

CKINVDCx5p33_ASAP7_75t_R g1940 ( 
.A(n_1577),
.Y(n_1940)
);

OR2x2_ASAP7_75t_L g1941 ( 
.A(n_1580),
.B(n_1587),
.Y(n_1941)
);

OAI22xp5_ASAP7_75t_L g1942 ( 
.A1(n_1605),
.A2(n_880),
.B1(n_877),
.B2(n_1028),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1739),
.B(n_1634),
.Y(n_1943)
);

AOI22xp33_ASAP7_75t_L g1944 ( 
.A1(n_1696),
.A2(n_877),
.B1(n_880),
.B2(n_1658),
.Y(n_1944)
);

AND2x4_ASAP7_75t_L g1945 ( 
.A(n_1582),
.B(n_1608),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1571),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1739),
.B(n_1634),
.Y(n_1947)
);

OAI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1605),
.A2(n_880),
.B1(n_877),
.B2(n_1028),
.Y(n_1948)
);

INVx4_ASAP7_75t_L g1949 ( 
.A(n_1715),
.Y(n_1949)
);

INVxp67_ASAP7_75t_L g1950 ( 
.A(n_1653),
.Y(n_1950)
);

OA21x2_ASAP7_75t_L g1951 ( 
.A1(n_1757),
.A2(n_1590),
.B(n_1613),
.Y(n_1951)
);

OAI221xp5_ASAP7_75t_L g1952 ( 
.A1(n_1584),
.A2(n_745),
.B1(n_1159),
.B2(n_891),
.C(n_1028),
.Y(n_1952)
);

AOI22xp33_ASAP7_75t_L g1953 ( 
.A1(n_1696),
.A2(n_877),
.B1(n_880),
.B2(n_1658),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1623),
.B(n_1699),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1571),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1739),
.B(n_1634),
.Y(n_1956)
);

OAI22xp33_ASAP7_75t_L g1957 ( 
.A1(n_1726),
.A2(n_1019),
.B1(n_1246),
.B2(n_611),
.Y(n_1957)
);

AND2x4_ASAP7_75t_L g1958 ( 
.A(n_1812),
.B(n_1821),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1941),
.B(n_1857),
.Y(n_1959)
);

HB1xp67_ASAP7_75t_L g1960 ( 
.A(n_1913),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1879),
.B(n_1863),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1777),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1879),
.B(n_1863),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1915),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1915),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1941),
.B(n_1857),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1918),
.Y(n_1967)
);

BUFx6f_ASAP7_75t_L g1968 ( 
.A(n_1805),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1925),
.B(n_1954),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1873),
.B(n_1803),
.Y(n_1970)
);

INVx3_ASAP7_75t_L g1971 ( 
.A(n_1812),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1806),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1879),
.B(n_1813),
.Y(n_1973)
);

INVx1_ASAP7_75t_SL g1974 ( 
.A(n_1836),
.Y(n_1974)
);

INVxp67_ASAP7_75t_SL g1975 ( 
.A(n_1890),
.Y(n_1975)
);

BUFx2_ASAP7_75t_L g1976 ( 
.A(n_1879),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1813),
.B(n_1872),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1815),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1819),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1872),
.B(n_1812),
.Y(n_1980)
);

OR2x2_ASAP7_75t_L g1981 ( 
.A(n_1823),
.B(n_1868),
.Y(n_1981)
);

HB1xp67_ASAP7_75t_L g1982 ( 
.A(n_1907),
.Y(n_1982)
);

CKINVDCx16_ASAP7_75t_R g1983 ( 
.A(n_1807),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1872),
.B(n_1821),
.Y(n_1984)
);

OR2x2_ASAP7_75t_L g1985 ( 
.A(n_1823),
.B(n_1876),
.Y(n_1985)
);

BUFx2_ASAP7_75t_L g1986 ( 
.A(n_1865),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1852),
.Y(n_1987)
);

NAND2x1_ASAP7_75t_L g1988 ( 
.A(n_1802),
.B(n_1845),
.Y(n_1988)
);

BUFx6f_ASAP7_75t_L g1989 ( 
.A(n_1881),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1821),
.B(n_1830),
.Y(n_1990)
);

INVx1_ASAP7_75t_SL g1991 ( 
.A(n_1809),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1885),
.Y(n_1992)
);

AND2x2_ASAP7_75t_SL g1993 ( 
.A(n_1921),
.B(n_1923),
.Y(n_1993)
);

BUFx2_ASAP7_75t_L g1994 ( 
.A(n_1865),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1938),
.B(n_1946),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1955),
.B(n_1826),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1907),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1931),
.B(n_1945),
.Y(n_1998)
);

BUFx3_ASAP7_75t_L g1999 ( 
.A(n_1779),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1945),
.B(n_1865),
.Y(n_2000)
);

OR2x2_ASAP7_75t_L g2001 ( 
.A(n_1876),
.B(n_1866),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1826),
.Y(n_2002)
);

INVx3_ASAP7_75t_L g2003 ( 
.A(n_1945),
.Y(n_2003)
);

INVx4_ASAP7_75t_L g2004 ( 
.A(n_1842),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1887),
.B(n_1896),
.Y(n_2005)
);

AND2x4_ASAP7_75t_SL g2006 ( 
.A(n_1842),
.B(n_1862),
.Y(n_2006)
);

OR2x2_ASAP7_75t_L g2007 ( 
.A(n_1919),
.B(n_1908),
.Y(n_2007)
);

INVxp67_ASAP7_75t_SL g2008 ( 
.A(n_1889),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1896),
.B(n_1894),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1791),
.B(n_1943),
.Y(n_2010)
);

AOI22xp33_ASAP7_75t_L g2011 ( 
.A1(n_1942),
.A2(n_1948),
.B1(n_1953),
.B2(n_1930),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1908),
.Y(n_2012)
);

AND2x4_ASAP7_75t_L g2013 ( 
.A(n_1825),
.B(n_1911),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1833),
.B(n_1886),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1791),
.B(n_1943),
.Y(n_2015)
);

BUFx3_ASAP7_75t_L g2016 ( 
.A(n_1779),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1916),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1916),
.Y(n_2018)
);

OR2x2_ASAP7_75t_L g2019 ( 
.A(n_1919),
.B(n_1947),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1900),
.Y(n_2020)
);

OR2x2_ASAP7_75t_L g2021 ( 
.A(n_1947),
.B(n_1956),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1904),
.B(n_1902),
.Y(n_2022)
);

INVx2_ASAP7_75t_SL g2023 ( 
.A(n_1911),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1956),
.B(n_1884),
.Y(n_2024)
);

BUFx6f_ASAP7_75t_L g2025 ( 
.A(n_1881),
.Y(n_2025)
);

AOI221xp5_ASAP7_75t_L g2026 ( 
.A1(n_1924),
.A2(n_1932),
.B1(n_1944),
.B2(n_1952),
.C(n_1922),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1904),
.Y(n_2027)
);

INVx3_ASAP7_75t_L g2028 ( 
.A(n_1927),
.Y(n_2028)
);

BUFx3_ASAP7_75t_L g2029 ( 
.A(n_1800),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1893),
.Y(n_2030)
);

INVx3_ASAP7_75t_L g2031 ( 
.A(n_1927),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1855),
.B(n_1880),
.Y(n_2032)
);

AND2x4_ASAP7_75t_L g2033 ( 
.A(n_1796),
.B(n_1797),
.Y(n_2033)
);

AND2x4_ASAP7_75t_SL g2034 ( 
.A(n_1842),
.B(n_1882),
.Y(n_2034)
);

INVx2_ASAP7_75t_SL g2035 ( 
.A(n_1796),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1880),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1880),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1912),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1864),
.B(n_1848),
.Y(n_2039)
);

AND2x4_ASAP7_75t_L g2040 ( 
.A(n_1797),
.B(n_1808),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_1856),
.B(n_1775),
.Y(n_2041)
);

OAI22xp33_ASAP7_75t_L g2042 ( 
.A1(n_1929),
.A2(n_1937),
.B1(n_1934),
.B2(n_1957),
.Y(n_2042)
);

OAI22xp5_ASAP7_75t_L g2043 ( 
.A1(n_1935),
.A2(n_1835),
.B1(n_1936),
.B2(n_1810),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1951),
.Y(n_2044)
);

AOI221xp5_ASAP7_75t_L g2045 ( 
.A1(n_1917),
.A2(n_1933),
.B1(n_1840),
.B2(n_1804),
.C(n_1853),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1914),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1951),
.Y(n_2047)
);

NOR2xp33_ASAP7_75t_L g2048 ( 
.A(n_1781),
.B(n_1926),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_1951),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1903),
.Y(n_2050)
);

HB1xp67_ASAP7_75t_L g2051 ( 
.A(n_1950),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1874),
.B(n_1844),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_1874),
.B(n_1877),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1827),
.Y(n_2054)
);

AOI222xp33_ASAP7_75t_L g2055 ( 
.A1(n_1837),
.A2(n_1843),
.B1(n_1838),
.B2(n_1867),
.C1(n_1939),
.C2(n_1859),
.Y(n_2055)
);

BUFx3_ASAP7_75t_L g2056 ( 
.A(n_1800),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1784),
.B(n_1789),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1892),
.Y(n_2058)
);

NOR2xp33_ASAP7_75t_L g2059 ( 
.A(n_1790),
.B(n_1816),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_SL g2060 ( 
.A(n_1854),
.B(n_1831),
.Y(n_2060)
);

HB1xp67_ASAP7_75t_L g2061 ( 
.A(n_1824),
.Y(n_2061)
);

INVxp67_ASAP7_75t_L g2062 ( 
.A(n_1878),
.Y(n_2062)
);

NOR2xp33_ASAP7_75t_L g2063 ( 
.A(n_1816),
.B(n_1841),
.Y(n_2063)
);

NAND2xp33_ASAP7_75t_R g2064 ( 
.A(n_1841),
.B(n_1940),
.Y(n_2064)
);

BUFx3_ASAP7_75t_L g2065 ( 
.A(n_1920),
.Y(n_2065)
);

AND2x4_ASAP7_75t_SL g2066 ( 
.A(n_1842),
.B(n_1807),
.Y(n_2066)
);

INVx1_ASAP7_75t_SL g2067 ( 
.A(n_1891),
.Y(n_2067)
);

NOR2xp33_ASAP7_75t_L g2068 ( 
.A(n_1940),
.B(n_1858),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1828),
.Y(n_2069)
);

AND2x4_ASAP7_75t_L g2070 ( 
.A(n_1808),
.B(n_1860),
.Y(n_2070)
);

OR2x2_ASAP7_75t_L g2071 ( 
.A(n_1792),
.B(n_1875),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_1783),
.B(n_1772),
.Y(n_2072)
);

OR2x2_ASAP7_75t_L g2073 ( 
.A(n_1959),
.B(n_1814),
.Y(n_2073)
);

BUFx3_ASAP7_75t_L g2074 ( 
.A(n_1999),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_1969),
.B(n_1871),
.Y(n_2075)
);

AOI221xp5_ASAP7_75t_L g2076 ( 
.A1(n_2043),
.A2(n_2042),
.B1(n_2045),
.B2(n_2011),
.C(n_2026),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1962),
.Y(n_2077)
);

NOR4xp25_ASAP7_75t_SL g2078 ( 
.A(n_2064),
.B(n_2060),
.C(n_2045),
.D(n_1870),
.Y(n_2078)
);

OAI33xp33_ASAP7_75t_L g2079 ( 
.A1(n_2043),
.A2(n_1883),
.A3(n_1939),
.B1(n_1785),
.B2(n_1794),
.B3(n_1780),
.Y(n_2079)
);

OAI33xp33_ASAP7_75t_L g2080 ( 
.A1(n_2042),
.A2(n_1861),
.A3(n_1798),
.B1(n_1906),
.B2(n_1898),
.B3(n_1909),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_1961),
.B(n_1778),
.Y(n_2081)
);

AOI31xp33_ASAP7_75t_L g2082 ( 
.A1(n_2026),
.A2(n_1846),
.A3(n_1776),
.B(n_1850),
.Y(n_2082)
);

AOI22xp33_ASAP7_75t_L g2083 ( 
.A1(n_1993),
.A2(n_1778),
.B1(n_1928),
.B2(n_1949),
.Y(n_2083)
);

OAI211xp5_ASAP7_75t_L g2084 ( 
.A1(n_2011),
.A2(n_1786),
.B(n_1773),
.C(n_1782),
.Y(n_2084)
);

INVx2_ASAP7_75t_L g2085 ( 
.A(n_1964),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1969),
.B(n_1778),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_1991),
.B(n_1778),
.Y(n_2087)
);

OAI22xp5_ASAP7_75t_L g2088 ( 
.A1(n_1993),
.A2(n_2071),
.B1(n_1851),
.B2(n_2068),
.Y(n_2088)
);

NOR2xp33_ASAP7_75t_L g2089 ( 
.A(n_2048),
.B(n_1949),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1962),
.Y(n_2090)
);

OAI33xp33_ASAP7_75t_L g2091 ( 
.A1(n_2062),
.A2(n_1897),
.A3(n_1834),
.B1(n_1949),
.B2(n_1839),
.B3(n_1928),
.Y(n_2091)
);

OR2x2_ASAP7_75t_L g2092 ( 
.A(n_1959),
.B(n_1799),
.Y(n_2092)
);

OAI22xp5_ASAP7_75t_L g2093 ( 
.A1(n_1993),
.A2(n_2071),
.B1(n_1928),
.B2(n_1839),
.Y(n_2093)
);

AOI33xp33_ASAP7_75t_L g2094 ( 
.A1(n_1991),
.A2(n_2054),
.A3(n_1974),
.B1(n_2070),
.B2(n_2038),
.B3(n_2053),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1972),
.Y(n_2095)
);

OAI22xp5_ASAP7_75t_L g2096 ( 
.A1(n_1983),
.A2(n_1839),
.B1(n_1787),
.B2(n_1807),
.Y(n_2096)
);

NAND4xp25_ASAP7_75t_SL g2097 ( 
.A(n_2055),
.B(n_2001),
.C(n_2052),
.D(n_2053),
.Y(n_2097)
);

BUFx2_ASAP7_75t_L g2098 ( 
.A(n_2013),
.Y(n_2098)
);

AO21x2_ASAP7_75t_L g2099 ( 
.A1(n_2037),
.A2(n_1824),
.B(n_1788),
.Y(n_2099)
);

AOI22xp33_ASAP7_75t_L g2100 ( 
.A1(n_2055),
.A2(n_1807),
.B1(n_1920),
.B2(n_1847),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1966),
.B(n_1834),
.Y(n_2101)
);

OAI211xp5_ASAP7_75t_SL g2102 ( 
.A1(n_2062),
.A2(n_1895),
.B(n_1901),
.C(n_1910),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_1966),
.B(n_1820),
.Y(n_2103)
);

AOI22xp5_ASAP7_75t_L g2104 ( 
.A1(n_2039),
.A2(n_1774),
.B1(n_1849),
.B2(n_1847),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1972),
.Y(n_2105)
);

BUFx3_ASAP7_75t_L g2106 ( 
.A(n_1999),
.Y(n_2106)
);

AOI221xp5_ASAP7_75t_L g2107 ( 
.A1(n_2054),
.A2(n_1801),
.B1(n_1793),
.B2(n_1817),
.C(n_1832),
.Y(n_2107)
);

AOI211xp5_ASAP7_75t_L g2108 ( 
.A1(n_2070),
.A2(n_1881),
.B(n_1869),
.C(n_1905),
.Y(n_2108)
);

INVx3_ASAP7_75t_SL g2109 ( 
.A(n_1983),
.Y(n_2109)
);

AOI22xp33_ASAP7_75t_L g2110 ( 
.A1(n_2039),
.A2(n_1847),
.B1(n_1849),
.B2(n_1899),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_1964),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_1961),
.B(n_1795),
.Y(n_2112)
);

INVxp67_ASAP7_75t_L g2113 ( 
.A(n_2051),
.Y(n_2113)
);

OAI221xp5_ASAP7_75t_L g2114 ( 
.A1(n_1988),
.A2(n_1888),
.B1(n_1849),
.B2(n_1818),
.C(n_1811),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_1964),
.Y(n_2115)
);

NAND4xp25_ASAP7_75t_L g2116 ( 
.A(n_2014),
.B(n_1829),
.C(n_1822),
.D(n_1869),
.Y(n_2116)
);

AOI221xp5_ASAP7_75t_L g2117 ( 
.A1(n_2069),
.A2(n_2014),
.B1(n_2070),
.B2(n_2051),
.C(n_2061),
.Y(n_2117)
);

INVxp67_ASAP7_75t_L g2118 ( 
.A(n_1974),
.Y(n_2118)
);

AOI22xp33_ASAP7_75t_L g2119 ( 
.A1(n_2041),
.A2(n_1881),
.B1(n_2057),
.B2(n_2072),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_1963),
.B(n_1977),
.Y(n_2120)
);

BUFx2_ASAP7_75t_L g2121 ( 
.A(n_2013),
.Y(n_2121)
);

OAI211xp5_ASAP7_75t_L g2122 ( 
.A1(n_1988),
.A2(n_2061),
.B(n_2001),
.C(n_2069),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_1963),
.B(n_1977),
.Y(n_2123)
);

OAI31xp33_ASAP7_75t_SL g2124 ( 
.A1(n_2052),
.A2(n_2070),
.A3(n_2057),
.B(n_2041),
.Y(n_2124)
);

AND2x4_ASAP7_75t_L g2125 ( 
.A(n_1976),
.B(n_2003),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1978),
.Y(n_2126)
);

AOI22xp33_ASAP7_75t_L g2127 ( 
.A1(n_2072),
.A2(n_2034),
.B1(n_2069),
.B2(n_2006),
.Y(n_2127)
);

HB1xp67_ASAP7_75t_L g2128 ( 
.A(n_1960),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_SL g2129 ( 
.A(n_1968),
.B(n_2058),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_1973),
.B(n_1976),
.Y(n_2130)
);

AOI22xp33_ASAP7_75t_SL g2131 ( 
.A1(n_2034),
.A2(n_2006),
.B1(n_2032),
.B2(n_1968),
.Y(n_2131)
);

INVx2_ASAP7_75t_SL g2132 ( 
.A(n_1999),
.Y(n_2132)
);

OAI22xp5_ASAP7_75t_L g2133 ( 
.A1(n_2034),
.A2(n_2006),
.B1(n_2058),
.B2(n_2005),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1978),
.Y(n_2134)
);

CKINVDCx5p33_ASAP7_75t_R g2135 ( 
.A(n_2059),
.Y(n_2135)
);

AOI221xp5_ASAP7_75t_L g2136 ( 
.A1(n_2050),
.A2(n_2032),
.B1(n_1975),
.B2(n_2046),
.C(n_2038),
.Y(n_2136)
);

OAI33xp33_ASAP7_75t_L g2137 ( 
.A1(n_2012),
.A2(n_2018),
.A3(n_2017),
.B1(n_2005),
.B2(n_1970),
.B3(n_2030),
.Y(n_2137)
);

OAI21xp5_ASAP7_75t_L g2138 ( 
.A1(n_2050),
.A2(n_2030),
.B(n_1975),
.Y(n_2138)
);

OAI221xp5_ASAP7_75t_L g2139 ( 
.A1(n_2063),
.A2(n_2046),
.B1(n_2008),
.B2(n_1968),
.C(n_2067),
.Y(n_2139)
);

OAI21x1_ASAP7_75t_L g2140 ( 
.A1(n_2028),
.A2(n_2031),
.B(n_2044),
.Y(n_2140)
);

OAI33xp33_ASAP7_75t_L g2141 ( 
.A1(n_2012),
.A2(n_2018),
.A3(n_2017),
.B1(n_1970),
.B2(n_1995),
.B3(n_1992),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1979),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_1973),
.B(n_1986),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_1986),
.B(n_1994),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_1979),
.Y(n_2145)
);

OAI31xp33_ASAP7_75t_L g2146 ( 
.A1(n_2040),
.A2(n_2066),
.A3(n_2067),
.B(n_2033),
.Y(n_2146)
);

OAI221xp5_ASAP7_75t_L g2147 ( 
.A1(n_2008),
.A2(n_1968),
.B1(n_1985),
.B2(n_2035),
.C(n_2004),
.Y(n_2147)
);

BUFx2_ASAP7_75t_L g2148 ( 
.A(n_2013),
.Y(n_2148)
);

INVxp67_ASAP7_75t_SL g2149 ( 
.A(n_1960),
.Y(n_2149)
);

NOR4xp25_ASAP7_75t_SL g2150 ( 
.A(n_1994),
.B(n_1992),
.C(n_1987),
.D(n_2002),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_1965),
.Y(n_2151)
);

AOI22xp5_ASAP7_75t_L g2152 ( 
.A1(n_2024),
.A2(n_2066),
.B1(n_1968),
.B2(n_2004),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_1965),
.Y(n_2153)
);

OR2x2_ASAP7_75t_L g2154 ( 
.A(n_1981),
.B(n_1985),
.Y(n_2154)
);

AOI22xp33_ASAP7_75t_L g2155 ( 
.A1(n_2024),
.A2(n_1968),
.B1(n_2040),
.B2(n_2033),
.Y(n_2155)
);

AOI221xp5_ASAP7_75t_L g2156 ( 
.A1(n_1987),
.A2(n_1995),
.B1(n_2040),
.B2(n_2010),
.C(n_2015),
.Y(n_2156)
);

AOI22xp33_ASAP7_75t_L g2157 ( 
.A1(n_2040),
.A2(n_2033),
.B1(n_1980),
.B2(n_1984),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_1965),
.Y(n_2158)
);

INVxp67_ASAP7_75t_L g2159 ( 
.A(n_1981),
.Y(n_2159)
);

OAI22xp5_ASAP7_75t_L g2160 ( 
.A1(n_2021),
.A2(n_2004),
.B1(n_2066),
.B2(n_2003),
.Y(n_2160)
);

OAI33xp33_ASAP7_75t_L g2161 ( 
.A1(n_2007),
.A2(n_1996),
.A3(n_1997),
.B1(n_2022),
.B2(n_2019),
.B3(n_2009),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_2128),
.B(n_2023),
.Y(n_2162)
);

NOR2x1_ASAP7_75t_L g2163 ( 
.A(n_2122),
.B(n_2065),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2077),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2077),
.Y(n_2165)
);

NOR2x1_ASAP7_75t_L g2166 ( 
.A(n_2147),
.B(n_2065),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_2159),
.B(n_2023),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_SL g2168 ( 
.A(n_2124),
.B(n_2094),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_2120),
.B(n_1982),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2090),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2090),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_2120),
.B(n_1982),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_2123),
.B(n_2007),
.Y(n_2173)
);

AND2x2_ASAP7_75t_L g2174 ( 
.A(n_2098),
.B(n_1980),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_2098),
.B(n_1984),
.Y(n_2175)
);

AND2x2_ASAP7_75t_L g2176 ( 
.A(n_2121),
.B(n_2036),
.Y(n_2176)
);

INVxp67_ASAP7_75t_SL g2177 ( 
.A(n_2149),
.Y(n_2177)
);

AND2x4_ASAP7_75t_L g2178 ( 
.A(n_2121),
.B(n_2013),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2095),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_2101),
.B(n_2023),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2095),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2105),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_2148),
.B(n_2036),
.Y(n_2183)
);

INVx1_ASAP7_75t_SL g2184 ( 
.A(n_2129),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_2148),
.B(n_2112),
.Y(n_2185)
);

NOR2x1_ASAP7_75t_L g2186 ( 
.A(n_2138),
.B(n_2065),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2112),
.B(n_2036),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_2143),
.B(n_1990),
.Y(n_2188)
);

INVx1_ASAP7_75t_SL g2189 ( 
.A(n_2144),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_2085),
.Y(n_2190)
);

NOR2xp67_ASAP7_75t_L g2191 ( 
.A(n_2139),
.B(n_2035),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2105),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2126),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2126),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_2154),
.B(n_2027),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_2154),
.B(n_2027),
.Y(n_2196)
);

BUFx2_ASAP7_75t_L g2197 ( 
.A(n_2125),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2134),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_2085),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_2130),
.B(n_2019),
.Y(n_2200)
);

NAND2x1p5_ASAP7_75t_L g2201 ( 
.A(n_2152),
.B(n_1971),
.Y(n_2201)
);

AND2x2_ASAP7_75t_SL g2202 ( 
.A(n_2107),
.B(n_1998),
.Y(n_2202)
);

BUFx2_ASAP7_75t_L g2203 ( 
.A(n_2109),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_2113),
.B(n_2002),
.Y(n_2204)
);

AND2x2_ASAP7_75t_L g2205 ( 
.A(n_2125),
.B(n_2049),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2134),
.Y(n_2206)
);

NOR2xp33_ASAP7_75t_L g2207 ( 
.A(n_2097),
.B(n_2021),
.Y(n_2207)
);

OAI22xp5_ASAP7_75t_L g2208 ( 
.A1(n_2076),
.A2(n_2015),
.B1(n_2010),
.B2(n_2004),
.Y(n_2208)
);

OR2x2_ASAP7_75t_L g2209 ( 
.A(n_2073),
.B(n_2092),
.Y(n_2209)
);

AND2x2_ASAP7_75t_L g2210 ( 
.A(n_2125),
.B(n_2049),
.Y(n_2210)
);

AND2x4_ASAP7_75t_L g2211 ( 
.A(n_2140),
.B(n_2003),
.Y(n_2211)
);

AND2x2_ASAP7_75t_L g2212 ( 
.A(n_2144),
.B(n_2099),
.Y(n_2212)
);

AND2x2_ASAP7_75t_L g2213 ( 
.A(n_2099),
.B(n_2047),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_2099),
.B(n_2047),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_2111),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2142),
.Y(n_2216)
);

OR2x2_ASAP7_75t_L g2217 ( 
.A(n_2073),
.B(n_2009),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2142),
.Y(n_2218)
);

AND2x4_ASAP7_75t_L g2219 ( 
.A(n_2140),
.B(n_2003),
.Y(n_2219)
);

BUFx2_ASAP7_75t_L g2220 ( 
.A(n_2109),
.Y(n_2220)
);

INVxp67_ASAP7_75t_L g2221 ( 
.A(n_2137),
.Y(n_2221)
);

AND2x4_ASAP7_75t_L g2222 ( 
.A(n_2115),
.B(n_1958),
.Y(n_2222)
);

OR2x2_ASAP7_75t_L g2223 ( 
.A(n_2092),
.B(n_1967),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_2151),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2145),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_2103),
.B(n_2020),
.Y(n_2226)
);

OR2x2_ASAP7_75t_L g2227 ( 
.A(n_2209),
.B(n_2118),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_2190),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_2180),
.B(n_2136),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2164),
.Y(n_2230)
);

INVx1_ASAP7_75t_SL g2231 ( 
.A(n_2203),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_2190),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2164),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2165),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2165),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_2185),
.B(n_2109),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2170),
.Y(n_2237)
);

HB1xp67_ASAP7_75t_L g2238 ( 
.A(n_2185),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_2190),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_2199),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_2180),
.B(n_2117),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2170),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2171),
.Y(n_2243)
);

AND2x2_ASAP7_75t_L g2244 ( 
.A(n_2185),
.B(n_2081),
.Y(n_2244)
);

OR2x2_ASAP7_75t_L g2245 ( 
.A(n_2209),
.B(n_2153),
.Y(n_2245)
);

INVx2_ASAP7_75t_L g2246 ( 
.A(n_2199),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2171),
.Y(n_2247)
);

OR3x2_ASAP7_75t_L g2248 ( 
.A(n_2209),
.B(n_2116),
.C(n_2078),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_2226),
.B(n_2075),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_2197),
.B(n_2081),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2226),
.B(n_2156),
.Y(n_2251)
);

HB1xp67_ASAP7_75t_L g2252 ( 
.A(n_2223),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2179),
.Y(n_2253)
);

OR2x2_ASAP7_75t_L g2254 ( 
.A(n_2223),
.B(n_2153),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2179),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_2221),
.B(n_2086),
.Y(n_2256)
);

OR2x6_ASAP7_75t_L g2257 ( 
.A(n_2163),
.B(n_2096),
.Y(n_2257)
);

NAND2x1p5_ASAP7_75t_L g2258 ( 
.A(n_2163),
.B(n_2074),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2221),
.B(n_2119),
.Y(n_2259)
);

OR2x2_ASAP7_75t_L g2260 ( 
.A(n_2223),
.B(n_2158),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_2197),
.B(n_2155),
.Y(n_2261)
);

AND2x2_ASAP7_75t_L g2262 ( 
.A(n_2197),
.B(n_2152),
.Y(n_2262)
);

AND2x4_ASAP7_75t_L g2263 ( 
.A(n_2178),
.B(n_2074),
.Y(n_2263)
);

NAND2xp33_ASAP7_75t_SL g2264 ( 
.A(n_2168),
.B(n_2100),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2217),
.B(n_2087),
.Y(n_2265)
);

OR2x2_ASAP7_75t_L g2266 ( 
.A(n_2217),
.B(n_2158),
.Y(n_2266)
);

OR2x2_ASAP7_75t_L g2267 ( 
.A(n_2217),
.B(n_2145),
.Y(n_2267)
);

OAI22xp5_ASAP7_75t_L g2268 ( 
.A1(n_2168),
.A2(n_2083),
.B1(n_2104),
.B2(n_2082),
.Y(n_2268)
);

OAI21xp33_ASAP7_75t_SL g2269 ( 
.A1(n_2186),
.A2(n_2146),
.B(n_2157),
.Y(n_2269)
);

INVx2_ASAP7_75t_L g2270 ( 
.A(n_2199),
.Y(n_2270)
);

NOR2xp67_ASAP7_75t_L g2271 ( 
.A(n_2191),
.B(n_2135),
.Y(n_2271)
);

OR2x2_ASAP7_75t_L g2272 ( 
.A(n_2195),
.B(n_2132),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_2167),
.B(n_2088),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_2167),
.B(n_2000),
.Y(n_2274)
);

AND2x4_ASAP7_75t_L g2275 ( 
.A(n_2178),
.B(n_2106),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2207),
.B(n_2000),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_2207),
.B(n_2132),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2181),
.Y(n_2278)
);

AND2x2_ASAP7_75t_L g2279 ( 
.A(n_2212),
.B(n_2131),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_2184),
.B(n_2033),
.Y(n_2280)
);

OR2x2_ASAP7_75t_L g2281 ( 
.A(n_2195),
.B(n_2022),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2181),
.Y(n_2282)
);

NAND4xp25_ASAP7_75t_L g2283 ( 
.A(n_2191),
.B(n_2102),
.C(n_2084),
.D(n_2127),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_2258),
.B(n_2212),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2256),
.B(n_2184),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2242),
.Y(n_2286)
);

AND2x2_ASAP7_75t_L g2287 ( 
.A(n_2258),
.B(n_2212),
.Y(n_2287)
);

NOR2xp33_ASAP7_75t_L g2288 ( 
.A(n_2259),
.B(n_2135),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2242),
.Y(n_2289)
);

INVx2_ASAP7_75t_SL g2290 ( 
.A(n_2258),
.Y(n_2290)
);

OR2x2_ASAP7_75t_L g2291 ( 
.A(n_2245),
.B(n_2196),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2243),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2243),
.Y(n_2293)
);

OR2x2_ASAP7_75t_L g2294 ( 
.A(n_2245),
.B(n_2196),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_2279),
.B(n_2203),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2229),
.B(n_2202),
.Y(n_2296)
);

OAI222xp33_ASAP7_75t_L g2297 ( 
.A1(n_2257),
.A2(n_2186),
.B1(n_2208),
.B2(n_2166),
.C1(n_2220),
.C2(n_2201),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2241),
.B(n_2202),
.Y(n_2298)
);

AND2x2_ASAP7_75t_L g2299 ( 
.A(n_2279),
.B(n_2220),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2247),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_2236),
.B(n_2166),
.Y(n_2301)
);

OR2x2_ASAP7_75t_L g2302 ( 
.A(n_2238),
.B(n_2267),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2247),
.Y(n_2303)
);

AOI22xp33_ASAP7_75t_L g2304 ( 
.A1(n_2248),
.A2(n_2079),
.B1(n_2202),
.B2(n_2080),
.Y(n_2304)
);

NOR2xp33_ASAP7_75t_L g2305 ( 
.A(n_2283),
.B(n_2089),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_2228),
.Y(n_2306)
);

AND2x2_ASAP7_75t_SL g2307 ( 
.A(n_2248),
.B(n_2202),
.Y(n_2307)
);

INVxp67_ASAP7_75t_L g2308 ( 
.A(n_2264),
.Y(n_2308)
);

NOR3xp33_ASAP7_75t_L g2309 ( 
.A(n_2264),
.B(n_2093),
.C(n_2091),
.Y(n_2309)
);

INVx1_ASAP7_75t_SL g2310 ( 
.A(n_2231),
.Y(n_2310)
);

NOR2x1_ASAP7_75t_L g2311 ( 
.A(n_2271),
.B(n_2208),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2278),
.Y(n_2312)
);

NAND2x1p5_ASAP7_75t_L g2313 ( 
.A(n_2236),
.B(n_2213),
.Y(n_2313)
);

AND2x4_ASAP7_75t_L g2314 ( 
.A(n_2262),
.B(n_2178),
.Y(n_2314)
);

BUFx3_ASAP7_75t_L g2315 ( 
.A(n_2227),
.Y(n_2315)
);

OAI21xp33_ASAP7_75t_L g2316 ( 
.A1(n_2269),
.A2(n_2201),
.B(n_2213),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2278),
.Y(n_2317)
);

INVx2_ASAP7_75t_SL g2318 ( 
.A(n_2263),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2282),
.Y(n_2319)
);

AND2x2_ASAP7_75t_L g2320 ( 
.A(n_2262),
.B(n_2201),
.Y(n_2320)
);

NOR2x1_ASAP7_75t_L g2321 ( 
.A(n_2257),
.B(n_2162),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2282),
.Y(n_2322)
);

AND2x2_ASAP7_75t_L g2323 ( 
.A(n_2263),
.B(n_2201),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2230),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_SL g2325 ( 
.A(n_2268),
.B(n_2133),
.Y(n_2325)
);

NAND2x1_ASAP7_75t_L g2326 ( 
.A(n_2257),
.B(n_2178),
.Y(n_2326)
);

NAND3xp33_ASAP7_75t_SL g2327 ( 
.A(n_2273),
.B(n_2150),
.C(n_2108),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2233),
.Y(n_2328)
);

AND2x2_ASAP7_75t_L g2329 ( 
.A(n_2263),
.B(n_2178),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2275),
.B(n_2173),
.Y(n_2330)
);

NOR3xp33_ASAP7_75t_L g2331 ( 
.A(n_2277),
.B(n_2114),
.C(n_2161),
.Y(n_2331)
);

OR2x2_ASAP7_75t_L g2332 ( 
.A(n_2267),
.B(n_2162),
.Y(n_2332)
);

NOR2xp67_ASAP7_75t_SL g2333 ( 
.A(n_2227),
.B(n_2016),
.Y(n_2333)
);

OAI31xp33_ASAP7_75t_L g2334 ( 
.A1(n_2261),
.A2(n_2160),
.A3(n_2213),
.B(n_2214),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_2249),
.B(n_2173),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_L g2336 ( 
.A(n_2251),
.B(n_2173),
.Y(n_2336)
);

AND2x2_ASAP7_75t_L g2337 ( 
.A(n_2275),
.B(n_2187),
.Y(n_2337)
);

NOR2xp33_ASAP7_75t_R g2338 ( 
.A(n_2276),
.B(n_2110),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2292),
.Y(n_2339)
);

O2A1O1Ixp33_ASAP7_75t_L g2340 ( 
.A1(n_2308),
.A2(n_2257),
.B(n_2252),
.C(n_2261),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_L g2341 ( 
.A(n_2298),
.B(n_2244),
.Y(n_2341)
);

AND2x2_ASAP7_75t_L g2342 ( 
.A(n_2295),
.B(n_2275),
.Y(n_2342)
);

OR2x2_ASAP7_75t_L g2343 ( 
.A(n_2302),
.B(n_2265),
.Y(n_2343)
);

NOR2xp33_ASAP7_75t_L g2344 ( 
.A(n_2307),
.B(n_2288),
.Y(n_2344)
);

AOI21xp33_ASAP7_75t_L g2345 ( 
.A1(n_2307),
.A2(n_2214),
.B(n_2177),
.Y(n_2345)
);

OAI22xp5_ASAP7_75t_L g2346 ( 
.A1(n_2304),
.A2(n_2189),
.B1(n_2250),
.B2(n_2244),
.Y(n_2346)
);

AOI322xp5_ASAP7_75t_L g2347 ( 
.A1(n_2331),
.A2(n_2177),
.A3(n_2250),
.B1(n_2214),
.B2(n_2189),
.C1(n_2169),
.C2(n_2172),
.Y(n_2347)
);

NAND2x1p5_ASAP7_75t_L g2348 ( 
.A(n_2321),
.B(n_2016),
.Y(n_2348)
);

INVxp67_ASAP7_75t_L g2349 ( 
.A(n_2295),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_2296),
.B(n_2281),
.Y(n_2350)
);

INVxp67_ASAP7_75t_SL g2351 ( 
.A(n_2311),
.Y(n_2351)
);

OR2x2_ASAP7_75t_L g2352 ( 
.A(n_2302),
.B(n_2281),
.Y(n_2352)
);

INVx1_ASAP7_75t_SL g2353 ( 
.A(n_2299),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2292),
.Y(n_2354)
);

OAI21xp33_ASAP7_75t_L g2355 ( 
.A1(n_2316),
.A2(n_2309),
.B(n_2325),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2300),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_SL g2357 ( 
.A(n_2338),
.B(n_2280),
.Y(n_2357)
);

INVxp67_ASAP7_75t_L g2358 ( 
.A(n_2299),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_L g2359 ( 
.A(n_2310),
.B(n_2305),
.Y(n_2359)
);

OAI22xp5_ASAP7_75t_L g2360 ( 
.A1(n_2326),
.A2(n_2274),
.B1(n_2272),
.B2(n_2266),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_2285),
.B(n_2272),
.Y(n_2361)
);

OAI21xp5_ASAP7_75t_L g2362 ( 
.A1(n_2297),
.A2(n_2204),
.B(n_2237),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_2313),
.Y(n_2363)
);

INVx1_ASAP7_75t_SL g2364 ( 
.A(n_2301),
.Y(n_2364)
);

INVxp67_ASAP7_75t_SL g2365 ( 
.A(n_2326),
.Y(n_2365)
);

AND2x2_ASAP7_75t_L g2366 ( 
.A(n_2301),
.B(n_2200),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_2313),
.Y(n_2367)
);

AOI221xp5_ASAP7_75t_L g2368 ( 
.A1(n_2327),
.A2(n_2141),
.B1(n_2255),
.B2(n_2253),
.C(n_2234),
.Y(n_2368)
);

OAI22xp5_ASAP7_75t_L g2369 ( 
.A1(n_2336),
.A2(n_2315),
.B1(n_2313),
.B2(n_2318),
.Y(n_2369)
);

O2A1O1Ixp33_ASAP7_75t_L g2370 ( 
.A1(n_2334),
.A2(n_2204),
.B(n_2270),
.C(n_2239),
.Y(n_2370)
);

AOI221xp5_ASAP7_75t_L g2371 ( 
.A1(n_2315),
.A2(n_2235),
.B1(n_2187),
.B2(n_2240),
.C(n_2246),
.Y(n_2371)
);

OAI22xp5_ASAP7_75t_L g2372 ( 
.A1(n_2318),
.A2(n_2266),
.B1(n_2187),
.B2(n_2200),
.Y(n_2372)
);

OAI21xp33_ASAP7_75t_SL g2373 ( 
.A1(n_2284),
.A2(n_2200),
.B(n_2260),
.Y(n_2373)
);

AND2x4_ASAP7_75t_L g2374 ( 
.A(n_2314),
.B(n_2228),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2300),
.Y(n_2375)
);

OAI221xp5_ASAP7_75t_SL g2376 ( 
.A1(n_2284),
.A2(n_2260),
.B1(n_2254),
.B2(n_2183),
.C(n_2176),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2303),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2303),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2322),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2335),
.B(n_2188),
.Y(n_2380)
);

AND2x2_ASAP7_75t_L g2381 ( 
.A(n_2342),
.B(n_2330),
.Y(n_2381)
);

XNOR2x2_ASAP7_75t_L g2382 ( 
.A(n_2344),
.B(n_2287),
.Y(n_2382)
);

INVxp67_ASAP7_75t_SL g2383 ( 
.A(n_2351),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2339),
.Y(n_2384)
);

INVx2_ASAP7_75t_L g2385 ( 
.A(n_2374),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_2374),
.Y(n_2386)
);

OAI21xp33_ASAP7_75t_L g2387 ( 
.A1(n_2355),
.A2(n_2287),
.B(n_2320),
.Y(n_2387)
);

AOI22xp33_ASAP7_75t_SL g2388 ( 
.A1(n_2344),
.A2(n_2320),
.B1(n_2323),
.B2(n_2290),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2354),
.Y(n_2389)
);

INVx2_ASAP7_75t_L g2390 ( 
.A(n_2374),
.Y(n_2390)
);

INVx1_ASAP7_75t_SL g2391 ( 
.A(n_2353),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2342),
.Y(n_2392)
);

AOI22xp5_ASAP7_75t_L g2393 ( 
.A1(n_2346),
.A2(n_2333),
.B1(n_2323),
.B2(n_2314),
.Y(n_2393)
);

OAI21xp33_ASAP7_75t_L g2394 ( 
.A1(n_2347),
.A2(n_2290),
.B(n_2314),
.Y(n_2394)
);

OR2x2_ASAP7_75t_L g2395 ( 
.A(n_2352),
.B(n_2332),
.Y(n_2395)
);

INVxp67_ASAP7_75t_L g2396 ( 
.A(n_2359),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2356),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2375),
.Y(n_2398)
);

AOI211x1_ASAP7_75t_SL g2399 ( 
.A1(n_2369),
.A2(n_2306),
.B(n_2239),
.C(n_2270),
.Y(n_2399)
);

AOI22xp33_ASAP7_75t_L g2400 ( 
.A1(n_2357),
.A2(n_2345),
.B1(n_2341),
.B2(n_2350),
.Y(n_2400)
);

AOI22xp5_ASAP7_75t_L g2401 ( 
.A1(n_2349),
.A2(n_2333),
.B1(n_2329),
.B2(n_2330),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2377),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2358),
.B(n_2337),
.Y(n_2403)
);

INVxp67_ASAP7_75t_L g2404 ( 
.A(n_2357),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2378),
.Y(n_2405)
);

AND2x2_ASAP7_75t_L g2406 ( 
.A(n_2366),
.B(n_2329),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2379),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_2364),
.B(n_2337),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2352),
.Y(n_2409)
);

OAI22xp5_ASAP7_75t_L g2410 ( 
.A1(n_2348),
.A2(n_2332),
.B1(n_2291),
.B2(n_2294),
.Y(n_2410)
);

AOI21xp5_ASAP7_75t_L g2411 ( 
.A1(n_2340),
.A2(n_2370),
.B(n_2362),
.Y(n_2411)
);

INVx1_ASAP7_75t_SL g2412 ( 
.A(n_2391),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2409),
.Y(n_2413)
);

NAND3xp33_ASAP7_75t_L g2414 ( 
.A(n_2411),
.B(n_2404),
.C(n_2383),
.Y(n_2414)
);

NOR4xp25_ASAP7_75t_SL g2415 ( 
.A(n_2394),
.B(n_2365),
.C(n_2376),
.D(n_2368),
.Y(n_2415)
);

AOI22xp5_ASAP7_75t_L g2416 ( 
.A1(n_2387),
.A2(n_2360),
.B1(n_2348),
.B2(n_2361),
.Y(n_2416)
);

INVxp67_ASAP7_75t_L g2417 ( 
.A(n_2382),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2409),
.Y(n_2418)
);

NAND2x1_ASAP7_75t_L g2419 ( 
.A(n_2401),
.B(n_2385),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2384),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2384),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_2381),
.B(n_2366),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_2396),
.B(n_2343),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_2392),
.B(n_2343),
.Y(n_2424)
);

NOR4xp25_ASAP7_75t_SL g2425 ( 
.A(n_2382),
.B(n_2371),
.C(n_2322),
.D(n_2328),
.Y(n_2425)
);

AND2x2_ASAP7_75t_L g2426 ( 
.A(n_2381),
.B(n_2363),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2389),
.Y(n_2427)
);

INVx2_ASAP7_75t_L g2428 ( 
.A(n_2392),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2389),
.Y(n_2429)
);

NAND4xp25_ASAP7_75t_L g2430 ( 
.A(n_2400),
.B(n_2367),
.C(n_2363),
.D(n_2372),
.Y(n_2430)
);

NAND2x1p5_ASAP7_75t_SL g2431 ( 
.A(n_2385),
.B(n_2386),
.Y(n_2431)
);

OAI22xp5_ASAP7_75t_L g2432 ( 
.A1(n_2393),
.A2(n_2388),
.B1(n_2408),
.B2(n_2403),
.Y(n_2432)
);

AND2x2_ASAP7_75t_L g2433 ( 
.A(n_2406),
.B(n_2367),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2386),
.B(n_2380),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_2412),
.B(n_2390),
.Y(n_2435)
);

NOR2xp33_ASAP7_75t_L g2436 ( 
.A(n_2414),
.B(n_2395),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2428),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_2417),
.B(n_2390),
.Y(n_2438)
);

OA21x2_ASAP7_75t_L g2439 ( 
.A1(n_2418),
.A2(n_2402),
.B(n_2407),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_SL g2440 ( 
.A(n_2423),
.B(n_2410),
.Y(n_2440)
);

AOI21xp5_ASAP7_75t_L g2441 ( 
.A1(n_2425),
.A2(n_2407),
.B(n_2398),
.Y(n_2441)
);

AND2x2_ASAP7_75t_L g2442 ( 
.A(n_2422),
.B(n_2406),
.Y(n_2442)
);

NOR3xp33_ASAP7_75t_L g2443 ( 
.A(n_2432),
.B(n_2405),
.C(n_2402),
.Y(n_2443)
);

AND2x2_ASAP7_75t_L g2444 ( 
.A(n_2422),
.B(n_2395),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2428),
.Y(n_2445)
);

OR2x2_ASAP7_75t_L g2446 ( 
.A(n_2431),
.B(n_2424),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_2426),
.B(n_2397),
.Y(n_2447)
);

NOR2xp33_ASAP7_75t_L g2448 ( 
.A(n_2419),
.B(n_2397),
.Y(n_2448)
);

NOR3xp33_ASAP7_75t_L g2449 ( 
.A(n_2419),
.B(n_2405),
.C(n_2398),
.Y(n_2449)
);

OAI211xp5_ASAP7_75t_SL g2450 ( 
.A1(n_2440),
.A2(n_2416),
.B(n_2413),
.C(n_2399),
.Y(n_2450)
);

AOI221xp5_ASAP7_75t_L g2451 ( 
.A1(n_2449),
.A2(n_2431),
.B1(n_2430),
.B2(n_2418),
.C(n_2429),
.Y(n_2451)
);

AOI221x1_ASAP7_75t_L g2452 ( 
.A1(n_2449),
.A2(n_2421),
.B1(n_2420),
.B2(n_2427),
.C(n_2434),
.Y(n_2452)
);

XNOR2x1_ASAP7_75t_L g2453 ( 
.A(n_2446),
.B(n_2415),
.Y(n_2453)
);

CKINVDCx16_ASAP7_75t_R g2454 ( 
.A(n_2436),
.Y(n_2454)
);

OAI221xp5_ASAP7_75t_L g2455 ( 
.A1(n_2443),
.A2(n_2426),
.B1(n_2433),
.B2(n_2373),
.C(n_2328),
.Y(n_2455)
);

OAI21xp33_ASAP7_75t_SL g2456 ( 
.A1(n_2448),
.A2(n_2433),
.B(n_2324),
.Y(n_2456)
);

AOI221xp5_ASAP7_75t_L g2457 ( 
.A1(n_2441),
.A2(n_2438),
.B1(n_2435),
.B2(n_2444),
.C(n_2447),
.Y(n_2457)
);

AOI221xp5_ASAP7_75t_L g2458 ( 
.A1(n_2441),
.A2(n_2324),
.B1(n_2319),
.B2(n_2317),
.C(n_2312),
.Y(n_2458)
);

AOI211xp5_ASAP7_75t_L g2459 ( 
.A1(n_2442),
.A2(n_2289),
.B(n_2286),
.C(n_2293),
.Y(n_2459)
);

AOI221xp5_ASAP7_75t_L g2460 ( 
.A1(n_2437),
.A2(n_2306),
.B1(n_2294),
.B2(n_2291),
.C(n_2246),
.Y(n_2460)
);

AOI21xp5_ASAP7_75t_L g2461 ( 
.A1(n_2439),
.A2(n_2240),
.B(n_2232),
.Y(n_2461)
);

AOI221x1_ASAP7_75t_L g2462 ( 
.A1(n_2445),
.A2(n_2232),
.B1(n_2192),
.B2(n_2193),
.C(n_2182),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2439),
.Y(n_2463)
);

AOI221xp5_ASAP7_75t_L g2464 ( 
.A1(n_2449),
.A2(n_2211),
.B1(n_2219),
.B2(n_2193),
.C(n_2216),
.Y(n_2464)
);

OAI21xp5_ASAP7_75t_L g2465 ( 
.A1(n_2453),
.A2(n_2211),
.B(n_2219),
.Y(n_2465)
);

NOR2xp33_ASAP7_75t_R g2466 ( 
.A(n_2454),
.B(n_2106),
.Y(n_2466)
);

NOR2xp33_ASAP7_75t_R g2467 ( 
.A(n_2463),
.B(n_2016),
.Y(n_2467)
);

NOR2x1_ASAP7_75t_L g2468 ( 
.A(n_2450),
.B(n_2254),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2456),
.Y(n_2469)
);

AOI22xp5_ASAP7_75t_L g2470 ( 
.A1(n_2451),
.A2(n_2219),
.B1(n_2211),
.B2(n_2035),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2452),
.Y(n_2471)
);

XOR2xp5_ASAP7_75t_L g2472 ( 
.A(n_2457),
.B(n_2056),
.Y(n_2472)
);

AND2x2_ASAP7_75t_SL g2473 ( 
.A(n_2458),
.B(n_2211),
.Y(n_2473)
);

OR2x2_ASAP7_75t_L g2474 ( 
.A(n_2469),
.B(n_2455),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2471),
.Y(n_2475)
);

HB1xp67_ASAP7_75t_L g2476 ( 
.A(n_2466),
.Y(n_2476)
);

NAND2x1p5_ASAP7_75t_L g2477 ( 
.A(n_2468),
.B(n_2461),
.Y(n_2477)
);

NAND4xp75_ASAP7_75t_L g2478 ( 
.A(n_2470),
.B(n_2462),
.C(n_2460),
.D(n_2464),
.Y(n_2478)
);

NAND4xp25_ASAP7_75t_L g2479 ( 
.A(n_2465),
.B(n_2459),
.C(n_2029),
.D(n_2056),
.Y(n_2479)
);

NOR2xp67_ASAP7_75t_L g2480 ( 
.A(n_2467),
.B(n_2225),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_SL g2481 ( 
.A(n_2473),
.B(n_2472),
.Y(n_2481)
);

AOI22xp5_ASAP7_75t_L g2482 ( 
.A1(n_2481),
.A2(n_2211),
.B1(n_2219),
.B2(n_2176),
.Y(n_2482)
);

AOI22xp5_ASAP7_75t_L g2483 ( 
.A1(n_2476),
.A2(n_2219),
.B1(n_2183),
.B2(n_2176),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2477),
.Y(n_2484)
);

NAND2xp5_ASAP7_75t_L g2485 ( 
.A(n_2475),
.B(n_2474),
.Y(n_2485)
);

AOI221xp5_ASAP7_75t_L g2486 ( 
.A1(n_2479),
.A2(n_2225),
.B1(n_2182),
.B2(n_2192),
.C(n_2194),
.Y(n_2486)
);

NOR3xp33_ASAP7_75t_SL g2487 ( 
.A(n_2478),
.B(n_2480),
.C(n_2206),
.Y(n_2487)
);

OAI221xp5_ASAP7_75t_L g2488 ( 
.A1(n_2477),
.A2(n_2029),
.B1(n_2056),
.B2(n_2218),
.C(n_2194),
.Y(n_2488)
);

AND3x4_ASAP7_75t_L g2489 ( 
.A(n_2487),
.B(n_2029),
.C(n_2222),
.Y(n_2489)
);

CKINVDCx5p33_ASAP7_75t_R g2490 ( 
.A(n_2484),
.Y(n_2490)
);

HB1xp67_ASAP7_75t_L g2491 ( 
.A(n_2485),
.Y(n_2491)
);

CKINVDCx5p33_ASAP7_75t_R g2492 ( 
.A(n_2482),
.Y(n_2492)
);

CKINVDCx16_ASAP7_75t_R g2493 ( 
.A(n_2483),
.Y(n_2493)
);

OAI211xp5_ASAP7_75t_L g2494 ( 
.A1(n_2491),
.A2(n_2488),
.B(n_2486),
.C(n_2174),
.Y(n_2494)
);

OAI21xp5_ASAP7_75t_L g2495 ( 
.A1(n_2490),
.A2(n_2175),
.B(n_2174),
.Y(n_2495)
);

OAI31xp33_ASAP7_75t_L g2496 ( 
.A1(n_2494),
.A2(n_2489),
.A3(n_2493),
.B(n_2492),
.Y(n_2496)
);

INVx1_ASAP7_75t_SL g2497 ( 
.A(n_2496),
.Y(n_2497)
);

INVx1_ASAP7_75t_SL g2498 ( 
.A(n_2496),
.Y(n_2498)
);

AOI222xp33_ASAP7_75t_L g2499 ( 
.A1(n_2497),
.A2(n_2495),
.B1(n_2489),
.B2(n_2218),
.C1(n_2198),
.C2(n_2206),
.Y(n_2499)
);

OAI22xp5_ASAP7_75t_L g2500 ( 
.A1(n_2498),
.A2(n_2198),
.B1(n_2216),
.B2(n_2224),
.Y(n_2500)
);

AOI22xp33_ASAP7_75t_L g2501 ( 
.A1(n_2499),
.A2(n_2183),
.B1(n_2025),
.B2(n_1989),
.Y(n_2501)
);

AOI221xp5_ASAP7_75t_L g2502 ( 
.A1(n_2500),
.A2(n_2224),
.B1(n_2215),
.B2(n_2174),
.C(n_2175),
.Y(n_2502)
);

AOI22xp5_ASAP7_75t_L g2503 ( 
.A1(n_2501),
.A2(n_2502),
.B1(n_2175),
.B2(n_2169),
.Y(n_2503)
);

OAI221xp5_ASAP7_75t_L g2504 ( 
.A1(n_2503),
.A2(n_2224),
.B1(n_2215),
.B2(n_2210),
.C(n_2205),
.Y(n_2504)
);

AOI211xp5_ASAP7_75t_L g2505 ( 
.A1(n_2504),
.A2(n_2205),
.B(n_2210),
.C(n_2025),
.Y(n_2505)
);


endmodule