module fake_ariane_1526_n_1891 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1891);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1891;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_899;
wire n_352;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_851;
wire n_212;
wire n_444;
wire n_355;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_1846;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

BUFx3_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_176),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_82),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_168),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_134),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_55),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_14),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_94),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_142),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_113),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_137),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_39),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_193),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_129),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_75),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_1),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_111),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_145),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_144),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_149),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_167),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_127),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_74),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_3),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_67),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_27),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_122),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_86),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_101),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_165),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_91),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_186),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_192),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_73),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_23),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_175),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_163),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_52),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_124),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_34),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_78),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_151),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_99),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_2),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_88),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_201),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_131),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_5),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_33),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_38),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_126),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_22),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_33),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_191),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_72),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_20),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_153),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_60),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_174),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_0),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_146),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_102),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_61),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_28),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_18),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_158),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_139),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_30),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_22),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_27),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_57),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_34),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_30),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_80),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_178),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_108),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_25),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_103),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_121),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_60),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_79),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_89),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_8),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_42),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_52),
.Y(n_287)
);

BUFx5_ASAP7_75t_L g288 ( 
.A(n_184),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_41),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_2),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_65),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_58),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_13),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_170),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_8),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_32),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_93),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_5),
.Y(n_298)
);

INVxp33_ASAP7_75t_L g299 ( 
.A(n_182),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_4),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_132),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_6),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_125),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_172),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_25),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_138),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_183),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_200),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_65),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_117),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_194),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_130),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_10),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_197),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_196),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_46),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_4),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_17),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_185),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_16),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_120),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_13),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_57),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_97),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_135),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_181),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_187),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_166),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_116),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_105),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_1),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_171),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_154),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_11),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_76),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_6),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_10),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_32),
.Y(n_338)
);

BUFx10_ASAP7_75t_L g339 ( 
.A(n_55),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_106),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_195),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_107),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_18),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_199),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_95),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_9),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_48),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_152),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_147),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_50),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_49),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_71),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_44),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_162),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_100),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_90),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_148),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_188),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_14),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_85),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_11),
.Y(n_361)
);

BUFx10_ASAP7_75t_L g362 ( 
.A(n_69),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_159),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_189),
.Y(n_364)
);

BUFx5_ASAP7_75t_L g365 ( 
.A(n_136),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_49),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_7),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_17),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_202),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_198),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_112),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_84),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_119),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_140),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_123),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_64),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_98),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_143),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_20),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_45),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_19),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_150),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_180),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_46),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_40),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_87),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_92),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_48),
.Y(n_388)
);

BUFx10_ASAP7_75t_L g389 ( 
.A(n_44),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_47),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_24),
.Y(n_391)
);

BUFx10_ASAP7_75t_L g392 ( 
.A(n_37),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_179),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_68),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_164),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_21),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_38),
.Y(n_397)
);

BUFx8_ASAP7_75t_SL g398 ( 
.A(n_77),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_62),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_56),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_0),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_128),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_45),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_66),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_279),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_279),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_279),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_279),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_205),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_203),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_246),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_388),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_215),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_219),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_246),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_353),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_221),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_353),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_279),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_300),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_300),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_339),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_308),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_300),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_339),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_395),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_300),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_339),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_300),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_239),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_368),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_368),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_368),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_368),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_269),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_236),
.Y(n_436)
);

INVxp67_ASAP7_75t_SL g437 ( 
.A(n_396),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_310),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_311),
.Y(n_439)
);

INVxp33_ASAP7_75t_L g440 ( 
.A(n_209),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_362),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_329),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_341),
.Y(n_443)
);

BUFx6f_ASAP7_75t_SL g444 ( 
.A(n_362),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_344),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_396),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_237),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_252),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_203),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_266),
.Y(n_450)
);

INVxp67_ASAP7_75t_SL g451 ( 
.A(n_368),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_362),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_208),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_260),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_208),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_260),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_267),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_211),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_348),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_285),
.Y(n_460)
);

INVxp33_ASAP7_75t_SL g461 ( 
.A(n_214),
.Y(n_461)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_389),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_256),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_286),
.Y(n_464)
);

INVxp67_ASAP7_75t_SL g465 ( 
.A(n_274),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_291),
.Y(n_466)
);

CKINVDCx14_ASAP7_75t_R g467 ( 
.A(n_378),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_305),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_211),
.Y(n_469)
);

BUFx2_ASAP7_75t_SL g470 ( 
.A(n_243),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_316),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_318),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_212),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_359),
.Y(n_474)
);

INVxp67_ASAP7_75t_SL g475 ( 
.A(n_274),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_361),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_212),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_255),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_376),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_389),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_256),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_214),
.Y(n_482)
);

CKINVDCx16_ASAP7_75t_R g483 ( 
.A(n_389),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_380),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_336),
.Y(n_485)
);

INVxp33_ASAP7_75t_SL g486 ( 
.A(n_218),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_218),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_398),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_381),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_385),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_309),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_309),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_323),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_340),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_217),
.Y(n_495)
);

INVxp67_ASAP7_75t_SL g496 ( 
.A(n_323),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_403),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_217),
.Y(n_498)
);

CKINVDCx14_ASAP7_75t_R g499 ( 
.A(n_392),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_403),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_392),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_220),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_220),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_222),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_222),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_206),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_206),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_434),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_410),
.B(n_340),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_R g510 ( 
.A(n_499),
.B(n_238),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_405),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g512 ( 
.A(n_412),
.B(n_455),
.Y(n_512)
);

INVx4_ASAP7_75t_L g513 ( 
.A(n_444),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_470),
.B(n_283),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_434),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_405),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_406),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_488),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_454),
.B(n_392),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_406),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_440),
.A2(n_228),
.B1(n_367),
.B2(n_226),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_407),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_407),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_470),
.B(n_437),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_467),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_409),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_465),
.B(n_299),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_408),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_408),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_419),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_419),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_455),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_475),
.B(n_391),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_410),
.B(n_204),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_420),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_449),
.B(n_243),
.Y(n_536)
);

BUFx2_ASAP7_75t_L g537 ( 
.A(n_482),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_449),
.B(n_463),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_463),
.B(n_207),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_420),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_421),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_436),
.A2(n_240),
.B1(n_254),
.B2(n_379),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_421),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_424),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_424),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_427),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_427),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_429),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_429),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_413),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_431),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_431),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_432),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_432),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_433),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_433),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_417),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_458),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_506),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_444),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_430),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_506),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_507),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_435),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_507),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_481),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_451),
.B(n_481),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_456),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_456),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_496),
.B(n_397),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_491),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_491),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_436),
.A2(n_401),
.B1(n_399),
.B2(n_390),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_438),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_492),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_478),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_492),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_493),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_494),
.B(n_210),
.Y(n_579)
);

AND2x6_ASAP7_75t_L g580 ( 
.A(n_494),
.B(n_225),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_493),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_411),
.B(n_307),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_415),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_497),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_416),
.B(n_307),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_497),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_500),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_500),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_418),
.B(n_213),
.Y(n_589)
);

AND2x6_ASAP7_75t_L g590 ( 
.A(n_519),
.B(n_225),
.Y(n_590)
);

AO22x2_ASAP7_75t_L g591 ( 
.A1(n_573),
.A2(n_425),
.B1(n_480),
.B2(n_422),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_516),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_511),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_516),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_565),
.Y(n_595)
);

OR2x2_ASAP7_75t_L g596 ( 
.A(n_537),
.B(n_512),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_543),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_SL g598 ( 
.A1(n_521),
.A2(n_444),
.B1(n_423),
.B2(n_414),
.Y(n_598)
);

INVx2_ASAP7_75t_SL g599 ( 
.A(n_527),
.Y(n_599)
);

INVx1_ASAP7_75t_SL g600 ( 
.A(n_576),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_511),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_516),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_516),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_520),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_517),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_558),
.B(n_458),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_558),
.B(n_469),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_527),
.B(n_482),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_520),
.Y(n_609)
);

OAI22xp33_ASAP7_75t_L g610 ( 
.A1(n_521),
.A2(n_426),
.B1(n_501),
.B2(n_452),
.Y(n_610)
);

BUFx6f_ASAP7_75t_SL g611 ( 
.A(n_513),
.Y(n_611)
);

INVxp67_ASAP7_75t_L g612 ( 
.A(n_537),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_543),
.Y(n_613)
);

BUFx8_ASAP7_75t_SL g614 ( 
.A(n_518),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_543),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_524),
.B(n_536),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_522),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_582),
.A2(n_486),
.B1(n_461),
.B2(n_453),
.Y(n_618)
);

INVx5_ASAP7_75t_L g619 ( 
.A(n_580),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_520),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_582),
.A2(n_487),
.B1(n_400),
.B2(n_452),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_523),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_523),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_528),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_528),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_530),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_520),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_530),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_536),
.B(n_441),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_510),
.B(n_469),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_529),
.Y(n_631)
);

INVx2_ASAP7_75t_SL g632 ( 
.A(n_509),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_514),
.B(n_426),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_543),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_513),
.B(n_473),
.Y(n_635)
);

INVxp67_ASAP7_75t_SL g636 ( 
.A(n_538),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_513),
.B(n_473),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_512),
.Y(n_638)
);

OR2x6_ASAP7_75t_L g639 ( 
.A(n_513),
.B(n_560),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_519),
.B(n_446),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_529),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_560),
.B(n_477),
.Y(n_642)
);

NAND2xp33_ASAP7_75t_SL g643 ( 
.A(n_560),
.B(n_477),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_531),
.Y(n_644)
);

NAND3xp33_ASAP7_75t_L g645 ( 
.A(n_589),
.B(n_498),
.C(n_495),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_560),
.B(n_495),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_536),
.B(n_441),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_531),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_567),
.B(n_498),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_536),
.B(n_502),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_529),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_535),
.Y(n_652)
);

NAND2xp33_ASAP7_75t_L g653 ( 
.A(n_580),
.B(n_502),
.Y(n_653)
);

INVx1_ASAP7_75t_SL g654 ( 
.A(n_526),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_509),
.B(n_503),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_535),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_509),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_535),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_547),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_540),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_547),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_509),
.B(n_503),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_567),
.B(n_582),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_582),
.B(n_504),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_540),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_547),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_585),
.B(n_566),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_554),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_541),
.Y(n_669)
);

INVx1_ASAP7_75t_SL g670 ( 
.A(n_550),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_554),
.Y(n_671)
);

AOI22xp33_ASAP7_75t_L g672 ( 
.A1(n_585),
.A2(n_448),
.B1(n_450),
.B2(n_447),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_554),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_585),
.B(n_504),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_565),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_541),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_583),
.B(n_505),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_571),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_543),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_545),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_585),
.B(n_566),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_543),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_566),
.B(n_505),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_544),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_544),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_545),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_546),
.Y(n_687)
);

NAND2xp33_ASAP7_75t_R g688 ( 
.A(n_525),
.B(n_439),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_565),
.Y(n_689)
);

OR2x6_ASAP7_75t_L g690 ( 
.A(n_589),
.B(n_457),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_565),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_565),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_573),
.A2(n_490),
.B1(n_464),
.B2(n_466),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_583),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_544),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_544),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_546),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_542),
.A2(n_228),
.B1(n_367),
.B2(n_226),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_566),
.B(n_428),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_544),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_548),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_544),
.Y(n_702)
);

NOR3xp33_ASAP7_75t_L g703 ( 
.A(n_532),
.B(n_338),
.C(n_258),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_548),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_565),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_549),
.Y(n_706)
);

OAI22xp33_ASAP7_75t_L g707 ( 
.A1(n_542),
.A2(n_483),
.B1(n_462),
.B2(n_384),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_583),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_559),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_533),
.A2(n_489),
.B1(n_484),
.B2(n_479),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_533),
.B(n_570),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_570),
.B(n_223),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_549),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_534),
.B(n_223),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_551),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_551),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_552),
.Y(n_717)
);

BUFx2_ASAP7_75t_L g718 ( 
.A(n_557),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_571),
.A2(n_468),
.B1(n_476),
.B2(n_474),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_552),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_553),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_539),
.B(n_460),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_553),
.Y(n_723)
);

OAI21xp33_ASAP7_75t_SL g724 ( 
.A1(n_559),
.A2(n_472),
.B(n_471),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_555),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_555),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_556),
.Y(n_727)
);

INVxp33_ASAP7_75t_L g728 ( 
.A(n_579),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_562),
.B(n_277),
.Y(n_729)
);

BUFx2_ASAP7_75t_L g730 ( 
.A(n_561),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_556),
.Y(n_731)
);

CKINVDCx6p67_ASAP7_75t_R g732 ( 
.A(n_580),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_571),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_563),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_562),
.B(n_442),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_563),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_563),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_581),
.B(n_588),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_581),
.B(n_588),
.Y(n_739)
);

INVx5_ASAP7_75t_L g740 ( 
.A(n_580),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_590),
.A2(n_580),
.B1(n_571),
.B2(n_572),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_649),
.B(n_581),
.Y(n_742)
);

A2O1A1Ixp33_ASAP7_75t_L g743 ( 
.A1(n_724),
.A2(n_588),
.B(n_581),
.C(n_569),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_590),
.A2(n_588),
.B1(n_580),
.B2(n_224),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_599),
.B(n_569),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_645),
.B(n_224),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_728),
.B(n_575),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_599),
.B(n_443),
.Y(n_748)
);

INVxp67_ASAP7_75t_L g749 ( 
.A(n_638),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_645),
.B(n_575),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_709),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_694),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_629),
.B(n_577),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_616),
.B(n_577),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_636),
.B(n_578),
.Y(n_755)
);

O2A1O1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_724),
.A2(n_587),
.B(n_586),
.C(n_578),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_596),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_722),
.B(n_586),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_677),
.B(n_587),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_678),
.B(n_229),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_709),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_590),
.B(n_571),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_590),
.A2(n_580),
.B1(n_304),
.B2(n_229),
.Y(n_763)
);

OAI22xp5_ASAP7_75t_L g764 ( 
.A1(n_650),
.A2(n_384),
.B1(n_390),
.B2(n_399),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_590),
.A2(n_580),
.B1(n_304),
.B2(n_234),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_596),
.Y(n_766)
);

BUFx2_ASAP7_75t_L g767 ( 
.A(n_638),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_614),
.Y(n_768)
);

OR2x6_ASAP7_75t_L g769 ( 
.A(n_718),
.B(n_730),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_590),
.B(n_571),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_678),
.B(n_230),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_647),
.B(n_572),
.Y(n_772)
);

INVx2_ASAP7_75t_SL g773 ( 
.A(n_608),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_709),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_590),
.B(n_572),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_683),
.B(n_572),
.Y(n_776)
);

OR2x6_ASAP7_75t_L g777 ( 
.A(n_718),
.B(n_564),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_711),
.B(n_572),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_593),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_664),
.B(n_572),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_631),
.Y(n_781)
);

INVx4_ASAP7_75t_L g782 ( 
.A(n_611),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_631),
.Y(n_783)
);

O2A1O1Ixp5_ASAP7_75t_L g784 ( 
.A1(n_595),
.A2(n_584),
.B(n_568),
.C(n_315),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_608),
.B(n_574),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_690),
.B(n_568),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_690),
.B(n_568),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_678),
.B(n_230),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_690),
.B(n_584),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_678),
.B(n_232),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_690),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_600),
.Y(n_792)
);

INVx5_ASAP7_75t_L g793 ( 
.A(n_639),
.Y(n_793)
);

NOR2x1p5_ASAP7_75t_L g794 ( 
.A(n_699),
.B(n_401),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_601),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_690),
.B(n_584),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_641),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_678),
.B(n_233),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_733),
.B(n_370),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_633),
.B(n_242),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_605),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_641),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_605),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_663),
.B(n_508),
.Y(n_804)
);

INVx4_ASAP7_75t_L g805 ( 
.A(n_611),
.Y(n_805)
);

NAND3xp33_ASAP7_75t_L g806 ( 
.A(n_698),
.B(n_251),
.C(n_250),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_641),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_739),
.B(n_508),
.Y(n_808)
);

OAI22xp5_ASAP7_75t_L g809 ( 
.A1(n_618),
.A2(n_320),
.B1(n_298),
.B2(n_296),
.Y(n_809)
);

OAI221xp5_ASAP7_75t_L g810 ( 
.A1(n_698),
.A2(n_275),
.B1(n_404),
.B2(n_262),
.C(n_265),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_655),
.B(n_270),
.Y(n_811)
);

BUFx2_ASAP7_75t_L g812 ( 
.A(n_612),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_651),
.Y(n_813)
);

O2A1O1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_738),
.A2(n_515),
.B(n_508),
.C(n_278),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_733),
.B(n_370),
.Y(n_815)
);

NOR2xp67_ASAP7_75t_L g816 ( 
.A(n_637),
.B(n_508),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_739),
.B(n_708),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_SL g818 ( 
.A(n_654),
.B(n_445),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_708),
.B(n_729),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_651),
.Y(n_820)
);

INVx2_ASAP7_75t_SL g821 ( 
.A(n_730),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_617),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_632),
.B(n_515),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_651),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_632),
.B(n_515),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_657),
.B(n_515),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_L g827 ( 
.A1(n_657),
.A2(n_272),
.B1(n_337),
.B2(n_343),
.Y(n_827)
);

AOI22x1_ASAP7_75t_R g828 ( 
.A1(n_617),
.A2(n_459),
.B1(n_485),
.B2(n_369),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_652),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_622),
.Y(n_830)
);

O2A1O1Ixp5_ASAP7_75t_L g831 ( 
.A1(n_595),
.A2(n_325),
.B(n_227),
.C(n_231),
.Y(n_831)
);

HB1xp67_ASAP7_75t_L g832 ( 
.A(n_670),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_622),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_652),
.Y(n_834)
);

INVxp67_ASAP7_75t_L g835 ( 
.A(n_735),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_606),
.A2(n_289),
.B1(n_313),
.B2(n_317),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_640),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_667),
.B(n_324),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_623),
.A2(n_235),
.B(n_216),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_623),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_681),
.B(n_364),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_598),
.A2(n_373),
.B1(n_386),
.B2(n_253),
.Y(n_842)
);

INVxp67_ASAP7_75t_L g843 ( 
.A(n_688),
.Y(n_843)
);

BUFx2_ASAP7_75t_L g844 ( 
.A(n_591),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_694),
.B(n_371),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_694),
.B(n_371),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_733),
.B(n_372),
.Y(n_847)
);

NOR3xp33_ASAP7_75t_L g848 ( 
.A(n_610),
.B(n_273),
.C(n_271),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_672),
.B(n_737),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_652),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_621),
.B(n_282),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_624),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_733),
.B(n_372),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_624),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_737),
.B(n_374),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_706),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_710),
.B(n_287),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_662),
.B(n_674),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_625),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_625),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_712),
.Y(n_861)
);

OAI22xp5_ASAP7_75t_L g862 ( 
.A1(n_607),
.A2(n_334),
.B1(n_290),
.B2(n_292),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_706),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_714),
.B(n_293),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_635),
.B(n_295),
.Y(n_865)
);

O2A1O1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_626),
.A2(n_248),
.B(n_244),
.C(n_280),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_592),
.B(n_374),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_693),
.B(n_302),
.Y(n_868)
);

INVx1_ASAP7_75t_SL g869 ( 
.A(n_630),
.Y(n_869)
);

OR2x2_ASAP7_75t_L g870 ( 
.A(n_707),
.B(n_322),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_706),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_713),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_733),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_592),
.B(n_375),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_642),
.B(n_646),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_713),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_594),
.B(n_602),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_594),
.B(n_375),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_602),
.B(n_377),
.Y(n_879)
);

INVx2_ASAP7_75t_SL g880 ( 
.A(n_591),
.Y(n_880)
);

NAND2xp33_ASAP7_75t_L g881 ( 
.A(n_620),
.B(n_377),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_603),
.B(n_382),
.Y(n_882)
);

INVxp33_ASAP7_75t_L g883 ( 
.A(n_703),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_595),
.B(n_331),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_597),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_603),
.B(n_382),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_591),
.B(n_719),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_604),
.B(n_387),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_604),
.B(n_387),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_626),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_SL g891 ( 
.A(n_611),
.B(n_346),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_595),
.B(n_347),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_609),
.B(n_393),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_591),
.B(n_350),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_620),
.B(n_393),
.Y(n_895)
);

NOR2x1p5_ASAP7_75t_L g896 ( 
.A(n_643),
.B(n_351),
.Y(n_896)
);

O2A1O1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_628),
.A2(n_284),
.B(n_297),
.C(n_303),
.Y(n_897)
);

NAND3xp33_ASAP7_75t_L g898 ( 
.A(n_653),
.B(n_366),
.C(n_402),
.Y(n_898)
);

BUFx2_ASAP7_75t_L g899 ( 
.A(n_639),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_713),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_609),
.B(n_394),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_620),
.B(n_394),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_627),
.B(n_402),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_627),
.B(n_327),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_716),
.Y(n_905)
);

NAND2x1p5_ASAP7_75t_L g906 ( 
.A(n_793),
.B(n_740),
.Y(n_906)
);

AOI22xp5_ASAP7_75t_L g907 ( 
.A1(n_800),
.A2(n_648),
.B1(n_665),
.B2(n_669),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_779),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_800),
.A2(n_648),
.B1(n_665),
.B2(n_669),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_781),
.Y(n_910)
);

BUFx2_ASAP7_75t_L g911 ( 
.A(n_767),
.Y(n_911)
);

NAND2x1p5_ASAP7_75t_L g912 ( 
.A(n_793),
.B(n_619),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_792),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_747),
.B(n_734),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_781),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_769),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_783),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_837),
.B(n_639),
.Y(n_918)
);

NOR2x2_ASAP7_75t_L g919 ( 
.A(n_769),
.B(n_639),
.Y(n_919)
);

INVxp67_ASAP7_75t_L g920 ( 
.A(n_812),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_749),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_793),
.B(n_627),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_747),
.B(n_759),
.Y(n_923)
);

INVx5_ASAP7_75t_L g924 ( 
.A(n_793),
.Y(n_924)
);

OAI22xp5_ASAP7_75t_L g925 ( 
.A1(n_817),
.A2(n_795),
.B1(n_803),
.B2(n_801),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_835),
.B(n_705),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_783),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_883),
.B(n_628),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_858),
.A2(n_687),
.B1(n_660),
.B2(n_644),
.Y(n_929)
);

NAND2x1p5_ASAP7_75t_L g930 ( 
.A(n_752),
.B(n_740),
.Y(n_930)
);

INVx1_ASAP7_75t_SL g931 ( 
.A(n_832),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_R g932 ( 
.A(n_768),
.B(n_732),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_769),
.B(n_644),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_758),
.B(n_734),
.Y(n_934)
);

INVx1_ASAP7_75t_SL g935 ( 
.A(n_785),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_757),
.B(n_766),
.Y(n_936)
);

INVx2_ASAP7_75t_SL g937 ( 
.A(n_821),
.Y(n_937)
);

CKINVDCx11_ASAP7_75t_R g938 ( 
.A(n_777),
.Y(n_938)
);

NAND3xp33_ASAP7_75t_L g939 ( 
.A(n_810),
.B(n_676),
.C(n_660),
.Y(n_939)
);

NOR2x1p5_ASAP7_75t_L g940 ( 
.A(n_870),
.B(n_732),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_753),
.B(n_736),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_858),
.A2(n_715),
.B1(n_687),
.B2(n_697),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_R g943 ( 
.A(n_818),
.B(n_597),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_797),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_753),
.B(n_736),
.Y(n_945)
);

CKINVDCx11_ASAP7_75t_R g946 ( 
.A(n_777),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_750),
.B(n_676),
.Y(n_947)
);

BUFx4f_ASAP7_75t_L g948 ( 
.A(n_777),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_773),
.B(n_680),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_797),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_750),
.B(n_680),
.Y(n_951)
);

NOR3xp33_ASAP7_75t_SL g952 ( 
.A(n_764),
.B(n_697),
.C(n_686),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_883),
.B(n_686),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_822),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_830),
.Y(n_955)
);

OR2x6_ASAP7_75t_L g956 ( 
.A(n_748),
.B(n_716),
.Y(n_956)
);

HB1xp67_ASAP7_75t_L g957 ( 
.A(n_748),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_802),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_861),
.B(n_701),
.Y(n_959)
);

OR2x6_ASAP7_75t_L g960 ( 
.A(n_880),
.B(n_716),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_868),
.B(n_721),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_752),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_877),
.A2(n_704),
.B(n_701),
.Y(n_963)
);

OAI22xp5_ASAP7_75t_L g964 ( 
.A1(n_833),
.A2(n_717),
.B1(n_715),
.B2(n_727),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_782),
.B(n_704),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_SL g966 ( 
.A1(n_842),
.A2(n_330),
.B1(n_332),
.B2(n_356),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_742),
.B(n_717),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_840),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_782),
.B(n_720),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_802),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_852),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_SL g972 ( 
.A(n_843),
.B(n_619),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_807),
.Y(n_973)
);

NOR3xp33_ASAP7_75t_SL g974 ( 
.A(n_746),
.B(n_723),
.C(n_720),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_SL g975 ( 
.A(n_805),
.B(n_619),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_745),
.B(n_723),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_819),
.B(n_725),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_754),
.B(n_725),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_873),
.B(n_705),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_778),
.B(n_727),
.Y(n_980)
);

INVx2_ASAP7_75t_SL g981 ( 
.A(n_794),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_807),
.Y(n_982)
);

NAND3xp33_ASAP7_75t_SL g983 ( 
.A(n_848),
.B(n_791),
.C(n_842),
.Y(n_983)
);

NOR3xp33_ASAP7_75t_SL g984 ( 
.A(n_746),
.B(n_261),
.C(n_241),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_854),
.Y(n_985)
);

AOI22xp33_ASAP7_75t_L g986 ( 
.A1(n_851),
.A2(n_731),
.B1(n_721),
.B2(n_726),
.Y(n_986)
);

AOI22xp33_ASAP7_75t_L g987 ( 
.A1(n_844),
.A2(n_731),
.B1(n_721),
.B2(n_726),
.Y(n_987)
);

HB1xp67_ASAP7_75t_L g988 ( 
.A(n_899),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_813),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_813),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_887),
.Y(n_991)
);

INVx5_ASAP7_75t_L g992 ( 
.A(n_873),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_820),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_869),
.B(n_726),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_873),
.B(n_705),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_859),
.Y(n_996)
);

INVx4_ASAP7_75t_L g997 ( 
.A(n_805),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_806),
.B(n_597),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_857),
.B(n_656),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_838),
.B(n_656),
.Y(n_1000)
);

INVx1_ASAP7_75t_SL g1001 ( 
.A(n_894),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_860),
.Y(n_1002)
);

AOI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_865),
.A2(n_864),
.B1(n_892),
.B2(n_884),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_873),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_841),
.B(n_658),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_890),
.B(n_658),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_SL g1007 ( 
.A1(n_811),
.A2(n_373),
.B1(n_386),
.B2(n_363),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_875),
.B(n_597),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_811),
.B(n_613),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_820),
.Y(n_1010)
);

INVx1_ASAP7_75t_SL g1011 ( 
.A(n_845),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_808),
.Y(n_1012)
);

AOI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_865),
.A2(n_675),
.B1(n_689),
.B2(n_691),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_751),
.A2(n_761),
.B1(n_774),
.B2(n_780),
.Y(n_1014)
);

BUFx3_ASAP7_75t_L g1015 ( 
.A(n_885),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_856),
.Y(n_1016)
);

INVx2_ASAP7_75t_SL g1017 ( 
.A(n_896),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_856),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_875),
.B(n_613),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_828),
.Y(n_1020)
);

AOI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_864),
.A2(n_675),
.B1(n_689),
.B2(n_691),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_755),
.B(n_613),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_863),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_884),
.B(n_659),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_828),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_892),
.B(n_659),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_885),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_905),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_863),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_772),
.B(n_661),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_871),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_772),
.B(n_849),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_824),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_871),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_824),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_809),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_829),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_872),
.Y(n_1038)
);

OR2x2_ASAP7_75t_L g1039 ( 
.A(n_827),
.B(n_661),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_804),
.B(n_666),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_776),
.A2(n_615),
.B(n_634),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_872),
.B(n_615),
.Y(n_1042)
);

BUFx4f_ASAP7_75t_L g1043 ( 
.A(n_876),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_786),
.B(n_666),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_787),
.B(n_668),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_876),
.A2(n_673),
.B1(n_668),
.B2(n_671),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_789),
.B(n_671),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_829),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_SL g1049 ( 
.A1(n_836),
.A2(n_342),
.B1(n_247),
.B2(n_249),
.Y(n_1049)
);

BUFx4f_ASAP7_75t_L g1050 ( 
.A(n_900),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_900),
.B(n_615),
.Y(n_1051)
);

INVxp67_ASAP7_75t_L g1052 ( 
.A(n_891),
.Y(n_1052)
);

AOI22xp33_ASAP7_75t_L g1053 ( 
.A1(n_905),
.A2(n_673),
.B1(n_692),
.B2(n_700),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_796),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_743),
.A2(n_855),
.B1(n_776),
.B2(n_889),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_862),
.B(n_692),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_834),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_756),
.Y(n_1058)
);

INVx2_ASAP7_75t_SL g1059 ( 
.A(n_895),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_834),
.Y(n_1060)
);

INVx2_ASAP7_75t_SL g1061 ( 
.A(n_895),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_743),
.B(n_634),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_850),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_846),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_850),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_823),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_744),
.B(n_634),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_816),
.B(n_634),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_867),
.B(n_679),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_874),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_878),
.B(n_679),
.Y(n_1071)
);

OR2x2_ASAP7_75t_L g1072 ( 
.A(n_879),
.B(n_679),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_825),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_763),
.B(n_679),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_765),
.B(n_685),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_882),
.B(n_685),
.Y(n_1076)
);

BUFx8_ASAP7_75t_L g1077 ( 
.A(n_866),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_826),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_886),
.B(n_685),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_904),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_897),
.A2(n_685),
.B(n_702),
.C(n_700),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_888),
.B(n_682),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_893),
.B(n_682),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_741),
.B(n_619),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_904),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_901),
.B(n_682),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_839),
.B(n_684),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_762),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_903),
.B(n_684),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_947),
.A2(n_951),
.B(n_978),
.Y(n_1090)
);

O2A1O1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_923),
.A2(n_881),
.B(n_760),
.C(n_788),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_941),
.A2(n_815),
.B(n_790),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_935),
.B(n_902),
.Y(n_1093)
);

AOI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_1036),
.A2(n_788),
.B1(n_853),
.B2(n_847),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_924),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_924),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_928),
.B(n_771),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_1003),
.A2(n_898),
.B1(n_853),
.B2(n_847),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_908),
.Y(n_1099)
);

O2A1O1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_953),
.A2(n_771),
.B(n_815),
.C(n_799),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_953),
.B(n_790),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_945),
.A2(n_799),
.B(n_798),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_910),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_994),
.B(n_798),
.Y(n_1104)
);

HB1xp67_ASAP7_75t_L g1105 ( 
.A(n_911),
.Y(n_1105)
);

AOI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_983),
.A2(n_770),
.B1(n_775),
.B2(n_741),
.Y(n_1106)
);

OR2x6_ASAP7_75t_L g1107 ( 
.A(n_956),
.B(n_814),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_1064),
.B(n_831),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_907),
.A2(n_702),
.B1(n_700),
.B2(n_696),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1055),
.A2(n_784),
.B(n_702),
.Y(n_1110)
);

NOR3xp33_ASAP7_75t_SL g1111 ( 
.A(n_1070),
.B(n_1025),
.C(n_1020),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_994),
.B(n_684),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_937),
.B(n_695),
.Y(n_1113)
);

OR2x6_ASAP7_75t_L g1114 ( 
.A(n_956),
.B(n_695),
.Y(n_1114)
);

BUFx4f_ASAP7_75t_L g1115 ( 
.A(n_933),
.Y(n_1115)
);

NAND3xp33_ASAP7_75t_SL g1116 ( 
.A(n_952),
.B(n_974),
.C(n_1007),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_961),
.B(n_695),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_933),
.B(n_696),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1011),
.B(n_696),
.Y(n_1119)
);

NAND2xp33_ASAP7_75t_L g1120 ( 
.A(n_952),
.B(n_619),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_909),
.A2(n_740),
.B1(n_619),
.B2(n_321),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_924),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_959),
.B(n_3),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_966),
.A2(n_740),
.B1(n_383),
.B2(n_352),
.Y(n_1124)
);

INVxp67_ASAP7_75t_L g1125 ( 
.A(n_921),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_959),
.B(n_7),
.Y(n_1126)
);

AOI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_936),
.A2(n_319),
.B1(n_257),
.B2(n_259),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_973),
.Y(n_1128)
);

AO32x1_ASAP7_75t_L g1129 ( 
.A1(n_1014),
.A2(n_9),
.A3(n_12),
.B1(n_15),
.B2(n_16),
.Y(n_1129)
);

AOI21x1_ASAP7_75t_L g1130 ( 
.A1(n_1024),
.A2(n_365),
.B(n_288),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_949),
.B(n_991),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_1009),
.A2(n_740),
.B(n_328),
.C(n_326),
.Y(n_1132)
);

BUFx3_ASAP7_75t_L g1133 ( 
.A(n_913),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_948),
.B(n_245),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_973),
.Y(n_1135)
);

INVxp67_ASAP7_75t_L g1136 ( 
.A(n_921),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_949),
.B(n_12),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_1009),
.A2(n_333),
.B(n_264),
.C(n_360),
.Y(n_1138)
);

CKINVDCx20_ASAP7_75t_R g1139 ( 
.A(n_938),
.Y(n_1139)
);

BUFx4f_ASAP7_75t_L g1140 ( 
.A(n_956),
.Y(n_1140)
);

O2A1O1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_920),
.A2(n_15),
.B(n_19),
.C(n_21),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_948),
.B(n_263),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_929),
.A2(n_335),
.B1(n_358),
.B2(n_357),
.Y(n_1143)
);

INVxp67_ASAP7_75t_SL g1144 ( 
.A(n_1028),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_R g1145 ( 
.A(n_938),
.B(n_268),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_974),
.A2(n_314),
.B(n_281),
.C(n_355),
.Y(n_1146)
);

AOI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1026),
.A2(n_365),
.B(n_288),
.Y(n_1147)
);

AOI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_999),
.A2(n_383),
.B1(n_352),
.B2(n_288),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_967),
.A2(n_312),
.B(n_354),
.Y(n_1149)
);

AOI22xp33_ASAP7_75t_L g1150 ( 
.A1(n_986),
.A2(n_383),
.B1(n_352),
.B2(n_365),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_946),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1012),
.B(n_23),
.Y(n_1152)
);

O2A1O1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_925),
.A2(n_926),
.B(n_976),
.C(n_977),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_931),
.B(n_306),
.Y(n_1154)
);

BUFx4f_ASAP7_75t_L g1155 ( 
.A(n_965),
.Y(n_1155)
);

AOI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1032),
.A2(n_365),
.B(n_288),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_SL g1157 ( 
.A1(n_1069),
.A2(n_998),
.B(n_1022),
.C(n_1027),
.Y(n_1157)
);

CKINVDCx8_ASAP7_75t_R g1158 ( 
.A(n_924),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_980),
.A2(n_349),
.B(n_345),
.Y(n_1159)
);

NOR3xp33_ASAP7_75t_SL g1160 ( 
.A(n_964),
.B(n_276),
.C(n_294),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_R g1161 ( 
.A(n_946),
.B(n_913),
.Y(n_1161)
);

AOI22xp33_ASAP7_75t_L g1162 ( 
.A1(n_986),
.A2(n_383),
.B1(n_352),
.B2(n_365),
.Y(n_1162)
);

INVx5_ASAP7_75t_L g1163 ( 
.A(n_960),
.Y(n_1163)
);

BUFx12f_ASAP7_75t_L g1164 ( 
.A(n_981),
.Y(n_1164)
);

CKINVDCx20_ASAP7_75t_R g1165 ( 
.A(n_932),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1054),
.B(n_24),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_934),
.A2(n_301),
.B(n_383),
.Y(n_1167)
);

OAI21xp5_ASAP7_75t_SL g1168 ( 
.A1(n_1052),
.A2(n_26),
.B(n_28),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_989),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_957),
.B(n_26),
.Y(n_1170)
);

O2A1O1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_926),
.A2(n_29),
.B(n_31),
.C(n_35),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_954),
.Y(n_1172)
);

AOI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_1077),
.A2(n_987),
.B1(n_914),
.B2(n_957),
.Y(n_1173)
);

BUFx12f_ASAP7_75t_L g1174 ( 
.A(n_916),
.Y(n_1174)
);

A2O1A1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_942),
.A2(n_352),
.B(n_365),
.C(n_288),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_963),
.A2(n_70),
.B(n_190),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_939),
.A2(n_365),
.B(n_288),
.C(n_35),
.Y(n_1177)
);

INVxp67_ASAP7_75t_L g1178 ( 
.A(n_988),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_990),
.Y(n_1179)
);

OAI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1022),
.A2(n_288),
.B(n_31),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_955),
.B(n_29),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_916),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_968),
.B(n_971),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_985),
.B(n_36),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_993),
.Y(n_1185)
);

OR2x2_ASAP7_75t_L g1186 ( 
.A(n_988),
.B(n_1001),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1030),
.A2(n_81),
.B(n_177),
.Y(n_1187)
);

OA22x2_ASAP7_75t_L g1188 ( 
.A1(n_1059),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_918),
.B(n_40),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1041),
.A2(n_83),
.B(n_173),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_996),
.B(n_1002),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1016),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_987),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_1193)
);

OR2x6_ASAP7_75t_L g1194 ( 
.A(n_940),
.B(n_43),
.Y(n_1194)
);

AOI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_918),
.A2(n_47),
.B1(n_50),
.B2(n_51),
.Y(n_1195)
);

OAI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1062),
.A2(n_51),
.B(n_53),
.Y(n_1196)
);

HB1xp67_ASAP7_75t_L g1197 ( 
.A(n_1028),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_1017),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1077),
.A2(n_1058),
.B1(n_1031),
.B2(n_1018),
.Y(n_1199)
);

INVx1_ASAP7_75t_SL g1200 ( 
.A(n_943),
.Y(n_1200)
);

AO21x1_ASAP7_75t_L g1201 ( 
.A1(n_998),
.A2(n_109),
.B(n_169),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_SL g1202 ( 
.A(n_997),
.B(n_53),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1068),
.A2(n_110),
.B(n_161),
.Y(n_1203)
);

AOI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_965),
.A2(n_54),
.B1(n_56),
.B2(n_58),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1068),
.A2(n_114),
.B(n_160),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_943),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_932),
.B(n_54),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_969),
.B(n_59),
.Y(n_1208)
);

A2O1A1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_1061),
.A2(n_59),
.B(n_61),
.C(n_62),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1076),
.A2(n_118),
.B(n_156),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_969),
.B(n_63),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_993),
.Y(n_1212)
);

A2O1A1Ixp33_ASAP7_75t_L g1213 ( 
.A1(n_1069),
.A2(n_63),
.B(n_64),
.C(n_66),
.Y(n_1213)
);

O2A1O1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1008),
.A2(n_96),
.B(n_104),
.C(n_115),
.Y(n_1214)
);

BUFx2_ASAP7_75t_L g1215 ( 
.A(n_919),
.Y(n_1215)
);

HB1xp67_ASAP7_75t_L g1216 ( 
.A(n_1060),
.Y(n_1216)
);

HB1xp67_ASAP7_75t_L g1217 ( 
.A(n_1060),
.Y(n_1217)
);

BUFx2_ASAP7_75t_L g1218 ( 
.A(n_1015),
.Y(n_1218)
);

BUFx4f_ASAP7_75t_SL g1219 ( 
.A(n_997),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1008),
.B(n_133),
.Y(n_1220)
);

BUFx3_ASAP7_75t_L g1221 ( 
.A(n_1015),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_SL g1222 ( 
.A(n_1043),
.B(n_141),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_1019),
.B(n_155),
.Y(n_1223)
);

INVx2_ASAP7_75t_SL g1224 ( 
.A(n_1050),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1049),
.A2(n_1080),
.B1(n_1078),
.B2(n_1073),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1066),
.B(n_1088),
.Y(n_1226)
);

CKINVDCx8_ASAP7_75t_R g1227 ( 
.A(n_992),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_962),
.Y(n_1228)
);

A2O1A1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_984),
.A2(n_1039),
.B(n_1056),
.C(n_1081),
.Y(n_1229)
);

BUFx3_ASAP7_75t_L g1230 ( 
.A(n_992),
.Y(n_1230)
);

O2A1O1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1081),
.A2(n_1079),
.B(n_984),
.C(n_1072),
.Y(n_1231)
);

CKINVDCx16_ASAP7_75t_R g1232 ( 
.A(n_975),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_1004),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1085),
.B(n_1029),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1042),
.A2(n_1051),
.B(n_1074),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1089),
.A2(n_1040),
.B(n_1086),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1000),
.B(n_1005),
.Y(n_1237)
);

BUFx3_ASAP7_75t_L g1238 ( 
.A(n_1133),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1099),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_1155),
.B(n_992),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1090),
.A2(n_1153),
.B(n_1236),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1157),
.A2(n_1067),
.B(n_1087),
.Y(n_1242)
);

INVx5_ASAP7_75t_L g1243 ( 
.A(n_1122),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1226),
.B(n_1023),
.Y(n_1244)
);

O2A1O1Ixp5_ASAP7_75t_SL g1245 ( 
.A1(n_1180),
.A2(n_979),
.B(n_995),
.C(n_1042),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1226),
.B(n_1034),
.Y(n_1246)
);

INVx5_ASAP7_75t_L g1247 ( 
.A(n_1122),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_1125),
.B(n_962),
.Y(n_1248)
);

CKINVDCx6p67_ASAP7_75t_R g1249 ( 
.A(n_1139),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1125),
.B(n_1136),
.Y(n_1250)
);

AOI211x1_ASAP7_75t_L g1251 ( 
.A1(n_1196),
.A2(n_1006),
.B(n_1051),
.C(n_1083),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1136),
.B(n_1093),
.Y(n_1252)
);

AO31x2_ASAP7_75t_L g1253 ( 
.A1(n_1229),
.A2(n_1082),
.A3(n_1037),
.B(n_1035),
.Y(n_1253)
);

NOR2xp67_ASAP7_75t_SL g1254 ( 
.A(n_1151),
.B(n_1004),
.Y(n_1254)
);

INVx3_ASAP7_75t_SL g1255 ( 
.A(n_1165),
.Y(n_1255)
);

OR2x2_ASAP7_75t_SL g1256 ( 
.A(n_1116),
.B(n_1004),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1092),
.A2(n_1067),
.B(n_1075),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1123),
.A2(n_1027),
.B1(n_1013),
.B2(n_1021),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1110),
.A2(n_995),
.B(n_979),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1093),
.B(n_1038),
.Y(n_1260)
);

AO31x2_ASAP7_75t_L g1261 ( 
.A1(n_1175),
.A2(n_1201),
.A3(n_1102),
.B(n_1098),
.Y(n_1261)
);

INVx2_ASAP7_75t_SL g1262 ( 
.A(n_1115),
.Y(n_1262)
);

BUFx2_ASAP7_75t_R g1263 ( 
.A(n_1227),
.Y(n_1263)
);

OR2x6_ASAP7_75t_L g1264 ( 
.A(n_1206),
.B(n_1084),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1130),
.A2(n_1063),
.B(n_1010),
.Y(n_1265)
);

AO31x2_ASAP7_75t_L g1266 ( 
.A1(n_1177),
.A2(n_1048),
.A3(n_1063),
.B(n_1010),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_SL g1267 ( 
.A(n_1155),
.B(n_1232),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1147),
.A2(n_1035),
.B(n_1037),
.Y(n_1268)
);

NOR3xp33_ASAP7_75t_SL g1269 ( 
.A(n_1168),
.B(n_922),
.C(n_1075),
.Y(n_1269)
);

AND2x4_ASAP7_75t_L g1270 ( 
.A(n_1221),
.B(n_1004),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_SL g1271 ( 
.A(n_1115),
.B(n_1038),
.Y(n_1271)
);

AOI21x1_ASAP7_75t_SL g1272 ( 
.A1(n_1126),
.A2(n_1071),
.B(n_1045),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1131),
.B(n_1048),
.Y(n_1273)
);

CKINVDCx20_ASAP7_75t_R g1274 ( 
.A(n_1145),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1156),
.A2(n_1047),
.B(n_1044),
.Y(n_1275)
);

NAND2xp33_ASAP7_75t_L g1276 ( 
.A(n_1160),
.B(n_1088),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1105),
.B(n_958),
.Y(n_1277)
);

AOI31xp67_ASAP7_75t_L g1278 ( 
.A1(n_1094),
.A2(n_1074),
.A3(n_922),
.B(n_915),
.Y(n_1278)
);

AO31x2_ASAP7_75t_L g1279 ( 
.A1(n_1237),
.A2(n_970),
.A3(n_1065),
.B(n_917),
.Y(n_1279)
);

INVx1_ASAP7_75t_SL g1280 ( 
.A(n_1200),
.Y(n_1280)
);

AO31x2_ASAP7_75t_L g1281 ( 
.A1(n_1103),
.A2(n_950),
.A3(n_1033),
.B(n_927),
.Y(n_1281)
);

AO31x2_ASAP7_75t_L g1282 ( 
.A1(n_1128),
.A2(n_982),
.A3(n_944),
.B(n_1053),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1120),
.A2(n_1084),
.B(n_1053),
.Y(n_1283)
);

OA21x2_ASAP7_75t_L g1284 ( 
.A1(n_1235),
.A2(n_1046),
.B(n_1057),
.Y(n_1284)
);

AOI221xp5_ASAP7_75t_L g1285 ( 
.A1(n_1116),
.A2(n_1046),
.B1(n_1057),
.B2(n_972),
.C(n_930),
.Y(n_1285)
);

NOR2xp67_ASAP7_75t_L g1286 ( 
.A(n_1095),
.B(n_906),
.Y(n_1286)
);

AO31x2_ASAP7_75t_L g1287 ( 
.A1(n_1135),
.A2(n_912),
.A3(n_1179),
.B(n_1169),
.Y(n_1287)
);

A2O1A1Ixp33_ASAP7_75t_L g1288 ( 
.A1(n_1100),
.A2(n_1091),
.B(n_1097),
.C(n_1101),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1190),
.A2(n_1176),
.B(n_1231),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_SL g1290 ( 
.A(n_1233),
.B(n_1225),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_SL g1291 ( 
.A1(n_1144),
.A2(n_1222),
.B(n_1223),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1105),
.B(n_1178),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1144),
.A2(n_1167),
.B(n_1210),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1187),
.A2(n_1109),
.B(n_1205),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1178),
.B(n_1208),
.Y(n_1295)
);

AO21x2_ASAP7_75t_L g1296 ( 
.A1(n_1112),
.A2(n_1104),
.B(n_1132),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_SL g1297 ( 
.A(n_1194),
.Y(n_1297)
);

AND2x4_ASAP7_75t_L g1298 ( 
.A(n_1182),
.B(n_1163),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1183),
.A2(n_1191),
.B(n_1152),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1170),
.B(n_1172),
.Y(n_1300)
);

O2A1O1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1213),
.A2(n_1141),
.B(n_1209),
.C(n_1211),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1170),
.B(n_1186),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1117),
.A2(n_1108),
.B(n_1138),
.Y(n_1303)
);

AO31x2_ASAP7_75t_L g1304 ( 
.A1(n_1185),
.A2(n_1212),
.A3(n_1192),
.B(n_1146),
.Y(n_1304)
);

HB1xp67_ASAP7_75t_L g1305 ( 
.A(n_1218),
.Y(n_1305)
);

OAI22x1_ASAP7_75t_L g1306 ( 
.A1(n_1195),
.A2(n_1204),
.B1(n_1215),
.B2(n_1189),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1173),
.B(n_1137),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_SL g1308 ( 
.A(n_1163),
.B(n_1199),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1173),
.B(n_1119),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1203),
.A2(n_1214),
.B(n_1096),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1199),
.B(n_1140),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_SL g1312 ( 
.A(n_1163),
.B(n_1158),
.Y(n_1312)
);

OA21x2_ASAP7_75t_L g1313 ( 
.A1(n_1150),
.A2(n_1162),
.B(n_1148),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1121),
.A2(n_1163),
.B(n_1166),
.Y(n_1314)
);

NAND2xp33_ASAP7_75t_SL g1315 ( 
.A(n_1160),
.B(n_1161),
.Y(n_1315)
);

INVx3_ASAP7_75t_L g1316 ( 
.A(n_1122),
.Y(n_1316)
);

A2O1A1Ixp33_ASAP7_75t_L g1317 ( 
.A1(n_1223),
.A2(n_1171),
.B(n_1184),
.C(n_1181),
.Y(n_1317)
);

AO31x2_ASAP7_75t_L g1318 ( 
.A1(n_1193),
.A2(n_1159),
.A3(n_1149),
.B(n_1143),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1150),
.A2(n_1162),
.B(n_1107),
.Y(n_1319)
);

INVx3_ASAP7_75t_L g1320 ( 
.A(n_1122),
.Y(n_1320)
);

OAI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1106),
.A2(n_1220),
.B(n_1148),
.Y(n_1321)
);

BUFx4f_ASAP7_75t_L g1322 ( 
.A(n_1194),
.Y(n_1322)
);

BUFx3_ASAP7_75t_L g1323 ( 
.A(n_1174),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1234),
.Y(n_1324)
);

AOI211x1_ASAP7_75t_L g1325 ( 
.A1(n_1113),
.A2(n_1118),
.B(n_1207),
.C(n_1142),
.Y(n_1325)
);

OAI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1188),
.A2(n_1107),
.B(n_1197),
.Y(n_1326)
);

INVx2_ASAP7_75t_SL g1327 ( 
.A(n_1219),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1230),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1194),
.B(n_1228),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1107),
.A2(n_1217),
.B(n_1197),
.Y(n_1330)
);

A2O1A1Ixp33_ASAP7_75t_L g1331 ( 
.A1(n_1124),
.A2(n_1224),
.B(n_1202),
.C(n_1127),
.Y(n_1331)
);

INVxp67_ASAP7_75t_SL g1332 ( 
.A(n_1216),
.Y(n_1332)
);

INVxp67_ASAP7_75t_SL g1333 ( 
.A(n_1134),
.Y(n_1333)
);

NAND2x1p5_ASAP7_75t_L g1334 ( 
.A(n_1198),
.B(n_1154),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1219),
.B(n_1111),
.Y(n_1335)
);

INVx5_ASAP7_75t_L g1336 ( 
.A(n_1114),
.Y(n_1336)
);

INVx4_ASAP7_75t_L g1337 ( 
.A(n_1164),
.Y(n_1337)
);

AO32x2_ASAP7_75t_L g1338 ( 
.A1(n_1129),
.A2(n_880),
.A3(n_1193),
.B1(n_1098),
.B2(n_1055),
.Y(n_1338)
);

OA21x2_ASAP7_75t_L g1339 ( 
.A1(n_1124),
.A2(n_1129),
.B(n_1111),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1114),
.B(n_1129),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1099),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1226),
.B(n_923),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1090),
.A2(n_1003),
.B(n_951),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1226),
.B(n_923),
.Y(n_1344)
);

AO31x2_ASAP7_75t_L g1345 ( 
.A1(n_1236),
.A2(n_1229),
.A3(n_1055),
.B(n_1175),
.Y(n_1345)
);

NAND2x1_ASAP7_75t_L g1346 ( 
.A(n_1095),
.B(n_1096),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1090),
.A2(n_1003),
.B(n_951),
.Y(n_1347)
);

INVx1_ASAP7_75t_SL g1348 ( 
.A(n_1200),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1130),
.A2(n_1147),
.B(n_1156),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1115),
.B(n_757),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1180),
.A2(n_1003),
.B(n_1090),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1090),
.A2(n_1003),
.B(n_951),
.Y(n_1352)
);

AO32x2_ASAP7_75t_L g1353 ( 
.A1(n_1193),
.A2(n_880),
.A3(n_1098),
.B1(n_1055),
.B2(n_966),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1090),
.A2(n_1003),
.B(n_951),
.Y(n_1354)
);

INVx6_ASAP7_75t_L g1355 ( 
.A(n_1174),
.Y(n_1355)
);

AO31x2_ASAP7_75t_L g1356 ( 
.A1(n_1236),
.A2(n_1229),
.A3(n_1055),
.B(n_1175),
.Y(n_1356)
);

AO21x2_ASAP7_75t_L g1357 ( 
.A1(n_1130),
.A2(n_1147),
.B(n_1156),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1226),
.B(n_923),
.Y(n_1358)
);

AO31x2_ASAP7_75t_L g1359 ( 
.A1(n_1236),
.A2(n_1229),
.A3(n_1055),
.B(n_1175),
.Y(n_1359)
);

AOI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1156),
.A2(n_1147),
.B(n_1130),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1226),
.B(n_923),
.Y(n_1361)
);

NAND2x1p5_ASAP7_75t_L g1362 ( 
.A(n_1115),
.B(n_1155),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1099),
.Y(n_1363)
);

NOR2xp67_ASAP7_75t_L g1364 ( 
.A(n_1095),
.B(n_992),
.Y(n_1364)
);

BUFx2_ASAP7_75t_L g1365 ( 
.A(n_1105),
.Y(n_1365)
);

OR2x6_ASAP7_75t_SL g1366 ( 
.A(n_1151),
.B(n_768),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1130),
.A2(n_1147),
.B(n_1156),
.Y(n_1367)
);

NOR2x1_ASAP7_75t_SL g1368 ( 
.A(n_1122),
.B(n_1163),
.Y(n_1368)
);

NOR2xp67_ASAP7_75t_L g1369 ( 
.A(n_1095),
.B(n_992),
.Y(n_1369)
);

INVx6_ASAP7_75t_L g1370 ( 
.A(n_1174),
.Y(n_1370)
);

NOR2xp67_ASAP7_75t_L g1371 ( 
.A(n_1095),
.B(n_992),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1226),
.B(n_923),
.Y(n_1372)
);

AOI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1116),
.A2(n_1036),
.B1(n_800),
.B2(n_983),
.Y(n_1373)
);

OAI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1180),
.A2(n_1003),
.B(n_1090),
.Y(n_1374)
);

BUFx6f_ASAP7_75t_L g1375 ( 
.A(n_1115),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_1161),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1221),
.B(n_1182),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1130),
.A2(n_1147),
.B(n_1156),
.Y(n_1378)
);

INVxp67_ASAP7_75t_SL g1379 ( 
.A(n_1144),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1090),
.A2(n_1003),
.B(n_951),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1180),
.A2(n_1003),
.B(n_1090),
.Y(n_1381)
);

INVx4_ASAP7_75t_L g1382 ( 
.A(n_1155),
.Y(n_1382)
);

OA21x2_ASAP7_75t_L g1383 ( 
.A1(n_1110),
.A2(n_1235),
.B(n_1229),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_SL g1384 ( 
.A(n_1155),
.B(n_1003),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1226),
.B(n_923),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_R g1386 ( 
.A(n_1165),
.B(n_768),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1155),
.B(n_1003),
.Y(n_1387)
);

BUFx8_ASAP7_75t_L g1388 ( 
.A(n_1164),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_1373),
.B(n_1384),
.Y(n_1389)
);

INVx2_ASAP7_75t_SL g1390 ( 
.A(n_1355),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1373),
.A2(n_1344),
.B1(n_1358),
.B2(n_1342),
.Y(n_1391)
);

AO31x2_ASAP7_75t_L g1392 ( 
.A1(n_1241),
.A2(n_1242),
.A3(n_1340),
.B(n_1258),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1295),
.B(n_1292),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1360),
.A2(n_1367),
.B(n_1349),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1378),
.A2(n_1289),
.B(n_1294),
.Y(n_1395)
);

INVxp67_ASAP7_75t_L g1396 ( 
.A(n_1332),
.Y(n_1396)
);

INVxp67_ASAP7_75t_SL g1397 ( 
.A(n_1379),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1361),
.B(n_1372),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1275),
.A2(n_1293),
.B(n_1268),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1321),
.A2(n_1307),
.B1(n_1319),
.B2(n_1313),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1351),
.A2(n_1381),
.B(n_1347),
.Y(n_1401)
);

AO31x2_ASAP7_75t_L g1402 ( 
.A1(n_1259),
.A2(n_1352),
.A3(n_1354),
.B(n_1380),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1321),
.A2(n_1313),
.B1(n_1297),
.B2(n_1306),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1265),
.A2(n_1310),
.B(n_1272),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1341),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1297),
.A2(n_1322),
.B1(n_1290),
.B2(n_1387),
.Y(n_1406)
);

INVx3_ASAP7_75t_L g1407 ( 
.A(n_1382),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1385),
.B(n_1252),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1322),
.A2(n_1309),
.B1(n_1302),
.B2(n_1324),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1300),
.B(n_1365),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1363),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1244),
.B(n_1246),
.Y(n_1412)
);

AND2x4_ASAP7_75t_L g1413 ( 
.A(n_1264),
.B(n_1336),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1269),
.A2(n_1256),
.B1(n_1301),
.B2(n_1331),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_SL g1415 ( 
.A1(n_1299),
.A2(n_1303),
.B(n_1311),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_SL g1416 ( 
.A1(n_1326),
.A2(n_1330),
.B(n_1335),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1283),
.A2(n_1291),
.B(n_1288),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1277),
.Y(n_1418)
);

AND2x4_ASAP7_75t_L g1419 ( 
.A(n_1264),
.B(n_1336),
.Y(n_1419)
);

INVx3_ASAP7_75t_L g1420 ( 
.A(n_1382),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1257),
.A2(n_1245),
.B(n_1314),
.Y(n_1421)
);

CKINVDCx11_ASAP7_75t_R g1422 ( 
.A(n_1366),
.Y(n_1422)
);

AND2x4_ASAP7_75t_L g1423 ( 
.A(n_1264),
.B(n_1336),
.Y(n_1423)
);

OAI221xp5_ASAP7_75t_L g1424 ( 
.A1(n_1333),
.A2(n_1315),
.B1(n_1276),
.B2(n_1334),
.C(n_1329),
.Y(n_1424)
);

BUFx10_ASAP7_75t_L g1425 ( 
.A(n_1376),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1284),
.A2(n_1383),
.B(n_1346),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1284),
.A2(n_1383),
.B(n_1326),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1250),
.A2(n_1248),
.B1(n_1305),
.B2(n_1251),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1260),
.B(n_1280),
.Y(n_1429)
);

BUFx4_ASAP7_75t_SL g1430 ( 
.A(n_1274),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1296),
.A2(n_1285),
.B(n_1357),
.Y(n_1431)
);

OAI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1339),
.A2(n_1348),
.B1(n_1353),
.B2(n_1362),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_1386),
.Y(n_1433)
);

CKINVDCx20_ASAP7_75t_R g1434 ( 
.A(n_1388),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1308),
.A2(n_1339),
.B1(n_1273),
.B2(n_1353),
.Y(n_1435)
);

INVx3_ASAP7_75t_L g1436 ( 
.A(n_1375),
.Y(n_1436)
);

O2A1O1Ixp33_ASAP7_75t_L g1437 ( 
.A1(n_1327),
.A2(n_1255),
.B(n_1267),
.C(n_1271),
.Y(n_1437)
);

AO31x2_ASAP7_75t_L g1438 ( 
.A1(n_1338),
.A2(n_1278),
.A3(n_1253),
.B(n_1279),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1251),
.A2(n_1325),
.B1(n_1263),
.B2(n_1350),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1353),
.A2(n_1375),
.B1(n_1262),
.B2(n_1355),
.Y(n_1440)
);

AOI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1240),
.A2(n_1312),
.B(n_1368),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1364),
.A2(n_1369),
.B(n_1371),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1377),
.B(n_1238),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1316),
.A2(n_1320),
.B(n_1328),
.Y(n_1444)
);

A2O1A1Ixp33_ASAP7_75t_L g1445 ( 
.A1(n_1338),
.A2(n_1286),
.B(n_1254),
.C(n_1371),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_SL g1446 ( 
.A1(n_1338),
.A2(n_1375),
.B1(n_1370),
.B2(n_1325),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1253),
.Y(n_1447)
);

CKINVDCx11_ASAP7_75t_R g1448 ( 
.A(n_1249),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1270),
.B(n_1298),
.Y(n_1449)
);

INVx3_ASAP7_75t_L g1450 ( 
.A(n_1243),
.Y(n_1450)
);

AO31x2_ASAP7_75t_L g1451 ( 
.A1(n_1261),
.A2(n_1266),
.A3(n_1359),
.B(n_1345),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_SL g1452 ( 
.A1(n_1337),
.A2(n_1261),
.B(n_1318),
.Y(n_1452)
);

OR2x6_ASAP7_75t_L g1453 ( 
.A(n_1298),
.B(n_1370),
.Y(n_1453)
);

INVxp67_ASAP7_75t_SL g1454 ( 
.A(n_1364),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1281),
.Y(n_1455)
);

NAND3xp33_ASAP7_75t_L g1456 ( 
.A(n_1243),
.B(n_1247),
.C(n_1270),
.Y(n_1456)
);

CKINVDCx20_ASAP7_75t_R g1457 ( 
.A(n_1388),
.Y(n_1457)
);

INVx1_ASAP7_75t_SL g1458 ( 
.A(n_1323),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_SL g1459 ( 
.A(n_1247),
.B(n_1356),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1345),
.A2(n_1356),
.B(n_1266),
.Y(n_1460)
);

OAI211xp5_ASAP7_75t_SL g1461 ( 
.A1(n_1318),
.A2(n_1304),
.B(n_1266),
.C(n_1287),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1281),
.Y(n_1462)
);

OAI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1304),
.A2(n_1282),
.B(n_1287),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1304),
.A2(n_1373),
.B1(n_1003),
.B2(n_800),
.Y(n_1464)
);

CKINVDCx20_ASAP7_75t_R g1465 ( 
.A(n_1282),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_L g1466 ( 
.A1(n_1360),
.A2(n_1367),
.B(n_1349),
.Y(n_1466)
);

OAI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1360),
.A2(n_1367),
.B(n_1349),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1373),
.A2(n_842),
.B1(n_894),
.B2(n_983),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1239),
.Y(n_1469)
);

A2O1A1Ixp33_ASAP7_75t_L g1470 ( 
.A1(n_1373),
.A2(n_1003),
.B(n_1374),
.C(n_1351),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1264),
.B(n_1336),
.Y(n_1471)
);

BUFx12f_ASAP7_75t_L g1472 ( 
.A(n_1388),
.Y(n_1472)
);

OAI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1373),
.A2(n_1003),
.B(n_800),
.Y(n_1473)
);

OA21x2_ASAP7_75t_L g1474 ( 
.A1(n_1241),
.A2(n_1242),
.B(n_1257),
.Y(n_1474)
);

OAI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1360),
.A2(n_1367),
.B(n_1349),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1295),
.B(n_1292),
.Y(n_1476)
);

BUFx2_ASAP7_75t_L g1477 ( 
.A(n_1365),
.Y(n_1477)
);

AOI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1360),
.A2(n_1242),
.B(n_1343),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1360),
.A2(n_1367),
.B(n_1349),
.Y(n_1479)
);

BUFx12f_ASAP7_75t_L g1480 ( 
.A(n_1388),
.Y(n_1480)
);

INVx3_ASAP7_75t_L g1481 ( 
.A(n_1382),
.Y(n_1481)
);

O2A1O1Ixp33_ASAP7_75t_L g1482 ( 
.A1(n_1317),
.A2(n_835),
.B(n_800),
.C(n_1351),
.Y(n_1482)
);

INVx4_ASAP7_75t_L g1483 ( 
.A(n_1255),
.Y(n_1483)
);

OAI22xp5_ASAP7_75t_SL g1484 ( 
.A1(n_1373),
.A2(n_598),
.B1(n_835),
.B2(n_1139),
.Y(n_1484)
);

NAND3x1_ASAP7_75t_L g1485 ( 
.A(n_1373),
.B(n_1374),
.C(n_1351),
.Y(n_1485)
);

OAI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1349),
.A2(n_1378),
.B(n_1367),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1373),
.A2(n_842),
.B1(n_894),
.B2(n_983),
.Y(n_1487)
);

OAI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1373),
.A2(n_1188),
.B1(n_1003),
.B2(n_1322),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_L g1489 ( 
.A1(n_1360),
.A2(n_1367),
.B(n_1349),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1373),
.B(n_1384),
.Y(n_1490)
);

INVxp67_ASAP7_75t_SL g1491 ( 
.A(n_1379),
.Y(n_1491)
);

BUFx2_ASAP7_75t_L g1492 ( 
.A(n_1365),
.Y(n_1492)
);

INVxp67_ASAP7_75t_L g1493 ( 
.A(n_1332),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_1264),
.B(n_1336),
.Y(n_1494)
);

OAI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1373),
.A2(n_1003),
.B1(n_800),
.B2(n_835),
.Y(n_1495)
);

OAI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1373),
.A2(n_1003),
.B(n_800),
.Y(n_1496)
);

OAI21x1_ASAP7_75t_L g1497 ( 
.A1(n_1360),
.A2(n_1367),
.B(n_1349),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1360),
.A2(n_1367),
.B(n_1349),
.Y(n_1498)
);

INVx3_ASAP7_75t_L g1499 ( 
.A(n_1382),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1239),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1302),
.B(n_1365),
.Y(n_1501)
);

OA21x2_ASAP7_75t_L g1502 ( 
.A1(n_1241),
.A2(n_1242),
.B(n_1257),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1360),
.A2(n_1367),
.B(n_1349),
.Y(n_1503)
);

AOI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1360),
.A2(n_1242),
.B(n_1343),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1393),
.B(n_1476),
.Y(n_1505)
);

BUFx3_ASAP7_75t_L g1506 ( 
.A(n_1443),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1412),
.B(n_1408),
.Y(n_1507)
);

NOR2xp67_ASAP7_75t_L g1508 ( 
.A(n_1483),
.B(n_1424),
.Y(n_1508)
);

BUFx10_ASAP7_75t_L g1509 ( 
.A(n_1433),
.Y(n_1509)
);

OA21x2_ASAP7_75t_L g1510 ( 
.A1(n_1431),
.A2(n_1421),
.B(n_1399),
.Y(n_1510)
);

O2A1O1Ixp5_ASAP7_75t_L g1511 ( 
.A1(n_1473),
.A2(n_1496),
.B(n_1470),
.C(n_1417),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1391),
.B(n_1398),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1397),
.Y(n_1513)
);

AOI21xp5_ASAP7_75t_SL g1514 ( 
.A1(n_1470),
.A2(n_1464),
.B(n_1482),
.Y(n_1514)
);

OA21x2_ASAP7_75t_L g1515 ( 
.A1(n_1395),
.A2(n_1401),
.B(n_1460),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1495),
.A2(n_1490),
.B1(n_1389),
.B2(n_1485),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1501),
.B(n_1410),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1477),
.B(n_1492),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1397),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1389),
.A2(n_1490),
.B1(n_1485),
.B2(n_1487),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1429),
.B(n_1418),
.Y(n_1521)
);

INVxp67_ASAP7_75t_L g1522 ( 
.A(n_1491),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1468),
.A2(n_1487),
.B1(n_1488),
.B2(n_1484),
.Y(n_1523)
);

BUFx3_ASAP7_75t_L g1524 ( 
.A(n_1433),
.Y(n_1524)
);

AOI21xp5_ASAP7_75t_SL g1525 ( 
.A1(n_1445),
.A2(n_1414),
.B(n_1491),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_1430),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1396),
.B(n_1493),
.Y(n_1527)
);

AND2x4_ASAP7_75t_L g1528 ( 
.A(n_1413),
.B(n_1419),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1396),
.B(n_1493),
.Y(n_1529)
);

AOI221x1_ASAP7_75t_SL g1530 ( 
.A1(n_1488),
.A2(n_1428),
.B1(n_1432),
.B2(n_1469),
.C(n_1500),
.Y(n_1530)
);

O2A1O1Ixp5_ASAP7_75t_L g1531 ( 
.A1(n_1459),
.A2(n_1432),
.B(n_1439),
.C(n_1478),
.Y(n_1531)
);

NAND2xp33_ASAP7_75t_SL g1532 ( 
.A(n_1434),
.B(n_1457),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_1430),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1405),
.B(n_1411),
.Y(n_1534)
);

O2A1O1Ixp5_ASAP7_75t_L g1535 ( 
.A1(n_1504),
.A2(n_1445),
.B(n_1454),
.C(n_1420),
.Y(n_1535)
);

INVx1_ASAP7_75t_SL g1536 ( 
.A(n_1458),
.Y(n_1536)
);

OA22x2_ASAP7_75t_L g1537 ( 
.A1(n_1416),
.A2(n_1452),
.B1(n_1449),
.B2(n_1415),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1409),
.B(n_1446),
.Y(n_1538)
);

AND2x4_ASAP7_75t_L g1539 ( 
.A(n_1413),
.B(n_1419),
.Y(n_1539)
);

O2A1O1Ixp5_ASAP7_75t_L g1540 ( 
.A1(n_1454),
.A2(n_1407),
.B(n_1420),
.C(n_1481),
.Y(n_1540)
);

O2A1O1Ixp33_ASAP7_75t_L g1541 ( 
.A1(n_1468),
.A2(n_1437),
.B(n_1403),
.C(n_1390),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1409),
.B(n_1446),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_SL g1543 ( 
.A1(n_1413),
.A2(n_1494),
.B(n_1423),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1440),
.B(n_1403),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1406),
.A2(n_1400),
.B1(n_1440),
.B2(n_1435),
.Y(n_1545)
);

OA21x2_ASAP7_75t_L g1546 ( 
.A1(n_1404),
.A2(n_1503),
.B(n_1498),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1400),
.B(n_1435),
.Y(n_1547)
);

OAI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1499),
.A2(n_1483),
.B1(n_1457),
.B2(n_1434),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1453),
.B(n_1451),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1444),
.B(n_1450),
.Y(n_1550)
);

O2A1O1Ixp5_ASAP7_75t_L g1551 ( 
.A1(n_1447),
.A2(n_1441),
.B(n_1436),
.C(n_1442),
.Y(n_1551)
);

OA21x2_ASAP7_75t_L g1552 ( 
.A1(n_1463),
.A2(n_1427),
.B(n_1479),
.Y(n_1552)
);

OA21x2_ASAP7_75t_L g1553 ( 
.A1(n_1394),
.A2(n_1489),
.B(n_1466),
.Y(n_1553)
);

O2A1O1Ixp33_ASAP7_75t_L g1554 ( 
.A1(n_1474),
.A2(n_1502),
.B(n_1447),
.C(n_1461),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1455),
.Y(n_1555)
);

CKINVDCx16_ASAP7_75t_R g1556 ( 
.A(n_1472),
.Y(n_1556)
);

AOI21xp5_ASAP7_75t_SL g1557 ( 
.A1(n_1423),
.A2(n_1471),
.B(n_1456),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_1472),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1451),
.B(n_1392),
.Y(n_1559)
);

AOI21x1_ASAP7_75t_SL g1560 ( 
.A1(n_1422),
.A2(n_1402),
.B(n_1448),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1462),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1422),
.B(n_1426),
.Y(n_1562)
);

OA21x2_ASAP7_75t_L g1563 ( 
.A1(n_1467),
.A2(n_1497),
.B(n_1475),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1448),
.B(n_1425),
.Y(n_1564)
);

NAND2xp33_ASAP7_75t_SL g1565 ( 
.A(n_1480),
.B(n_1425),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1438),
.B(n_1465),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1486),
.B(n_1393),
.Y(n_1567)
);

BUFx8_ASAP7_75t_SL g1568 ( 
.A(n_1472),
.Y(n_1568)
);

OAI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1473),
.A2(n_1373),
.B1(n_1496),
.B2(n_1495),
.Y(n_1569)
);

O2A1O1Ixp33_ASAP7_75t_L g1570 ( 
.A1(n_1495),
.A2(n_1496),
.B(n_1473),
.C(n_1470),
.Y(n_1570)
);

AOI21xp5_ASAP7_75t_L g1571 ( 
.A1(n_1473),
.A2(n_1496),
.B(n_1401),
.Y(n_1571)
);

O2A1O1Ixp33_ASAP7_75t_L g1572 ( 
.A1(n_1495),
.A2(n_1496),
.B(n_1473),
.C(n_1470),
.Y(n_1572)
);

A2O1A1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_1473),
.A2(n_1496),
.B(n_1373),
.C(n_1003),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_SL g1574 ( 
.A1(n_1484),
.A2(n_1434),
.B1(n_1457),
.B2(n_1389),
.Y(n_1574)
);

A2O1A1Ixp33_ASAP7_75t_L g1575 ( 
.A1(n_1473),
.A2(n_1496),
.B(n_1373),
.C(n_1003),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_1430),
.Y(n_1576)
);

INVx1_ASAP7_75t_SL g1577 ( 
.A(n_1443),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1412),
.B(n_1408),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1412),
.B(n_1408),
.Y(n_1579)
);

AOI211xp5_ASAP7_75t_L g1580 ( 
.A1(n_1495),
.A2(n_1484),
.B(n_1488),
.C(n_1473),
.Y(n_1580)
);

O2A1O1Ixp5_ASAP7_75t_L g1581 ( 
.A1(n_1473),
.A2(n_1496),
.B(n_1470),
.C(n_1417),
.Y(n_1581)
);

OAI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1473),
.A2(n_1373),
.B1(n_1496),
.B2(n_1495),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1412),
.B(n_1408),
.Y(n_1583)
);

NOR2xp67_ASAP7_75t_L g1584 ( 
.A(n_1483),
.B(n_1424),
.Y(n_1584)
);

AOI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1473),
.A2(n_1496),
.B(n_1401),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1412),
.B(n_1408),
.Y(n_1586)
);

INVx4_ASAP7_75t_L g1587 ( 
.A(n_1407),
.Y(n_1587)
);

O2A1O1Ixp5_ASAP7_75t_L g1588 ( 
.A1(n_1473),
.A2(n_1496),
.B(n_1470),
.C(n_1417),
.Y(n_1588)
);

AOI221x1_ASAP7_75t_SL g1589 ( 
.A1(n_1495),
.A2(n_1391),
.B1(n_521),
.B2(n_252),
.C(n_266),
.Y(n_1589)
);

AOI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1473),
.A2(n_1496),
.B(n_1401),
.Y(n_1590)
);

AOI221xp5_ASAP7_75t_L g1591 ( 
.A1(n_1495),
.A2(n_810),
.B1(n_800),
.B2(n_1488),
.C(n_1464),
.Y(n_1591)
);

O2A1O1Ixp33_ASAP7_75t_L g1592 ( 
.A1(n_1495),
.A2(n_1496),
.B(n_1473),
.C(n_1470),
.Y(n_1592)
);

CKINVDCx6p67_ASAP7_75t_R g1593 ( 
.A(n_1556),
.Y(n_1593)
);

NOR2x1_ASAP7_75t_L g1594 ( 
.A(n_1525),
.B(n_1514),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1512),
.B(n_1507),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1526),
.B(n_1533),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1513),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1567),
.B(n_1505),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1555),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1561),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1519),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1578),
.B(n_1579),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1583),
.B(n_1586),
.Y(n_1603)
);

AND2x4_ASAP7_75t_L g1604 ( 
.A(n_1550),
.B(n_1562),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1522),
.B(n_1517),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_SL g1606 ( 
.A(n_1576),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1559),
.Y(n_1607)
);

INVx3_ASAP7_75t_L g1608 ( 
.A(n_1552),
.Y(n_1608)
);

NAND2x1p5_ASAP7_75t_L g1609 ( 
.A(n_1508),
.B(n_1584),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1534),
.Y(n_1610)
);

OA21x2_ASAP7_75t_L g1611 ( 
.A1(n_1531),
.A2(n_1581),
.B(n_1511),
.Y(n_1611)
);

NOR2x1_ASAP7_75t_R g1612 ( 
.A(n_1558),
.B(n_1524),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1527),
.B(n_1529),
.Y(n_1613)
);

HB1xp67_ASAP7_75t_L g1614 ( 
.A(n_1518),
.Y(n_1614)
);

BUFx3_ASAP7_75t_L g1615 ( 
.A(n_1506),
.Y(n_1615)
);

OAI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1573),
.A2(n_1575),
.B(n_1588),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1547),
.B(n_1566),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1571),
.B(n_1585),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1548),
.B(n_1574),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1528),
.B(n_1539),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1549),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1521),
.Y(n_1622)
);

AO21x2_ASAP7_75t_L g1623 ( 
.A1(n_1590),
.A2(n_1554),
.B(n_1523),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1537),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1537),
.Y(n_1625)
);

AO21x2_ASAP7_75t_L g1626 ( 
.A1(n_1520),
.A2(n_1545),
.B(n_1575),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1516),
.B(n_1510),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1510),
.B(n_1515),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1510),
.B(n_1515),
.Y(n_1629)
);

AOI221xp5_ASAP7_75t_L g1630 ( 
.A1(n_1589),
.A2(n_1530),
.B1(n_1591),
.B2(n_1580),
.C(n_1569),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1551),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1540),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1511),
.B(n_1581),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1540),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1588),
.B(n_1538),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1598),
.B(n_1563),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1599),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1600),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1618),
.B(n_1553),
.Y(n_1639)
);

AND2x4_ASAP7_75t_SL g1640 ( 
.A(n_1620),
.B(n_1587),
.Y(n_1640)
);

NAND3xp33_ASAP7_75t_SL g1641 ( 
.A(n_1630),
.B(n_1573),
.C(n_1570),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1597),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1635),
.B(n_1592),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1627),
.B(n_1546),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1627),
.B(n_1582),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1628),
.B(n_1592),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1601),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1628),
.B(n_1570),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1629),
.B(n_1572),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_L g1650 ( 
.A(n_1594),
.B(n_1572),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1629),
.B(n_1535),
.Y(n_1651)
);

NOR2xp67_ASAP7_75t_L g1652 ( 
.A(n_1632),
.B(n_1542),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1608),
.B(n_1544),
.Y(n_1653)
);

BUFx3_ASAP7_75t_L g1654 ( 
.A(n_1609),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1635),
.B(n_1577),
.Y(n_1655)
);

INVx1_ASAP7_75t_SL g1656 ( 
.A(n_1615),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1608),
.B(n_1543),
.Y(n_1657)
);

INVxp67_ASAP7_75t_L g1658 ( 
.A(n_1632),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1637),
.Y(n_1659)
);

NAND3xp33_ASAP7_75t_SL g1660 ( 
.A(n_1643),
.B(n_1650),
.C(n_1616),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1637),
.Y(n_1661)
);

NOR3xp33_ASAP7_75t_L g1662 ( 
.A(n_1641),
.B(n_1594),
.C(n_1616),
.Y(n_1662)
);

AOI21x1_ASAP7_75t_L g1663 ( 
.A1(n_1651),
.A2(n_1634),
.B(n_1631),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1643),
.B(n_1605),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1637),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1645),
.B(n_1614),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1645),
.B(n_1605),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1645),
.B(n_1604),
.Y(n_1668)
);

AOI221xp5_ASAP7_75t_L g1669 ( 
.A1(n_1641),
.A2(n_1626),
.B1(n_1623),
.B2(n_1633),
.C(n_1619),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_R g1670 ( 
.A(n_1650),
.B(n_1565),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1645),
.B(n_1595),
.Y(n_1671)
);

INVx1_ASAP7_75t_SL g1672 ( 
.A(n_1656),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1653),
.B(n_1604),
.Y(n_1673)
);

AND2x4_ASAP7_75t_L g1674 ( 
.A(n_1657),
.B(n_1604),
.Y(n_1674)
);

INVxp67_ASAP7_75t_L g1675 ( 
.A(n_1655),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1657),
.B(n_1620),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_R g1677 ( 
.A(n_1656),
.B(n_1532),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1642),
.Y(n_1678)
);

NOR5xp2_ASAP7_75t_SL g1679 ( 
.A(n_1658),
.B(n_1560),
.C(n_1593),
.D(n_1612),
.E(n_1623),
.Y(n_1679)
);

NOR3xp33_ASAP7_75t_L g1680 ( 
.A(n_1658),
.B(n_1633),
.C(n_1634),
.Y(n_1680)
);

OAI221xp5_ASAP7_75t_L g1681 ( 
.A1(n_1652),
.A2(n_1541),
.B1(n_1611),
.B2(n_1617),
.C(n_1622),
.Y(n_1681)
);

OAI31xp33_ASAP7_75t_L g1682 ( 
.A1(n_1646),
.A2(n_1541),
.A3(n_1609),
.B(n_1625),
.Y(n_1682)
);

OR2x2_ASAP7_75t_L g1683 ( 
.A(n_1646),
.B(n_1613),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1646),
.B(n_1612),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1642),
.Y(n_1685)
);

AOI211xp5_ASAP7_75t_L g1686 ( 
.A1(n_1646),
.A2(n_1624),
.B(n_1625),
.C(n_1631),
.Y(n_1686)
);

OAI222xp33_ASAP7_75t_L g1687 ( 
.A1(n_1648),
.A2(n_1617),
.B1(n_1621),
.B2(n_1624),
.C1(n_1626),
.C2(n_1607),
.Y(n_1687)
);

CKINVDCx20_ASAP7_75t_R g1688 ( 
.A(n_1640),
.Y(n_1688)
);

AOI221xp5_ASAP7_75t_L g1689 ( 
.A1(n_1648),
.A2(n_1626),
.B1(n_1623),
.B2(n_1610),
.C(n_1622),
.Y(n_1689)
);

AOI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1652),
.A2(n_1611),
.B1(n_1648),
.B2(n_1649),
.Y(n_1690)
);

AND2x4_ASAP7_75t_L g1691 ( 
.A(n_1657),
.B(n_1620),
.Y(n_1691)
);

OAI221xp5_ASAP7_75t_L g1692 ( 
.A1(n_1648),
.A2(n_1611),
.B1(n_1610),
.B2(n_1603),
.C(n_1602),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1690),
.B(n_1636),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_SL g1694 ( 
.A(n_1669),
.B(n_1649),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1683),
.B(n_1649),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1678),
.Y(n_1696)
);

OAI21xp5_ASAP7_75t_L g1697 ( 
.A1(n_1662),
.A2(n_1611),
.B(n_1651),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1659),
.Y(n_1698)
);

OA21x2_ASAP7_75t_L g1699 ( 
.A1(n_1689),
.A2(n_1663),
.B(n_1687),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1659),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1668),
.B(n_1636),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1668),
.B(n_1673),
.Y(n_1702)
);

NAND3xp33_ASAP7_75t_SL g1703 ( 
.A(n_1692),
.B(n_1651),
.C(n_1644),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1661),
.Y(n_1704)
);

INVx3_ASAP7_75t_L g1705 ( 
.A(n_1663),
.Y(n_1705)
);

BUFx3_ASAP7_75t_L g1706 ( 
.A(n_1688),
.Y(n_1706)
);

BUFx3_ASAP7_75t_L g1707 ( 
.A(n_1688),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1671),
.B(n_1638),
.Y(n_1708)
);

BUFx2_ASAP7_75t_L g1709 ( 
.A(n_1685),
.Y(n_1709)
);

BUFx3_ASAP7_75t_L g1710 ( 
.A(n_1672),
.Y(n_1710)
);

INVx4_ASAP7_75t_SL g1711 ( 
.A(n_1691),
.Y(n_1711)
);

BUFx6f_ASAP7_75t_L g1712 ( 
.A(n_1660),
.Y(n_1712)
);

OR2x6_ASAP7_75t_L g1713 ( 
.A(n_1674),
.B(n_1557),
.Y(n_1713)
);

HB1xp67_ASAP7_75t_L g1714 ( 
.A(n_1665),
.Y(n_1714)
);

INVxp67_ASAP7_75t_L g1715 ( 
.A(n_1681),
.Y(n_1715)
);

INVx3_ASAP7_75t_L g1716 ( 
.A(n_1674),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1664),
.B(n_1683),
.Y(n_1717)
);

INVx4_ASAP7_75t_SL g1718 ( 
.A(n_1691),
.Y(n_1718)
);

AND4x1_ASAP7_75t_L g1719 ( 
.A(n_1682),
.B(n_1596),
.C(n_1564),
.D(n_1593),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1664),
.B(n_1647),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1714),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1694),
.B(n_1666),
.Y(n_1722)
);

AND2x4_ASAP7_75t_L g1723 ( 
.A(n_1711),
.B(n_1674),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1714),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1717),
.B(n_1680),
.Y(n_1725)
);

INVx1_ASAP7_75t_SL g1726 ( 
.A(n_1706),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1698),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1695),
.B(n_1667),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1717),
.B(n_1667),
.Y(n_1729)
);

INVx1_ASAP7_75t_SL g1730 ( 
.A(n_1706),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1711),
.B(n_1718),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1698),
.Y(n_1732)
);

AND3x1_ASAP7_75t_L g1733 ( 
.A(n_1697),
.B(n_1684),
.C(n_1686),
.Y(n_1733)
);

NOR3xp33_ASAP7_75t_SL g1734 ( 
.A(n_1703),
.B(n_1679),
.C(n_1606),
.Y(n_1734)
);

NAND2x1_ASAP7_75t_L g1735 ( 
.A(n_1716),
.B(n_1693),
.Y(n_1735)
);

OR2x6_ASAP7_75t_L g1736 ( 
.A(n_1697),
.B(n_1713),
.Y(n_1736)
);

INVx4_ASAP7_75t_L g1737 ( 
.A(n_1712),
.Y(n_1737)
);

INVx4_ASAP7_75t_L g1738 ( 
.A(n_1712),
.Y(n_1738)
);

NAND3xp33_ASAP7_75t_L g1739 ( 
.A(n_1712),
.B(n_1651),
.C(n_1639),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1700),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1720),
.B(n_1675),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1696),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1700),
.Y(n_1743)
);

NAND2x1p5_ASAP7_75t_L g1744 ( 
.A(n_1719),
.B(n_1654),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1718),
.B(n_1702),
.Y(n_1745)
);

INVx1_ASAP7_75t_SL g1746 ( 
.A(n_1706),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1704),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1718),
.B(n_1676),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1716),
.B(n_1693),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1702),
.B(n_1676),
.Y(n_1750)
);

INVx2_ASAP7_75t_SL g1751 ( 
.A(n_1731),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1729),
.B(n_1720),
.Y(n_1752)
);

NAND2x1_ASAP7_75t_L g1753 ( 
.A(n_1731),
.B(n_1716),
.Y(n_1753)
);

AOI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1733),
.A2(n_1712),
.B1(n_1715),
.B2(n_1703),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1745),
.B(n_1750),
.Y(n_1755)
);

INVxp67_ASAP7_75t_SL g1756 ( 
.A(n_1744),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1726),
.B(n_1712),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1729),
.B(n_1720),
.Y(n_1758)
);

AND2x2_ASAP7_75t_SL g1759 ( 
.A(n_1733),
.B(n_1712),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1726),
.B(n_1712),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1730),
.B(n_1715),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1742),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1742),
.Y(n_1763)
);

AND2x4_ASAP7_75t_L g1764 ( 
.A(n_1745),
.B(n_1707),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1749),
.Y(n_1765)
);

INVxp67_ASAP7_75t_L g1766 ( 
.A(n_1730),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1746),
.B(n_1710),
.Y(n_1767)
);

NOR2x1_ASAP7_75t_L g1768 ( 
.A(n_1737),
.B(n_1707),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1749),
.Y(n_1769)
);

INVx3_ASAP7_75t_L g1770 ( 
.A(n_1735),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1728),
.B(n_1696),
.Y(n_1771)
);

OR2x2_ASAP7_75t_L g1772 ( 
.A(n_1728),
.B(n_1708),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1749),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1727),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1727),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1732),
.Y(n_1776)
);

NAND2xp33_ASAP7_75t_SL g1777 ( 
.A(n_1734),
.B(n_1677),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1746),
.B(n_1710),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1750),
.B(n_1702),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1744),
.B(n_1716),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1732),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1725),
.B(n_1710),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1740),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1744),
.B(n_1701),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1749),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1725),
.B(n_1709),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1741),
.B(n_1708),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_SL g1788 ( 
.A(n_1759),
.B(n_1744),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1759),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1754),
.B(n_1721),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1766),
.B(n_1721),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1762),
.B(n_1724),
.Y(n_1792)
);

NOR2x1_ASAP7_75t_L g1793 ( 
.A(n_1768),
.B(n_1737),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1779),
.B(n_1723),
.Y(n_1794)
);

INVx1_ASAP7_75t_SL g1795 ( 
.A(n_1767),
.Y(n_1795)
);

INVx3_ASAP7_75t_SL g1796 ( 
.A(n_1764),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1779),
.B(n_1734),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1774),
.Y(n_1798)
);

INVx1_ASAP7_75t_SL g1799 ( 
.A(n_1778),
.Y(n_1799)
);

NAND2xp33_ASAP7_75t_R g1800 ( 
.A(n_1757),
.B(n_1670),
.Y(n_1800)
);

AOI22xp33_ASAP7_75t_L g1801 ( 
.A1(n_1784),
.A2(n_1699),
.B1(n_1739),
.B2(n_1736),
.Y(n_1801)
);

AND2x4_ASAP7_75t_L g1802 ( 
.A(n_1755),
.B(n_1723),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1755),
.B(n_1723),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1765),
.Y(n_1804)
);

INVx1_ASAP7_75t_SL g1805 ( 
.A(n_1761),
.Y(n_1805)
);

HB1xp67_ASAP7_75t_L g1806 ( 
.A(n_1782),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1765),
.Y(n_1807)
);

NAND2xp33_ASAP7_75t_L g1808 ( 
.A(n_1777),
.B(n_1760),
.Y(n_1808)
);

INVx1_ASAP7_75t_SL g1809 ( 
.A(n_1764),
.Y(n_1809)
);

INVxp67_ASAP7_75t_SL g1810 ( 
.A(n_1786),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1763),
.B(n_1724),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1764),
.B(n_1723),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1769),
.Y(n_1813)
);

HB1xp67_ASAP7_75t_L g1814 ( 
.A(n_1775),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1776),
.Y(n_1815)
);

AOI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1801),
.A2(n_1699),
.B1(n_1739),
.B2(n_1737),
.Y(n_1816)
);

OA21x2_ASAP7_75t_SL g1817 ( 
.A1(n_1805),
.A2(n_1777),
.B(n_1722),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1814),
.Y(n_1818)
);

OAI21xp33_ASAP7_75t_L g1819 ( 
.A1(n_1797),
.A2(n_1773),
.B(n_1769),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1805),
.B(n_1806),
.Y(n_1820)
);

AOI221xp5_ASAP7_75t_L g1821 ( 
.A1(n_1790),
.A2(n_1737),
.B1(n_1738),
.B2(n_1756),
.C(n_1705),
.Y(n_1821)
);

NAND3xp33_ASAP7_75t_L g1822 ( 
.A(n_1790),
.B(n_1738),
.C(n_1773),
.Y(n_1822)
);

OAI21xp5_ASAP7_75t_L g1823 ( 
.A1(n_1810),
.A2(n_1738),
.B(n_1722),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1796),
.B(n_1751),
.Y(n_1824)
);

OAI22xp33_ASAP7_75t_SL g1825 ( 
.A1(n_1789),
.A2(n_1738),
.B1(n_1736),
.B2(n_1735),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1794),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1794),
.Y(n_1827)
);

NOR2x1_ASAP7_75t_L g1828 ( 
.A(n_1793),
.B(n_1770),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1814),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1806),
.B(n_1785),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1796),
.B(n_1751),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1810),
.B(n_1781),
.Y(n_1832)
);

OAI22xp5_ASAP7_75t_L g1833 ( 
.A1(n_1795),
.A2(n_1799),
.B1(n_1788),
.B2(n_1797),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1804),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1796),
.B(n_1785),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1834),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1826),
.B(n_1812),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1818),
.Y(n_1838)
);

OR2x2_ASAP7_75t_L g1839 ( 
.A(n_1820),
.B(n_1795),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1829),
.B(n_1799),
.Y(n_1840)
);

NOR3xp33_ASAP7_75t_L g1841 ( 
.A(n_1833),
.B(n_1789),
.C(n_1808),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1827),
.B(n_1812),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1832),
.B(n_1809),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1824),
.B(n_1809),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1830),
.Y(n_1845)
);

NOR2xp33_ASAP7_75t_L g1846 ( 
.A(n_1831),
.B(n_1568),
.Y(n_1846)
);

AOI221xp5_ASAP7_75t_L g1847 ( 
.A1(n_1841),
.A2(n_1833),
.B1(n_1816),
.B2(n_1789),
.C(n_1822),
.Y(n_1847)
);

NOR2xp67_ASAP7_75t_L g1848 ( 
.A(n_1846),
.B(n_1770),
.Y(n_1848)
);

AOI22xp5_ASAP7_75t_L g1849 ( 
.A1(n_1844),
.A2(n_1699),
.B1(n_1797),
.B2(n_1819),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_SL g1850 ( 
.A(n_1839),
.B(n_1825),
.Y(n_1850)
);

AOI211xp5_ASAP7_75t_L g1851 ( 
.A1(n_1840),
.A2(n_1823),
.B(n_1817),
.C(n_1821),
.Y(n_1851)
);

NOR4xp25_ASAP7_75t_L g1852 ( 
.A(n_1840),
.B(n_1832),
.C(n_1823),
.D(n_1835),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1837),
.B(n_1804),
.Y(n_1853)
);

AOI31xp33_ASAP7_75t_L g1854 ( 
.A1(n_1843),
.A2(n_1828),
.A3(n_1793),
.B(n_1791),
.Y(n_1854)
);

AOI21xp5_ASAP7_75t_SL g1855 ( 
.A1(n_1843),
.A2(n_1791),
.B(n_1792),
.Y(n_1855)
);

AOI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1842),
.A2(n_1811),
.B(n_1792),
.Y(n_1856)
);

AOI221xp5_ASAP7_75t_L g1857 ( 
.A1(n_1852),
.A2(n_1836),
.B1(n_1845),
.B2(n_1838),
.C(n_1798),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_SL g1858 ( 
.A(n_1847),
.B(n_1770),
.Y(n_1858)
);

OAI21xp33_ASAP7_75t_L g1859 ( 
.A1(n_1849),
.A2(n_1803),
.B(n_1802),
.Y(n_1859)
);

BUFx2_ASAP7_75t_L g1860 ( 
.A(n_1853),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_SL g1861 ( 
.A(n_1851),
.B(n_1802),
.Y(n_1861)
);

OAI211xp5_ASAP7_75t_SL g1862 ( 
.A1(n_1850),
.A2(n_1811),
.B(n_1807),
.C(n_1813),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1860),
.Y(n_1863)
);

CKINVDCx16_ASAP7_75t_R g1864 ( 
.A(n_1861),
.Y(n_1864)
);

NAND3xp33_ASAP7_75t_L g1865 ( 
.A(n_1857),
.B(n_1862),
.C(n_1854),
.Y(n_1865)
);

NAND3xp33_ASAP7_75t_L g1866 ( 
.A(n_1858),
.B(n_1855),
.C(n_1856),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1859),
.Y(n_1867)
);

INVx3_ASAP7_75t_L g1868 ( 
.A(n_1860),
.Y(n_1868)
);

OAI32xp33_ASAP7_75t_L g1869 ( 
.A1(n_1862),
.A2(n_1804),
.A3(n_1807),
.B1(n_1813),
.B2(n_1815),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1868),
.Y(n_1870)
);

AOI221xp5_ASAP7_75t_SL g1871 ( 
.A1(n_1867),
.A2(n_1813),
.B1(n_1807),
.B2(n_1815),
.C(n_1798),
.Y(n_1871)
);

AOI211xp5_ASAP7_75t_L g1872 ( 
.A1(n_1865),
.A2(n_1848),
.B(n_1780),
.C(n_1784),
.Y(n_1872)
);

CKINVDCx20_ASAP7_75t_R g1873 ( 
.A(n_1864),
.Y(n_1873)
);

NOR2x1_ASAP7_75t_L g1874 ( 
.A(n_1866),
.B(n_1802),
.Y(n_1874)
);

XNOR2xp5_ASAP7_75t_SL g1875 ( 
.A(n_1870),
.B(n_1863),
.Y(n_1875)
);

AND2x4_ASAP7_75t_L g1876 ( 
.A(n_1873),
.B(n_1802),
.Y(n_1876)
);

OAI21xp5_ASAP7_75t_L g1877 ( 
.A1(n_1874),
.A2(n_1869),
.B(n_1780),
.Y(n_1877)
);

NAND4xp75_ASAP7_75t_L g1878 ( 
.A(n_1877),
.B(n_1871),
.C(n_1872),
.D(n_1803),
.Y(n_1878)
);

OAI221xp5_ASAP7_75t_L g1879 ( 
.A1(n_1878),
.A2(n_1875),
.B1(n_1800),
.B2(n_1736),
.C(n_1753),
.Y(n_1879)
);

CKINVDCx20_ASAP7_75t_R g1880 ( 
.A(n_1879),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1879),
.Y(n_1881)
);

OAI321xp33_ASAP7_75t_L g1882 ( 
.A1(n_1881),
.A2(n_1876),
.A3(n_1736),
.B1(n_1783),
.B2(n_1771),
.C(n_1787),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1880),
.Y(n_1883)
);

OAI22x1_ASAP7_75t_SL g1884 ( 
.A1(n_1883),
.A2(n_1882),
.B1(n_1536),
.B2(n_1509),
.Y(n_1884)
);

OAI22xp5_ASAP7_75t_L g1885 ( 
.A1(n_1883),
.A2(n_1752),
.B1(n_1758),
.B2(n_1771),
.Y(n_1885)
);

OAI311xp33_ASAP7_75t_L g1886 ( 
.A1(n_1884),
.A2(n_1758),
.A3(n_1752),
.B1(n_1787),
.C1(n_1772),
.Y(n_1886)
);

OAI21xp5_ASAP7_75t_L g1887 ( 
.A1(n_1886),
.A2(n_1885),
.B(n_1753),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1887),
.B(n_1705),
.Y(n_1888)
);

AOI22xp33_ASAP7_75t_L g1889 ( 
.A1(n_1888),
.A2(n_1736),
.B1(n_1705),
.B2(n_1772),
.Y(n_1889)
);

AOI221xp5_ASAP7_75t_L g1890 ( 
.A1(n_1889),
.A2(n_1705),
.B1(n_1740),
.B2(n_1743),
.C(n_1747),
.Y(n_1890)
);

AOI211xp5_ASAP7_75t_L g1891 ( 
.A1(n_1890),
.A2(n_1509),
.B(n_1707),
.C(n_1748),
.Y(n_1891)
);


endmodule