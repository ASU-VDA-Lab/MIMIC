module fake_ariane_1664_n_1808 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1808);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1808;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_677;
wire n_604;
wire n_439;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1777;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1252;
wire n_1129;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_31),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_109),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_120),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_22),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_48),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_4),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_116),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_160),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_75),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_28),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_84),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_8),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_3),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_137),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_85),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_143),
.Y(n_185)
);

BUFx10_ASAP7_75t_L g186 ( 
.A(n_76),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_61),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_130),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_127),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_114),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_11),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_72),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_50),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_47),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_86),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_95),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_128),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_112),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_65),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_122),
.Y(n_200)
);

BUFx2_ASAP7_75t_SL g201 ( 
.A(n_60),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_7),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_101),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_45),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_38),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_49),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_159),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_7),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_110),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_111),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_106),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_88),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_48),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_102),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_15),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_99),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_119),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_83),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_78),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_133),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_92),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_140),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_124),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_161),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_32),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_53),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_64),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_18),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_42),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_113),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_59),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_165),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_70),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_3),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_93),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_90),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_163),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_117),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_52),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_164),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_69),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_15),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_82),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_162),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_63),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_10),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_16),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_60),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_25),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_132),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_10),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_45),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_100),
.Y(n_253)
);

BUFx8_ASAP7_75t_SL g254 ( 
.A(n_87),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_126),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_156),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_0),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_42),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_36),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_18),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_9),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_1),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_50),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_157),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_134),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_68),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_68),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_61),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_4),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_142),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_13),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_55),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_36),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_64),
.Y(n_274)
);

BUFx2_ASAP7_75t_SL g275 ( 
.A(n_6),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_2),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_31),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_148),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_16),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_158),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_69),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_138),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_29),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_33),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_8),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_34),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_141),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_34),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_54),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_51),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_27),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_12),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_118),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_52),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_37),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_107),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_149),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_11),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_97),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_103),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_13),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_9),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_58),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_65),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_56),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_62),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_58),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_44),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_125),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_81),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_30),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_136),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_44),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_38),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_104),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_2),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_150),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_32),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_39),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_129),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_62),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_96),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_94),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_145),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_26),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_74),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_27),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_29),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_108),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_59),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_30),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_228),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_228),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_228),
.Y(n_334)
);

INVxp33_ASAP7_75t_SL g335 ( 
.A(n_194),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_228),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_183),
.B(n_168),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_168),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_291),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_260),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_170),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_254),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_194),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_183),
.B(n_0),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_230),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_182),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_170),
.B(n_1),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_174),
.B(n_5),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_174),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_188),
.Y(n_350)
);

INVxp33_ASAP7_75t_SL g351 ( 
.A(n_201),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_189),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_250),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_177),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_270),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_177),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_226),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_226),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_279),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_279),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_167),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_172),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_184),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_173),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_291),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_178),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_184),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_190),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_190),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_192),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_180),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_181),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_187),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_191),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_192),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_196),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_196),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_229),
.Y(n_378)
);

NOR2xp67_ASAP7_75t_L g379 ( 
.A(n_246),
.B(n_5),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_269),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_202),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_204),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_197),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_197),
.B(n_6),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_198),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_198),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_207),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_284),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_313),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_207),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_239),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_210),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_210),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_211),
.B(n_12),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_211),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_242),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_193),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_245),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_212),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_212),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_247),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_195),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_214),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_230),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_214),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_224),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_221),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_195),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_221),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_256),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_223),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_193),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_223),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_235),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_235),
.Y(n_415)
);

BUFx2_ASAP7_75t_SL g416 ( 
.A(n_186),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_238),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_195),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_238),
.B(n_14),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_332),
.Y(n_420)
);

AND2x6_ASAP7_75t_L g421 ( 
.A(n_338),
.B(n_209),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_337),
.B(n_264),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_416),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_397),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_397),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_397),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_332),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_333),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_333),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_365),
.B(n_291),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_357),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_346),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_412),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_334),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_334),
.B(n_336),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_336),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_338),
.Y(n_437)
);

INVx2_ASAP7_75t_SL g438 ( 
.A(n_402),
.Y(n_438)
);

INVx5_ASAP7_75t_L g439 ( 
.A(n_412),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_402),
.B(n_264),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_412),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_341),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_341),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_349),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_349),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_416),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_365),
.B(n_227),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_344),
.B(n_193),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_358),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_354),
.B(n_227),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_402),
.B(n_287),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_408),
.B(n_227),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_408),
.B(n_287),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_345),
.B(n_379),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_354),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_345),
.B(n_186),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_408),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_356),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_356),
.B(n_328),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_363),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_359),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_363),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_367),
.B(n_368),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_367),
.B(n_328),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_368),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_369),
.B(n_299),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_369),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_370),
.B(n_328),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_370),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_375),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_375),
.B(n_246),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_376),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_376),
.B(n_193),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_377),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_377),
.Y(n_475)
);

AND2x4_ASAP7_75t_L g476 ( 
.A(n_383),
.B(n_193),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_383),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_385),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_385),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_386),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_350),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_386),
.Y(n_482)
);

INVx4_ASAP7_75t_L g483 ( 
.A(n_387),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_418),
.B(n_186),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_387),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_390),
.B(n_299),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_390),
.B(n_392),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_392),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_393),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_393),
.Y(n_490)
);

OA21x2_ASAP7_75t_L g491 ( 
.A1(n_395),
.A2(n_317),
.B(n_315),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_395),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_399),
.B(n_315),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_399),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_400),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_400),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_403),
.Y(n_497)
);

AND2x2_ASAP7_75t_SL g498 ( 
.A(n_456),
.B(n_219),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_430),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_469),
.Y(n_500)
);

INVx5_ASAP7_75t_L g501 ( 
.A(n_421),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_423),
.B(n_362),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_457),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_457),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_459),
.B(n_468),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_469),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_425),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_469),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_457),
.Y(n_509)
);

AOI22xp33_ASAP7_75t_L g510 ( 
.A1(n_422),
.A2(n_335),
.B1(n_456),
.B2(n_448),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_457),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_430),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_469),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_457),
.Y(n_514)
);

INVx1_ASAP7_75t_SL g515 ( 
.A(n_432),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_469),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_425),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_469),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_423),
.B(n_364),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_469),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_425),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_457),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_457),
.Y(n_523)
);

AND2x6_ASAP7_75t_L g524 ( 
.A(n_473),
.B(n_219),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_484),
.B(n_186),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_469),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_457),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_446),
.B(n_366),
.Y(n_528)
);

OAI22x1_ASAP7_75t_L g529 ( 
.A1(n_432),
.A2(n_481),
.B1(n_343),
.B2(n_360),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_446),
.A2(n_351),
.B1(n_394),
.B2(n_347),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_472),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_422),
.B(n_339),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_448),
.A2(n_384),
.B1(n_348),
.B2(n_379),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_431),
.Y(n_534)
);

AND2x6_ASAP7_75t_L g535 ( 
.A(n_473),
.B(n_476),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_425),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_454),
.B(n_371),
.Y(n_537)
);

BUFx8_ASAP7_75t_SL g538 ( 
.A(n_481),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_433),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_472),
.Y(n_540)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_430),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_461),
.B(n_361),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_433),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_433),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_472),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_433),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_454),
.B(n_373),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_438),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_431),
.B(n_374),
.Y(n_549)
);

OR2x6_ASAP7_75t_L g550 ( 
.A(n_471),
.B(n_419),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_472),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_483),
.B(n_381),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_483),
.B(n_382),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_472),
.Y(n_554)
);

OAI22xp33_ASAP7_75t_L g555 ( 
.A1(n_484),
.A2(n_171),
.B1(n_277),
.B2(n_268),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_441),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_472),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_441),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_431),
.A2(n_449),
.B1(n_306),
.B2(n_307),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_467),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_472),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_472),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_449),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_490),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_490),
.Y(n_565)
);

INVx1_ASAP7_75t_SL g566 ( 
.A(n_449),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_441),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_447),
.Y(n_568)
);

INVx4_ASAP7_75t_SL g569 ( 
.A(n_421),
.Y(n_569)
);

AND3x2_ASAP7_75t_L g570 ( 
.A(n_447),
.B(n_391),
.C(n_372),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_490),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_490),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_483),
.B(n_405),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_471),
.A2(n_257),
.B1(n_318),
.B2(n_252),
.Y(n_574)
);

INVx1_ASAP7_75t_SL g575 ( 
.A(n_447),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_421),
.Y(n_576)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_459),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_483),
.B(n_405),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_441),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_490),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_490),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_490),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_471),
.B(n_396),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_490),
.Y(n_584)
);

NAND3xp33_ASAP7_75t_L g585 ( 
.A(n_437),
.B(n_409),
.C(n_407),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_471),
.B(n_398),
.Y(n_586)
);

BUFx8_ASAP7_75t_SL g587 ( 
.A(n_450),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_495),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_495),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_495),
.Y(n_590)
);

CKINVDCx11_ASAP7_75t_R g591 ( 
.A(n_471),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_495),
.Y(n_592)
);

OR2x2_ASAP7_75t_L g593 ( 
.A(n_463),
.B(n_352),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_495),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_495),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_467),
.B(n_407),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_467),
.B(n_401),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_495),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_463),
.B(n_353),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_495),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_459),
.B(n_409),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_497),
.Y(n_602)
);

AND2x6_ASAP7_75t_L g603 ( 
.A(n_473),
.B(n_219),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_497),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_L g605 ( 
.A1(n_487),
.A2(n_288),
.B1(n_259),
.B2(n_261),
.Y(n_605)
);

OAI22xp33_ASAP7_75t_L g606 ( 
.A1(n_466),
.A2(n_283),
.B1(n_286),
.B2(n_298),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_497),
.Y(n_607)
);

NOR3xp33_ASAP7_75t_L g608 ( 
.A(n_487),
.B(n_205),
.C(n_199),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_497),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_468),
.B(n_411),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_497),
.Y(n_611)
);

INVx5_ASAP7_75t_L g612 ( 
.A(n_421),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_497),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_497),
.Y(n_614)
);

OAI22xp33_ASAP7_75t_L g615 ( 
.A1(n_466),
.A2(n_404),
.B1(n_342),
.B2(n_263),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_467),
.B(n_411),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_497),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_443),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_467),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_464),
.A2(n_281),
.B1(n_316),
.B2(n_262),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_482),
.B(n_406),
.Y(n_621)
);

INVx5_ASAP7_75t_L g622 ( 
.A(n_421),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_424),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_443),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_443),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_482),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_424),
.Y(n_627)
);

BUFx4f_ASAP7_75t_L g628 ( 
.A(n_421),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_482),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_482),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_443),
.Y(n_631)
);

INVx1_ASAP7_75t_SL g632 ( 
.A(n_440),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_452),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_482),
.B(n_410),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_444),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_488),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_468),
.B(n_413),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_488),
.B(n_413),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_488),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_452),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_452),
.Y(n_641)
);

NOR2x1p5_ASAP7_75t_L g642 ( 
.A(n_435),
.B(n_199),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_452),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_488),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_488),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_420),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_420),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_632),
.B(n_437),
.Y(n_648)
);

NAND2xp33_ASAP7_75t_SL g649 ( 
.A(n_532),
.B(n_442),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_618),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_618),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_566),
.B(n_486),
.Y(n_652)
);

NAND2x1_ASAP7_75t_L g653 ( 
.A(n_576),
.B(n_421),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_624),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_646),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_537),
.B(n_440),
.Y(n_656)
);

INVx5_ASAP7_75t_L g657 ( 
.A(n_576),
.Y(n_657)
);

BUFx2_ASAP7_75t_L g658 ( 
.A(n_534),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_538),
.Y(n_659)
);

O2A1O1Ixp33_ASAP7_75t_L g660 ( 
.A1(n_499),
.A2(n_435),
.B(n_445),
.C(n_442),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_563),
.B(n_340),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_647),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_499),
.B(n_452),
.Y(n_663)
);

NOR2x1p5_ASAP7_75t_L g664 ( 
.A(n_593),
.B(n_599),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_547),
.B(n_451),
.Y(n_665)
);

A2O1A1Ixp33_ASAP7_75t_L g666 ( 
.A1(n_498),
.A2(n_455),
.B(n_458),
.C(n_444),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_498),
.A2(n_491),
.B1(n_421),
.B2(n_450),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_629),
.Y(n_668)
);

AND2x2_ASAP7_75t_SL g669 ( 
.A(n_498),
.B(n_491),
.Y(n_669)
);

INVx8_ASAP7_75t_L g670 ( 
.A(n_535),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_624),
.Y(n_671)
);

AOI22xp33_ASAP7_75t_L g672 ( 
.A1(n_524),
.A2(n_491),
.B1(n_421),
.B2(n_450),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_577),
.B(n_445),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_575),
.B(n_355),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_629),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_577),
.B(n_462),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_576),
.B(n_462),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_552),
.B(n_475),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_576),
.B(n_475),
.Y(n_679)
);

INVx2_ASAP7_75t_SL g680 ( 
.A(n_593),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_636),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_553),
.B(n_478),
.Y(n_682)
);

INVxp33_ASAP7_75t_L g683 ( 
.A(n_542),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_625),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_633),
.Y(n_685)
);

AO22x2_ASAP7_75t_L g686 ( 
.A1(n_575),
.A2(n_201),
.B1(n_275),
.B2(n_414),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_510),
.A2(n_480),
.B1(n_494),
.B2(n_478),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_636),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_507),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_599),
.B(n_451),
.Y(n_690)
);

NAND2xp33_ASAP7_75t_SL g691 ( 
.A(n_512),
.B(n_479),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_601),
.B(n_479),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_525),
.B(n_453),
.Y(n_693)
);

INVxp67_ASAP7_75t_L g694 ( 
.A(n_515),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_525),
.B(n_453),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_628),
.B(n_480),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_507),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_512),
.B(n_489),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_639),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_639),
.Y(n_700)
);

INVxp67_ASAP7_75t_L g701 ( 
.A(n_542),
.Y(n_701)
);

INVx5_ASAP7_75t_L g702 ( 
.A(n_524),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_601),
.B(n_489),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_610),
.B(n_494),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_610),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_644),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_560),
.Y(n_707)
);

OR2x2_ASAP7_75t_L g708 ( 
.A(n_559),
.B(n_486),
.Y(n_708)
);

OR2x6_ASAP7_75t_L g709 ( 
.A(n_541),
.B(n_529),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_626),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_541),
.B(n_464),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_637),
.B(n_464),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_626),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_568),
.B(n_378),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_633),
.B(n_427),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_628),
.B(n_444),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_560),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_530),
.A2(n_421),
.B1(n_464),
.B2(n_450),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_637),
.B(n_464),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_505),
.B(n_444),
.Y(n_720)
);

A2O1A1Ixp33_ASAP7_75t_L g721 ( 
.A1(n_585),
.A2(n_496),
.B(n_455),
.C(n_492),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_625),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_628),
.B(n_455),
.Y(n_723)
);

BUFx5_ASAP7_75t_L g724 ( 
.A(n_535),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_501),
.B(n_455),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_505),
.B(n_458),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_501),
.B(n_458),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_642),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_630),
.Y(n_729)
);

OAI221xp5_ASAP7_75t_L g730 ( 
.A1(n_620),
.A2(n_205),
.B1(n_311),
.B2(n_206),
.C(n_314),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_597),
.B(n_502),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_630),
.B(n_645),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_630),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_524),
.A2(n_491),
.B1(n_421),
.B2(n_450),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_631),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_645),
.B(n_458),
.Y(n_736)
);

NOR3xp33_ASAP7_75t_L g737 ( 
.A(n_549),
.B(n_213),
.C(n_206),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_620),
.B(n_380),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_640),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_640),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_641),
.B(n_460),
.Y(n_741)
);

OAI21xp33_ASAP7_75t_L g742 ( 
.A1(n_533),
.A2(n_428),
.B(n_427),
.Y(n_742)
);

INVx8_ASAP7_75t_L g743 ( 
.A(n_535),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_550),
.A2(n_535),
.B1(n_643),
.B2(n_641),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_643),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_501),
.B(n_460),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_535),
.B(n_460),
.Y(n_747)
);

OAI22xp5_ASAP7_75t_L g748 ( 
.A1(n_550),
.A2(n_436),
.B1(n_428),
.B2(n_429),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_560),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_519),
.B(n_429),
.Y(n_750)
);

BUFx2_ASAP7_75t_L g751 ( 
.A(n_587),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_619),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_535),
.B(n_460),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_535),
.B(n_465),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_517),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_L g756 ( 
.A1(n_550),
.A2(n_436),
.B1(n_434),
.B2(n_493),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_642),
.B(n_573),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_501),
.B(n_465),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_528),
.B(n_434),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_529),
.B(n_388),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_578),
.B(n_465),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_550),
.A2(n_450),
.B1(n_493),
.B2(n_492),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_635),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_569),
.B(n_473),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_619),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_635),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_583),
.B(n_470),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_596),
.B(n_470),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_524),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_501),
.B(n_470),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_616),
.B(n_474),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_638),
.B(n_474),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_517),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_569),
.B(n_473),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_521),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_521),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_501),
.B(n_474),
.Y(n_777)
);

OR2x2_ASAP7_75t_L g778 ( 
.A(n_574),
.B(n_389),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_536),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_536),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_550),
.B(n_474),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_548),
.B(n_477),
.Y(n_782)
);

INVxp67_ASAP7_75t_L g783 ( 
.A(n_586),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_539),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_548),
.B(n_477),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_524),
.A2(n_492),
.B1(n_485),
.B2(n_477),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_612),
.B(n_477),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_591),
.B(n_485),
.Y(n_788)
);

NAND3xp33_ASAP7_75t_L g789 ( 
.A(n_605),
.B(n_496),
.C(n_485),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_524),
.A2(n_491),
.B1(n_415),
.B2(n_417),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_539),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_543),
.Y(n_792)
);

OR2x6_ASAP7_75t_L g793 ( 
.A(n_621),
.B(n_634),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_543),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_544),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_548),
.B(n_496),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_L g797 ( 
.A1(n_602),
.A2(n_266),
.B1(n_267),
.B2(n_271),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_544),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_546),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_555),
.B(n_292),
.Y(n_800)
);

NOR2xp67_ASAP7_75t_L g801 ( 
.A(n_585),
.B(n_414),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_546),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_556),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_524),
.B(n_473),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_570),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_603),
.B(n_476),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_603),
.A2(n_491),
.B1(n_329),
.B2(n_324),
.Y(n_807)
);

OAI22xp5_ASAP7_75t_L g808 ( 
.A1(n_571),
.A2(n_330),
.B1(n_295),
.B2(n_301),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_670),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_690),
.B(n_603),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_690),
.B(n_603),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_656),
.B(n_603),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_782),
.A2(n_522),
.B(n_503),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_780),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_785),
.A2(n_527),
.B(n_523),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_796),
.A2(n_527),
.B(n_523),
.Y(n_816)
);

A2O1A1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_656),
.A2(n_584),
.B(n_617),
.C(n_571),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_665),
.B(n_603),
.Y(n_818)
);

AOI21xp33_ASAP7_75t_L g819 ( 
.A1(n_800),
.A2(n_606),
.B(n_615),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_677),
.A2(n_527),
.B(n_523),
.Y(n_820)
);

OAI21xp5_ASAP7_75t_L g821 ( 
.A1(n_747),
.A2(n_506),
.B(n_500),
.Y(n_821)
);

NOR2x1_ASAP7_75t_L g822 ( 
.A(n_652),
.B(n_664),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_724),
.B(n_545),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_665),
.B(n_608),
.Y(n_824)
);

BUFx12f_ASAP7_75t_L g825 ( 
.A(n_659),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_648),
.B(n_571),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_674),
.B(n_476),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_714),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_788),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_715),
.B(n_584),
.Y(n_830)
);

O2A1O1Ixp33_ASAP7_75t_SL g831 ( 
.A1(n_666),
.A2(n_513),
.B(n_516),
.C(n_508),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_753),
.A2(n_518),
.B(n_516),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_715),
.B(n_584),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_751),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_650),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_698),
.B(n_617),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_698),
.B(n_617),
.Y(n_837)
);

BUFx4f_ASAP7_75t_L g838 ( 
.A(n_793),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_679),
.A2(n_732),
.B(n_736),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_693),
.B(n_556),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_655),
.Y(n_841)
);

OAI22xp33_ASAP7_75t_L g842 ( 
.A1(n_708),
.A2(n_417),
.B1(n_415),
.B2(n_302),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_693),
.B(n_558),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_695),
.B(n_558),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_680),
.B(n_518),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_800),
.A2(n_581),
.B1(n_520),
.B2(n_526),
.Y(n_846)
);

INVxp67_ASAP7_75t_L g847 ( 
.A(n_658),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_695),
.B(n_567),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_673),
.B(n_567),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_685),
.B(n_520),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_679),
.A2(n_531),
.B(n_526),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_L g852 ( 
.A1(n_754),
.A2(n_540),
.B(n_531),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_761),
.A2(n_551),
.B(n_540),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_676),
.B(n_705),
.Y(n_854)
);

BUFx12f_ASAP7_75t_L g855 ( 
.A(n_805),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_685),
.B(n_551),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_696),
.A2(n_557),
.B(n_554),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_669),
.A2(n_476),
.B1(n_579),
.B2(n_231),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_696),
.A2(n_557),
.B(n_554),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_711),
.B(n_579),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_L g861 ( 
.A1(n_678),
.A2(n_588),
.B1(n_561),
.B2(n_614),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_716),
.A2(n_562),
.B(n_561),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_768),
.A2(n_564),
.B(n_562),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_744),
.A2(n_580),
.B1(n_572),
.B2(n_564),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_724),
.B(n_545),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_771),
.A2(n_572),
.B(n_565),
.Y(n_866)
);

INVx11_ASAP7_75t_L g867 ( 
.A(n_694),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_783),
.B(n_565),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_711),
.B(n_476),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_772),
.A2(n_581),
.B(n_580),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_682),
.A2(n_588),
.B(n_582),
.Y(n_871)
);

NAND2x1p5_ASAP7_75t_L g872 ( 
.A(n_769),
.B(n_612),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_724),
.B(n_545),
.Y(n_873)
);

A2O1A1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_750),
.A2(n_594),
.B(n_595),
.C(n_592),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_662),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_692),
.B(n_476),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_793),
.B(n_582),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_703),
.B(n_589),
.Y(n_878)
);

INVx3_ASAP7_75t_L g879 ( 
.A(n_670),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_651),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_738),
.B(n_275),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_701),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_704),
.B(n_589),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_661),
.B(n_213),
.Y(n_884)
);

NOR2xp67_ASAP7_75t_L g885 ( 
.A(n_778),
.B(n_594),
.Y(n_885)
);

OAI21xp5_ASAP7_75t_L g886 ( 
.A1(n_716),
.A2(n_598),
.B(n_590),
.Y(n_886)
);

AND2x2_ASAP7_75t_SL g887 ( 
.A(n_669),
.B(n_240),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_723),
.A2(n_609),
.B(n_600),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_670),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_723),
.A2(n_609),
.B(n_600),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_712),
.B(n_595),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_719),
.B(n_604),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_789),
.A2(n_614),
.B(n_611),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_793),
.B(n_611),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_L g895 ( 
.A1(n_667),
.A2(n_743),
.B1(n_740),
.B2(n_739),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_663),
.B(n_604),
.Y(n_896)
);

NOR2xp67_ASAP7_75t_L g897 ( 
.A(n_728),
.B(n_607),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_657),
.B(n_613),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_668),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_657),
.A2(n_726),
.B(n_720),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_663),
.B(n_607),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_743),
.A2(n_613),
.B1(n_569),
.B2(n_329),
.Y(n_902)
);

NOR2xp67_ASAP7_75t_L g903 ( 
.A(n_731),
.B(n_612),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_657),
.A2(n_511),
.B(n_509),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_657),
.B(n_613),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_675),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_654),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_649),
.A2(n_653),
.B(n_741),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_731),
.B(n_757),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_750),
.B(n_613),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_654),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_759),
.B(n_509),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_681),
.A2(n_511),
.B(n_509),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_743),
.Y(n_914)
);

NOR2x1_ASAP7_75t_L g915 ( 
.A(n_709),
.B(n_511),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_683),
.B(n_215),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_688),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_759),
.B(n_767),
.Y(n_918)
);

INVx4_ASAP7_75t_L g919 ( 
.A(n_702),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_699),
.A2(n_706),
.B(n_700),
.Y(n_920)
);

O2A1O1Ixp5_ASAP7_75t_L g921 ( 
.A1(n_691),
.A2(n_303),
.B(n_208),
.C(n_314),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_702),
.B(n_623),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_767),
.B(n_745),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_687),
.B(n_762),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_710),
.B(n_713),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_769),
.Y(n_926)
);

A2O1A1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_666),
.A2(n_660),
.B(n_730),
.C(n_781),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_683),
.B(n_215),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_702),
.B(n_623),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_721),
.A2(n_514),
.B(n_612),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_L g931 ( 
.A1(n_667),
.A2(n_308),
.B1(n_305),
.B2(n_321),
.Y(n_931)
);

OAI21xp33_ASAP7_75t_L g932 ( 
.A1(n_797),
.A2(n_808),
.B(n_752),
.Y(n_932)
);

BUFx2_ASAP7_75t_L g933 ( 
.A(n_764),
.Y(n_933)
);

O2A1O1Ixp5_ASAP7_75t_L g934 ( 
.A1(n_756),
.A2(n_303),
.B(n_208),
.C(n_331),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_764),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_729),
.A2(n_504),
.B(n_623),
.Y(n_936)
);

AND2x4_ASAP7_75t_L g937 ( 
.A(n_774),
.B(n_569),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_790),
.A2(n_327),
.B1(n_612),
.B2(n_622),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_702),
.B(n_672),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_671),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_672),
.B(n_623),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_733),
.B(n_504),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_801),
.B(n_623),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_671),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_790),
.B(n_627),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_749),
.B(n_765),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_684),
.A2(n_627),
.B(n_622),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_734),
.B(n_627),
.Y(n_948)
);

NAND3xp33_ASAP7_75t_L g949 ( 
.A(n_737),
.B(n_622),
.C(n_323),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_766),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_686),
.B(n_627),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_686),
.B(n_225),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_760),
.B(n_225),
.Y(n_953)
);

AND2x2_ASAP7_75t_SL g954 ( 
.A(n_734),
.B(n_240),
.Y(n_954)
);

AOI22xp5_ASAP7_75t_L g955 ( 
.A1(n_686),
.A2(n_317),
.B1(n_323),
.B2(n_324),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_718),
.B(n_231),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_707),
.B(n_717),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_722),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_774),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_707),
.B(n_424),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_717),
.B(n_742),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_735),
.B(n_234),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_763),
.B(n_234),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_773),
.Y(n_964)
);

A2O1A1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_807),
.A2(n_249),
.B(n_274),
.C(n_285),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_748),
.A2(n_185),
.B(n_175),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_806),
.B(n_241),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_804),
.B(n_241),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_775),
.Y(n_969)
);

O2A1O1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_776),
.A2(n_803),
.B(n_802),
.C(n_799),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_784),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_791),
.B(n_248),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_792),
.A2(n_179),
.B(n_176),
.Y(n_973)
);

AOI22xp33_ASAP7_75t_L g974 ( 
.A1(n_795),
.A2(n_274),
.B1(n_248),
.B2(n_249),
.Y(n_974)
);

INVx4_ASAP7_75t_L g975 ( 
.A(n_689),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_697),
.A2(n_169),
.B(n_216),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_909),
.B(n_755),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_814),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_918),
.A2(n_798),
.B(n_794),
.Y(n_979)
);

CKINVDCx20_ASAP7_75t_R g980 ( 
.A(n_825),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_841),
.Y(n_981)
);

AOI22xp33_ASAP7_75t_L g982 ( 
.A1(n_954),
.A2(n_779),
.B1(n_770),
.B2(n_787),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_812),
.A2(n_787),
.B(n_725),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_818),
.A2(n_746),
.B(n_777),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_824),
.A2(n_786),
.B1(n_294),
.B2(n_290),
.Y(n_985)
);

O2A1O1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_819),
.A2(n_294),
.B(n_251),
.C(n_258),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_909),
.B(n_725),
.Y(n_987)
);

HB1xp67_ASAP7_75t_L g988 ( 
.A(n_847),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_935),
.Y(n_989)
);

NAND2xp33_ASAP7_75t_SL g990 ( 
.A(n_935),
.B(n_727),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_916),
.B(n_928),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_900),
.A2(n_777),
.B(n_770),
.Y(n_992)
);

NOR3xp33_ASAP7_75t_SL g993 ( 
.A(n_834),
.B(n_285),
.C(n_251),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_935),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_881),
.B(n_258),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_854),
.B(n_727),
.Y(n_996)
);

NOR3xp33_ASAP7_75t_L g997 ( 
.A(n_842),
.B(n_290),
.C(n_289),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_822),
.B(n_758),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_884),
.B(n_272),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_R g1000 ( 
.A(n_882),
.B(n_218),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_SL g1001 ( 
.A1(n_887),
.A2(n_273),
.B1(n_272),
.B2(n_331),
.Y(n_1001)
);

BUFx4f_ASAP7_75t_L g1002 ( 
.A(n_935),
.Y(n_1002)
);

AND2x2_ASAP7_75t_SL g1003 ( 
.A(n_954),
.B(n_240),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_SL g1004 ( 
.A(n_855),
.B(n_220),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_867),
.B(n_273),
.Y(n_1005)
);

BUFx3_ASAP7_75t_L g1006 ( 
.A(n_828),
.Y(n_1006)
);

NAND2x1_ASAP7_75t_L g1007 ( 
.A(n_879),
.B(n_424),
.Y(n_1007)
);

NOR2x1_ASAP7_75t_L g1008 ( 
.A(n_809),
.B(n_200),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_959),
.Y(n_1009)
);

AND2x4_ASAP7_75t_L g1010 ( 
.A(n_937),
.B(n_276),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_956),
.B(n_276),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_953),
.B(n_289),
.Y(n_1012)
);

BUFx3_ASAP7_75t_L g1013 ( 
.A(n_838),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_933),
.B(n_304),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_827),
.B(n_304),
.Y(n_1015)
);

BUFx2_ASAP7_75t_L g1016 ( 
.A(n_829),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_830),
.A2(n_255),
.B(n_203),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_833),
.A2(n_255),
.B(n_203),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_959),
.B(n_222),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_838),
.B(n_311),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_959),
.B(n_319),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_959),
.B(n_319),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_924),
.A2(n_209),
.B(n_217),
.C(n_243),
.Y(n_1023)
);

OAI22x1_ASAP7_75t_L g1024 ( 
.A1(n_955),
.A2(n_325),
.B1(n_209),
.B2(n_326),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_839),
.A2(n_209),
.B(n_325),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_937),
.Y(n_1026)
);

INVx4_ASAP7_75t_L g1027 ( 
.A(n_926),
.Y(n_1027)
);

AOI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_887),
.A2(n_280),
.B1(n_233),
.B2(n_236),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_L g1029 ( 
.A1(n_936),
.A2(n_426),
.B(n_424),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_875),
.Y(n_1030)
);

CKINVDCx8_ASAP7_75t_R g1031 ( 
.A(n_926),
.Y(n_1031)
);

BUFx3_ASAP7_75t_L g1032 ( 
.A(n_926),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_810),
.B(n_232),
.Y(n_1033)
);

O2A1O1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_927),
.A2(n_200),
.B(n_217),
.C(n_243),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_908),
.A2(n_426),
.B(n_424),
.Y(n_1035)
);

OR2x2_ASAP7_75t_L g1036 ( 
.A(n_931),
.B(n_424),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_811),
.A2(n_200),
.B(n_217),
.C(n_243),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_885),
.B(n_14),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_850),
.A2(n_193),
.B1(n_237),
.B2(n_244),
.Y(n_1039)
);

AO32x1_ASAP7_75t_L g1040 ( 
.A1(n_861),
.A2(n_424),
.A3(n_426),
.B1(n_20),
.B2(n_21),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_974),
.B(n_17),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_923),
.A2(n_17),
.B(n_19),
.C(n_20),
.Y(n_1042)
);

O2A1O1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_876),
.A2(n_19),
.B(n_21),
.C(n_22),
.Y(n_1043)
);

O2A1O1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_932),
.A2(n_23),
.B(n_24),
.C(n_25),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_850),
.B(n_23),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_SL g1046 ( 
.A1(n_856),
.A2(n_26),
.B(n_28),
.C(n_33),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_926),
.B(n_809),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_899),
.Y(n_1048)
);

NAND2xp33_ASAP7_75t_R g1049 ( 
.A(n_951),
.B(n_253),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_965),
.A2(n_35),
.B(n_37),
.C(n_39),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_831),
.A2(n_426),
.B(n_439),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_835),
.Y(n_1052)
);

BUFx3_ASAP7_75t_L g1053 ( 
.A(n_906),
.Y(n_1053)
);

BUFx12f_ASAP7_75t_L g1054 ( 
.A(n_919),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_831),
.A2(n_426),
.B(n_439),
.Y(n_1055)
);

AOI22xp33_ASAP7_75t_L g1056 ( 
.A1(n_952),
.A2(n_939),
.B1(n_858),
.B2(n_969),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_856),
.B(n_300),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_877),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_858),
.A2(n_265),
.B1(n_278),
.B2(n_282),
.Y(n_1059)
);

AOI21x1_ASAP7_75t_L g1060 ( 
.A1(n_840),
.A2(n_426),
.B(n_439),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_868),
.A2(n_310),
.B(n_322),
.C(n_320),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_845),
.B(n_35),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_974),
.B(n_40),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_817),
.A2(n_312),
.B(n_309),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_836),
.A2(n_439),
.B(n_297),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_868),
.A2(n_296),
.B(n_293),
.C(n_439),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_845),
.B(n_40),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_879),
.B(n_439),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_837),
.A2(n_439),
.B(n_43),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_878),
.A2(n_41),
.B(n_43),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_R g1071 ( 
.A(n_889),
.B(n_89),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_883),
.A2(n_41),
.B(n_46),
.Y(n_1072)
);

OAI22x1_ASAP7_75t_L g1073 ( 
.A1(n_915),
.A2(n_46),
.B1(n_47),
.B2(n_51),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_917),
.B(n_53),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_889),
.B(n_54),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_895),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_1076)
);

O2A1O1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_826),
.A2(n_57),
.B(n_63),
.C(n_66),
.Y(n_1077)
);

OAI22x1_ASAP7_75t_L g1078 ( 
.A1(n_877),
.A2(n_66),
.B1(n_67),
.B2(n_71),
.Y(n_1078)
);

HB1xp67_ASAP7_75t_L g1079 ( 
.A(n_894),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_910),
.A2(n_67),
.B1(n_73),
.B2(n_77),
.Y(n_1080)
);

OR2x6_ASAP7_75t_L g1081 ( 
.A(n_939),
.B(n_79),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_914),
.B(n_80),
.Y(n_1082)
);

AOI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_894),
.A2(n_91),
.B1(n_98),
.B2(n_105),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_914),
.B(n_115),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_950),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_846),
.A2(n_121),
.B1(n_123),
.B2(n_131),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_964),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_975),
.B(n_135),
.Y(n_1088)
);

AOI22xp33_ASAP7_75t_L g1089 ( 
.A1(n_971),
.A2(n_139),
.B1(n_146),
.B2(n_147),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_934),
.A2(n_152),
.B(n_153),
.C(n_154),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_967),
.B(n_166),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_968),
.B(n_869),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_871),
.A2(n_813),
.B(n_816),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_919),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_962),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_920),
.A2(n_925),
.B(n_852),
.C(n_832),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_975),
.B(n_957),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_815),
.A2(n_853),
.B(n_866),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_963),
.Y(n_1099)
);

NAND2xp33_ASAP7_75t_L g1100 ( 
.A(n_912),
.B(n_891),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_897),
.B(n_860),
.Y(n_1101)
);

AO22x1_ASAP7_75t_L g1102 ( 
.A1(n_946),
.A2(n_925),
.B1(n_972),
.B2(n_938),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_849),
.B(n_843),
.Y(n_1103)
);

NOR2xp67_ASAP7_75t_L g1104 ( 
.A(n_949),
.B(n_966),
.Y(n_1104)
);

NAND2xp33_ASAP7_75t_R g1105 ( 
.A(n_945),
.B(n_961),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_844),
.B(n_848),
.Y(n_1106)
);

O2A1O1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_892),
.A2(n_874),
.B(n_921),
.C(n_946),
.Y(n_1107)
);

BUFx4f_ASAP7_75t_L g1108 ( 
.A(n_872),
.Y(n_1108)
);

O2A1O1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_957),
.A2(n_893),
.B(n_970),
.C(n_896),
.Y(n_1109)
);

OR2x2_ASAP7_75t_L g1110 ( 
.A(n_901),
.B(n_907),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_SL g1111 ( 
.A(n_872),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_880),
.B(n_907),
.Y(n_1112)
);

O2A1O1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_862),
.A2(n_886),
.B(n_821),
.C(n_960),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_880),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_SL g1115 ( 
.A(n_903),
.B(n_911),
.Y(n_1115)
);

INVxp67_ASAP7_75t_L g1116 ( 
.A(n_940),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_944),
.Y(n_1117)
);

INVx4_ASAP7_75t_L g1118 ( 
.A(n_944),
.Y(n_1118)
);

OA22x2_ASAP7_75t_L g1119 ( 
.A1(n_864),
.A2(n_941),
.B1(n_948),
.B2(n_958),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_943),
.B(n_960),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_942),
.B(n_948),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1100),
.A2(n_823),
.B(n_873),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_991),
.B(n_973),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_1006),
.Y(n_1124)
);

BUFx3_ASAP7_75t_L g1125 ( 
.A(n_1016),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1003),
.A2(n_941),
.B1(n_942),
.B2(n_902),
.Y(n_1126)
);

AO31x2_ASAP7_75t_L g1127 ( 
.A1(n_1098),
.A2(n_913),
.A3(n_863),
.B(n_870),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_1035),
.A2(n_890),
.B(n_888),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_SL g1129 ( 
.A1(n_1081),
.A2(n_929),
.B(n_922),
.Y(n_1129)
);

AO31x2_ASAP7_75t_L g1130 ( 
.A1(n_1098),
.A2(n_947),
.A3(n_859),
.B(n_857),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_988),
.B(n_976),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_1044),
.A2(n_987),
.B(n_1034),
.C(n_997),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_1001),
.A2(n_851),
.B1(n_930),
.B2(n_820),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_1108),
.B(n_922),
.Y(n_1134)
);

INVx4_ASAP7_75t_L g1135 ( 
.A(n_1002),
.Y(n_1135)
);

OA21x2_ASAP7_75t_L g1136 ( 
.A1(n_1093),
.A2(n_865),
.B(n_873),
.Y(n_1136)
);

BUFx10_ASAP7_75t_L g1137 ( 
.A(n_1005),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_1000),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_999),
.B(n_898),
.Y(n_1139)
);

NOR2xp67_ASAP7_75t_L g1140 ( 
.A(n_1027),
.B(n_905),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1012),
.B(n_904),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1045),
.A2(n_1067),
.B1(n_1062),
.B2(n_1011),
.Y(n_1142)
);

AOI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1102),
.A2(n_1060),
.B(n_1025),
.Y(n_1143)
);

INVxp67_ASAP7_75t_SL g1144 ( 
.A(n_1053),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_995),
.B(n_1058),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_1079),
.B(n_998),
.Y(n_1146)
);

AO21x1_ASAP7_75t_L g1147 ( 
.A1(n_1076),
.A2(n_1034),
.B(n_1042),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_980),
.Y(n_1148)
);

AO32x2_ASAP7_75t_L g1149 ( 
.A1(n_1080),
.A2(n_985),
.A3(n_1118),
.B1(n_1039),
.B2(n_1086),
.Y(n_1149)
);

BUFx8_ASAP7_75t_L g1150 ( 
.A(n_1020),
.Y(n_1150)
);

O2A1O1Ixp5_ASAP7_75t_SL g1151 ( 
.A1(n_1075),
.A2(n_1038),
.B(n_1085),
.C(n_1087),
.Y(n_1151)
);

AOI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1041),
.A2(n_1063),
.B1(n_1022),
.B2(n_1024),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_977),
.B(n_1014),
.Y(n_1153)
);

AOI22xp33_ASAP7_75t_L g1154 ( 
.A1(n_1081),
.A2(n_1119),
.B1(n_1010),
.B2(n_1099),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1096),
.A2(n_1106),
.B(n_1103),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_1050),
.A2(n_1092),
.B(n_1042),
.C(n_1109),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_SL g1157 ( 
.A1(n_1109),
.A2(n_1113),
.B(n_1107),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1113),
.A2(n_1091),
.B(n_1107),
.Y(n_1158)
);

O2A1O1Ixp33_ASAP7_75t_SL g1159 ( 
.A1(n_1057),
.A2(n_1061),
.B(n_1084),
.C(n_1066),
.Y(n_1159)
);

O2A1O1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_1046),
.A2(n_1050),
.B(n_1043),
.C(n_1077),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_1026),
.Y(n_1161)
);

AOI22xp33_ASAP7_75t_L g1162 ( 
.A1(n_1081),
.A2(n_1119),
.B1(n_1010),
.B2(n_1095),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_992),
.A2(n_979),
.B(n_1055),
.Y(n_1163)
);

CKINVDCx11_ASAP7_75t_R g1164 ( 
.A(n_1054),
.Y(n_1164)
);

AOI221x1_ASAP7_75t_L g1165 ( 
.A1(n_1078),
.A2(n_1073),
.B1(n_1070),
.B2(n_1072),
.C(n_1023),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1021),
.B(n_993),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_1026),
.B(n_1013),
.Y(n_1167)
);

INVx4_ASAP7_75t_L g1168 ( 
.A(n_1002),
.Y(n_1168)
);

O2A1O1Ixp33_ASAP7_75t_SL g1169 ( 
.A1(n_1033),
.A2(n_1074),
.B(n_1007),
.C(n_1090),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_989),
.B(n_994),
.Y(n_1170)
);

BUFx2_ASAP7_75t_L g1171 ( 
.A(n_989),
.Y(n_1171)
);

BUFx10_ASAP7_75t_L g1172 ( 
.A(n_1082),
.Y(n_1172)
);

NAND2x1p5_ASAP7_75t_L g1173 ( 
.A(n_1108),
.B(n_989),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_SL g1174 ( 
.A(n_1031),
.B(n_1111),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_983),
.A2(n_984),
.B(n_1121),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_994),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_979),
.A2(n_1055),
.B(n_1051),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1051),
.A2(n_1025),
.B(n_983),
.Y(n_1178)
);

AOI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1056),
.A2(n_1015),
.B1(n_990),
.B2(n_1028),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1065),
.A2(n_984),
.B(n_1115),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1030),
.B(n_1048),
.Y(n_1181)
);

NAND2xp33_ASAP7_75t_L g1182 ( 
.A(n_1094),
.B(n_1071),
.Y(n_1182)
);

INVx1_ASAP7_75t_SL g1183 ( 
.A(n_994),
.Y(n_1183)
);

OA21x2_ASAP7_75t_L g1184 ( 
.A1(n_1017),
.A2(n_1018),
.B(n_1065),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1120),
.A2(n_1017),
.B(n_1018),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1104),
.A2(n_1036),
.B(n_1068),
.Y(n_1186)
);

AOI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1059),
.A2(n_1097),
.B1(n_1004),
.B2(n_996),
.Y(n_1187)
);

OAI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1083),
.A2(n_1072),
.B1(n_1070),
.B2(n_1049),
.Y(n_1188)
);

OAI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1037),
.A2(n_1069),
.B(n_982),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1088),
.A2(n_1040),
.B(n_1082),
.Y(n_1190)
);

AOI221xp5_ASAP7_75t_SL g1191 ( 
.A1(n_1043),
.A2(n_1077),
.B1(n_1064),
.B2(n_1019),
.C(n_1089),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1040),
.A2(n_1047),
.B(n_1101),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1040),
.A2(n_1118),
.B(n_1112),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1114),
.A2(n_1110),
.B(n_1116),
.Y(n_1194)
);

OAI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1009),
.A2(n_1105),
.B1(n_1027),
.B2(n_1094),
.Y(n_1195)
);

OR2x2_ASAP7_75t_L g1196 ( 
.A(n_1009),
.B(n_1117),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1009),
.B(n_1052),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1032),
.B(n_1008),
.Y(n_1198)
);

AND2x6_ASAP7_75t_L g1199 ( 
.A(n_1094),
.B(n_1114),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_991),
.B(n_909),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1100),
.A2(n_1096),
.B(n_1098),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_991),
.B(n_909),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_SL g1203 ( 
.A1(n_1081),
.A2(n_918),
.B(n_1088),
.Y(n_1203)
);

AOI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1003),
.A2(n_1001),
.B1(n_525),
.B2(n_954),
.Y(n_1204)
);

AO32x2_ASAP7_75t_L g1205 ( 
.A1(n_1076),
.A2(n_1001),
.A3(n_1080),
.B1(n_756),
.B2(n_985),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1096),
.A2(n_818),
.B(n_812),
.Y(n_1206)
);

INVx2_ASAP7_75t_SL g1207 ( 
.A(n_1013),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1100),
.A2(n_1096),
.B(n_1098),
.Y(n_1208)
);

HB1xp67_ASAP7_75t_L g1209 ( 
.A(n_988),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_978),
.Y(n_1210)
);

OAI22x1_ASAP7_75t_L g1211 ( 
.A1(n_1041),
.A2(n_955),
.B1(n_542),
.B2(n_800),
.Y(n_1211)
);

INVx2_ASAP7_75t_SL g1212 ( 
.A(n_1013),
.Y(n_1212)
);

INVx2_ASAP7_75t_SL g1213 ( 
.A(n_1013),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_988),
.B(n_515),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_981),
.Y(n_1215)
);

O2A1O1Ixp33_ASAP7_75t_SL g1216 ( 
.A1(n_1096),
.A2(n_824),
.B(n_1045),
.C(n_818),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_991),
.B(n_674),
.Y(n_1217)
);

AO32x2_ASAP7_75t_L g1218 ( 
.A1(n_1076),
.A2(n_1001),
.A3(n_1080),
.B1(n_756),
.B2(n_985),
.Y(n_1218)
);

INVxp67_ASAP7_75t_L g1219 ( 
.A(n_988),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_1031),
.Y(n_1220)
);

A2O1A1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1003),
.A2(n_819),
.B(n_909),
.C(n_665),
.Y(n_1221)
);

A2O1A1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1003),
.A2(n_819),
.B(n_909),
.C(n_665),
.Y(n_1222)
);

BUFx3_ASAP7_75t_L g1223 ( 
.A(n_1006),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1100),
.A2(n_1096),
.B(n_1098),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_991),
.B(n_909),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1026),
.B(n_1013),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_981),
.Y(n_1227)
);

NAND3x1_ASAP7_75t_L g1228 ( 
.A(n_1020),
.B(n_800),
.C(n_760),
.Y(n_1228)
);

BUFx4_ASAP7_75t_SL g1229 ( 
.A(n_980),
.Y(n_1229)
);

AO31x2_ASAP7_75t_L g1230 ( 
.A1(n_1098),
.A2(n_1093),
.A3(n_1096),
.B(n_1023),
.Y(n_1230)
);

CKINVDCx11_ASAP7_75t_R g1231 ( 
.A(n_980),
.Y(n_1231)
);

CKINVDCx11_ASAP7_75t_R g1232 ( 
.A(n_980),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1100),
.A2(n_1096),
.B(n_1098),
.Y(n_1233)
);

OAI22x1_ASAP7_75t_L g1234 ( 
.A1(n_1041),
.A2(n_955),
.B1(n_542),
.B2(n_800),
.Y(n_1234)
);

AO21x1_ASAP7_75t_L g1235 ( 
.A1(n_1044),
.A2(n_1076),
.B(n_986),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1100),
.A2(n_1096),
.B(n_1098),
.Y(n_1236)
);

BUFx2_ASAP7_75t_R g1237 ( 
.A(n_1013),
.Y(n_1237)
);

NAND3xp33_ASAP7_75t_SL g1238 ( 
.A(n_997),
.B(n_481),
.C(n_432),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_988),
.B(n_515),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_981),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_981),
.Y(n_1241)
);

BUFx8_ASAP7_75t_L g1242 ( 
.A(n_1016),
.Y(n_1242)
);

AOI221x1_ASAP7_75t_L g1243 ( 
.A1(n_1076),
.A2(n_1078),
.B1(n_819),
.B2(n_1024),
.C(n_1001),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1029),
.A2(n_1035),
.B(n_1093),
.Y(n_1244)
);

OAI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1096),
.A2(n_818),
.B(n_812),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_981),
.Y(n_1246)
);

BUFx3_ASAP7_75t_L g1247 ( 
.A(n_1006),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1026),
.B(n_1013),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_987),
.B(n_918),
.Y(n_1249)
);

AO32x2_ASAP7_75t_L g1250 ( 
.A1(n_1076),
.A2(n_1001),
.A3(n_1080),
.B1(n_756),
.B2(n_985),
.Y(n_1250)
);

AO31x2_ASAP7_75t_L g1251 ( 
.A1(n_1098),
.A2(n_1093),
.A3(n_1096),
.B(n_1023),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_981),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1029),
.A2(n_1035),
.B(n_1093),
.Y(n_1253)
);

OAI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1045),
.A2(n_525),
.B1(n_456),
.B2(n_484),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1029),
.A2(n_1035),
.B(n_1093),
.Y(n_1255)
);

AOI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1003),
.A2(n_1001),
.B1(n_525),
.B2(n_954),
.Y(n_1256)
);

OR2x6_ASAP7_75t_L g1257 ( 
.A(n_1013),
.B(n_1081),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_988),
.B(n_515),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_981),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1211),
.A2(n_1234),
.B1(n_1204),
.B2(n_1256),
.Y(n_1260)
);

INVx4_ASAP7_75t_L g1261 ( 
.A(n_1135),
.Y(n_1261)
);

AOI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1204),
.A2(n_1256),
.B1(n_1238),
.B2(n_1254),
.Y(n_1262)
);

BUFx12f_ASAP7_75t_L g1263 ( 
.A(n_1231),
.Y(n_1263)
);

BUFx2_ASAP7_75t_SL g1264 ( 
.A(n_1220),
.Y(n_1264)
);

BUFx4f_ASAP7_75t_SL g1265 ( 
.A(n_1242),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_1232),
.Y(n_1266)
);

AOI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1214),
.A2(n_1239),
.B1(n_1258),
.B2(n_1137),
.Y(n_1267)
);

CKINVDCx11_ASAP7_75t_R g1268 ( 
.A(n_1164),
.Y(n_1268)
);

NAND2x1p5_ASAP7_75t_L g1269 ( 
.A(n_1135),
.B(n_1168),
.Y(n_1269)
);

INVx1_ASAP7_75t_SL g1270 ( 
.A(n_1138),
.Y(n_1270)
);

AOI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1137),
.A2(n_1152),
.B1(n_1166),
.B2(n_1179),
.Y(n_1271)
);

INVx6_ASAP7_75t_L g1272 ( 
.A(n_1168),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_SL g1273 ( 
.A1(n_1257),
.A2(n_1148),
.B1(n_1152),
.B2(n_1225),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1235),
.A2(n_1142),
.B1(n_1217),
.B2(n_1257),
.Y(n_1274)
);

CKINVDCx20_ASAP7_75t_R g1275 ( 
.A(n_1150),
.Y(n_1275)
);

OAI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1243),
.A2(n_1179),
.B1(n_1200),
.B2(n_1202),
.Y(n_1276)
);

BUFx6f_ASAP7_75t_L g1277 ( 
.A(n_1172),
.Y(n_1277)
);

BUFx2_ASAP7_75t_L g1278 ( 
.A(n_1144),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1215),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1227),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1221),
.A2(n_1222),
.B1(n_1142),
.B2(n_1203),
.Y(n_1281)
);

CKINVDCx6p67_ASAP7_75t_R g1282 ( 
.A(n_1124),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1220),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_1229),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1210),
.Y(n_1285)
);

INVx1_ASAP7_75t_SL g1286 ( 
.A(n_1237),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1240),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1241),
.Y(n_1288)
);

BUFx2_ASAP7_75t_SL g1289 ( 
.A(n_1223),
.Y(n_1289)
);

INVx6_ASAP7_75t_L g1290 ( 
.A(n_1172),
.Y(n_1290)
);

CKINVDCx11_ASAP7_75t_R g1291 ( 
.A(n_1247),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1153),
.B(n_1249),
.Y(n_1292)
);

INVx6_ASAP7_75t_L g1293 ( 
.A(n_1242),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1246),
.Y(n_1294)
);

INVx3_ASAP7_75t_L g1295 ( 
.A(n_1173),
.Y(n_1295)
);

BUFx12f_ASAP7_75t_L g1296 ( 
.A(n_1150),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1257),
.A2(n_1147),
.B1(n_1162),
.B2(n_1154),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1145),
.A2(n_1188),
.B1(n_1126),
.B2(n_1123),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1126),
.A2(n_1157),
.B1(n_1139),
.B2(n_1190),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_1125),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1155),
.A2(n_1189),
.B1(n_1252),
.B2(n_1259),
.Y(n_1301)
);

OAI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1187),
.A2(n_1165),
.B1(n_1174),
.B2(n_1141),
.Y(n_1302)
);

INVx2_ASAP7_75t_SL g1303 ( 
.A(n_1207),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1189),
.A2(n_1158),
.B1(n_1133),
.B2(n_1187),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1209),
.B(n_1219),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1133),
.A2(n_1131),
.B1(n_1206),
.B2(n_1245),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1196),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1206),
.A2(n_1245),
.B1(n_1250),
.B2(n_1205),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1197),
.Y(n_1309)
);

OAI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1174),
.A2(n_1205),
.B1(n_1250),
.B2(n_1218),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1132),
.A2(n_1156),
.B1(n_1160),
.B2(n_1201),
.Y(n_1311)
);

INVxp67_ASAP7_75t_SL g1312 ( 
.A(n_1208),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1205),
.A2(n_1218),
.B1(n_1250),
.B2(n_1228),
.Y(n_1313)
);

AOI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1182),
.A2(n_1191),
.B1(n_1213),
.B2(n_1212),
.Y(n_1314)
);

HB1xp67_ASAP7_75t_L g1315 ( 
.A(n_1230),
.Y(n_1315)
);

CKINVDCx11_ASAP7_75t_R g1316 ( 
.A(n_1176),
.Y(n_1316)
);

CKINVDCx20_ASAP7_75t_R g1317 ( 
.A(n_1167),
.Y(n_1317)
);

INVx2_ASAP7_75t_SL g1318 ( 
.A(n_1226),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_SL g1319 ( 
.A1(n_1224),
.A2(n_1236),
.B(n_1233),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1171),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1161),
.B(n_1248),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1218),
.A2(n_1198),
.B1(n_1248),
.B2(n_1195),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1194),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1176),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1183),
.Y(n_1325)
);

BUFx4f_ASAP7_75t_SL g1326 ( 
.A(n_1161),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1183),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1173),
.Y(n_1328)
);

BUFx4_ASAP7_75t_R g1329 ( 
.A(n_1129),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1170),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1199),
.Y(n_1331)
);

BUFx6f_ASAP7_75t_L g1332 ( 
.A(n_1199),
.Y(n_1332)
);

BUFx12f_ASAP7_75t_L g1333 ( 
.A(n_1199),
.Y(n_1333)
);

BUFx12f_ASAP7_75t_L g1334 ( 
.A(n_1151),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1175),
.A2(n_1193),
.B1(n_1192),
.B2(n_1191),
.Y(n_1335)
);

NAND2x1p5_ASAP7_75t_L g1336 ( 
.A(n_1134),
.B(n_1140),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1180),
.A2(n_1185),
.B1(n_1184),
.B2(n_1186),
.Y(n_1337)
);

CKINVDCx20_ASAP7_75t_R g1338 ( 
.A(n_1184),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1216),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1149),
.B(n_1251),
.Y(n_1340)
);

INVx6_ASAP7_75t_L g1341 ( 
.A(n_1159),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_SL g1342 ( 
.A1(n_1122),
.A2(n_1149),
.B(n_1143),
.Y(n_1342)
);

INVx4_ASAP7_75t_SL g1343 ( 
.A(n_1251),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1136),
.B(n_1178),
.Y(n_1344)
);

BUFx10_ASAP7_75t_L g1345 ( 
.A(n_1149),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1136),
.B(n_1169),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1177),
.A2(n_1163),
.B1(n_1130),
.B2(n_1127),
.Y(n_1347)
);

BUFx3_ASAP7_75t_L g1348 ( 
.A(n_1128),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_SL g1349 ( 
.A1(n_1244),
.A2(n_1253),
.B(n_1255),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1181),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1200),
.B(n_1202),
.Y(n_1351)
);

CKINVDCx11_ASAP7_75t_R g1352 ( 
.A(n_1231),
.Y(n_1352)
);

BUFx2_ASAP7_75t_SL g1353 ( 
.A(n_1220),
.Y(n_1353)
);

INVx1_ASAP7_75t_SL g1354 ( 
.A(n_1138),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1181),
.Y(n_1355)
);

NAND2x1p5_ASAP7_75t_L g1356 ( 
.A(n_1135),
.B(n_1108),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1211),
.A2(n_1234),
.B1(n_1001),
.B2(n_1003),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1181),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1217),
.B(n_1146),
.Y(n_1359)
);

OAI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1204),
.A2(n_1256),
.B1(n_1152),
.B2(n_525),
.Y(n_1360)
);

INVx5_ASAP7_75t_L g1361 ( 
.A(n_1257),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1211),
.A2(n_1234),
.B1(n_1001),
.B2(n_1003),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_1144),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1204),
.A2(n_1256),
.B1(n_1003),
.B2(n_1222),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_1231),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1181),
.Y(n_1366)
);

AOI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1204),
.A2(n_1256),
.B1(n_525),
.B2(n_1001),
.Y(n_1367)
);

BUFx3_ASAP7_75t_L g1368 ( 
.A(n_1220),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_1229),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1181),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_SL g1371 ( 
.A1(n_1142),
.A2(n_1003),
.B1(n_954),
.B2(n_887),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_SL g1372 ( 
.A(n_1150),
.Y(n_1372)
);

BUFx10_ASAP7_75t_L g1373 ( 
.A(n_1148),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1181),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_SL g1375 ( 
.A1(n_1142),
.A2(n_1003),
.B1(n_954),
.B2(n_887),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1340),
.B(n_1345),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1345),
.B(n_1313),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_1284),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1278),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1350),
.B(n_1355),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1347),
.A2(n_1337),
.B(n_1344),
.Y(n_1381)
);

CKINVDCx6p67_ASAP7_75t_R g1382 ( 
.A(n_1296),
.Y(n_1382)
);

AOI21xp33_ASAP7_75t_L g1383 ( 
.A1(n_1360),
.A2(n_1281),
.B(n_1302),
.Y(n_1383)
);

AND2x4_ASAP7_75t_L g1384 ( 
.A(n_1361),
.B(n_1343),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_SL g1385 ( 
.A(n_1372),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1323),
.Y(n_1386)
);

INVx2_ASAP7_75t_SL g1387 ( 
.A(n_1363),
.Y(n_1387)
);

INVx2_ASAP7_75t_SL g1388 ( 
.A(n_1361),
.Y(n_1388)
);

AND2x4_ASAP7_75t_L g1389 ( 
.A(n_1361),
.B(n_1343),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1305),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1279),
.Y(n_1391)
);

OR2x2_ASAP7_75t_L g1392 ( 
.A(n_1313),
.B(n_1310),
.Y(n_1392)
);

OR2x2_ASAP7_75t_L g1393 ( 
.A(n_1310),
.B(n_1308),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1280),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1287),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1288),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1294),
.Y(n_1397)
);

INVx2_ASAP7_75t_SL g1398 ( 
.A(n_1361),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1320),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1325),
.Y(n_1400)
);

BUFx2_ASAP7_75t_L g1401 ( 
.A(n_1338),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1308),
.B(n_1306),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1315),
.Y(n_1403)
);

OAI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1367),
.A2(n_1262),
.B1(n_1364),
.B2(n_1271),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_SL g1405 ( 
.A(n_1369),
.B(n_1286),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1315),
.Y(n_1406)
);

INVx3_ASAP7_75t_L g1407 ( 
.A(n_1348),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1312),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1312),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1306),
.B(n_1304),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1346),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1327),
.Y(n_1412)
);

BUFx2_ASAP7_75t_L g1413 ( 
.A(n_1343),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1301),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1301),
.Y(n_1415)
);

AO21x2_ASAP7_75t_L g1416 ( 
.A1(n_1360),
.A2(n_1302),
.B(n_1342),
.Y(n_1416)
);

OA21x2_ASAP7_75t_L g1417 ( 
.A1(n_1319),
.A2(n_1337),
.B(n_1335),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1349),
.A2(n_1311),
.B(n_1335),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1309),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1339),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1358),
.Y(n_1421)
);

AOI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1304),
.A2(n_1375),
.B(n_1371),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1351),
.B(n_1270),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1299),
.B(n_1298),
.Y(n_1424)
);

INVxp67_ASAP7_75t_L g1425 ( 
.A(n_1359),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1366),
.Y(n_1426)
);

OA21x2_ASAP7_75t_L g1427 ( 
.A1(n_1299),
.A2(n_1298),
.B(n_1274),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1370),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1374),
.Y(n_1429)
);

INVx3_ASAP7_75t_L g1430 ( 
.A(n_1341),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1285),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1274),
.B(n_1260),
.Y(n_1432)
);

OR2x6_ASAP7_75t_L g1433 ( 
.A(n_1333),
.B(n_1332),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1307),
.Y(n_1434)
);

BUFx2_ASAP7_75t_L g1435 ( 
.A(n_1334),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1341),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1260),
.B(n_1330),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1331),
.A2(n_1336),
.B(n_1297),
.Y(n_1438)
);

INVx1_ASAP7_75t_SL g1439 ( 
.A(n_1317),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1324),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1322),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1322),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1276),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1292),
.B(n_1276),
.Y(n_1444)
);

INVx2_ASAP7_75t_SL g1445 ( 
.A(n_1290),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1336),
.A2(n_1297),
.B(n_1295),
.Y(n_1446)
);

INVxp33_ASAP7_75t_L g1447 ( 
.A(n_1291),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1273),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1329),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1329),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1314),
.Y(n_1451)
);

BUFx12f_ASAP7_75t_L g1452 ( 
.A(n_1268),
.Y(n_1452)
);

INVxp67_ASAP7_75t_L g1453 ( 
.A(n_1267),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1321),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1354),
.B(n_1300),
.Y(n_1455)
);

BUFx8_ASAP7_75t_L g1456 ( 
.A(n_1263),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1283),
.B(n_1368),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1283),
.B(n_1368),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1426),
.Y(n_1459)
);

AOI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1404),
.A2(n_1375),
.B1(n_1371),
.B2(n_1362),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1429),
.B(n_1264),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1401),
.B(n_1289),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1401),
.B(n_1303),
.Y(n_1463)
);

NOR2xp33_ASAP7_75t_L g1464 ( 
.A(n_1405),
.B(n_1282),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1379),
.B(n_1387),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1402),
.B(n_1353),
.Y(n_1466)
);

AOI221xp5_ASAP7_75t_L g1467 ( 
.A1(n_1422),
.A2(n_1357),
.B1(n_1362),
.B2(n_1275),
.C(n_1277),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1390),
.B(n_1387),
.Y(n_1468)
);

A2O1A1Ixp33_ASAP7_75t_L g1469 ( 
.A1(n_1383),
.A2(n_1357),
.B(n_1328),
.C(n_1318),
.Y(n_1469)
);

OAI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1410),
.A2(n_1356),
.B(n_1269),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1413),
.B(n_1384),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1402),
.B(n_1316),
.Y(n_1472)
);

NOR2x1_ASAP7_75t_SL g1473 ( 
.A(n_1449),
.B(n_1261),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1376),
.B(n_1293),
.Y(n_1474)
);

O2A1O1Ixp33_ASAP7_75t_L g1475 ( 
.A1(n_1410),
.A2(n_1356),
.B(n_1266),
.C(n_1365),
.Y(n_1475)
);

NOR2x1_ASAP7_75t_L g1476 ( 
.A(n_1457),
.B(n_1265),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_SL g1477 ( 
.A(n_1430),
.B(n_1326),
.Y(n_1477)
);

O2A1O1Ixp33_ASAP7_75t_L g1478 ( 
.A1(n_1453),
.A2(n_1326),
.B(n_1265),
.C(n_1272),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1411),
.B(n_1290),
.Y(n_1479)
);

INVxp67_ASAP7_75t_L g1480 ( 
.A(n_1411),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1425),
.B(n_1293),
.Y(n_1481)
);

AND2x4_ASAP7_75t_L g1482 ( 
.A(n_1413),
.B(n_1293),
.Y(n_1482)
);

INVxp67_ASAP7_75t_L g1483 ( 
.A(n_1400),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1439),
.B(n_1352),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1399),
.B(n_1373),
.Y(n_1485)
);

A2O1A1Ixp33_ASAP7_75t_L g1486 ( 
.A1(n_1432),
.A2(n_1272),
.B(n_1373),
.C(n_1443),
.Y(n_1486)
);

NAND4xp25_ASAP7_75t_L g1487 ( 
.A(n_1435),
.B(n_1444),
.C(n_1424),
.D(n_1432),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_SL g1488 ( 
.A1(n_1424),
.A2(n_1427),
.B1(n_1416),
.B2(n_1393),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1414),
.B(n_1415),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1447),
.B(n_1378),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1414),
.B(n_1415),
.Y(n_1491)
);

INVx5_ASAP7_75t_SL g1492 ( 
.A(n_1382),
.Y(n_1492)
);

OAI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1427),
.A2(n_1451),
.B(n_1418),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_SL g1494 ( 
.A1(n_1458),
.A2(n_1445),
.B(n_1450),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1386),
.B(n_1421),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1391),
.B(n_1412),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1423),
.B(n_1377),
.Y(n_1497)
);

O2A1O1Ixp33_ASAP7_75t_L g1498 ( 
.A1(n_1451),
.A2(n_1416),
.B(n_1427),
.C(n_1448),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1386),
.B(n_1421),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1384),
.B(n_1389),
.Y(n_1500)
);

AOI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1416),
.A2(n_1448),
.B1(n_1427),
.B2(n_1437),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1428),
.B(n_1408),
.Y(n_1502)
);

BUFx3_ASAP7_75t_L g1503 ( 
.A(n_1456),
.Y(n_1503)
);

OR2x6_ASAP7_75t_L g1504 ( 
.A(n_1449),
.B(n_1450),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1428),
.B(n_1408),
.Y(n_1505)
);

CKINVDCx20_ASAP7_75t_R g1506 ( 
.A(n_1456),
.Y(n_1506)
);

OAI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1392),
.A2(n_1393),
.B1(n_1441),
.B2(n_1442),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1394),
.B(n_1395),
.Y(n_1508)
);

AO32x2_ASAP7_75t_L g1509 ( 
.A1(n_1388),
.A2(n_1398),
.A3(n_1445),
.B1(n_1392),
.B2(n_1434),
.Y(n_1509)
);

NOR2x1_ASAP7_75t_SL g1510 ( 
.A(n_1433),
.B(n_1436),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1440),
.Y(n_1511)
);

OAI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1418),
.A2(n_1417),
.B(n_1420),
.Y(n_1512)
);

A2O1A1Ixp33_ASAP7_75t_L g1513 ( 
.A1(n_1441),
.A2(n_1442),
.B(n_1446),
.C(n_1438),
.Y(n_1513)
);

AND2x4_ASAP7_75t_L g1514 ( 
.A(n_1500),
.B(n_1407),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1502),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1500),
.B(n_1407),
.Y(n_1516)
);

INVx2_ASAP7_75t_SL g1517 ( 
.A(n_1468),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1496),
.B(n_1403),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1512),
.B(n_1417),
.Y(n_1519)
);

INVx1_ASAP7_75t_SL g1520 ( 
.A(n_1465),
.Y(n_1520)
);

BUFx3_ASAP7_75t_L g1521 ( 
.A(n_1494),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1480),
.B(n_1409),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1483),
.B(n_1459),
.Y(n_1523)
);

INVxp67_ASAP7_75t_SL g1524 ( 
.A(n_1480),
.Y(n_1524)
);

NOR2x1_ASAP7_75t_L g1525 ( 
.A(n_1461),
.B(n_1479),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1512),
.B(n_1417),
.Y(n_1526)
);

INVx2_ASAP7_75t_SL g1527 ( 
.A(n_1482),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1502),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1509),
.B(n_1417),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1505),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1460),
.A2(n_1430),
.B1(n_1420),
.B2(n_1436),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1505),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1509),
.B(n_1381),
.Y(n_1533)
);

OAI221xp5_ASAP7_75t_SL g1534 ( 
.A1(n_1467),
.A2(n_1409),
.B1(n_1382),
.B2(n_1435),
.C(n_1430),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_SL g1535 ( 
.A1(n_1507),
.A2(n_1452),
.B1(n_1430),
.B2(n_1446),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1509),
.B(n_1381),
.Y(n_1536)
);

BUFx2_ASAP7_75t_L g1537 ( 
.A(n_1509),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1488),
.A2(n_1454),
.B1(n_1438),
.B2(n_1431),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1483),
.B(n_1396),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1508),
.B(n_1397),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1511),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1464),
.B(n_1452),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1495),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1495),
.Y(n_1544)
);

INVxp67_ASAP7_75t_L g1545 ( 
.A(n_1466),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1499),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1499),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1489),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1521),
.Y(n_1549)
);

HB1xp67_ASAP7_75t_L g1550 ( 
.A(n_1541),
.Y(n_1550)
);

AOI221xp5_ASAP7_75t_L g1551 ( 
.A1(n_1537),
.A2(n_1498),
.B1(n_1467),
.B2(n_1487),
.C(n_1501),
.Y(n_1551)
);

NOR2xp33_ASAP7_75t_L g1552 ( 
.A(n_1521),
.B(n_1472),
.Y(n_1552)
);

NAND2x1_ASAP7_75t_L g1553 ( 
.A(n_1525),
.B(n_1462),
.Y(n_1553)
);

OAI221xp5_ASAP7_75t_L g1554 ( 
.A1(n_1537),
.A2(n_1488),
.B1(n_1498),
.B2(n_1493),
.C(n_1469),
.Y(n_1554)
);

INVx5_ASAP7_75t_L g1555 ( 
.A(n_1529),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1541),
.Y(n_1556)
);

OAI21xp5_ASAP7_75t_SL g1557 ( 
.A1(n_1529),
.A2(n_1475),
.B(n_1478),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1520),
.B(n_1497),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_SL g1559 ( 
.A(n_1529),
.B(n_1466),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1520),
.B(n_1474),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1521),
.B(n_1471),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1545),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1546),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1522),
.Y(n_1564)
);

BUFx2_ASAP7_75t_L g1565 ( 
.A(n_1527),
.Y(n_1565)
);

NAND3xp33_ASAP7_75t_L g1566 ( 
.A(n_1525),
.B(n_1493),
.C(n_1479),
.Y(n_1566)
);

INVxp67_ASAP7_75t_SL g1567 ( 
.A(n_1524),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1522),
.Y(n_1568)
);

AOI221xp5_ASAP7_75t_L g1569 ( 
.A1(n_1519),
.A2(n_1507),
.B1(n_1475),
.B2(n_1489),
.C(n_1491),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1524),
.B(n_1461),
.Y(n_1570)
);

OAI322xp33_ASAP7_75t_L g1571 ( 
.A1(n_1531),
.A2(n_1472),
.A3(n_1491),
.B1(n_1463),
.B2(n_1440),
.C1(n_1380),
.C2(n_1434),
.Y(n_1571)
);

OAI221xp5_ASAP7_75t_L g1572 ( 
.A1(n_1534),
.A2(n_1486),
.B1(n_1470),
.B2(n_1513),
.C(n_1419),
.Y(n_1572)
);

AOI21xp5_ASAP7_75t_L g1573 ( 
.A1(n_1534),
.A2(n_1478),
.B(n_1470),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1517),
.B(n_1485),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1546),
.Y(n_1575)
);

OAI211xp5_ASAP7_75t_SL g1576 ( 
.A1(n_1523),
.A2(n_1476),
.B(n_1455),
.C(n_1484),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1514),
.B(n_1516),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1518),
.B(n_1523),
.Y(n_1578)
);

INVxp67_ASAP7_75t_L g1579 ( 
.A(n_1539),
.Y(n_1579)
);

INVx2_ASAP7_75t_SL g1580 ( 
.A(n_1518),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1546),
.B(n_1403),
.Y(n_1581)
);

INVx3_ASAP7_75t_L g1582 ( 
.A(n_1514),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1543),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1548),
.B(n_1406),
.Y(n_1584)
);

AOI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1531),
.A2(n_1473),
.B(n_1510),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1539),
.B(n_1481),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1543),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1533),
.B(n_1504),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1540),
.B(n_1406),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1544),
.Y(n_1590)
);

OAI21xp33_ASAP7_75t_L g1591 ( 
.A1(n_1551),
.A2(n_1526),
.B(n_1519),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1555),
.B(n_1533),
.Y(n_1592)
);

INVx1_ASAP7_75t_SL g1593 ( 
.A(n_1553),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1555),
.B(n_1582),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1564),
.B(n_1515),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1579),
.B(n_1515),
.Y(n_1596)
);

BUFx2_ASAP7_75t_L g1597 ( 
.A(n_1555),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1581),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1568),
.B(n_1528),
.Y(n_1599)
);

BUFx3_ASAP7_75t_L g1600 ( 
.A(n_1549),
.Y(n_1600)
);

INVxp67_ASAP7_75t_L g1601 ( 
.A(n_1550),
.Y(n_1601)
);

AND2x4_ASAP7_75t_L g1602 ( 
.A(n_1577),
.B(n_1533),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1581),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1555),
.B(n_1536),
.Y(n_1604)
);

NAND2x1p5_ASAP7_75t_L g1605 ( 
.A(n_1555),
.B(n_1536),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1582),
.B(n_1536),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1583),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1563),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1582),
.B(n_1519),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_SL g1610 ( 
.A(n_1585),
.B(n_1527),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1587),
.Y(n_1611)
);

HB1xp67_ASAP7_75t_L g1612 ( 
.A(n_1562),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_SL g1613 ( 
.A(n_1561),
.B(n_1527),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1577),
.B(n_1526),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1556),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1577),
.B(n_1526),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1565),
.B(n_1528),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1590),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1563),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1567),
.B(n_1530),
.Y(n_1620)
);

HB1xp67_ASAP7_75t_L g1621 ( 
.A(n_1584),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1580),
.B(n_1530),
.Y(n_1622)
);

AND2x6_ASAP7_75t_SL g1623 ( 
.A(n_1552),
.B(n_1542),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1549),
.B(n_1514),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1578),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1578),
.B(n_1532),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1559),
.B(n_1532),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1575),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1614),
.B(n_1549),
.Y(n_1629)
);

INVx2_ASAP7_75t_SL g1630 ( 
.A(n_1600),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1607),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1607),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1607),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1611),
.Y(n_1634)
);

NOR2x1_ASAP7_75t_L g1635 ( 
.A(n_1597),
.B(n_1506),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1625),
.B(n_1580),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1614),
.B(n_1561),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1625),
.B(n_1589),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1621),
.B(n_1544),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1612),
.B(n_1569),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1605),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1605),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1614),
.B(n_1561),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1616),
.B(n_1552),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1621),
.B(n_1591),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1611),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1616),
.B(n_1574),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1615),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1591),
.B(n_1620),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1611),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1591),
.B(n_1547),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1618),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1618),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1618),
.Y(n_1654)
);

NAND2x1p5_ASAP7_75t_L g1655 ( 
.A(n_1597),
.B(n_1482),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1616),
.B(n_1574),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1605),
.B(n_1602),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1605),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1620),
.B(n_1547),
.Y(n_1659)
);

AOI32xp33_ASAP7_75t_L g1660 ( 
.A1(n_1592),
.A2(n_1554),
.A3(n_1576),
.B1(n_1559),
.B2(n_1572),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1625),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1599),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1605),
.B(n_1560),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1602),
.B(n_1560),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1620),
.B(n_1558),
.Y(n_1665)
);

AOI21xp33_ASAP7_75t_L g1666 ( 
.A1(n_1612),
.A2(n_1557),
.B(n_1566),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1615),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1626),
.B(n_1570),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1599),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1602),
.B(n_1592),
.Y(n_1670)
);

OAI31xp33_ASAP7_75t_L g1671 ( 
.A1(n_1592),
.A2(n_1573),
.A3(n_1588),
.B(n_1538),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1644),
.B(n_1593),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1635),
.B(n_1597),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1631),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1644),
.B(n_1593),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1647),
.B(n_1602),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1647),
.B(n_1602),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1640),
.B(n_1601),
.Y(n_1678)
);

OAI21xp33_ASAP7_75t_L g1679 ( 
.A1(n_1649),
.A2(n_1604),
.B(n_1610),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1670),
.Y(n_1680)
);

INVx2_ASAP7_75t_SL g1681 ( 
.A(n_1635),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1631),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1632),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1656),
.B(n_1602),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1660),
.B(n_1601),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1632),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1660),
.B(n_1627),
.Y(n_1687)
);

NAND4xp75_ASAP7_75t_L g1688 ( 
.A(n_1671),
.B(n_1649),
.C(n_1666),
.D(n_1645),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1648),
.B(n_1667),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1638),
.B(n_1626),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1638),
.B(n_1626),
.Y(n_1691)
);

O2A1O1Ixp33_ASAP7_75t_L g1692 ( 
.A1(n_1666),
.A2(n_1610),
.B(n_1604),
.C(n_1571),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1645),
.B(n_1596),
.Y(n_1693)
);

AOI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1671),
.A2(n_1613),
.B(n_1596),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1656),
.B(n_1604),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1651),
.B(n_1598),
.Y(n_1696)
);

INVxp67_ASAP7_75t_L g1697 ( 
.A(n_1630),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1637),
.B(n_1624),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1637),
.B(n_1624),
.Y(n_1699)
);

NAND2xp33_ASAP7_75t_SL g1700 ( 
.A(n_1657),
.B(n_1594),
.Y(n_1700)
);

OAI21xp33_ASAP7_75t_L g1701 ( 
.A1(n_1651),
.A2(n_1609),
.B(n_1606),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1633),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1665),
.B(n_1662),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1633),
.Y(n_1704)
);

AND2x4_ASAP7_75t_L g1705 ( 
.A(n_1643),
.B(n_1600),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1670),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1634),
.Y(n_1707)
);

INVxp67_ASAP7_75t_SL g1708 ( 
.A(n_1685),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1674),
.Y(n_1709)
);

A2O1A1Ixp33_ASAP7_75t_L g1710 ( 
.A1(n_1687),
.A2(n_1657),
.B(n_1658),
.C(n_1641),
.Y(n_1710)
);

AOI32xp33_ASAP7_75t_L g1711 ( 
.A1(n_1678),
.A2(n_1642),
.A3(n_1641),
.B1(n_1658),
.B2(n_1663),
.Y(n_1711)
);

AOI222xp33_ASAP7_75t_L g1712 ( 
.A1(n_1679),
.A2(n_1688),
.B1(n_1701),
.B2(n_1681),
.C1(n_1703),
.C2(n_1689),
.Y(n_1712)
);

NAND3xp33_ASAP7_75t_L g1713 ( 
.A(n_1692),
.B(n_1661),
.C(n_1630),
.Y(n_1713)
);

NOR3xp33_ASAP7_75t_L g1714 ( 
.A(n_1688),
.B(n_1642),
.C(n_1641),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1680),
.Y(n_1715)
);

INVxp67_ASAP7_75t_L g1716 ( 
.A(n_1681),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1674),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1690),
.B(n_1665),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1697),
.B(n_1662),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1690),
.B(n_1669),
.Y(n_1720)
);

NAND3x2_ASAP7_75t_L g1721 ( 
.A(n_1693),
.B(n_1663),
.C(n_1629),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1680),
.Y(n_1722)
);

AO22x1_ASAP7_75t_L g1723 ( 
.A1(n_1673),
.A2(n_1456),
.B1(n_1600),
.B2(n_1503),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1691),
.B(n_1669),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1691),
.B(n_1661),
.Y(n_1725)
);

HAxp5_ASAP7_75t_SL g1726 ( 
.A(n_1694),
.B(n_1456),
.CON(n_1726),
.SN(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1706),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1672),
.B(n_1643),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1672),
.B(n_1675),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_SL g1730 ( 
.A(n_1673),
.B(n_1655),
.Y(n_1730)
);

A2O1A1Ixp33_ASAP7_75t_L g1731 ( 
.A1(n_1693),
.A2(n_1658),
.B(n_1642),
.C(n_1623),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1682),
.Y(n_1732)
);

AOI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1675),
.A2(n_1535),
.B1(n_1664),
.B2(n_1629),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1715),
.Y(n_1734)
);

NOR2xp67_ASAP7_75t_L g1735 ( 
.A(n_1729),
.B(n_1706),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1715),
.Y(n_1736)
);

XNOR2xp5_ASAP7_75t_L g1737 ( 
.A(n_1729),
.B(n_1385),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1728),
.B(n_1705),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1728),
.B(n_1705),
.Y(n_1739)
);

NAND3xp33_ASAP7_75t_L g1740 ( 
.A(n_1712),
.B(n_1673),
.C(n_1704),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1722),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1716),
.B(n_1705),
.Y(n_1742)
);

NOR2x1_ASAP7_75t_L g1743 ( 
.A(n_1713),
.B(n_1682),
.Y(n_1743)
);

AOI33xp33_ASAP7_75t_L g1744 ( 
.A1(n_1709),
.A2(n_1707),
.A3(n_1702),
.B1(n_1683),
.B2(n_1686),
.B3(n_1695),
.Y(n_1744)
);

AOI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1708),
.A2(n_1684),
.B1(n_1676),
.B2(n_1677),
.Y(n_1745)
);

OAI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1731),
.A2(n_1655),
.B1(n_1684),
.B2(n_1677),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_SL g1747 ( 
.A(n_1731),
.B(n_1700),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1722),
.B(n_1676),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1727),
.Y(n_1749)
);

NOR2x1_ASAP7_75t_L g1750 ( 
.A(n_1730),
.B(n_1683),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1727),
.B(n_1695),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1717),
.Y(n_1752)
);

OAI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1710),
.A2(n_1702),
.B(n_1686),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_SL g1754 ( 
.A(n_1737),
.B(n_1714),
.Y(n_1754)
);

AOI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1740),
.A2(n_1733),
.B1(n_1710),
.B2(n_1721),
.Y(n_1755)
);

OAI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1747),
.A2(n_1718),
.B1(n_1726),
.B2(n_1730),
.Y(n_1756)
);

INVxp67_ASAP7_75t_L g1757 ( 
.A(n_1742),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1749),
.Y(n_1758)
);

O2A1O1Ixp33_ASAP7_75t_L g1759 ( 
.A1(n_1747),
.A2(n_1743),
.B(n_1750),
.C(n_1753),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1735),
.B(n_1720),
.Y(n_1760)
);

A2O1A1Ixp33_ASAP7_75t_SL g1761 ( 
.A1(n_1746),
.A2(n_1711),
.B(n_1732),
.C(n_1719),
.Y(n_1761)
);

O2A1O1Ixp33_ASAP7_75t_L g1762 ( 
.A1(n_1734),
.A2(n_1741),
.B(n_1736),
.C(n_1749),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1748),
.B(n_1724),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1738),
.B(n_1623),
.Y(n_1764)
);

AOI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1748),
.A2(n_1725),
.B1(n_1723),
.B2(n_1726),
.Y(n_1765)
);

AOI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1759),
.A2(n_1751),
.B(n_1742),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1757),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1758),
.Y(n_1768)
);

NAND2xp33_ASAP7_75t_SL g1769 ( 
.A(n_1763),
.B(n_1738),
.Y(n_1769)
);

NOR3xp33_ASAP7_75t_L g1770 ( 
.A(n_1754),
.B(n_1752),
.C(n_1744),
.Y(n_1770)
);

NOR2xp33_ASAP7_75t_L g1771 ( 
.A(n_1764),
.B(n_1739),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1760),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1755),
.B(n_1739),
.Y(n_1773)
);

NAND4xp25_ASAP7_75t_L g1774 ( 
.A(n_1761),
.B(n_1745),
.C(n_1744),
.D(n_1698),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1756),
.B(n_1664),
.Y(n_1775)
);

AOI322xp5_ASAP7_75t_L g1776 ( 
.A1(n_1770),
.A2(n_1765),
.A3(n_1762),
.B1(n_1707),
.B2(n_1659),
.C1(n_1606),
.C2(n_1646),
.Y(n_1776)
);

AOI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1766),
.A2(n_1696),
.B(n_1634),
.Y(n_1777)
);

O2A1O1Ixp33_ASAP7_75t_L g1778 ( 
.A1(n_1774),
.A2(n_1696),
.B(n_1646),
.C(n_1650),
.Y(n_1778)
);

AOI221xp5_ASAP7_75t_L g1779 ( 
.A1(n_1773),
.A2(n_1652),
.B1(n_1653),
.B2(n_1654),
.C(n_1650),
.Y(n_1779)
);

AOI322xp5_ASAP7_75t_L g1780 ( 
.A1(n_1772),
.A2(n_1659),
.A3(n_1606),
.B1(n_1652),
.B2(n_1654),
.C1(n_1653),
.C2(n_1609),
.Y(n_1780)
);

OAI211xp5_ASAP7_75t_SL g1781 ( 
.A1(n_1775),
.A2(n_1613),
.B(n_1636),
.C(n_1668),
.Y(n_1781)
);

AOI221xp5_ASAP7_75t_L g1782 ( 
.A1(n_1778),
.A2(n_1768),
.B1(n_1769),
.B2(n_1771),
.C(n_1767),
.Y(n_1782)
);

AOI221xp5_ASAP7_75t_SL g1783 ( 
.A1(n_1777),
.A2(n_1699),
.B1(n_1698),
.B2(n_1594),
.C(n_1490),
.Y(n_1783)
);

A2O1A1Ixp33_ASAP7_75t_L g1784 ( 
.A1(n_1776),
.A2(n_1600),
.B(n_1699),
.C(n_1594),
.Y(n_1784)
);

O2A1O1Ixp33_ASAP7_75t_L g1785 ( 
.A1(n_1781),
.A2(n_1655),
.B(n_1668),
.C(n_1639),
.Y(n_1785)
);

NOR3xp33_ASAP7_75t_L g1786 ( 
.A(n_1779),
.B(n_1639),
.C(n_1636),
.Y(n_1786)
);

AOI211xp5_ASAP7_75t_L g1787 ( 
.A1(n_1780),
.A2(n_1492),
.B(n_1609),
.C(n_1627),
.Y(n_1787)
);

OAI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1778),
.A2(n_1622),
.B1(n_1603),
.B2(n_1598),
.Y(n_1788)
);

AND2x2_ASAP7_75t_SL g1789 ( 
.A(n_1782),
.B(n_1492),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1784),
.A2(n_1492),
.B1(n_1598),
.B2(n_1603),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1786),
.B(n_1624),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1788),
.Y(n_1792)
);

NAND4xp75_ASAP7_75t_L g1793 ( 
.A(n_1783),
.B(n_1627),
.C(n_1623),
.D(n_1603),
.Y(n_1793)
);

AND2x4_ASAP7_75t_L g1794 ( 
.A(n_1791),
.B(n_1624),
.Y(n_1794)
);

INVx2_ASAP7_75t_SL g1795 ( 
.A(n_1789),
.Y(n_1795)
);

NAND3xp33_ASAP7_75t_SL g1796 ( 
.A(n_1792),
.B(n_1785),
.C(n_1787),
.Y(n_1796)
);

XNOR2xp5_ASAP7_75t_L g1797 ( 
.A(n_1796),
.B(n_1793),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1797),
.Y(n_1798)
);

INVx4_ASAP7_75t_L g1799 ( 
.A(n_1798),
.Y(n_1799)
);

INVx3_ASAP7_75t_SL g1800 ( 
.A(n_1798),
.Y(n_1800)
);

OAI22xp5_ASAP7_75t_L g1801 ( 
.A1(n_1800),
.A2(n_1795),
.B1(n_1790),
.B2(n_1794),
.Y(n_1801)
);

OAI22x1_ASAP7_75t_L g1802 ( 
.A1(n_1799),
.A2(n_1791),
.B1(n_1624),
.B2(n_1617),
.Y(n_1802)
);

AOI21xp5_ASAP7_75t_L g1803 ( 
.A1(n_1801),
.A2(n_1622),
.B(n_1595),
.Y(n_1803)
);

AOI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1803),
.A2(n_1802),
.B(n_1595),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1804),
.B(n_1608),
.Y(n_1805)
);

XNOR2xp5_ASAP7_75t_L g1806 ( 
.A(n_1805),
.B(n_1433),
.Y(n_1806)
);

AOI221xp5_ASAP7_75t_L g1807 ( 
.A1(n_1806),
.A2(n_1628),
.B1(n_1608),
.B2(n_1619),
.C(n_1586),
.Y(n_1807)
);

AOI211xp5_ASAP7_75t_L g1808 ( 
.A1(n_1807),
.A2(n_1477),
.B(n_1617),
.C(n_1586),
.Y(n_1808)
);


endmodule