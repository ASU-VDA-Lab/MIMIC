module fake_netlist_5_505_n_1488 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_1488);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1488;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_150;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_709;
wire n_317;
wire n_1236;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_297;
wire n_156;
wire n_1078;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1284;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_184;
wire n_446;
wire n_1064;
wire n_144;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1233;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_1468;
wire n_689;
wire n_738;
wire n_640;
wire n_252;
wire n_624;
wire n_1380;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_456;
wire n_959;
wire n_535;
wire n_152;
wire n_940;
wire n_1445;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_256;
wire n_950;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_146;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_153;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1470;
wire n_1096;
wire n_234;
wire n_833;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1419;
wire n_338;
wire n_149;
wire n_693;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_151;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1335;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_754;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_791;
wire n_732;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_148;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_147;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_733;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_145;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_499;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_236;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1220;
wire n_229;
wire n_437;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_246;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_64),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_55),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_88),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_4),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_78),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_97),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_51),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_92),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_94),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_123),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_103),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_89),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_107),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_108),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_98),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_18),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_71),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_63),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_13),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_57),
.Y(n_165)
);

BUFx10_ASAP7_75t_L g166 ( 
.A(n_42),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_134),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_20),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_122),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_102),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_53),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_26),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_5),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_101),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_132),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_74),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_32),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_128),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_24),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_45),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_22),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_110),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_14),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_49),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_139),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_19),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_19),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_129),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_113),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_44),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_99),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_116),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_66),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_4),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_10),
.Y(n_195)
);

BUFx10_ASAP7_75t_L g196 ( 
.A(n_12),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_11),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_75),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_67),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_38),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_82),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_105),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_69),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_77),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_93),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_83),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_76),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_16),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_28),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_137),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_25),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_39),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_125),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_68),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_80),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_136),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_81),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_34),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_7),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_141),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_42),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_73),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_117),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_54),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_40),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_38),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_65),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_124),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_115),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_100),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_35),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_16),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_29),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_135),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_26),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_70),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_138),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_31),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_37),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_3),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_17),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_46),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_133),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_44),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_22),
.Y(n_245)
);

BUFx10_ASAP7_75t_L g246 ( 
.A(n_131),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_3),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_119),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_111),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_18),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_118),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_84),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_41),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_120),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_29),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_11),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_34),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_5),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_2),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_61),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_28),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_95),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_121),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_30),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_79),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_36),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_59),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_142),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_62),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_96),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_47),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_90),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_112),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_33),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_23),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_2),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_60),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_114),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_12),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_17),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_6),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_58),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_31),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_126),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_21),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_85),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_10),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_143),
.Y(n_288)
);

BUFx10_ASAP7_75t_L g289 ( 
.A(n_20),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_146),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_240),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_240),
.Y(n_292)
);

NOR2xp67_ASAP7_75t_L g293 ( 
.A(n_186),
.B(n_0),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_240),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_155),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_240),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_240),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_149),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_255),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_201),
.B(n_271),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_255),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_255),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_151),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_255),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_153),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_149),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_255),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_154),
.Y(n_308)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_222),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_216),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_201),
.B(n_0),
.Y(n_311)
);

INVxp33_ASAP7_75t_SL g312 ( 
.A(n_160),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_156),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_175),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_162),
.B(n_1),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_216),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_228),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_228),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_176),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_183),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_204),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_183),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_218),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_178),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_182),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_184),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_188),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_193),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_218),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_221),
.Y(n_330)
);

NOR2xp67_ASAP7_75t_L g331 ( 
.A(n_186),
.B(n_1),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_221),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_198),
.Y(n_333)
);

INVxp33_ASAP7_75t_SL g334 ( 
.A(n_160),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_164),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_172),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_204),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_202),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_203),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_251),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_148),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_226),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_205),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_251),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_173),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_232),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_206),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_207),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_263),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_210),
.Y(n_350)
);

NOR2xp67_ASAP7_75t_L g351 ( 
.A(n_200),
.B(n_6),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_190),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_194),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_215),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_233),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_263),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_217),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_166),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_286),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_165),
.B(n_174),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_168),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_223),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_227),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_286),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_290),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_292),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_303),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_305),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_308),
.Y(n_369)
);

INVx5_ASAP7_75t_L g370 ( 
.A(n_309),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_341),
.B(n_269),
.Y(n_371)
);

OA21x2_ASAP7_75t_L g372 ( 
.A1(n_360),
.A2(n_174),
.B(n_165),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_337),
.B(n_144),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_309),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_298),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_313),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_292),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_314),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_294),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_309),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_294),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_361),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_296),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_319),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_324),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_300),
.B(n_325),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_296),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_309),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_306),
.Y(n_389)
);

NAND2xp33_ASAP7_75t_R g390 ( 
.A(n_312),
.B(n_144),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_291),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_326),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_301),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_327),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_342),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_297),
.B(n_145),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_297),
.B(n_145),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_299),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_328),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_333),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_299),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_302),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_338),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_339),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_295),
.B(n_246),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_310),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_302),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_304),
.B(n_242),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_304),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_307),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_343),
.Y(n_411)
);

NOR2xp67_ASAP7_75t_L g412 ( 
.A(n_307),
.B(n_150),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_316),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_322),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_322),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_320),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_347),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_348),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_321),
.B(n_157),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_321),
.B(n_200),
.Y(n_420)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_295),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_311),
.B(n_242),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_354),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_320),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_335),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_357),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_335),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_362),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_323),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_336),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_336),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_386),
.B(n_363),
.Y(n_432)
);

OR2x2_ASAP7_75t_L g433 ( 
.A(n_371),
.B(n_350),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_371),
.B(n_350),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_380),
.Y(n_435)
);

INVx5_ASAP7_75t_L g436 ( 
.A(n_380),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_390),
.A2(n_334),
.B1(n_288),
.B2(n_315),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_420),
.B(n_323),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_425),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_L g440 ( 
.A1(n_422),
.A2(n_346),
.B1(n_293),
.B2(n_331),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_373),
.B(n_358),
.Y(n_441)
);

OAI21xp33_ASAP7_75t_SL g442 ( 
.A1(n_420),
.A2(n_331),
.B(n_293),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_373),
.B(n_317),
.Y(n_443)
);

BUFx10_ASAP7_75t_L g444 ( 
.A(n_365),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_422),
.B(n_260),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_422),
.B(n_230),
.Y(n_446)
);

OAI22xp33_ASAP7_75t_L g447 ( 
.A1(n_395),
.A2(n_187),
.B1(n_225),
.B2(n_285),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_419),
.B(n_260),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_395),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_427),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_393),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_396),
.B(n_222),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_393),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_430),
.B(n_345),
.Y(n_454)
);

NAND2xp33_ASAP7_75t_SL g455 ( 
.A(n_405),
.B(n_288),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_391),
.Y(n_456)
);

INVx2_ASAP7_75t_SL g457 ( 
.A(n_382),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_430),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_431),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_431),
.B(n_329),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_366),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_396),
.B(n_234),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_375),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_L g464 ( 
.A1(n_372),
.A2(n_351),
.B1(n_266),
.B2(n_280),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_397),
.B(n_237),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_389),
.Y(n_466)
);

INVx2_ASAP7_75t_SL g467 ( 
.A(n_397),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_377),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_377),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_374),
.B(n_248),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_372),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_367),
.B(n_222),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_368),
.B(n_318),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_406),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_408),
.B(n_345),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_379),
.Y(n_476)
);

INVx1_ASAP7_75t_SL g477 ( 
.A(n_413),
.Y(n_477)
);

NAND2xp33_ASAP7_75t_L g478 ( 
.A(n_391),
.B(n_222),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_421),
.Y(n_479)
);

AND3x2_ASAP7_75t_L g480 ( 
.A(n_385),
.B(n_400),
.C(n_399),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_369),
.B(n_340),
.Y(n_481)
);

INVx5_ASAP7_75t_L g482 ( 
.A(n_391),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_374),
.Y(n_483)
);

AND2x2_ASAP7_75t_SL g484 ( 
.A(n_421),
.B(n_222),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_379),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_381),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_L g487 ( 
.A1(n_372),
.A2(n_351),
.B1(n_266),
.B2(n_258),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_376),
.B(n_344),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_381),
.Y(n_489)
);

INVx5_ASAP7_75t_L g490 ( 
.A(n_374),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_374),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_383),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_383),
.B(n_252),
.Y(n_493)
);

INVx5_ASAP7_75t_L g494 ( 
.A(n_402),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_378),
.Y(n_495)
);

INVx1_ASAP7_75t_SL g496 ( 
.A(n_384),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_387),
.Y(n_497)
);

OR2x2_ASAP7_75t_SL g498 ( 
.A(n_418),
.B(n_257),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_392),
.B(n_349),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_394),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_403),
.B(n_356),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_398),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_404),
.B(n_352),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_372),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_429),
.B(n_330),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_401),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_L g507 ( 
.A1(n_408),
.A2(n_259),
.B1(n_279),
.B2(n_287),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_411),
.B(n_359),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_429),
.B(n_330),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_401),
.B(n_262),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_429),
.B(n_332),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_408),
.B(n_352),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_415),
.Y(n_513)
);

AND2x6_ASAP7_75t_L g514 ( 
.A(n_408),
.B(n_152),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_407),
.Y(n_515)
);

BUFx8_ASAP7_75t_SL g516 ( 
.A(n_417),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_409),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_423),
.B(n_159),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_426),
.A2(n_212),
.B1(n_211),
.B2(n_209),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_410),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g521 ( 
.A(n_429),
.B(n_353),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_412),
.B(n_353),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_428),
.Y(n_523)
);

OAI22xp33_ASAP7_75t_L g524 ( 
.A1(n_424),
.A2(n_195),
.B1(n_219),
.B2(n_197),
.Y(n_524)
);

AND2x2_ASAP7_75t_SL g525 ( 
.A(n_416),
.B(n_163),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_402),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g527 ( 
.A(n_412),
.B(n_147),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_402),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_416),
.B(n_170),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_L g530 ( 
.A1(n_416),
.A2(n_261),
.B1(n_264),
.B2(n_275),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_402),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_388),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_414),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_424),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_414),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_424),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_414),
.B(n_364),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_414),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_370),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_370),
.Y(n_540)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_370),
.Y(n_541)
);

INVxp33_ASAP7_75t_SL g542 ( 
.A(n_370),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_380),
.Y(n_543)
);

CKINVDCx16_ASAP7_75t_R g544 ( 
.A(n_421),
.Y(n_544)
);

BUFx10_ASAP7_75t_L g545 ( 
.A(n_386),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_390),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_420),
.B(n_332),
.Y(n_547)
);

BUFx4f_ASAP7_75t_L g548 ( 
.A(n_422),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_420),
.B(n_355),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_SL g550 ( 
.A(n_365),
.B(n_147),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_515),
.Y(n_551)
);

NAND2xp33_ASAP7_75t_L g552 ( 
.A(n_467),
.B(n_267),
.Y(n_552)
);

AOI221xp5_ASAP7_75t_L g553 ( 
.A1(n_447),
.A2(n_208),
.B1(n_181),
.B2(n_283),
.C(n_281),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_432),
.B(n_180),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_441),
.B(n_185),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_434),
.B(n_157),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_548),
.B(n_189),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_433),
.B(n_158),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_538),
.B(n_191),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_548),
.B(n_192),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_443),
.A2(n_268),
.B1(n_270),
.B2(n_272),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_462),
.B(n_465),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_515),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_484),
.B(n_199),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_520),
.B(n_213),
.Y(n_565)
);

BUFx6f_ASAP7_75t_SL g566 ( 
.A(n_444),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_503),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_484),
.B(n_214),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_464),
.B(n_220),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_549),
.B(n_166),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_R g571 ( 
.A(n_546),
.B(n_158),
.Y(n_571)
);

NAND2xp33_ASAP7_75t_L g572 ( 
.A(n_514),
.B(n_273),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_487),
.B(n_224),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_439),
.B(n_229),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_483),
.Y(n_575)
);

INVx8_ASAP7_75t_L g576 ( 
.A(n_516),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_527),
.B(n_236),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_517),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_549),
.B(n_166),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_450),
.B(n_243),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_445),
.A2(n_208),
.B1(n_181),
.B2(n_254),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_460),
.Y(n_582)
);

A2O1A1Ixp33_ASAP7_75t_L g583 ( 
.A1(n_442),
.A2(n_355),
.B(n_282),
.C(n_249),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_438),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_L g585 ( 
.A1(n_470),
.A2(n_265),
.B(n_284),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_458),
.B(n_161),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_SL g587 ( 
.A(n_516),
.B(n_246),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_460),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_459),
.B(n_161),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_483),
.Y(n_590)
);

OR2x2_ASAP7_75t_L g591 ( 
.A(n_449),
.B(n_168),
.Y(n_591)
);

NAND3xp33_ASAP7_75t_L g592 ( 
.A(n_440),
.B(n_245),
.C(n_177),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_545),
.B(n_167),
.Y(n_593)
);

O2A1O1Ixp33_ASAP7_75t_L g594 ( 
.A1(n_448),
.A2(n_169),
.B(n_284),
.C(n_171),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_457),
.B(n_283),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_455),
.A2(n_169),
.B1(n_171),
.B2(n_278),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_545),
.B(n_277),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_461),
.B(n_277),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_444),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_468),
.B(n_179),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_SL g601 ( 
.A(n_496),
.B(n_246),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_491),
.B(n_247),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_495),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_491),
.B(n_244),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_469),
.B(n_231),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_525),
.A2(n_276),
.B1(n_281),
.B2(n_289),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_476),
.B(n_235),
.Y(n_607)
);

AND3x1_ASAP7_75t_L g608 ( 
.A(n_437),
.B(n_289),
.C(n_196),
.Y(n_608)
);

NOR3xp33_ASAP7_75t_L g609 ( 
.A(n_455),
.B(n_537),
.C(n_519),
.Y(n_609)
);

OR2x2_ASAP7_75t_L g610 ( 
.A(n_457),
.B(n_276),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_485),
.B(n_238),
.Y(n_611)
);

BUFx6f_ASAP7_75t_SL g612 ( 
.A(n_444),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_446),
.A2(n_471),
.B1(n_504),
.B2(n_546),
.Y(n_613)
);

NOR2x1p5_ASAP7_75t_L g614 ( 
.A(n_438),
.B(n_250),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_517),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_491),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_518),
.A2(n_274),
.B1(n_256),
.B2(n_253),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_486),
.B(n_239),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_489),
.B(n_241),
.Y(n_619)
);

OAI221xp5_ASAP7_75t_L g620 ( 
.A1(n_530),
.A2(n_289),
.B1(n_196),
.B2(n_9),
.C(n_13),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_492),
.B(n_497),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_521),
.Y(n_622)
);

OAI21xp33_ASAP7_75t_L g623 ( 
.A1(n_547),
.A2(n_196),
.B(n_8),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_502),
.B(n_506),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_545),
.B(n_518),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_525),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_521),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_505),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_472),
.B(n_14),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_505),
.Y(n_630)
);

NAND2xp33_ASAP7_75t_L g631 ( 
.A(n_514),
.B(n_130),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_509),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_531),
.B(n_526),
.Y(n_633)
);

AO221x1_ASAP7_75t_L g634 ( 
.A1(n_524),
.A2(n_15),
.B1(n_21),
.B2(n_23),
.C(n_24),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_509),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_L g636 ( 
.A1(n_471),
.A2(n_127),
.B(n_106),
.Y(n_636)
);

NAND2xp33_ASAP7_75t_L g637 ( 
.A(n_514),
.B(n_104),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_533),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_547),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_534),
.B(n_91),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_531),
.B(n_87),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_550),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_528),
.B(n_86),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_490),
.B(n_72),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_536),
.B(n_56),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_504),
.A2(n_52),
.B1(n_50),
.B2(n_48),
.Y(n_646)
);

INVx1_ASAP7_75t_SL g647 ( 
.A(n_466),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_490),
.B(n_15),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_511),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_454),
.Y(n_650)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_479),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_500),
.B(n_25),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_533),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_472),
.B(n_27),
.Y(n_654)
);

O2A1O1Ixp5_ASAP7_75t_L g655 ( 
.A1(n_448),
.A2(n_27),
.B(n_30),
.C(n_32),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_454),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_493),
.B(n_33),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_490),
.B(n_35),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_510),
.B(n_498),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_536),
.B(n_36),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_490),
.B(n_37),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_490),
.B(n_39),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_454),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_475),
.B(n_40),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_475),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_475),
.B(n_41),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_512),
.Y(n_667)
);

OR2x6_ASAP7_75t_L g668 ( 
.A(n_463),
.B(n_43),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_512),
.B(n_43),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_452),
.B(n_522),
.Y(n_670)
);

AOI22xp5_ASAP7_75t_L g671 ( 
.A1(n_514),
.A2(n_522),
.B1(n_529),
.B2(n_544),
.Y(n_671)
);

AND3x1_ASAP7_75t_L g672 ( 
.A(n_473),
.B(n_508),
.C(n_499),
.Y(n_672)
);

AOI21xp5_ASAP7_75t_L g673 ( 
.A1(n_542),
.A2(n_541),
.B(n_539),
.Y(n_673)
);

OAI22xp5_ASAP7_75t_SL g674 ( 
.A1(n_477),
.A2(n_474),
.B1(n_488),
.B2(n_501),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_535),
.Y(n_675)
);

OAI22xp5_ASAP7_75t_L g676 ( 
.A1(n_562),
.A2(n_523),
.B1(n_507),
.B2(n_481),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_551),
.Y(n_677)
);

A2O1A1Ixp33_ASAP7_75t_L g678 ( 
.A1(n_556),
.A2(n_529),
.B(n_456),
.C(n_513),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_638),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_638),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_622),
.B(n_514),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_627),
.B(n_435),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_638),
.Y(n_683)
);

BUFx4f_ASAP7_75t_L g684 ( 
.A(n_576),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_551),
.Y(n_685)
);

A2O1A1Ixp33_ASAP7_75t_L g686 ( 
.A1(n_657),
.A2(n_540),
.B(n_451),
.C(n_453),
.Y(n_686)
);

NOR2x1_ASAP7_75t_R g687 ( 
.A(n_599),
.B(n_480),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_628),
.B(n_435),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_563),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_563),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_625),
.B(n_435),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_630),
.B(n_543),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_570),
.B(n_532),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_632),
.B(n_635),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_649),
.B(n_543),
.Y(n_695)
);

INVxp67_ASAP7_75t_L g696 ( 
.A(n_567),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_578),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_615),
.Y(n_698)
);

OAI21xp5_ASAP7_75t_L g699 ( 
.A1(n_569),
.A2(n_478),
.B(n_494),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_566),
.Y(n_700)
);

CKINVDCx8_ASAP7_75t_R g701 ( 
.A(n_576),
.Y(n_701)
);

OAI21xp5_ASAP7_75t_L g702 ( 
.A1(n_583),
.A2(n_494),
.B(n_436),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_593),
.B(n_494),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_615),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_R g705 ( 
.A(n_603),
.B(n_566),
.Y(n_705)
);

INVx2_ASAP7_75t_SL g706 ( 
.A(n_603),
.Y(n_706)
);

O2A1O1Ixp33_ASAP7_75t_L g707 ( 
.A1(n_664),
.A2(n_564),
.B(n_568),
.C(n_654),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_593),
.B(n_436),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_590),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_591),
.B(n_482),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_597),
.B(n_482),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_579),
.B(n_482),
.Y(n_712)
);

OAI22xp5_ASAP7_75t_L g713 ( 
.A1(n_581),
.A2(n_656),
.B1(n_663),
.B2(n_650),
.Y(n_713)
);

NOR2xp67_ASAP7_75t_L g714 ( 
.A(n_651),
.B(n_597),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_582),
.B(n_588),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_L g716 ( 
.A1(n_581),
.A2(n_626),
.B1(n_573),
.B2(n_659),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_L g717 ( 
.A1(n_626),
.A2(n_665),
.B1(n_667),
.B2(n_575),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_558),
.B(n_595),
.Y(n_718)
);

OAI21xp33_ASAP7_75t_L g719 ( 
.A1(n_606),
.A2(n_617),
.B(n_553),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_558),
.B(n_610),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_621),
.B(n_624),
.Y(n_721)
);

OAI21xp33_ASAP7_75t_L g722 ( 
.A1(n_606),
.A2(n_601),
.B(n_571),
.Y(n_722)
);

A2O1A1Ixp33_ASAP7_75t_L g723 ( 
.A1(n_657),
.A2(n_654),
.B(n_629),
.C(n_577),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_560),
.A2(n_633),
.B(n_673),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_671),
.B(n_666),
.Y(n_725)
);

HB1xp67_ASAP7_75t_L g726 ( 
.A(n_666),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_642),
.B(n_647),
.Y(n_727)
);

O2A1O1Ixp33_ASAP7_75t_L g728 ( 
.A1(n_664),
.A2(n_564),
.B(n_568),
.C(n_629),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_669),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_636),
.A2(n_631),
.B(n_637),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_616),
.A2(n_572),
.B(n_602),
.Y(n_731)
);

AOI21xp5_ASAP7_75t_L g732 ( 
.A1(n_602),
.A2(n_604),
.B(n_559),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_604),
.A2(n_640),
.B(n_645),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_571),
.B(n_652),
.Y(n_734)
);

AO21x1_ASAP7_75t_L g735 ( 
.A1(n_646),
.A2(n_577),
.B(n_643),
.Y(n_735)
);

A2O1A1Ixp33_ASAP7_75t_L g736 ( 
.A1(n_583),
.A2(n_594),
.B(n_623),
.C(n_675),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_614),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_552),
.A2(n_565),
.B1(n_600),
.B2(n_605),
.Y(n_738)
);

INVx4_ASAP7_75t_L g739 ( 
.A(n_638),
.Y(n_739)
);

O2A1O1Ixp33_ASAP7_75t_L g740 ( 
.A1(n_648),
.A2(n_662),
.B(n_661),
.C(n_658),
.Y(n_740)
);

O2A1O1Ixp33_ASAP7_75t_L g741 ( 
.A1(n_648),
.A2(n_662),
.B(n_661),
.C(n_658),
.Y(n_741)
);

NOR2x1_ASAP7_75t_L g742 ( 
.A(n_592),
.B(n_644),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_574),
.B(n_580),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_596),
.B(n_674),
.Y(n_744)
);

A2O1A1Ixp33_ASAP7_75t_L g745 ( 
.A1(n_655),
.A2(n_611),
.B(n_618),
.C(n_619),
.Y(n_745)
);

NAND2x1p5_ASAP7_75t_L g746 ( 
.A(n_653),
.B(n_644),
.Y(n_746)
);

A2O1A1Ixp33_ASAP7_75t_L g747 ( 
.A1(n_607),
.A2(n_561),
.B(n_598),
.C(n_589),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_653),
.Y(n_748)
);

BUFx12f_ASAP7_75t_L g749 ( 
.A(n_668),
.Y(n_749)
);

INVx3_ASAP7_75t_L g750 ( 
.A(n_660),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_668),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_586),
.A2(n_672),
.B1(n_585),
.B2(n_643),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_641),
.Y(n_753)
);

AOI22xp5_ASAP7_75t_L g754 ( 
.A1(n_608),
.A2(n_641),
.B1(n_634),
.B2(n_620),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_668),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_587),
.B(n_576),
.Y(n_756)
);

BUFx4f_ASAP7_75t_L g757 ( 
.A(n_612),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_612),
.A2(n_548),
.B(n_670),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_638),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_562),
.B(n_467),
.Y(n_760)
);

INVx4_ASAP7_75t_L g761 ( 
.A(n_638),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_562),
.B(n_467),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_562),
.B(n_467),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_670),
.A2(n_548),
.B(n_504),
.Y(n_764)
);

O2A1O1Ixp5_ASAP7_75t_L g765 ( 
.A1(n_557),
.A2(n_560),
.B(n_554),
.C(n_555),
.Y(n_765)
);

OAI21xp5_ASAP7_75t_L g766 ( 
.A1(n_613),
.A2(n_504),
.B(n_471),
.Y(n_766)
);

A2O1A1Ixp33_ASAP7_75t_L g767 ( 
.A1(n_556),
.A2(n_562),
.B(n_657),
.C(n_554),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_659),
.A2(n_562),
.B1(n_609),
.B2(n_467),
.Y(n_768)
);

AND2x6_ASAP7_75t_L g769 ( 
.A(n_562),
.B(n_629),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_562),
.B(n_467),
.Y(n_770)
);

NAND2x1p5_ASAP7_75t_L g771 ( 
.A(n_638),
.B(n_548),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_562),
.B(n_467),
.Y(n_772)
);

INVx3_ASAP7_75t_L g773 ( 
.A(n_638),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_562),
.B(n_467),
.Y(n_774)
);

OAI21xp5_ASAP7_75t_L g775 ( 
.A1(n_613),
.A2(n_504),
.B(n_471),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_625),
.B(n_546),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_625),
.B(n_484),
.Y(n_777)
);

NOR2x1p5_ASAP7_75t_SL g778 ( 
.A(n_590),
.B(n_616),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_659),
.A2(n_562),
.B1(n_609),
.B2(n_467),
.Y(n_779)
);

A2O1A1Ixp33_ASAP7_75t_L g780 ( 
.A1(n_556),
.A2(n_562),
.B(n_657),
.C(n_554),
.Y(n_780)
);

A2O1A1Ixp33_ASAP7_75t_L g781 ( 
.A1(n_556),
.A2(n_562),
.B(n_657),
.C(n_554),
.Y(n_781)
);

OAI21xp5_ASAP7_75t_L g782 ( 
.A1(n_613),
.A2(n_504),
.B(n_471),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_562),
.B(n_467),
.Y(n_783)
);

AO21x1_ASAP7_75t_L g784 ( 
.A1(n_636),
.A2(n_613),
.B(n_629),
.Y(n_784)
);

AOI33xp33_ASAP7_75t_L g785 ( 
.A1(n_581),
.A2(n_447),
.A3(n_553),
.B1(n_606),
.B2(n_626),
.B3(n_457),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_562),
.B(n_467),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_625),
.B(n_546),
.Y(n_787)
);

AND2x6_ASAP7_75t_L g788 ( 
.A(n_562),
.B(n_629),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_613),
.A2(n_504),
.B(n_471),
.Y(n_789)
);

A2O1A1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_556),
.A2(n_562),
.B(n_657),
.C(n_554),
.Y(n_790)
);

OAI21xp5_ASAP7_75t_L g791 ( 
.A1(n_613),
.A2(n_504),
.B(n_471),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_551),
.Y(n_792)
);

BUFx4f_ASAP7_75t_SL g793 ( 
.A(n_603),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_562),
.B(n_467),
.Y(n_794)
);

INVx1_ASAP7_75t_SL g795 ( 
.A(n_647),
.Y(n_795)
);

NAND2x1p5_ASAP7_75t_L g796 ( 
.A(n_638),
.B(n_548),
.Y(n_796)
);

NOR2xp67_ASAP7_75t_L g797 ( 
.A(n_599),
.B(n_500),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_584),
.B(n_639),
.Y(n_798)
);

BUFx2_ASAP7_75t_L g799 ( 
.A(n_603),
.Y(n_799)
);

NAND2x1p5_ASAP7_75t_L g800 ( 
.A(n_638),
.B(n_548),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_562),
.B(n_467),
.Y(n_801)
);

OAI21xp5_ASAP7_75t_L g802 ( 
.A1(n_613),
.A2(n_504),
.B(n_471),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_562),
.B(n_467),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_562),
.B(n_467),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_638),
.Y(n_805)
);

OA22x2_ASAP7_75t_L g806 ( 
.A1(n_634),
.A2(n_623),
.B1(n_639),
.B2(n_584),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_705),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_793),
.Y(n_808)
);

O2A1O1Ixp5_ASAP7_75t_L g809 ( 
.A1(n_784),
.A2(n_780),
.B(n_790),
.C(n_781),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_760),
.B(n_762),
.Y(n_810)
);

AO21x2_ASAP7_75t_L g811 ( 
.A1(n_766),
.A2(n_782),
.B(n_775),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_676),
.B(n_763),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_770),
.B(n_772),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_774),
.B(n_783),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_786),
.B(n_794),
.Y(n_815)
);

INVxp67_ASAP7_75t_SL g816 ( 
.A(n_683),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_801),
.B(n_803),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_804),
.B(n_721),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_685),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_677),
.Y(n_820)
);

AND2x2_ASAP7_75t_SL g821 ( 
.A(n_785),
.B(n_744),
.Y(n_821)
);

OAI22x1_ASAP7_75t_L g822 ( 
.A1(n_776),
.A2(n_787),
.B1(n_754),
.B2(n_779),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_722),
.B(n_795),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_769),
.B(n_788),
.Y(n_824)
);

BUFx2_ASAP7_75t_L g825 ( 
.A(n_795),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_718),
.B(n_720),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_768),
.B(n_769),
.Y(n_827)
);

OAI21xp33_ASAP7_75t_SL g828 ( 
.A1(n_725),
.A2(n_777),
.B(n_753),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_769),
.B(n_788),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_683),
.Y(n_830)
);

NAND3xp33_ASAP7_75t_L g831 ( 
.A(n_719),
.B(n_716),
.C(n_707),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_766),
.A2(n_775),
.B(n_789),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_769),
.B(n_788),
.Y(n_833)
);

A2O1A1Ixp33_ASAP7_75t_L g834 ( 
.A1(n_728),
.A2(n_740),
.B(n_741),
.C(n_765),
.Y(n_834)
);

O2A1O1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_734),
.A2(n_736),
.B(n_729),
.C(n_747),
.Y(n_835)
);

OA21x2_ASAP7_75t_L g836 ( 
.A1(n_782),
.A2(n_791),
.B(n_789),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_788),
.B(n_693),
.Y(n_837)
);

BUFx2_ASAP7_75t_L g838 ( 
.A(n_799),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_727),
.B(n_696),
.Y(n_839)
);

AO31x2_ASAP7_75t_L g840 ( 
.A1(n_745),
.A2(n_678),
.A3(n_717),
.B(n_724),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_743),
.B(n_694),
.Y(n_841)
);

NAND2x1_ASAP7_75t_L g842 ( 
.A(n_739),
.B(n_761),
.Y(n_842)
);

AOI21x1_ASAP7_75t_L g843 ( 
.A1(n_731),
.A2(n_732),
.B(n_733),
.Y(n_843)
);

OA22x2_ASAP7_75t_L g844 ( 
.A1(n_755),
.A2(n_751),
.B1(n_798),
.B2(n_706),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_726),
.B(n_798),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_714),
.B(n_715),
.Y(n_846)
);

OAI21x1_ASAP7_75t_SL g847 ( 
.A1(n_758),
.A2(n_702),
.B(n_681),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_689),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_802),
.A2(n_712),
.B(n_691),
.Y(n_849)
);

BUFx4_ASAP7_75t_SL g850 ( 
.A(n_700),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_690),
.Y(n_851)
);

BUFx2_ASAP7_75t_L g852 ( 
.A(n_749),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_750),
.B(n_738),
.Y(n_853)
);

AND2x6_ASAP7_75t_L g854 ( 
.A(n_742),
.B(n_752),
.Y(n_854)
);

INVx1_ASAP7_75t_SL g855 ( 
.A(n_710),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_L g856 ( 
.A1(n_806),
.A2(n_713),
.B1(n_746),
.B2(n_750),
.Y(n_856)
);

INVx4_ASAP7_75t_L g857 ( 
.A(n_683),
.Y(n_857)
);

BUFx2_ASAP7_75t_L g858 ( 
.A(n_806),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_701),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_682),
.B(n_703),
.Y(n_860)
);

AO31x2_ASAP7_75t_L g861 ( 
.A1(n_711),
.A2(n_708),
.A3(n_792),
.B(n_698),
.Y(n_861)
);

INVx4_ASAP7_75t_L g862 ( 
.A(n_748),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_748),
.Y(n_863)
);

OA21x2_ASAP7_75t_L g864 ( 
.A1(n_702),
.A2(n_699),
.B(n_692),
.Y(n_864)
);

AND2x4_ASAP7_75t_L g865 ( 
.A(n_737),
.B(n_739),
.Y(n_865)
);

OAI21x1_ASAP7_75t_L g866 ( 
.A1(n_771),
.A2(n_800),
.B(n_796),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_797),
.B(n_757),
.Y(n_867)
);

OAI21xp33_ASAP7_75t_SL g868 ( 
.A1(n_709),
.A2(n_695),
.B(n_688),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_757),
.B(n_684),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_748),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_679),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_761),
.B(n_679),
.Y(n_872)
);

NOR2x1_ASAP7_75t_L g873 ( 
.A(n_756),
.B(n_680),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_684),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_SL g875 ( 
.A1(n_746),
.A2(n_697),
.B(n_704),
.Y(n_875)
);

OAI21xp5_ASAP7_75t_L g876 ( 
.A1(n_759),
.A2(n_773),
.B(n_805),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_778),
.B(n_687),
.Y(n_877)
);

INVx1_ASAP7_75t_SL g878 ( 
.A(n_795),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_718),
.B(n_720),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_760),
.B(n_762),
.Y(n_880)
);

AO31x2_ASAP7_75t_L g881 ( 
.A1(n_784),
.A2(n_735),
.A3(n_723),
.B(n_686),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_730),
.A2(n_548),
.B(n_764),
.Y(n_882)
);

AO31x2_ASAP7_75t_L g883 ( 
.A1(n_784),
.A2(n_735),
.A3(n_723),
.B(n_686),
.Y(n_883)
);

AOI21xp33_ASAP7_75t_L g884 ( 
.A1(n_716),
.A2(n_719),
.B(n_707),
.Y(n_884)
);

INVx2_ASAP7_75t_SL g885 ( 
.A(n_795),
.Y(n_885)
);

AO31x2_ASAP7_75t_L g886 ( 
.A1(n_784),
.A2(n_735),
.A3(n_723),
.B(n_686),
.Y(n_886)
);

O2A1O1Ixp5_ASAP7_75t_L g887 ( 
.A1(n_784),
.A2(n_554),
.B(n_780),
.C(n_767),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_760),
.B(n_762),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_760),
.B(n_762),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_760),
.B(n_762),
.Y(n_890)
);

OAI22xp5_ASAP7_75t_L g891 ( 
.A1(n_723),
.A2(n_626),
.B1(n_780),
.B2(n_767),
.Y(n_891)
);

OAI21xp5_ASAP7_75t_L g892 ( 
.A1(n_723),
.A2(n_775),
.B(n_766),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_760),
.B(n_762),
.Y(n_893)
);

OAI21xp5_ASAP7_75t_L g894 ( 
.A1(n_723),
.A2(n_775),
.B(n_766),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_SL g895 ( 
.A1(n_730),
.A2(n_723),
.B(n_636),
.Y(n_895)
);

A2O1A1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_767),
.A2(n_781),
.B(n_790),
.C(n_780),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_718),
.B(n_720),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_718),
.B(n_720),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_683),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_776),
.B(n_787),
.Y(n_900)
);

AO21x1_ASAP7_75t_L g901 ( 
.A1(n_730),
.A2(n_728),
.B(n_707),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_683),
.Y(n_902)
);

BUFx2_ASAP7_75t_L g903 ( 
.A(n_795),
.Y(n_903)
);

BUFx4_ASAP7_75t_R g904 ( 
.A(n_701),
.Y(n_904)
);

AO31x2_ASAP7_75t_L g905 ( 
.A1(n_784),
.A2(n_735),
.A3(n_723),
.B(n_686),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_676),
.B(n_760),
.Y(n_906)
);

OAI22xp5_ASAP7_75t_L g907 ( 
.A1(n_723),
.A2(n_626),
.B1(n_780),
.B2(n_767),
.Y(n_907)
);

OAI22xp5_ASAP7_75t_L g908 ( 
.A1(n_723),
.A2(n_626),
.B1(n_780),
.B2(n_767),
.Y(n_908)
);

OAI21xp5_ASAP7_75t_L g909 ( 
.A1(n_723),
.A2(n_775),
.B(n_766),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_865),
.B(n_845),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_865),
.B(n_845),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_895),
.A2(n_849),
.B(n_882),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_818),
.B(n_841),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_819),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_820),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_818),
.B(n_841),
.Y(n_916)
);

INVx5_ASAP7_75t_L g917 ( 
.A(n_830),
.Y(n_917)
);

OR2x2_ASAP7_75t_L g918 ( 
.A(n_878),
.B(n_826),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_878),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_825),
.Y(n_920)
);

INVx4_ASAP7_75t_L g921 ( 
.A(n_904),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_879),
.B(n_897),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_900),
.A2(n_823),
.B1(n_821),
.B2(n_898),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_848),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_851),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_877),
.B(n_874),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_817),
.B(n_880),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_877),
.B(n_869),
.Y(n_928)
);

BUFx2_ASAP7_75t_L g929 ( 
.A(n_903),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_846),
.B(n_839),
.Y(n_930)
);

BUFx8_ASAP7_75t_L g931 ( 
.A(n_852),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_885),
.B(n_855),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_838),
.Y(n_933)
);

O2A1O1Ixp5_ASAP7_75t_L g934 ( 
.A1(n_891),
.A2(n_908),
.B(n_907),
.C(n_909),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_817),
.B(n_880),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_888),
.B(n_889),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_888),
.B(n_889),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_855),
.B(n_858),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_890),
.B(n_810),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_813),
.B(n_814),
.Y(n_940)
);

NAND2x1_ASAP7_75t_L g941 ( 
.A(n_875),
.B(n_857),
.Y(n_941)
);

BUFx3_ASAP7_75t_L g942 ( 
.A(n_808),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_873),
.B(n_867),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_871),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_890),
.B(n_815),
.Y(n_945)
);

INVx6_ASAP7_75t_SL g946 ( 
.A(n_850),
.Y(n_946)
);

AOI221xp5_ASAP7_75t_L g947 ( 
.A1(n_891),
.A2(n_908),
.B1(n_907),
.B2(n_884),
.C(n_831),
.Y(n_947)
);

HB1xp67_ASAP7_75t_L g948 ( 
.A(n_830),
.Y(n_948)
);

BUFx4f_ASAP7_75t_L g949 ( 
.A(n_830),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_L g950 ( 
.A1(n_893),
.A2(n_896),
.B1(n_831),
.B2(n_853),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_860),
.A2(n_909),
.B1(n_892),
.B2(n_894),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_822),
.B(n_835),
.Y(n_952)
);

INVx2_ASAP7_75t_SL g953 ( 
.A(n_844),
.Y(n_953)
);

CKINVDCx20_ASAP7_75t_R g954 ( 
.A(n_807),
.Y(n_954)
);

INVx1_ASAP7_75t_SL g955 ( 
.A(n_859),
.Y(n_955)
);

CKINVDCx6p67_ASAP7_75t_R g956 ( 
.A(n_902),
.Y(n_956)
);

OA21x2_ASAP7_75t_L g957 ( 
.A1(n_892),
.A2(n_894),
.B(n_809),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_844),
.B(n_863),
.Y(n_958)
);

AOI22xp33_ASAP7_75t_L g959 ( 
.A1(n_884),
.A2(n_906),
.B1(n_812),
.B2(n_854),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_854),
.B(n_834),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_856),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_870),
.B(n_899),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_870),
.B(n_899),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_854),
.B(n_828),
.Y(n_964)
);

INVx2_ASAP7_75t_SL g965 ( 
.A(n_871),
.Y(n_965)
);

BUFx3_ASAP7_75t_L g966 ( 
.A(n_902),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_816),
.B(n_827),
.Y(n_967)
);

HB1xp67_ASAP7_75t_L g968 ( 
.A(n_902),
.Y(n_968)
);

NAND2x1p5_ASAP7_75t_L g969 ( 
.A(n_857),
.B(n_862),
.Y(n_969)
);

AND2x6_ASAP7_75t_L g970 ( 
.A(n_824),
.B(n_829),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_854),
.B(n_837),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_887),
.A2(n_832),
.B(n_868),
.C(n_901),
.Y(n_972)
);

INVx2_ASAP7_75t_SL g973 ( 
.A(n_862),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_876),
.Y(n_974)
);

INVxp67_ASAP7_75t_L g975 ( 
.A(n_833),
.Y(n_975)
);

AOI21xp33_ASAP7_75t_SL g976 ( 
.A1(n_872),
.A2(n_866),
.B(n_832),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_842),
.Y(n_977)
);

CKINVDCx20_ASAP7_75t_R g978 ( 
.A(n_864),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_881),
.B(n_905),
.Y(n_979)
);

AOI22xp33_ASAP7_75t_L g980 ( 
.A1(n_811),
.A2(n_836),
.B1(n_864),
.B2(n_847),
.Y(n_980)
);

INVx4_ASAP7_75t_L g981 ( 
.A(n_811),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_881),
.B(n_886),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_883),
.B(n_886),
.Y(n_983)
);

CKINVDCx8_ASAP7_75t_R g984 ( 
.A(n_883),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_883),
.B(n_840),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_840),
.B(n_861),
.Y(n_986)
);

INVx3_ASAP7_75t_SL g987 ( 
.A(n_861),
.Y(n_987)
);

BUFx12f_ASAP7_75t_L g988 ( 
.A(n_843),
.Y(n_988)
);

BUFx2_ASAP7_75t_SL g989 ( 
.A(n_885),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_818),
.B(n_841),
.Y(n_990)
);

INVx2_ASAP7_75t_SL g991 ( 
.A(n_885),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_818),
.B(n_841),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_900),
.A2(n_818),
.B1(n_841),
.B2(n_760),
.Y(n_993)
);

INVx2_ASAP7_75t_SL g994 ( 
.A(n_885),
.Y(n_994)
);

BUFx12f_ASAP7_75t_L g995 ( 
.A(n_808),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_878),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_826),
.B(n_879),
.Y(n_997)
);

AOI22xp33_ASAP7_75t_L g998 ( 
.A1(n_821),
.A2(n_719),
.B1(n_716),
.B2(n_891),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_904),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_865),
.B(n_845),
.Y(n_1000)
);

BUFx12f_ASAP7_75t_L g1001 ( 
.A(n_808),
.Y(n_1001)
);

INVxp67_ASAP7_75t_L g1002 ( 
.A(n_825),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_820),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_878),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_826),
.B(n_879),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_871),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_818),
.B(n_841),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_904),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_820),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_819),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_819),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_900),
.B(n_776),
.Y(n_1012)
);

OA21x2_ASAP7_75t_L g1013 ( 
.A1(n_892),
.A2(n_909),
.B(n_894),
.Y(n_1013)
);

INVx4_ASAP7_75t_L g1014 ( 
.A(n_904),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_878),
.Y(n_1015)
);

INVx5_ASAP7_75t_L g1016 ( 
.A(n_830),
.Y(n_1016)
);

BUFx12f_ASAP7_75t_L g1017 ( 
.A(n_808),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_830),
.Y(n_1018)
);

INVx1_ASAP7_75t_SL g1019 ( 
.A(n_878),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_900),
.B(n_776),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_895),
.A2(n_730),
.B(n_849),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_900),
.A2(n_818),
.B1(n_841),
.B2(n_760),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_830),
.Y(n_1023)
);

AOI22xp33_ASAP7_75t_L g1024 ( 
.A1(n_821),
.A2(n_719),
.B1(n_716),
.B2(n_891),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_895),
.A2(n_730),
.B(n_849),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_900),
.B(n_776),
.Y(n_1026)
);

AO32x2_ASAP7_75t_L g1027 ( 
.A1(n_891),
.A2(n_907),
.A3(n_908),
.B1(n_856),
.B2(n_716),
.Y(n_1027)
);

NAND2x1p5_ASAP7_75t_L g1028 ( 
.A(n_917),
.B(n_1016),
.Y(n_1028)
);

BUFx12f_ASAP7_75t_L g1029 ( 
.A(n_999),
.Y(n_1029)
);

BUFx2_ASAP7_75t_L g1030 ( 
.A(n_933),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_940),
.B(n_998),
.Y(n_1031)
);

HB1xp67_ASAP7_75t_L g1032 ( 
.A(n_919),
.Y(n_1032)
);

BUFx2_ASAP7_75t_SL g1033 ( 
.A(n_954),
.Y(n_1033)
);

OAI22xp33_ASAP7_75t_L g1034 ( 
.A1(n_1012),
.A2(n_1020),
.B1(n_1026),
.B2(n_923),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_SL g1035 ( 
.A1(n_1012),
.A2(n_1020),
.B1(n_1026),
.B2(n_930),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_913),
.B(n_916),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_919),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_925),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_990),
.B(n_992),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_914),
.Y(n_1040)
);

OR2x6_ASAP7_75t_L g1041 ( 
.A(n_1021),
.B(n_1025),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_998),
.B(n_1024),
.Y(n_1042)
);

OAI22xp33_ASAP7_75t_L g1043 ( 
.A1(n_939),
.A2(n_945),
.B1(n_1007),
.B2(n_937),
.Y(n_1043)
);

INVx3_ASAP7_75t_L g1044 ( 
.A(n_988),
.Y(n_1044)
);

BUFx8_ASAP7_75t_L g1045 ( 
.A(n_995),
.Y(n_1045)
);

BUFx3_ASAP7_75t_L g1046 ( 
.A(n_933),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1010),
.Y(n_1047)
);

BUFx2_ASAP7_75t_R g1048 ( 
.A(n_1008),
.Y(n_1048)
);

INVx1_ASAP7_75t_SL g1049 ( 
.A(n_1019),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1011),
.Y(n_1050)
);

AOI22xp5_ASAP7_75t_SL g1051 ( 
.A1(n_928),
.A2(n_926),
.B1(n_935),
.B2(n_936),
.Y(n_1051)
);

HB1xp67_ASAP7_75t_L g1052 ( 
.A(n_996),
.Y(n_1052)
);

HB1xp67_ASAP7_75t_L g1053 ( 
.A(n_996),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_915),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1003),
.Y(n_1055)
);

AOI22xp33_ASAP7_75t_L g1056 ( 
.A1(n_1024),
.A2(n_952),
.B1(n_947),
.B2(n_959),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1009),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_927),
.A2(n_993),
.B1(n_1022),
.B2(n_959),
.Y(n_1058)
);

AOI22xp33_ASAP7_75t_L g1059 ( 
.A1(n_960),
.A2(n_950),
.B1(n_1013),
.B2(n_951),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_928),
.B(n_943),
.Y(n_1060)
);

HB1xp67_ASAP7_75t_L g1061 ( 
.A(n_1004),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_1015),
.Y(n_1062)
);

AOI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_1013),
.A2(n_997),
.B1(n_1005),
.B2(n_922),
.Y(n_1063)
);

INVx2_ASAP7_75t_SL g1064 ( 
.A(n_949),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_926),
.A2(n_943),
.B1(n_911),
.B2(n_1000),
.Y(n_1065)
);

BUFx2_ASAP7_75t_R g1066 ( 
.A(n_942),
.Y(n_1066)
);

BUFx2_ASAP7_75t_R g1067 ( 
.A(n_942),
.Y(n_1067)
);

AOI22xp33_ASAP7_75t_SL g1068 ( 
.A1(n_989),
.A2(n_964),
.B1(n_1013),
.B2(n_938),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_949),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_918),
.B(n_932),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_958),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_946),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_970),
.Y(n_1073)
);

BUFx2_ASAP7_75t_L g1074 ( 
.A(n_975),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_948),
.Y(n_1075)
);

BUFx3_ASAP7_75t_L g1076 ( 
.A(n_920),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_968),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_929),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_970),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_967),
.B(n_1027),
.Y(n_1080)
);

BUFx4f_ASAP7_75t_SL g1081 ( 
.A(n_946),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_1002),
.B(n_971),
.Y(n_1082)
);

AND2x4_ASAP7_75t_SL g1083 ( 
.A(n_910),
.B(n_1000),
.Y(n_1083)
);

AOI22xp33_ASAP7_75t_L g1084 ( 
.A1(n_953),
.A2(n_975),
.B1(n_970),
.B2(n_961),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_SL g1085 ( 
.A1(n_912),
.A2(n_921),
.B1(n_1014),
.B2(n_957),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_1018),
.Y(n_1086)
);

INVx2_ASAP7_75t_SL g1087 ( 
.A(n_966),
.Y(n_1087)
);

BUFx2_ASAP7_75t_L g1088 ( 
.A(n_970),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_966),
.Y(n_1089)
);

OA21x2_ASAP7_75t_L g1090 ( 
.A1(n_934),
.A2(n_986),
.B(n_980),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_962),
.Y(n_1091)
);

BUFx2_ASAP7_75t_L g1092 ( 
.A(n_970),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_972),
.A2(n_941),
.B(n_985),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_963),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_957),
.Y(n_1095)
);

BUFx2_ASAP7_75t_L g1096 ( 
.A(n_1002),
.Y(n_1096)
);

HB1xp67_ASAP7_75t_L g1097 ( 
.A(n_991),
.Y(n_1097)
);

CKINVDCx20_ASAP7_75t_R g1098 ( 
.A(n_954),
.Y(n_1098)
);

NAND2x1p5_ASAP7_75t_L g1099 ( 
.A(n_977),
.B(n_944),
.Y(n_1099)
);

BUFx10_ASAP7_75t_L g1100 ( 
.A(n_994),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_974),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_974),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_SL g1103 ( 
.A1(n_921),
.A2(n_1014),
.B1(n_978),
.B2(n_931),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_944),
.Y(n_1104)
);

AOI22xp33_ASAP7_75t_L g1105 ( 
.A1(n_978),
.A2(n_987),
.B1(n_981),
.B2(n_983),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_979),
.A2(n_982),
.B(n_969),
.Y(n_1106)
);

OAI21xp5_ASAP7_75t_SL g1107 ( 
.A1(n_955),
.A2(n_976),
.B(n_1027),
.Y(n_1107)
);

OAI21xp5_ASAP7_75t_SL g1108 ( 
.A1(n_1027),
.A2(n_969),
.B(n_973),
.Y(n_1108)
);

BUFx3_ASAP7_75t_L g1109 ( 
.A(n_956),
.Y(n_1109)
);

INVx3_ASAP7_75t_L g1110 ( 
.A(n_1006),
.Y(n_1110)
);

BUFx8_ASAP7_75t_SL g1111 ( 
.A(n_1001),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_1027),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1023),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1023),
.Y(n_1114)
);

BUFx2_ASAP7_75t_L g1115 ( 
.A(n_987),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_SL g1116 ( 
.A1(n_1023),
.A2(n_984),
.B(n_965),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_931),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1017),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_940),
.B(n_821),
.Y(n_1119)
);

AOI22xp33_ASAP7_75t_L g1120 ( 
.A1(n_1012),
.A2(n_1020),
.B1(n_1026),
.B2(n_744),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_924),
.Y(n_1121)
);

BUFx2_ASAP7_75t_L g1122 ( 
.A(n_919),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_924),
.Y(n_1123)
);

OAI221xp5_ASAP7_75t_L g1124 ( 
.A1(n_1120),
.A2(n_1035),
.B1(n_1056),
.B2(n_1058),
.C(n_1085),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_1073),
.B(n_1079),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1080),
.B(n_1101),
.Y(n_1126)
);

BUFx3_ASAP7_75t_L g1127 ( 
.A(n_1115),
.Y(n_1127)
);

HB1xp67_ASAP7_75t_L g1128 ( 
.A(n_1062),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_1115),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1036),
.B(n_1043),
.Y(n_1130)
);

INVxp67_ASAP7_75t_SL g1131 ( 
.A(n_1032),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1095),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_1080),
.B(n_1102),
.Y(n_1133)
);

AOI22xp33_ASAP7_75t_L g1134 ( 
.A1(n_1034),
.A2(n_1042),
.B1(n_1031),
.B2(n_1119),
.Y(n_1134)
);

HB1xp67_ASAP7_75t_SL g1135 ( 
.A(n_1066),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_1073),
.B(n_1079),
.Y(n_1136)
);

HB1xp67_ASAP7_75t_L g1137 ( 
.A(n_1062),
.Y(n_1137)
);

INVx5_ASAP7_75t_SL g1138 ( 
.A(n_1041),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1119),
.B(n_1031),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_1088),
.B(n_1092),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1112),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_1106),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_1098),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_1042),
.B(n_1071),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1090),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_1088),
.B(n_1092),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1090),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1090),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1059),
.B(n_1063),
.Y(n_1149)
);

INVx3_ASAP7_75t_L g1150 ( 
.A(n_1041),
.Y(n_1150)
);

CKINVDCx20_ASAP7_75t_R g1151 ( 
.A(n_1098),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_1106),
.B(n_1060),
.Y(n_1152)
);

AO21x2_ASAP7_75t_L g1153 ( 
.A1(n_1093),
.A2(n_1108),
.B(n_1107),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1041),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_1060),
.B(n_1041),
.Y(n_1155)
);

AO21x1_ASAP7_75t_SL g1156 ( 
.A1(n_1105),
.A2(n_1084),
.B(n_1116),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_1122),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_1070),
.B(n_1049),
.Y(n_1158)
);

HB1xp67_ASAP7_75t_L g1159 ( 
.A(n_1122),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1040),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_1116),
.A2(n_1044),
.B(n_1050),
.Y(n_1161)
);

CKINVDCx20_ASAP7_75t_R g1162 ( 
.A(n_1081),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1047),
.Y(n_1163)
);

INVxp67_ASAP7_75t_L g1164 ( 
.A(n_1078),
.Y(n_1164)
);

BUFx4f_ASAP7_75t_SL g1165 ( 
.A(n_1029),
.Y(n_1165)
);

INVx2_ASAP7_75t_SL g1166 ( 
.A(n_1037),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_1044),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1074),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1038),
.Y(n_1169)
);

INVx3_ASAP7_75t_L g1170 ( 
.A(n_1044),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_1060),
.Y(n_1171)
);

OA21x2_ASAP7_75t_L g1172 ( 
.A1(n_1082),
.A2(n_1123),
.B(n_1121),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1082),
.B(n_1036),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1054),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1039),
.B(n_1061),
.Y(n_1175)
);

INVxp67_ASAP7_75t_SL g1176 ( 
.A(n_1052),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1091),
.B(n_1094),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1055),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1057),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_1068),
.A2(n_1076),
.B1(n_1033),
.B2(n_1103),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_1053),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1141),
.Y(n_1182)
);

INVx5_ASAP7_75t_L g1183 ( 
.A(n_1138),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1126),
.B(n_1051),
.Y(n_1184)
);

HB1xp67_ASAP7_75t_L g1185 ( 
.A(n_1172),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1126),
.B(n_1077),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1133),
.B(n_1075),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1124),
.A2(n_1096),
.B1(n_1076),
.B2(n_1117),
.Y(n_1188)
);

AO21x2_ASAP7_75t_L g1189 ( 
.A1(n_1145),
.A2(n_1148),
.B(n_1147),
.Y(n_1189)
);

OAI221xp5_ASAP7_75t_L g1190 ( 
.A1(n_1130),
.A2(n_1065),
.B1(n_1097),
.B2(n_1030),
.C(n_1118),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1153),
.B(n_1114),
.Y(n_1191)
);

AND3x1_ASAP7_75t_L g1192 ( 
.A(n_1130),
.B(n_1118),
.C(n_1087),
.Y(n_1192)
);

INVx6_ASAP7_75t_L g1193 ( 
.A(n_1155),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1153),
.B(n_1132),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1173),
.B(n_1110),
.Y(n_1195)
);

HB1xp67_ASAP7_75t_L g1196 ( 
.A(n_1172),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1153),
.B(n_1113),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1153),
.B(n_1110),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1168),
.B(n_1046),
.Y(n_1199)
);

OR2x2_ASAP7_75t_L g1200 ( 
.A(n_1147),
.B(n_1046),
.Y(n_1200)
);

OR2x6_ASAP7_75t_L g1201 ( 
.A(n_1154),
.B(n_1099),
.Y(n_1201)
);

INVx1_ASAP7_75t_SL g1202 ( 
.A(n_1181),
.Y(n_1202)
);

NOR2x1p5_ASAP7_75t_L g1203 ( 
.A(n_1170),
.B(n_1109),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1154),
.B(n_1104),
.Y(n_1204)
);

AND2x4_ASAP7_75t_L g1205 ( 
.A(n_1154),
.B(n_1150),
.Y(n_1205)
);

AOI221xp5_ASAP7_75t_L g1206 ( 
.A1(n_1134),
.A2(n_1149),
.B1(n_1164),
.B2(n_1158),
.C(n_1180),
.Y(n_1206)
);

OR2x2_ASAP7_75t_L g1207 ( 
.A(n_1148),
.B(n_1087),
.Y(n_1207)
);

BUFx2_ASAP7_75t_L g1208 ( 
.A(n_1142),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1150),
.B(n_1138),
.Y(n_1209)
);

BUFx3_ASAP7_75t_L g1210 ( 
.A(n_1152),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1150),
.B(n_1086),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_SL g1212 ( 
.A(n_1192),
.B(n_1167),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1210),
.B(n_1152),
.Y(n_1213)
);

OAI221xp5_ASAP7_75t_SL g1214 ( 
.A1(n_1188),
.A2(n_1149),
.B1(n_1175),
.B2(n_1139),
.C(n_1144),
.Y(n_1214)
);

NAND3xp33_ASAP7_75t_L g1215 ( 
.A(n_1188),
.B(n_1157),
.C(n_1159),
.Y(n_1215)
);

OAI221xp5_ASAP7_75t_L g1216 ( 
.A1(n_1206),
.A2(n_1170),
.B1(n_1143),
.B2(n_1167),
.C(n_1131),
.Y(n_1216)
);

NOR3xp33_ASAP7_75t_L g1217 ( 
.A(n_1190),
.B(n_1161),
.C(n_1170),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_1195),
.B(n_1151),
.Y(n_1218)
);

AND4x1_ASAP7_75t_L g1219 ( 
.A(n_1206),
.B(n_1135),
.C(n_1067),
.D(n_1178),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1190),
.A2(n_1155),
.B1(n_1156),
.B2(n_1152),
.Y(n_1220)
);

NAND3xp33_ASAP7_75t_L g1221 ( 
.A(n_1192),
.B(n_1137),
.C(n_1128),
.Y(n_1221)
);

NAND4xp25_ASAP7_75t_L g1222 ( 
.A(n_1202),
.B(n_1181),
.C(n_1169),
.D(n_1177),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1202),
.B(n_1176),
.Y(n_1223)
);

NAND3xp33_ASAP7_75t_L g1224 ( 
.A(n_1199),
.B(n_1166),
.C(n_1169),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1199),
.B(n_1166),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1186),
.B(n_1187),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1186),
.B(n_1139),
.Y(n_1227)
);

NAND3xp33_ASAP7_75t_L g1228 ( 
.A(n_1200),
.B(n_1179),
.C(n_1178),
.Y(n_1228)
);

OAI221xp5_ASAP7_75t_L g1229 ( 
.A1(n_1201),
.A2(n_1170),
.B1(n_1167),
.B2(n_1064),
.C(n_1127),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1210),
.B(n_1152),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1193),
.A2(n_1155),
.B1(n_1171),
.B2(n_1140),
.Y(n_1231)
);

OAI21xp5_ASAP7_75t_SL g1232 ( 
.A1(n_1184),
.A2(n_1155),
.B(n_1083),
.Y(n_1232)
);

OAI221xp5_ASAP7_75t_SL g1233 ( 
.A1(n_1184),
.A2(n_1144),
.B1(n_1177),
.B2(n_1129),
.C(n_1127),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1193),
.A2(n_1171),
.B1(n_1140),
.B2(n_1146),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1210),
.B(n_1191),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_SL g1236 ( 
.A(n_1183),
.B(n_1167),
.Y(n_1236)
);

NAND3xp33_ASAP7_75t_L g1237 ( 
.A(n_1200),
.B(n_1179),
.C(n_1174),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1191),
.B(n_1140),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1203),
.A2(n_1167),
.B1(n_1138),
.B2(n_1146),
.Y(n_1239)
);

OAI221xp5_ASAP7_75t_SL g1240 ( 
.A1(n_1191),
.A2(n_1197),
.B1(n_1198),
.B2(n_1201),
.C(n_1194),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1197),
.B(n_1146),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1182),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1204),
.B(n_1160),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1197),
.B(n_1146),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1198),
.B(n_1138),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1193),
.A2(n_1171),
.B1(n_1167),
.B2(n_1205),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1193),
.A2(n_1171),
.B1(n_1136),
.B2(n_1125),
.Y(n_1247)
);

NAND3xp33_ASAP7_75t_L g1248 ( 
.A(n_1200),
.B(n_1174),
.C(n_1163),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1242),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1235),
.B(n_1194),
.Y(n_1250)
);

NOR2xp67_ASAP7_75t_L g1251 ( 
.A(n_1221),
.B(n_1185),
.Y(n_1251)
);

BUFx2_ASAP7_75t_L g1252 ( 
.A(n_1213),
.Y(n_1252)
);

INVx2_ASAP7_75t_SL g1253 ( 
.A(n_1213),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1238),
.B(n_1198),
.Y(n_1254)
);

OR2x2_ASAP7_75t_L g1255 ( 
.A(n_1240),
.B(n_1185),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1242),
.Y(n_1256)
);

BUFx2_ASAP7_75t_L g1257 ( 
.A(n_1230),
.Y(n_1257)
);

INVx3_ASAP7_75t_L g1258 ( 
.A(n_1230),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1238),
.B(n_1196),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1248),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1241),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1244),
.B(n_1189),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1248),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1244),
.B(n_1189),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1245),
.B(n_1189),
.Y(n_1265)
);

AND2x2_ASAP7_75t_SL g1266 ( 
.A(n_1219),
.B(n_1208),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1245),
.B(n_1189),
.Y(n_1267)
);

OR2x2_ASAP7_75t_L g1268 ( 
.A(n_1243),
.B(n_1189),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1228),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1226),
.B(n_1205),
.Y(n_1270)
);

INVx6_ASAP7_75t_L g1271 ( 
.A(n_1232),
.Y(n_1271)
);

AND2x4_ASAP7_75t_SL g1272 ( 
.A(n_1217),
.B(n_1201),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1228),
.Y(n_1273)
);

INVx2_ASAP7_75t_SL g1274 ( 
.A(n_1236),
.Y(n_1274)
);

OR2x2_ASAP7_75t_L g1275 ( 
.A(n_1223),
.B(n_1207),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1237),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1275),
.B(n_1225),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1275),
.B(n_1227),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1249),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1271),
.B(n_1165),
.Y(n_1280)
);

NAND3xp33_ASAP7_75t_L g1281 ( 
.A(n_1276),
.B(n_1219),
.C(n_1215),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1249),
.Y(n_1282)
);

HB1xp67_ASAP7_75t_L g1283 ( 
.A(n_1276),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_L g1284 ( 
.A(n_1271),
.B(n_1218),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1258),
.B(n_1246),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1258),
.B(n_1209),
.Y(n_1286)
);

AOI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1266),
.A2(n_1216),
.B1(n_1215),
.B2(n_1221),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1256),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1258),
.B(n_1209),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1258),
.B(n_1209),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1258),
.B(n_1193),
.Y(n_1291)
);

OR2x2_ASAP7_75t_L g1292 ( 
.A(n_1255),
.B(n_1222),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1275),
.B(n_1224),
.Y(n_1293)
);

OR2x2_ASAP7_75t_L g1294 ( 
.A(n_1255),
.B(n_1222),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1254),
.B(n_1193),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1256),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1260),
.Y(n_1297)
);

OR2x2_ASAP7_75t_L g1298 ( 
.A(n_1255),
.B(n_1224),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1254),
.B(n_1193),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1261),
.Y(n_1300)
);

NAND2x1_ASAP7_75t_L g1301 ( 
.A(n_1251),
.B(n_1237),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1261),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1254),
.B(n_1231),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1250),
.B(n_1211),
.Y(n_1304)
);

INVx6_ASAP7_75t_L g1305 ( 
.A(n_1266),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1260),
.B(n_1220),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1263),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1263),
.B(n_1269),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1269),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1271),
.B(n_1111),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1259),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1266),
.A2(n_1214),
.B1(n_1233),
.B2(n_1234),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1250),
.B(n_1211),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1273),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1306),
.B(n_1273),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1295),
.B(n_1262),
.Y(n_1316)
);

INVxp67_ASAP7_75t_L g1317 ( 
.A(n_1308),
.Y(n_1317)
);

INVxp33_ASAP7_75t_L g1318 ( 
.A(n_1310),
.Y(n_1318)
);

OR2x2_ASAP7_75t_L g1319 ( 
.A(n_1298),
.B(n_1268),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1279),
.Y(n_1320)
);

NAND2x1_ASAP7_75t_L g1321 ( 
.A(n_1305),
.B(n_1271),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1288),
.Y(n_1322)
);

INVxp67_ASAP7_75t_L g1323 ( 
.A(n_1283),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1295),
.B(n_1262),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1279),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1299),
.B(n_1262),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1293),
.B(n_1270),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1282),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1299),
.B(n_1264),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1298),
.B(n_1270),
.Y(n_1330)
);

OR2x6_ASAP7_75t_L g1331 ( 
.A(n_1301),
.B(n_1271),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1282),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1296),
.Y(n_1333)
);

NAND2x1_ASAP7_75t_L g1334 ( 
.A(n_1305),
.B(n_1271),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1285),
.B(n_1264),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1292),
.B(n_1294),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1296),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1288),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1297),
.B(n_1274),
.Y(n_1339)
);

HB1xp67_ASAP7_75t_L g1340 ( 
.A(n_1297),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1305),
.A2(n_1251),
.B1(n_1229),
.B2(n_1212),
.Y(n_1341)
);

OR2x2_ASAP7_75t_L g1342 ( 
.A(n_1292),
.B(n_1268),
.Y(n_1342)
);

INVxp67_ASAP7_75t_L g1343 ( 
.A(n_1284),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1307),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1304),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1304),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1313),
.Y(n_1347)
);

AOI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1281),
.A2(n_1239),
.B1(n_1272),
.B2(n_1274),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1285),
.B(n_1264),
.Y(n_1349)
);

INVx1_ASAP7_75t_SL g1350 ( 
.A(n_1305),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1294),
.B(n_1270),
.Y(n_1351)
);

AOI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1281),
.A2(n_1272),
.B1(n_1274),
.B2(n_1265),
.Y(n_1352)
);

INVx1_ASAP7_75t_SL g1353 ( 
.A(n_1280),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1307),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1313),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1309),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1340),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1344),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1331),
.B(n_1303),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1354),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1356),
.Y(n_1361)
);

AOI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1331),
.A2(n_1287),
.B1(n_1350),
.B2(n_1343),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1336),
.B(n_1309),
.Y(n_1363)
);

INVxp67_ASAP7_75t_SL g1364 ( 
.A(n_1321),
.Y(n_1364)
);

OR2x2_ASAP7_75t_L g1365 ( 
.A(n_1330),
.B(n_1314),
.Y(n_1365)
);

OR2x2_ASAP7_75t_L g1366 ( 
.A(n_1342),
.B(n_1314),
.Y(n_1366)
);

INVx1_ASAP7_75t_SL g1367 ( 
.A(n_1353),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1339),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1339),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1315),
.B(n_1303),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1342),
.B(n_1301),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1339),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1331),
.B(n_1311),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1351),
.B(n_1311),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1320),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1325),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1328),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1331),
.Y(n_1378)
);

OR2x2_ASAP7_75t_L g1379 ( 
.A(n_1323),
.B(n_1311),
.Y(n_1379)
);

CKINVDCx16_ASAP7_75t_R g1380 ( 
.A(n_1348),
.Y(n_1380)
);

BUFx2_ASAP7_75t_L g1381 ( 
.A(n_1321),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1345),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1332),
.Y(n_1383)
);

BUFx2_ASAP7_75t_L g1384 ( 
.A(n_1334),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1333),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1317),
.B(n_1287),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1337),
.Y(n_1387)
);

NOR3xp33_ASAP7_75t_L g1388 ( 
.A(n_1334),
.B(n_1312),
.C(n_1277),
.Y(n_1388)
);

BUFx3_ASAP7_75t_L g1389 ( 
.A(n_1322),
.Y(n_1389)
);

CKINVDCx16_ASAP7_75t_R g1390 ( 
.A(n_1352),
.Y(n_1390)
);

INVx1_ASAP7_75t_SL g1391 ( 
.A(n_1318),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1375),
.Y(n_1392)
);

CKINVDCx16_ASAP7_75t_R g1393 ( 
.A(n_1380),
.Y(n_1393)
);

AND2x4_ASAP7_75t_L g1394 ( 
.A(n_1367),
.B(n_1364),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1375),
.Y(n_1395)
);

INVxp67_ASAP7_75t_L g1396 ( 
.A(n_1391),
.Y(n_1396)
);

AOI211xp5_ASAP7_75t_L g1397 ( 
.A1(n_1386),
.A2(n_1341),
.B(n_1318),
.C(n_1319),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1359),
.B(n_1335),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1390),
.A2(n_1319),
.B(n_1327),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1362),
.B(n_1335),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1359),
.B(n_1349),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1370),
.B(n_1345),
.Y(n_1402)
);

OAI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1371),
.A2(n_1355),
.B1(n_1346),
.B2(n_1347),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1358),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1378),
.Y(n_1405)
);

OA21x2_ASAP7_75t_L g1406 ( 
.A1(n_1381),
.A2(n_1322),
.B(n_1338),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1363),
.B(n_1346),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1388),
.B(n_1349),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1360),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1361),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1376),
.Y(n_1411)
);

INVxp67_ASAP7_75t_SL g1412 ( 
.A(n_1389),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1377),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1383),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1385),
.Y(n_1415)
);

A2O1A1Ixp33_ASAP7_75t_L g1416 ( 
.A1(n_1378),
.A2(n_1272),
.B(n_1072),
.C(n_1267),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1396),
.B(n_1363),
.Y(n_1417)
);

INVx1_ASAP7_75t_SL g1418 ( 
.A(n_1393),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1397),
.A2(n_1371),
.B1(n_1381),
.B2(n_1384),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1394),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1412),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1394),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1412),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1398),
.B(n_1384),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1396),
.B(n_1408),
.Y(n_1425)
);

NAND3xp33_ASAP7_75t_L g1426 ( 
.A(n_1399),
.B(n_1357),
.C(n_1368),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1405),
.B(n_1357),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_L g1428 ( 
.A(n_1400),
.B(n_1111),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1401),
.A2(n_1374),
.B1(n_1373),
.B2(n_1382),
.Y(n_1429)
);

NAND2xp33_ASAP7_75t_SL g1430 ( 
.A(n_1405),
.B(n_1072),
.Y(n_1430)
);

AND2x4_ASAP7_75t_L g1431 ( 
.A(n_1404),
.B(n_1368),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1409),
.B(n_1369),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1402),
.B(n_1407),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1410),
.B(n_1387),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1411),
.B(n_1162),
.Y(n_1435)
);

O2A1O1Ixp33_ASAP7_75t_SL g1436 ( 
.A1(n_1419),
.A2(n_1403),
.B(n_1416),
.C(n_1395),
.Y(n_1436)
);

OAI222xp33_ASAP7_75t_L g1437 ( 
.A1(n_1419),
.A2(n_1403),
.B1(n_1373),
.B2(n_1379),
.C1(n_1372),
.C2(n_1369),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1418),
.A2(n_1382),
.B1(n_1372),
.B2(n_1374),
.Y(n_1438)
);

NAND4xp25_ASAP7_75t_SL g1439 ( 
.A(n_1426),
.B(n_1416),
.C(n_1415),
.D(n_1413),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1425),
.A2(n_1414),
.B1(n_1365),
.B2(n_1389),
.Y(n_1440)
);

AOI211xp5_ASAP7_75t_L g1441 ( 
.A1(n_1417),
.A2(n_1392),
.B(n_1365),
.C(n_1379),
.Y(n_1441)
);

OAI21xp33_ASAP7_75t_L g1442 ( 
.A1(n_1424),
.A2(n_1422),
.B(n_1420),
.Y(n_1442)
);

AOI211xp5_ASAP7_75t_L g1443 ( 
.A1(n_1430),
.A2(n_1366),
.B(n_1347),
.C(n_1355),
.Y(n_1443)
);

AOI211xp5_ASAP7_75t_L g1444 ( 
.A1(n_1428),
.A2(n_1366),
.B(n_1406),
.C(n_1316),
.Y(n_1444)
);

OAI21xp33_ASAP7_75t_L g1445 ( 
.A1(n_1429),
.A2(n_1324),
.B(n_1316),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1427),
.A2(n_1406),
.B(n_1278),
.Y(n_1446)
);

AOI221x1_ASAP7_75t_L g1447 ( 
.A1(n_1421),
.A2(n_1406),
.B1(n_1324),
.B2(n_1329),
.C(n_1326),
.Y(n_1447)
);

AOI211xp5_ASAP7_75t_L g1448 ( 
.A1(n_1436),
.A2(n_1423),
.B(n_1427),
.C(n_1432),
.Y(n_1448)
);

AND2x4_ASAP7_75t_L g1449 ( 
.A(n_1438),
.B(n_1435),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_SL g1450 ( 
.A(n_1444),
.B(n_1433),
.Y(n_1450)
);

NOR2x1_ASAP7_75t_L g1451 ( 
.A(n_1437),
.B(n_1439),
.Y(n_1451)
);

NAND3xp33_ASAP7_75t_L g1452 ( 
.A(n_1442),
.B(n_1431),
.C(n_1434),
.Y(n_1452)
);

NOR3xp33_ASAP7_75t_L g1453 ( 
.A(n_1441),
.B(n_1434),
.C(n_1431),
.Y(n_1453)
);

NOR3x1_ASAP7_75t_L g1454 ( 
.A(n_1440),
.B(n_1045),
.C(n_1064),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1445),
.B(n_1045),
.Y(n_1455)
);

NOR4xp75_ASAP7_75t_L g1456 ( 
.A(n_1447),
.B(n_1329),
.C(n_1326),
.D(n_1045),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1443),
.B(n_1265),
.Y(n_1457)
);

AOI211xp5_ASAP7_75t_L g1458 ( 
.A1(n_1448),
.A2(n_1446),
.B(n_1109),
.C(n_1069),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1449),
.B(n_1300),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_SL g1460 ( 
.A(n_1451),
.B(n_1029),
.Y(n_1460)
);

NOR4xp25_ASAP7_75t_SL g1461 ( 
.A(n_1450),
.B(n_1252),
.C(n_1257),
.D(n_1048),
.Y(n_1461)
);

NOR2x1_ASAP7_75t_L g1462 ( 
.A(n_1452),
.B(n_1069),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1459),
.Y(n_1463)
);

AOI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1460),
.A2(n_1455),
.B1(n_1453),
.B2(n_1457),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1462),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1461),
.A2(n_1456),
.B1(n_1454),
.B2(n_1203),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1458),
.Y(n_1467)
);

NOR3xp33_ASAP7_75t_L g1468 ( 
.A(n_1460),
.B(n_1161),
.C(n_1286),
.Y(n_1468)
);

NOR2x1_ASAP7_75t_L g1469 ( 
.A(n_1465),
.B(n_1069),
.Y(n_1469)
);

OAI211xp5_ASAP7_75t_L g1470 ( 
.A1(n_1464),
.A2(n_1069),
.B(n_1089),
.C(n_1289),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1463),
.Y(n_1471)
);

CKINVDCx20_ASAP7_75t_R g1472 ( 
.A(n_1467),
.Y(n_1472)
);

NOR5xp2_ASAP7_75t_L g1473 ( 
.A(n_1466),
.B(n_1100),
.C(n_1286),
.D(n_1289),
.E(n_1290),
.Y(n_1473)
);

INVx3_ASAP7_75t_L g1474 ( 
.A(n_1469),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1471),
.Y(n_1475)
);

NAND2x1p5_ASAP7_75t_L g1476 ( 
.A(n_1472),
.B(n_1089),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1474),
.Y(n_1477)
);

NAND5xp2_ASAP7_75t_L g1478 ( 
.A(n_1477),
.B(n_1475),
.C(n_1470),
.D(n_1476),
.E(n_1468),
.Y(n_1478)
);

O2A1O1Ixp5_ASAP7_75t_L g1479 ( 
.A1(n_1478),
.A2(n_1474),
.B(n_1476),
.C(n_1473),
.Y(n_1479)
);

OAI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1478),
.A2(n_1302),
.B1(n_1300),
.B2(n_1253),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1479),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1480),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1481),
.B(n_1100),
.Y(n_1483)
);

AOI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1482),
.A2(n_1302),
.B(n_1290),
.Y(n_1484)
);

OAI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1483),
.A2(n_1291),
.B(n_1267),
.Y(n_1485)
);

AOI22xp5_ASAP7_75t_SL g1486 ( 
.A1(n_1485),
.A2(n_1484),
.B1(n_1100),
.B2(n_1028),
.Y(n_1486)
);

OAI221xp5_ASAP7_75t_R g1487 ( 
.A1(n_1486),
.A2(n_1247),
.B1(n_1291),
.B2(n_1257),
.C(n_1252),
.Y(n_1487)
);

AOI211xp5_ASAP7_75t_L g1488 ( 
.A1(n_1487),
.A2(n_1086),
.B(n_1267),
.C(n_1265),
.Y(n_1488)
);


endmodule