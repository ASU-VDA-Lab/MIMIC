module fake_netlist_1_7488_n_17 (n_1, n_2, n_0, n_17);
input n_1;
input n_2;
input n_0;
output n_17;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
NOR2xp33_ASAP7_75t_SL g3 ( .A(n_0), .B(n_1), .Y(n_3) );
INVx1_ASAP7_75t_L g4 ( .A(n_0), .Y(n_4) );
AND2x6_ASAP7_75t_L g5 ( .A(n_0), .B(n_2), .Y(n_5) );
AND2x2_ASAP7_75t_L g6 ( .A(n_0), .B(n_1), .Y(n_6) );
AND2x2_ASAP7_75t_L g7 ( .A(n_6), .B(n_1), .Y(n_7) );
INVx2_ASAP7_75t_L g8 ( .A(n_4), .Y(n_8) );
OAI21x1_ASAP7_75t_L g9 ( .A1(n_4), .A2(n_2), .B(n_6), .Y(n_9) );
AND2x2_ASAP7_75t_L g10 ( .A(n_7), .B(n_5), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_8), .Y(n_11) );
OAI22xp5_ASAP7_75t_L g12 ( .A1(n_10), .A2(n_8), .B1(n_3), .B2(n_9), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_11), .B(n_9), .Y(n_13) );
NAND4xp75_ASAP7_75t_L g14 ( .A(n_13), .B(n_2), .C(n_5), .D(n_12), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_13), .Y(n_15) );
NAND2xp5_ASAP7_75t_SL g16 ( .A(n_15), .B(n_5), .Y(n_16) );
AOI22xp5_ASAP7_75t_L g17 ( .A1(n_16), .A2(n_5), .B1(n_14), .B2(n_10), .Y(n_17) );
endmodule