module fake_jpeg_840_n_178 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_178);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_13),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_9),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_16),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_0),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_61),
.Y(n_72)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_51),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_68),
.B(n_70),
.Y(n_73)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_44),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_62),
.B1(n_46),
.B2(n_52),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_71),
.A2(n_55),
.B1(n_74),
.B2(n_59),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_60),
.Y(n_92)
);

CKINVDCx9p33_ASAP7_75t_R g77 ( 
.A(n_69),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g89 ( 
.A(n_77),
.Y(n_89)
);

CKINVDCx12_ASAP7_75t_R g78 ( 
.A(n_63),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_78),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_53),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_80),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_46),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_58),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_R g86 ( 
.A(n_81),
.B(n_52),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_81),
.A2(n_62),
.B1(n_65),
.B2(n_67),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_91),
.B1(n_95),
.B2(n_98),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_88),
.Y(n_106)
);

NAND2xp33_ASAP7_75t_SL g88 ( 
.A(n_76),
.B(n_69),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

OA21x2_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_83),
.B(n_82),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_99),
.Y(n_103)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_60),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_97),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_56),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_74),
.A2(n_50),
.B1(n_56),
.B2(n_48),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_48),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_91),
.Y(n_119)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_76),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_108),
.B(n_109),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_50),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_1),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_117),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_45),
.C(n_24),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_115),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_1),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_2),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_45),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_118),
.B(n_21),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_106),
.A2(n_47),
.B(n_89),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_120),
.A2(n_122),
.B(n_30),
.Y(n_148)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_123),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_2),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_124),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_144)
);

XNOR2x2_ASAP7_75t_SL g125 ( 
.A(n_118),
.B(n_3),
.Y(n_125)
);

OAI32xp33_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_31),
.A3(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_4),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_127),
.B(n_129),
.Y(n_154)
);

AND2x6_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_28),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_132),
.Y(n_143)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_131),
.Y(n_151)
);

AND2x6_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_43),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_135),
.A2(n_114),
.B1(n_11),
.B2(n_12),
.Y(n_142)
);

NOR2x1_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_6),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_137),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_8),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_101),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_145),
.C(n_130),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_153),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_144),
.A2(n_146),
.B1(n_147),
.B2(n_123),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_128),
.C(n_119),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_126),
.A2(n_15),
.B1(n_18),
.B2(n_19),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_137),
.A2(n_15),
.B1(n_25),
.B2(n_27),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_147),
.Y(n_160)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_149),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_160),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_138),
.Y(n_159)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_159),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_162),
.C(n_154),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_37),
.C(n_38),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_163),
.A2(n_164),
.B1(n_162),
.B2(n_140),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_161),
.A2(n_152),
.B1(n_157),
.B2(n_156),
.Y(n_164)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_166),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_169),
.Y(n_171)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_164),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_169),
.B(n_167),
.Y(n_172)
);

AOI322xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_166),
.A3(n_167),
.B1(n_170),
.B2(n_152),
.C1(n_165),
.C2(n_141),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_173),
.A2(n_165),
.B(n_171),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_174),
.Y(n_175)
);

AOI322xp5_ASAP7_75t_L g176 ( 
.A1(n_175),
.A2(n_166),
.A3(n_143),
.B1(n_163),
.B2(n_151),
.C1(n_41),
.C2(n_42),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_151),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_39),
.Y(n_178)
);


endmodule