module real_aes_8791_n_350 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_350);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_350;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_979;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_900;
wire n_841;
wire n_718;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_555;
wire n_421;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_593;
wire n_460;
wire n_937;
wire n_989;
wire n_773;
wire n_401;
wire n_538;
wire n_353;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_537;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_1021;
wire n_700;
wire n_677;
wire n_958;
wire n_1046;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_1040;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_994;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_875;
wire n_467;
wire n_951;
wire n_992;
wire n_774;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_962;
wire n_693;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_755;
wire n_1025;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_725;
wire n_973;
wire n_455;
wire n_504;
wire n_671;
wire n_960;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_940;
wire n_770;
wire n_808;
wire n_722;
wire n_745;
wire n_867;
wire n_398;
wire n_688;
wire n_609;
wire n_425;
wire n_1042;
wire n_879;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_676;
wire n_658;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_1031;
wire n_880;
wire n_1037;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_999;
wire n_490;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_985;
wire n_777;
wire n_488;
wire n_501;
wire n_1041;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_756;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_1028;
wire n_366;
wire n_727;
wire n_1014;
wire n_397;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_354;
wire n_720;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_365;
wire n_653;
wire n_526;
wire n_928;
wire n_637;
wire n_899;
wire n_692;
wire n_789;
wire n_544;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_959;
wire n_715;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_721;
wire n_446;
wire n_681;
wire n_982;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_587;
wire n_546;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_968;
wire n_650;
wire n_646;
wire n_710;
wire n_743;
wire n_393;
wire n_652;
wire n_703;
wire n_823;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1024;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_0), .A2(n_182), .B1(n_486), .B2(n_973), .Y(n_972) );
INVx1_ASAP7_75t_L g854 ( .A(n_1), .Y(n_854) );
AOI22xp33_ASAP7_75t_SL g1042 ( .A1(n_2), .A2(n_139), .B1(n_423), .B2(n_428), .Y(n_1042) );
AOI222xp33_ASAP7_75t_L g431 ( .A1(n_3), .A2(n_172), .B1(n_306), .B2(n_432), .C1(n_434), .C2(n_438), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_4), .A2(n_239), .B1(n_524), .B2(n_647), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_5), .A2(n_104), .B1(n_650), .B2(n_708), .Y(n_707) );
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_6), .A2(n_302), .B1(n_650), .B2(n_688), .C(n_689), .Y(n_687) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_7), .Y(n_733) );
AOI22xp33_ASAP7_75t_SL g517 ( .A1(n_8), .A2(n_155), .B1(n_518), .B2(n_519), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_9), .A2(n_95), .B1(n_522), .B2(n_564), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_10), .A2(n_80), .B1(n_438), .B2(n_613), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_11), .B(n_510), .Y(n_509) );
AO22x2_ASAP7_75t_L g381 ( .A1(n_12), .A2(n_210), .B1(n_373), .B2(n_378), .Y(n_381) );
INVx1_ASAP7_75t_L g1000 ( .A(n_12), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_13), .A2(n_166), .B1(n_402), .B2(n_405), .Y(n_401) );
AOI22xp33_ASAP7_75t_SL g813 ( .A1(n_14), .A2(n_330), .B1(n_423), .B2(n_460), .Y(n_813) );
AOI222xp33_ASAP7_75t_L g1046 ( .A1(n_15), .A2(n_301), .B1(n_307), .B2(n_589), .C1(n_591), .C2(n_964), .Y(n_1046) );
AOI22xp5_ASAP7_75t_L g952 ( .A1(n_16), .A2(n_152), .B1(n_526), .B2(n_620), .Y(n_952) );
CKINVDCx20_ASAP7_75t_R g919 ( .A(n_17), .Y(n_919) );
CKINVDCx20_ASAP7_75t_R g930 ( .A(n_18), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_19), .A2(n_188), .B1(n_507), .B2(n_667), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_20), .A2(n_235), .B1(n_585), .B2(n_620), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_21), .A2(n_295), .B1(n_489), .B2(n_561), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_22), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_23), .A2(n_296), .B1(n_494), .B2(n_735), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_24), .A2(n_220), .B1(n_493), .B2(n_494), .Y(n_492) );
AOI222xp33_ASAP7_75t_L g588 ( .A1(n_25), .A2(n_67), .B1(n_262), .B2(n_460), .C1(n_589), .C2(n_591), .Y(n_588) );
AOI22xp5_ASAP7_75t_SL g800 ( .A1(n_26), .A2(n_233), .B1(n_526), .B2(n_801), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g940 ( .A(n_27), .Y(n_940) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_28), .A2(n_39), .B1(n_507), .B2(n_696), .C(n_697), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_29), .A2(n_151), .B1(n_526), .B2(n_791), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_30), .A2(n_334), .B1(n_519), .B2(n_587), .Y(n_953) );
CKINVDCx20_ASAP7_75t_R g913 ( .A(n_31), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_32), .A2(n_231), .B1(n_405), .B2(n_522), .Y(n_670) );
AO22x2_ASAP7_75t_L g383 ( .A1(n_33), .A2(n_118), .B1(n_373), .B2(n_374), .Y(n_383) );
INVx1_ASAP7_75t_L g451 ( .A(n_34), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_35), .A2(n_170), .B1(n_396), .B2(n_409), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g593 ( .A(n_36), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g958 ( .A1(n_37), .A2(n_959), .B1(n_979), .B2(n_980), .Y(n_958) );
INVx1_ASAP7_75t_L g980 ( .A(n_37), .Y(n_980) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_38), .A2(n_56), .B1(n_479), .B2(n_522), .Y(n_782) );
CKINVDCx20_ASAP7_75t_R g549 ( .A(n_40), .Y(n_549) );
AOI22xp33_ASAP7_75t_SL g673 ( .A1(n_41), .A2(n_61), .B1(n_390), .B2(n_402), .Y(n_673) );
INVx1_ASAP7_75t_L g832 ( .A(n_42), .Y(n_832) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_43), .A2(n_271), .B1(n_438), .B2(n_663), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g1009 ( .A1(n_44), .A2(n_63), .B1(n_367), .B2(n_404), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_45), .A2(n_159), .B1(n_405), .B2(n_791), .Y(n_899) );
INVx1_ASAP7_75t_L g693 ( .A(n_46), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_47), .A2(n_281), .B1(n_650), .B2(n_654), .Y(n_977) );
INVx1_ASAP7_75t_L g895 ( .A(n_48), .Y(n_895) );
AOI22xp5_ASAP7_75t_L g830 ( .A1(n_49), .A2(n_199), .B1(n_428), .B2(n_439), .Y(n_830) );
AOI222xp33_ASAP7_75t_L g700 ( .A1(n_50), .A2(n_132), .B1(n_140), .B2(n_432), .C1(n_458), .C2(n_463), .Y(n_700) );
AOI222xp33_ASAP7_75t_L g722 ( .A1(n_51), .A2(n_279), .B1(n_294), .B2(n_639), .C1(n_723), .C2(n_724), .Y(n_722) );
AOI22xp5_ASAP7_75t_SL g799 ( .A1(n_52), .A2(n_291), .B1(n_524), .B2(n_616), .Y(n_799) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_53), .Y(n_441) );
AOI22xp5_ASAP7_75t_SL g1008 ( .A1(n_54), .A2(n_209), .B1(n_616), .B2(n_620), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g1037 ( .A1(n_55), .A2(n_90), .B1(n_519), .B2(n_616), .Y(n_1037) );
CKINVDCx20_ASAP7_75t_R g917 ( .A(n_57), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_58), .A2(n_303), .B1(n_512), .B2(n_582), .Y(n_581) );
CKINVDCx16_ASAP7_75t_R g909 ( .A(n_59), .Y(n_909) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_60), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g1041 ( .A(n_62), .B(n_667), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_64), .B(n_724), .Y(n_776) );
CKINVDCx20_ASAP7_75t_R g675 ( .A(n_65), .Y(n_675) );
AOI22xp33_ASAP7_75t_SL g876 ( .A1(n_66), .A2(n_232), .B1(n_877), .B2(n_879), .Y(n_876) );
AOI22xp5_ASAP7_75t_L g896 ( .A1(n_68), .A2(n_94), .B1(n_438), .B2(n_512), .Y(n_896) );
INVx1_ASAP7_75t_L g461 ( .A(n_69), .Y(n_461) );
AOI22xp33_ASAP7_75t_SL g514 ( .A1(n_70), .A2(n_125), .B1(n_515), .B2(n_516), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_71), .A2(n_322), .B1(n_402), .B2(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g851 ( .A(n_72), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_73), .A2(n_142), .B1(n_408), .B2(n_789), .Y(n_788) );
NAND2xp5_ASAP7_75t_SL g841 ( .A(n_74), .B(n_805), .Y(n_841) );
CKINVDCx20_ASAP7_75t_R g962 ( .A(n_75), .Y(n_962) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_76), .A2(n_93), .B1(n_644), .B2(n_645), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_77), .A2(n_206), .B1(n_508), .B2(n_667), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g950 ( .A(n_78), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_79), .A2(n_217), .B1(n_555), .B2(n_556), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_81), .A2(n_99), .B1(n_647), .B2(n_784), .Y(n_783) );
AOI22xp33_ASAP7_75t_SL g881 ( .A1(n_82), .A2(n_215), .B1(n_577), .B2(n_882), .Y(n_881) );
AOI22xp5_ASAP7_75t_SL g1011 ( .A1(n_83), .A2(n_100), .B1(n_522), .B2(n_882), .Y(n_1011) );
AO22x2_ASAP7_75t_L g377 ( .A1(n_84), .A2(n_243), .B1(n_373), .B2(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g997 ( .A(n_84), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_85), .A2(n_252), .B1(n_396), .B2(n_587), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_86), .A2(n_325), .B1(n_591), .B2(n_946), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_87), .A2(n_323), .B1(n_411), .B2(n_791), .Y(n_955) );
AOI211xp5_ASAP7_75t_L g350 ( .A1(n_88), .A2(n_351), .B(n_359), .C(n_1002), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_89), .A2(n_339), .B1(n_793), .B2(n_794), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_91), .A2(n_275), .B1(n_580), .B2(n_719), .Y(n_966) );
AOI22xp5_ASAP7_75t_L g963 ( .A1(n_92), .A2(n_203), .B1(n_724), .B2(n_964), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_96), .A2(n_268), .B1(n_493), .B2(n_494), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_97), .A2(n_287), .B1(n_367), .B2(n_516), .Y(n_954) );
OA22x2_ASAP7_75t_L g703 ( .A1(n_98), .A2(n_704), .B1(n_705), .B2(n_725), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_98), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g900 ( .A1(n_101), .A2(n_114), .B1(n_515), .B2(n_522), .Y(n_900) );
AOI22xp33_ASAP7_75t_SL g1012 ( .A1(n_102), .A2(n_194), .B1(n_654), .B2(n_805), .Y(n_1012) );
AOI22xp33_ASAP7_75t_SL g665 ( .A1(n_103), .A2(n_107), .B1(n_423), .B2(n_639), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_105), .A2(n_124), .B1(n_566), .B2(n_975), .Y(n_974) );
AOI22xp33_ASAP7_75t_SL g867 ( .A1(n_106), .A2(n_154), .B1(n_721), .B2(n_868), .Y(n_867) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_108), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g809 ( .A(n_109), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g840 ( .A(n_110), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_111), .B(n_891), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_112), .A2(n_136), .B1(n_489), .B2(n_491), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g833 ( .A(n_113), .Y(n_833) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_115), .A2(n_261), .B1(n_577), .B2(n_616), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_116), .A2(n_258), .B1(n_516), .B2(n_975), .Y(n_1044) );
INVx1_ASAP7_75t_L g611 ( .A(n_117), .Y(n_611) );
INVx1_ASAP7_75t_L g1001 ( .A(n_118), .Y(n_1001) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_119), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_120), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_121), .A2(n_191), .B1(n_424), .B2(n_609), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_122), .A2(n_126), .B1(n_618), .B2(n_654), .Y(n_903) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_123), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g1015 ( .A(n_127), .Y(n_1015) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_128), .Y(n_745) );
AOI211xp5_ASAP7_75t_L g911 ( .A1(n_129), .A2(n_723), .B(n_912), .C(n_916), .Y(n_911) );
INVx1_ASAP7_75t_L g623 ( .A(n_130), .Y(n_623) );
CKINVDCx20_ASAP7_75t_R g837 ( .A(n_131), .Y(n_837) );
INVx1_ASAP7_75t_L g904 ( .A(n_133), .Y(n_904) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_134), .A2(n_169), .B1(n_384), .B2(n_515), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_135), .A2(n_310), .B1(n_622), .B2(n_652), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g1019 ( .A1(n_137), .A2(n_242), .B1(n_427), .B2(n_865), .Y(n_1019) );
AOI22xp33_ASAP7_75t_SL g478 ( .A1(n_138), .A2(n_228), .B1(n_479), .B2(n_482), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_141), .A2(n_332), .B1(n_423), .B2(n_460), .Y(n_893) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_143), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_144), .A2(n_248), .B1(n_561), .B2(n_562), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_145), .A2(n_178), .B1(n_390), .B2(n_396), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_146), .A2(n_331), .B1(n_721), .B2(n_868), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_147), .A2(n_283), .B1(n_405), .B2(n_411), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_148), .A2(n_255), .B1(n_428), .B2(n_721), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_149), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g978 ( .A1(n_150), .A2(n_222), .B1(n_493), .B2(n_879), .Y(n_978) );
AND2x6_ASAP7_75t_L g353 ( .A(n_153), .B(n_354), .Y(n_353) );
HB1xp67_ASAP7_75t_L g994 ( .A(n_153), .Y(n_994) );
CKINVDCx20_ASAP7_75t_R g835 ( .A(n_156), .Y(n_835) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_157), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g1021 ( .A(n_158), .Y(n_1021) );
AOI22xp33_ASAP7_75t_SL g902 ( .A1(n_160), .A2(n_327), .B1(n_390), .B2(n_786), .Y(n_902) );
AOI22xp5_ASAP7_75t_L g811 ( .A1(n_161), .A2(n_227), .B1(n_428), .B2(n_438), .Y(n_811) );
CKINVDCx20_ASAP7_75t_R g1032 ( .A(n_162), .Y(n_1032) );
AOI22xp33_ASAP7_75t_SL g521 ( .A1(n_163), .A2(n_340), .B1(n_405), .B2(n_522), .Y(n_521) );
AO22x1_ASAP7_75t_L g685 ( .A1(n_164), .A2(n_174), .B1(n_491), .B2(n_686), .Y(n_685) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_165), .Y(n_527) );
AOI221xp5_ASAP7_75t_L g684 ( .A1(n_167), .A2(n_309), .B1(n_524), .B2(n_647), .C(n_685), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_168), .A2(n_250), .B1(n_711), .B2(n_713), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_171), .A2(n_347), .B1(n_464), .B2(n_613), .Y(n_612) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_173), .Y(n_741) );
AOI22xp33_ASAP7_75t_SL g617 ( .A1(n_175), .A2(n_179), .B1(n_408), .B2(n_618), .Y(n_617) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_176), .Y(n_778) );
AO22x2_ASAP7_75t_L g372 ( .A1(n_177), .A2(n_234), .B1(n_373), .B2(n_374), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g998 ( .A(n_177), .B(n_999), .Y(n_998) );
CKINVDCx20_ASAP7_75t_R g1039 ( .A(n_180), .Y(n_1039) );
CKINVDCx20_ASAP7_75t_R g941 ( .A(n_181), .Y(n_941) );
AOI22xp33_ASAP7_75t_SL g523 ( .A1(n_183), .A2(n_249), .B1(n_524), .B2(n_526), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_184), .A2(n_236), .B1(n_367), .B2(n_384), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_185), .A2(n_285), .B1(n_864), .B2(n_865), .Y(n_863) );
AOI22xp33_ASAP7_75t_SL g619 ( .A1(n_186), .A2(n_320), .B1(n_384), .B2(n_620), .Y(n_619) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_187), .Y(n_545) );
AOI22xp5_ASAP7_75t_SL g803 ( .A1(n_189), .A2(n_257), .B1(n_804), .B2(n_805), .Y(n_803) );
CKINVDCx20_ASAP7_75t_R g637 ( .A(n_190), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_192), .A2(n_224), .B1(n_405), .B2(n_411), .Y(n_575) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_193), .Y(n_768) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_195), .A2(n_315), .B1(n_396), .B2(n_652), .Y(n_651) );
CKINVDCx20_ASAP7_75t_R g655 ( .A(n_196), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_197), .B(n_419), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_198), .A2(n_729), .B1(n_760), .B2(n_761), .Y(n_728) );
INVx1_ASAP7_75t_L g760 ( .A(n_198), .Y(n_760) );
XOR2xp5_ASAP7_75t_L g1003 ( .A(n_200), .B(n_1004), .Y(n_1003) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_201), .Y(n_774) );
AOI22xp33_ASAP7_75t_SL g649 ( .A1(n_202), .A2(n_341), .B1(n_616), .B2(n_650), .Y(n_649) );
CKINVDCx20_ASAP7_75t_R g926 ( .A(n_204), .Y(n_926) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_205), .A2(n_681), .B1(n_682), .B2(n_701), .Y(n_680) );
INVx1_ASAP7_75t_L g701 ( .A(n_205), .Y(n_701) );
INVx1_ASAP7_75t_L g456 ( .A(n_207), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g943 ( .A(n_208), .Y(n_943) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_211), .A2(n_534), .B1(n_567), .B2(n_568), .Y(n_533) );
INVx1_ASAP7_75t_L g567 ( .A(n_211), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_212), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_213), .A2(n_226), .B1(n_402), .B2(n_688), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_214), .A2(n_328), .B1(n_622), .B2(n_652), .Y(n_923) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_216), .B(n_507), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_218), .A2(n_277), .B1(n_868), .B2(n_968), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_219), .A2(n_336), .B1(n_408), .B2(n_411), .Y(n_407) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_221), .Y(n_815) );
AOI22xp33_ASAP7_75t_SL g874 ( .A1(n_223), .A2(n_253), .B1(n_804), .B2(n_875), .Y(n_874) );
AOI22xp5_ASAP7_75t_SL g443 ( .A1(n_225), .A2(n_444), .B1(n_495), .B2(n_496), .Y(n_443) );
INVx1_ASAP7_75t_L g496 ( .A(n_225), .Y(n_496) );
INVx2_ASAP7_75t_L g358 ( .A(n_229), .Y(n_358) );
AOI22xp33_ASAP7_75t_SL g504 ( .A1(n_230), .A2(n_300), .B1(n_439), .B2(n_460), .Y(n_504) );
INVx1_ASAP7_75t_L g447 ( .A(n_237), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_238), .A2(n_247), .B1(n_524), .B2(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g471 ( .A(n_240), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_241), .A2(n_290), .B1(n_515), .B2(n_585), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_244), .A2(n_289), .B1(n_518), .B2(n_879), .Y(n_924) );
INVx1_ASAP7_75t_L g829 ( .A(n_245), .Y(n_829) );
CKINVDCx20_ASAP7_75t_R g862 ( .A(n_246), .Y(n_862) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_251), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_254), .A2(n_293), .B1(n_696), .B2(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_256), .B(n_507), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g849 ( .A(n_259), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_260), .A2(n_335), .B1(n_507), .B2(n_580), .Y(n_579) );
AOI22xp33_ASAP7_75t_SL g883 ( .A1(n_263), .A2(n_349), .B1(n_644), .B2(n_647), .Y(n_883) );
CKINVDCx20_ASAP7_75t_R g1016 ( .A(n_264), .Y(n_1016) );
INVx1_ASAP7_75t_L g373 ( .A(n_265), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_265), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_266), .A2(n_270), .B1(n_696), .B2(n_871), .Y(n_870) );
INVx1_ASAP7_75t_L g632 ( .A(n_267), .Y(n_632) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_269), .Y(n_769) );
CKINVDCx20_ASAP7_75t_R g843 ( .A(n_272), .Y(n_843) );
CKINVDCx20_ASAP7_75t_R g847 ( .A(n_273), .Y(n_847) );
CKINVDCx20_ASAP7_75t_R g698 ( .A(n_274), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_276), .A2(n_313), .B1(n_515), .B2(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g630 ( .A(n_278), .Y(n_630) );
CKINVDCx20_ASAP7_75t_R g1023 ( .A(n_280), .Y(n_1023) );
AOI22xp33_ASAP7_75t_SL g511 ( .A1(n_282), .A2(n_321), .B1(n_424), .B2(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_284), .B(n_463), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g948 ( .A(n_286), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_288), .A2(n_314), .B1(n_423), .B2(n_427), .Y(n_422) );
AO22x2_ASAP7_75t_L g936 ( .A1(n_292), .A2(n_937), .B1(n_956), .B2(n_957), .Y(n_936) );
CKINVDCx20_ASAP7_75t_R g957 ( .A(n_292), .Y(n_957) );
CKINVDCx20_ASAP7_75t_R g858 ( .A(n_297), .Y(n_858) );
INVx1_ASAP7_75t_L g357 ( .A(n_298), .Y(n_357) );
INVx1_ASAP7_75t_L g354 ( .A(n_299), .Y(n_354) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_304), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_305), .B(n_419), .Y(n_892) );
INVx1_ASAP7_75t_L g855 ( .A(n_308), .Y(n_855) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_311), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_312), .B(n_580), .Y(n_914) );
CKINVDCx20_ASAP7_75t_R g844 ( .A(n_316), .Y(n_844) );
CKINVDCx20_ASAP7_75t_R g1018 ( .A(n_317), .Y(n_1018) );
CKINVDCx20_ASAP7_75t_R g415 ( .A(n_318), .Y(n_415) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_319), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g640 ( .A(n_324), .Y(n_640) );
INVx1_ASAP7_75t_L g932 ( .A(n_326), .Y(n_932) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_329), .B(n_419), .Y(n_606) );
CKINVDCx20_ASAP7_75t_R g928 ( .A(n_333), .Y(n_928) );
INVx1_ASAP7_75t_L g466 ( .A(n_337), .Y(n_466) );
INVx1_ASAP7_75t_L g690 ( .A(n_338), .Y(n_690) );
CKINVDCx20_ASAP7_75t_R g634 ( .A(n_342), .Y(n_634) );
OA22x2_ASAP7_75t_L g763 ( .A1(n_343), .A2(n_764), .B1(n_765), .B2(n_795), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_343), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g699 ( .A(n_344), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_345), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_346), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g661 ( .A(n_348), .Y(n_661) );
INVx2_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_SL g352 ( .A(n_353), .B(n_355), .Y(n_352) );
HB1xp67_ASAP7_75t_L g993 ( .A(n_354), .Y(n_993) );
OA21x2_ASAP7_75t_L g1030 ( .A1(n_355), .A2(n_992), .B(n_1031), .Y(n_1030) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .Y(n_355) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AOI221xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_596), .B1(n_987), .B2(n_988), .C(n_989), .Y(n_359) );
INVx1_ASAP7_75t_L g988 ( .A(n_360), .Y(n_988) );
AOI22xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_530), .B1(n_594), .B2(n_595), .Y(n_360) );
INVx1_ASAP7_75t_L g594 ( .A(n_361), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_363), .B1(n_442), .B2(n_529), .Y(n_361) );
INVx2_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
XOR2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_441), .Y(n_363) );
NAND4xp75_ASAP7_75t_L g364 ( .A(n_365), .B(n_400), .C(n_414), .D(n_431), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_389), .Y(n_365) );
INVx3_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx3_ASAP7_75t_L g515 ( .A(n_368), .Y(n_515) );
OAI22xp5_ASAP7_75t_SL g842 ( .A1(n_368), .A2(n_403), .B1(n_843), .B2(n_844), .Y(n_842) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_369), .Y(n_490) );
BUFx2_ASAP7_75t_SL g801 ( .A(n_369), .Y(n_801) );
BUFx2_ASAP7_75t_SL g975 ( .A(n_369), .Y(n_975) );
AND2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_379), .Y(n_369) );
AND2x6_ASAP7_75t_L g386 ( .A(n_370), .B(n_387), .Y(n_386) );
AND2x4_ASAP7_75t_L g404 ( .A(n_370), .B(n_395), .Y(n_404) );
AND2x6_ASAP7_75t_L g433 ( .A(n_370), .B(n_430), .Y(n_433) );
AND2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_376), .Y(n_370) );
AND2x2_ASAP7_75t_L g410 ( .A(n_371), .B(n_377), .Y(n_410) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g393 ( .A(n_372), .B(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_372), .B(n_377), .Y(n_399) );
AND2x2_ASAP7_75t_L g426 ( .A(n_372), .B(n_381), .Y(n_426) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g378 ( .A(n_375), .Y(n_378) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g394 ( .A(n_377), .Y(n_394) );
INVx1_ASAP7_75t_L g437 ( .A(n_377), .Y(n_437) );
AND2x2_ASAP7_75t_L g406 ( .A(n_379), .B(n_393), .Y(n_406) );
AND2x4_ASAP7_75t_L g409 ( .A(n_379), .B(n_410), .Y(n_409) );
AND2x4_ASAP7_75t_L g412 ( .A(n_379), .B(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_379), .B(n_393), .Y(n_852) );
AND2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
OR2x2_ASAP7_75t_L g388 ( .A(n_380), .B(n_383), .Y(n_388) );
AND2x2_ASAP7_75t_L g395 ( .A(n_380), .B(n_383), .Y(n_395) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g430 ( .A(n_381), .B(n_383), .Y(n_430) );
AND2x2_ASAP7_75t_L g436 ( .A(n_382), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g470 ( .A(n_382), .Y(n_470) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g398 ( .A(n_383), .Y(n_398) );
INVx5_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g486 ( .A(n_385), .Y(n_486) );
INVx2_ASAP7_75t_SL g791 ( .A(n_385), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g853 ( .A(n_385), .B(n_854), .Y(n_853) );
INVx11_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx11_ASAP7_75t_L g525 ( .A(n_386), .Y(n_525) );
AND2x4_ASAP7_75t_L g421 ( .A(n_387), .B(n_410), .Y(n_421) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OR2x2_ASAP7_75t_L g449 ( .A(n_388), .B(n_450), .Y(n_449) );
BUFx6f_ASAP7_75t_L g493 ( .A(n_390), .Y(n_493) );
BUFx2_ASAP7_75t_L g793 ( .A(n_390), .Y(n_793) );
INVx5_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g518 ( .A(n_391), .Y(n_518) );
INVx2_ASAP7_75t_L g587 ( .A(n_391), .Y(n_587) );
INVx3_ASAP7_75t_L g616 ( .A(n_391), .Y(n_616) );
INVx4_ASAP7_75t_L g712 ( .A(n_391), .Y(n_712) );
INVx8_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_395), .Y(n_392) );
NAND2xp5_ASAP7_75t_SL g692 ( .A(n_393), .B(n_395), .Y(n_692) );
INVx1_ASAP7_75t_L g429 ( .A(n_394), .Y(n_429) );
NAND2x1p5_ASAP7_75t_L g417 ( .A(n_395), .B(n_410), .Y(n_417) );
AND2x6_ASAP7_75t_L g508 ( .A(n_395), .B(n_410), .Y(n_508) );
BUFx4f_ASAP7_75t_SL g494 ( .A(n_396), .Y(n_494) );
BUFx2_ASAP7_75t_L g519 ( .A(n_396), .Y(n_519) );
BUFx2_ASAP7_75t_L g713 ( .A(n_396), .Y(n_713) );
INVx6_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g618 ( .A(n_397), .Y(n_618) );
INVx1_ASAP7_75t_L g794 ( .A(n_397), .Y(n_794) );
INVx1_ASAP7_75t_SL g879 ( .A(n_397), .Y(n_879) );
OR2x6_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
INVx1_ASAP7_75t_L g425 ( .A(n_398), .Y(n_425) );
INVx1_ASAP7_75t_L g413 ( .A(n_399), .Y(n_413) );
AND2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_407), .Y(n_400) );
INVx3_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g562 ( .A(n_403), .Y(n_562) );
INVx2_ASAP7_75t_L g577 ( .A(n_403), .Y(n_577) );
INVx2_ASAP7_75t_L g650 ( .A(n_403), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g925 ( .A1(n_403), .A2(n_926), .B1(n_927), .B2(n_928), .Y(n_925) );
INVx6_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx3_ASAP7_75t_L g526 ( .A(n_404), .Y(n_526) );
BUFx3_ASAP7_75t_L g786 ( .A(n_404), .Y(n_786) );
BUFx3_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx3_ASAP7_75t_L g481 ( .A(n_406), .Y(n_481) );
BUFx3_ASAP7_75t_L g566 ( .A(n_406), .Y(n_566) );
BUFx3_ASAP7_75t_L g620 ( .A(n_406), .Y(n_620) );
BUFx2_ASAP7_75t_L g491 ( .A(n_408), .Y(n_491) );
BUFx3_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx3_ASAP7_75t_L g516 ( .A(n_409), .Y(n_516) );
INVx2_ASAP7_75t_L g557 ( .A(n_409), .Y(n_557) );
BUFx3_ASAP7_75t_L g585 ( .A(n_409), .Y(n_585) );
BUFx6f_ASAP7_75t_L g654 ( .A(n_409), .Y(n_654) );
INVx1_ASAP7_75t_L g450 ( .A(n_410), .Y(n_450) );
BUFx3_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx3_ASAP7_75t_L g484 ( .A(n_412), .Y(n_484) );
BUFx3_ASAP7_75t_L g522 ( .A(n_412), .Y(n_522) );
BUFx2_ASAP7_75t_L g622 ( .A(n_412), .Y(n_622) );
BUFx2_ASAP7_75t_SL g645 ( .A(n_412), .Y(n_645) );
BUFx3_ASAP7_75t_L g804 ( .A(n_412), .Y(n_804) );
INVx1_ASAP7_75t_L g848 ( .A(n_412), .Y(n_848) );
BUFx2_ASAP7_75t_SL g973 ( .A(n_412), .Y(n_973) );
AND2x2_ASAP7_75t_L g805 ( .A(n_413), .B(n_470), .Y(n_805) );
OA211x2_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_416), .B(n_418), .C(n_422), .Y(n_414) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_416), .A2(n_537), .B1(n_538), .B2(n_540), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_416), .A2(n_630), .B1(n_631), .B2(n_632), .Y(n_629) );
INVx2_ASAP7_75t_L g771 ( .A(n_416), .Y(n_771) );
OAI22xp5_ASAP7_75t_L g831 ( .A1(n_416), .A2(n_469), .B1(n_832), .B2(n_833), .Y(n_831) );
BUFx3_ASAP7_75t_L g1040 ( .A(n_416), .Y(n_1040) );
BUFx3_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g453 ( .A(n_417), .Y(n_453) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g510 ( .A(n_420), .Y(n_510) );
INVx2_ASAP7_75t_L g580 ( .A(n_420), .Y(n_580) );
INVx5_ASAP7_75t_L g667 ( .A(n_420), .Y(n_667) );
INVx4_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx3_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
BUFx2_ASAP7_75t_L g582 ( .A(n_424), .Y(n_582) );
BUFx2_ASAP7_75t_L g721 ( .A(n_424), .Y(n_721) );
INVx1_ASAP7_75t_L g969 ( .A(n_424), .Y(n_969) );
AND2x4_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
AND2x4_ASAP7_75t_L g435 ( .A(n_426), .B(n_436), .Y(n_435) );
AND2x4_ASAP7_75t_L g439 ( .A(n_426), .B(n_440), .Y(n_439) );
NAND2x1p5_ASAP7_75t_L g469 ( .A(n_426), .B(n_470), .Y(n_469) );
INVx1_ASAP7_75t_SL g869 ( .A(n_427), .Y(n_869) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx3_ASAP7_75t_L g512 ( .A(n_428), .Y(n_512) );
BUFx2_ASAP7_75t_SL g613 ( .A(n_428), .Y(n_613) );
BUFx2_ASAP7_75t_SL g663 ( .A(n_428), .Y(n_663) );
AND2x4_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx1_ASAP7_75t_L g475 ( .A(n_429), .Y(n_475) );
INVx1_ASAP7_75t_L g474 ( .A(n_430), .Y(n_474) );
INVx2_ASAP7_75t_SL g455 ( .A(n_432), .Y(n_455) );
INVx2_ASAP7_75t_L g752 ( .A(n_432), .Y(n_752) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g502 ( .A(n_433), .Y(n_502) );
INVx4_ASAP7_75t_L g590 ( .A(n_433), .Y(n_590) );
BUFx3_ASAP7_75t_L g723 ( .A(n_433), .Y(n_723) );
INVx2_ASAP7_75t_L g810 ( .A(n_433), .Y(n_810) );
INVx2_ASAP7_75t_SL g836 ( .A(n_433), .Y(n_836) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_434), .Y(n_750) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_435), .Y(n_460) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_435), .Y(n_609) );
BUFx4f_ASAP7_75t_SL g639 ( .A(n_435), .Y(n_639) );
BUFx2_ASAP7_75t_L g946 ( .A(n_435), .Y(n_946) );
INVx1_ASAP7_75t_L g440 ( .A(n_437), .Y(n_440) );
INVx2_ASAP7_75t_L g592 ( .A(n_438), .Y(n_592) );
BUFx4f_ASAP7_75t_SL g724 ( .A(n_438), .Y(n_724) );
BUFx12f_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_439), .Y(n_464) );
BUFx6f_ASAP7_75t_L g865 ( .A(n_439), .Y(n_865) );
INVx2_ASAP7_75t_SL g529 ( .A(n_442), .Y(n_529) );
OA22x2_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_497), .B1(n_498), .B2(n_528), .Y(n_442) );
INVx1_ASAP7_75t_L g528 ( .A(n_443), .Y(n_528) );
INVx2_ASAP7_75t_SL g495 ( .A(n_444), .Y(n_495) );
AND2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_476), .Y(n_444) );
NOR3xp33_ASAP7_75t_L g445 ( .A(n_446), .B(n_454), .C(n_465), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_448), .B1(n_451), .B2(n_452), .Y(n_446) );
OAI21xp5_ASAP7_75t_SL g1017 ( .A1(n_448), .A2(n_1018), .B(n_1019), .Y(n_1017) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g539 ( .A(n_449), .Y(n_539) );
OAI21xp5_ASAP7_75t_L g828 ( .A1(n_449), .A2(n_829), .B(n_830), .Y(n_828) );
INVx1_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g748 ( .A(n_453), .Y(n_748) );
OAI221xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_456), .B1(n_457), .B2(n_461), .C(n_462), .Y(n_454) );
OAI222xp33_ASAP7_75t_L g541 ( .A1(n_455), .A2(n_459), .B1(n_542), .B2(n_543), .C1(n_544), .C2(n_545), .Y(n_541) );
OAI21xp33_ASAP7_75t_L g633 ( .A1(n_455), .A2(n_634), .B(n_635), .Y(n_633) );
OAI221xp5_ASAP7_75t_L g772 ( .A1(n_457), .A2(n_773), .B1(n_774), .B2(n_775), .C(n_776), .Y(n_772) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g834 ( .A1(n_459), .A2(n_835), .B1(n_836), .B2(n_837), .Y(n_834) );
INVx4_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
BUFx2_ASAP7_75t_L g864 ( .A(n_460), .Y(n_864) );
INVx2_ASAP7_75t_L g1022 ( .A(n_460), .Y(n_1022) );
INVx2_ASAP7_75t_L g754 ( .A(n_463), .Y(n_754) );
BUFx3_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g544 ( .A(n_464), .Y(n_544) );
OAI22xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_467), .B1(n_471), .B2(n_472), .Y(n_465) );
OAI22xp5_ASAP7_75t_SL g1014 ( .A1(n_467), .A2(n_748), .B1(n_1015), .B2(n_1016), .Y(n_1014) );
INVx3_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g949 ( .A(n_468), .Y(n_949) );
INVx4_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_469), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_469), .A2(n_550), .B1(n_698), .B2(n_699), .Y(n_697) );
BUFx3_ASAP7_75t_L g758 ( .A(n_469), .Y(n_758) );
OAI22xp5_ASAP7_75t_L g777 ( .A1(n_472), .A2(n_758), .B1(n_778), .B2(n_779), .Y(n_777) );
BUFx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
CKINVDCx16_ASAP7_75t_R g551 ( .A(n_473), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g947 ( .A1(n_473), .A2(n_948), .B1(n_949), .B2(n_950), .Y(n_947) );
OR2x6_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_477), .B(n_487), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_485), .Y(n_477) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
BUFx4f_ASAP7_75t_SL g644 ( .A(n_481), .Y(n_644) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OAI221xp5_ASAP7_75t_SL g731 ( .A1(n_483), .A2(n_525), .B1(n_732), .B2(n_733), .C(n_734), .Y(n_731) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_484), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_488), .B(n_492), .Y(n_487) );
BUFx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx3_ASAP7_75t_L g555 ( .A(n_490), .Y(n_555) );
BUFx6f_ASAP7_75t_L g647 ( .A(n_490), .Y(n_647) );
INVx3_ASAP7_75t_L g737 ( .A(n_490), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g694 ( .A(n_494), .Y(n_694) );
AO22x2_ASAP7_75t_L g570 ( .A1(n_497), .A2(n_498), .B1(n_571), .B2(n_572), .Y(n_570) );
INVx4_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
XOR2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_527), .Y(n_498) );
NAND3x1_ASAP7_75t_L g499 ( .A(n_500), .B(n_513), .C(n_520), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_501), .B(n_505), .Y(n_500) );
OAI21xp5_ASAP7_75t_SL g501 ( .A1(n_502), .A2(n_503), .B(n_504), .Y(n_501) );
OAI21xp5_ASAP7_75t_L g610 ( .A1(n_502), .A2(n_611), .B(n_612), .Y(n_610) );
OAI21xp5_ASAP7_75t_L g660 ( .A1(n_502), .A2(n_661), .B(n_662), .Y(n_660) );
OAI21xp5_ASAP7_75t_SL g894 ( .A1(n_502), .A2(n_895), .B(n_896), .Y(n_894) );
OAI21xp5_ASAP7_75t_SL g961 ( .A1(n_502), .A2(n_962), .B(n_963), .Y(n_961) );
NAND3xp33_ASAP7_75t_L g505 ( .A(n_506), .B(n_509), .C(n_511), .Y(n_505) );
BUFx4f_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx2_ASAP7_75t_L g719 ( .A(n_508), .Y(n_719) );
INVx1_ASAP7_75t_SL g872 ( .A(n_508), .Y(n_872) );
BUFx2_ASAP7_75t_L g891 ( .A(n_508), .Y(n_891) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_517), .Y(n_513) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_523), .Y(n_520) );
INVx1_ASAP7_75t_L g927 ( .A(n_524), .Y(n_927) );
INVx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_SL g561 ( .A(n_525), .Y(n_561) );
INVx4_ASAP7_75t_L g882 ( .A(n_525), .Y(n_882) );
INVx3_ASAP7_75t_L g595 ( .A(n_530), .Y(n_595) );
BUFx3_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .B1(n_569), .B2(n_570), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g568 ( .A(n_534), .Y(n_568) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_552), .Y(n_534) );
NOR3xp33_ASAP7_75t_L g535 ( .A(n_536), .B(n_541), .C(n_546), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g939 ( .A1(n_538), .A2(n_748), .B1(n_940), .B2(n_941), .Y(n_939) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_SL g631 ( .A(n_539), .Y(n_631) );
INVx2_ASAP7_75t_L g746 ( .A(n_539), .Y(n_746) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_548), .B1(n_549), .B2(n_550), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_548), .A2(n_637), .B1(n_638), .B2(n_640), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_550), .A2(n_757), .B1(n_758), .B2(n_759), .Y(n_756) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_553), .B(n_559), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_558), .Y(n_553) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
OAI21xp5_ASAP7_75t_SL g839 ( .A1(n_557), .A2(n_840), .B(n_841), .Y(n_839) );
INVx2_ASAP7_75t_L g875 ( .A(n_557), .Y(n_875) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_560), .B(n_563), .Y(n_559) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
XOR2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_593), .Y(n_572) );
NAND4xp75_ASAP7_75t_L g573 ( .A(n_574), .B(n_578), .C(n_583), .D(n_588), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
AND2x2_ASAP7_75t_SL g578 ( .A(n_579), .B(n_581), .Y(n_578) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_586), .Y(n_583) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_585), .Y(n_740) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_587), .Y(n_735) );
INVx4_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
BUFx2_ASAP7_75t_L g773 ( .A(n_590), .Y(n_773) );
OAI22xp5_ASAP7_75t_SL g1020 ( .A1(n_590), .A2(n_1021), .B1(n_1022), .B2(n_1023), .Y(n_1020) );
INVx1_ASAP7_75t_L g920 ( .A(n_591), .Y(n_920) );
INVx3_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g987 ( .A(n_596), .Y(n_987) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_820), .B1(n_985), .B2(n_986), .Y(n_596) );
INVx1_ASAP7_75t_L g985 ( .A(n_597), .Y(n_985) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_599), .B1(n_677), .B2(n_819), .Y(n_597) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
OA22x2_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B1(n_624), .B2(n_676), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
XOR2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_623), .Y(n_602) );
NAND4xp75_ASAP7_75t_SL g603 ( .A(n_604), .B(n_614), .C(n_619), .D(n_621), .Y(n_603) );
NOR2xp67_ASAP7_75t_SL g604 ( .A(n_605), .B(n_610), .Y(n_604) );
NAND3xp33_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .C(n_608), .Y(n_605) );
INVx1_ASAP7_75t_L g918 ( .A(n_609), .Y(n_918) );
BUFx6f_ASAP7_75t_L g964 ( .A(n_609), .Y(n_964) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_617), .Y(n_614) );
BUFx2_ASAP7_75t_L g688 ( .A(n_620), .Y(n_688) );
INVx1_ASAP7_75t_L g709 ( .A(n_620), .Y(n_709) );
INVx1_ASAP7_75t_L g676 ( .A(n_624), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_626), .B1(n_656), .B2(n_657), .Y(n_624) );
INVx1_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
XNOR2x1_ASAP7_75t_L g626 ( .A(n_627), .B(n_655), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_641), .Y(n_627) );
NOR3xp33_ASAP7_75t_L g628 ( .A(n_629), .B(n_633), .C(n_636), .Y(n_628) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_642), .B(n_648), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_646), .Y(n_642) );
INVx1_ASAP7_75t_SL g931 ( .A(n_647), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_651), .Y(n_648) );
INVx3_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx4_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx3_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
XOR2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_675), .Y(n_657) );
NAND2xp5_ASAP7_75t_SL g658 ( .A(n_659), .B(n_668), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_660), .B(n_664), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
BUFx6f_ASAP7_75t_L g696 ( .A(n_667), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_669), .B(n_672), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
INVx1_ASAP7_75t_L g819 ( .A(n_677), .Y(n_819) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_726), .B1(n_817), .B2(n_818), .Y(n_677) );
INVx1_ASAP7_75t_L g817 ( .A(n_678), .Y(n_817) );
OAI22xp5_ASAP7_75t_SL g678 ( .A1(n_679), .A2(n_680), .B1(n_702), .B2(n_703), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AND4x1_ASAP7_75t_L g683 ( .A(n_684), .B(n_687), .C(n_695), .D(n_700), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_691), .B1(n_693), .B2(n_694), .Y(n_689) );
BUFx2_ASAP7_75t_R g691 ( .A(n_692), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g846 ( .A1(n_692), .A2(n_847), .B1(n_848), .B2(n_849), .Y(n_846) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_SL g725 ( .A(n_705), .Y(n_725) );
NAND4xp75_ASAP7_75t_L g705 ( .A(n_706), .B(n_714), .C(n_717), .D(n_722), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_710), .Y(n_706) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
BUFx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g878 ( .A(n_712), .Y(n_878) );
AND2x2_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
AND2x2_ASAP7_75t_SL g717 ( .A(n_718), .B(n_720), .Y(n_717) );
INVx3_ASAP7_75t_L g944 ( .A(n_723), .Y(n_944) );
INVx1_ASAP7_75t_L g818 ( .A(n_726), .Y(n_818) );
XOR2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_762), .Y(n_726) );
BUFx3_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g761 ( .A(n_729), .Y(n_761) );
AND2x2_ASAP7_75t_SL g729 ( .A(n_730), .B(n_743), .Y(n_729) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_731), .B(n_736), .Y(n_730) );
OAI221xp5_ASAP7_75t_SL g736 ( .A1(n_737), .A2(n_738), .B1(n_739), .B2(n_741), .C(n_742), .Y(n_736) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
NOR3xp33_ASAP7_75t_L g743 ( .A(n_744), .B(n_749), .C(n_756), .Y(n_743) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_746), .B1(n_747), .B2(n_748), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_746), .A2(n_768), .B1(n_769), .B2(n_770), .Y(n_767) );
OAI222xp33_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_751), .B1(n_752), .B2(n_753), .C1(n_754), .C2(n_755), .Y(n_749) );
OAI21xp5_ASAP7_75t_SL g861 ( .A1(n_752), .A2(n_862), .B(n_863), .Y(n_861) );
OAI22xp5_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_796), .B1(n_797), .B2(n_816), .Y(n_762) );
INVx1_ASAP7_75t_L g816 ( .A(n_763), .Y(n_816) );
INVx1_ASAP7_75t_L g795 ( .A(n_765), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_766), .B(n_780), .Y(n_765) );
NOR3xp33_ASAP7_75t_L g766 ( .A(n_767), .B(n_772), .C(n_777), .Y(n_766) );
OAI211xp5_ASAP7_75t_L g912 ( .A1(n_770), .A2(n_913), .B(n_914), .C(n_915), .Y(n_912) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
NOR2xp67_ASAP7_75t_L g780 ( .A(n_781), .B(n_787), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_782), .B(n_783), .Y(n_781) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_788), .B(n_792), .Y(n_787) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx2_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
XOR2x2_ASAP7_75t_L g856 ( .A(n_797), .B(n_857), .Y(n_856) );
XOR2x2_ASAP7_75t_L g797 ( .A(n_798), .B(n_815), .Y(n_797) );
NAND4xp75_ASAP7_75t_SL g798 ( .A(n_799), .B(n_800), .C(n_802), .D(n_807), .Y(n_798) );
AND2x2_ASAP7_75t_L g802 ( .A(n_803), .B(n_806), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g807 ( .A(n_808), .B(n_812), .Y(n_807) );
OAI21xp5_ASAP7_75t_L g808 ( .A1(n_809), .A2(n_810), .B(n_811), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .Y(n_812) );
INVx1_ASAP7_75t_L g986 ( .A(n_820), .Y(n_986) );
AOI22xp5_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_884), .B1(n_983), .B2(n_984), .Y(n_820) );
INVx1_ASAP7_75t_SL g983 ( .A(n_821), .Y(n_983) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
XNOR2xp5_ASAP7_75t_L g823 ( .A(n_824), .B(n_856), .Y(n_823) );
BUFx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
XNOR2x1_ASAP7_75t_L g825 ( .A(n_826), .B(n_855), .Y(n_825) );
AND3x2_ASAP7_75t_L g826 ( .A(n_827), .B(n_838), .C(n_845), .Y(n_826) );
NOR3xp33_ASAP7_75t_L g827 ( .A(n_828), .B(n_831), .C(n_834), .Y(n_827) );
NOR2xp33_ASAP7_75t_L g838 ( .A(n_839), .B(n_842), .Y(n_838) );
NOR3xp33_ASAP7_75t_L g845 ( .A(n_846), .B(n_850), .C(n_853), .Y(n_845) );
NOR2xp33_ASAP7_75t_L g850 ( .A(n_851), .B(n_852), .Y(n_850) );
INVx1_ASAP7_75t_L g934 ( .A(n_852), .Y(n_934) );
XNOR2xp5_ASAP7_75t_L g857 ( .A(n_858), .B(n_859), .Y(n_857) );
NAND3xp33_ASAP7_75t_L g859 ( .A(n_860), .B(n_873), .C(n_880), .Y(n_859) );
NOR2xp33_ASAP7_75t_L g860 ( .A(n_861), .B(n_866), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_867), .B(n_870), .Y(n_866) );
INVx2_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx1_ASAP7_75t_SL g871 ( .A(n_872), .Y(n_871) );
AND2x2_ASAP7_75t_L g873 ( .A(n_874), .B(n_876), .Y(n_873) );
INVx3_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
AND2x2_ASAP7_75t_L g880 ( .A(n_881), .B(n_883), .Y(n_880) );
INVx1_ASAP7_75t_L g984 ( .A(n_884), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_885), .A2(n_886), .B1(n_905), .B2(n_982), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
XOR2x2_ASAP7_75t_SL g886 ( .A(n_887), .B(n_904), .Y(n_886) );
NAND2x1p5_ASAP7_75t_L g887 ( .A(n_888), .B(n_897), .Y(n_887) );
NOR2xp33_ASAP7_75t_L g888 ( .A(n_889), .B(n_894), .Y(n_888) );
NAND3xp33_ASAP7_75t_L g889 ( .A(n_890), .B(n_892), .C(n_893), .Y(n_889) );
NOR2x1_ASAP7_75t_L g897 ( .A(n_898), .B(n_901), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_899), .B(n_900), .Y(n_898) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_902), .B(n_903), .Y(n_901) );
INVx2_ASAP7_75t_SL g982 ( .A(n_905), .Y(n_982) );
AOI22xp5_ASAP7_75t_L g905 ( .A1(n_906), .A2(n_907), .B1(n_935), .B2(n_981), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
INVx2_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
XNOR2xp5_ASAP7_75t_L g908 ( .A(n_909), .B(n_910), .Y(n_908) );
AND2x2_ASAP7_75t_L g910 ( .A(n_911), .B(n_921), .Y(n_910) );
OAI22xp5_ASAP7_75t_L g916 ( .A1(n_917), .A2(n_918), .B1(n_919), .B2(n_920), .Y(n_916) );
NOR3xp33_ASAP7_75t_L g921 ( .A(n_922), .B(n_925), .C(n_929), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_923), .B(n_924), .Y(n_922) );
OAI22xp5_ASAP7_75t_L g929 ( .A1(n_930), .A2(n_931), .B1(n_932), .B2(n_933), .Y(n_929) );
INVx1_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
INVx2_ASAP7_75t_L g981 ( .A(n_935), .Y(n_981) );
XNOR2x2_ASAP7_75t_L g935 ( .A(n_936), .B(n_958), .Y(n_935) );
INVx1_ASAP7_75t_SL g956 ( .A(n_937), .Y(n_956) );
AND2x2_ASAP7_75t_SL g937 ( .A(n_938), .B(n_951), .Y(n_937) );
NOR3xp33_ASAP7_75t_L g938 ( .A(n_939), .B(n_942), .C(n_947), .Y(n_938) );
OAI21xp33_ASAP7_75t_L g942 ( .A1(n_943), .A2(n_944), .B(n_945), .Y(n_942) );
AND4x1_ASAP7_75t_L g951 ( .A(n_952), .B(n_953), .C(n_954), .D(n_955), .Y(n_951) );
INVx2_ASAP7_75t_SL g979 ( .A(n_959), .Y(n_979) );
AND2x2_ASAP7_75t_L g959 ( .A(n_960), .B(n_970), .Y(n_959) );
NOR2xp33_ASAP7_75t_L g960 ( .A(n_961), .B(n_965), .Y(n_960) );
NAND2xp5_ASAP7_75t_SL g965 ( .A(n_966), .B(n_967), .Y(n_965) );
INVx1_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
NOR2xp33_ASAP7_75t_L g970 ( .A(n_971), .B(n_976), .Y(n_970) );
NAND2xp5_ASAP7_75t_L g971 ( .A(n_972), .B(n_974), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g976 ( .A(n_977), .B(n_978), .Y(n_976) );
INVx1_ASAP7_75t_SL g989 ( .A(n_990), .Y(n_989) );
NOR2x1_ASAP7_75t_L g990 ( .A(n_991), .B(n_995), .Y(n_990) );
OR2x2_ASAP7_75t_SL g1049 ( .A(n_991), .B(n_996), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g991 ( .A(n_992), .B(n_994), .Y(n_991) );
CKINVDCx20_ASAP7_75t_R g1025 ( .A(n_992), .Y(n_1025) );
INVx1_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
NAND2xp5_ASAP7_75t_L g1031 ( .A(n_993), .B(n_1029), .Y(n_1031) );
CKINVDCx16_ASAP7_75t_R g1029 ( .A(n_994), .Y(n_1029) );
CKINVDCx20_ASAP7_75t_R g995 ( .A(n_996), .Y(n_995) );
NAND2xp5_ASAP7_75t_L g996 ( .A(n_997), .B(n_998), .Y(n_996) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1001), .Y(n_999) );
OAI322xp33_ASAP7_75t_L g1002 ( .A1(n_1003), .A2(n_1024), .A3(n_1026), .B1(n_1030), .B2(n_1032), .C1(n_1033), .C2(n_1047), .Y(n_1002) );
CKINVDCx20_ASAP7_75t_R g1004 ( .A(n_1005), .Y(n_1004) );
HB1xp67_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
NAND3x1_ASAP7_75t_SL g1006 ( .A(n_1007), .B(n_1010), .C(n_1013), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1009), .Y(n_1007) );
AND2x2_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1012), .Y(n_1010) );
NOR3xp33_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1017), .C(n_1020), .Y(n_1013) );
HB1xp67_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
HB1xp67_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
HB1xp67_ASAP7_75t_L g1027 ( .A(n_1028), .Y(n_1027) );
INVx1_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
XOR2x2_ASAP7_75t_L g1033 ( .A(n_1032), .B(n_1034), .Y(n_1033) );
NAND4xp75_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1038), .C(n_1043), .D(n_1046), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_1036), .B(n_1037), .Y(n_1035) );
OA211x2_ASAP7_75t_L g1038 ( .A1(n_1039), .A2(n_1040), .B(n_1041), .C(n_1042), .Y(n_1038) );
AND2x2_ASAP7_75t_L g1043 ( .A(n_1044), .B(n_1045), .Y(n_1043) );
CKINVDCx20_ASAP7_75t_R g1047 ( .A(n_1048), .Y(n_1047) );
CKINVDCx20_ASAP7_75t_R g1048 ( .A(n_1049), .Y(n_1048) );
endmodule