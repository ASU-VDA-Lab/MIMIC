module fake_jpeg_3399_n_204 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_204);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_2),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_25),
.B(n_45),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_4),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_20),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_23),
.Y(n_71)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

BUFx4f_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_64),
.Y(n_73)
);

CKINVDCx6p67_ASAP7_75t_R g83 ( 
.A(n_73),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_0),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_79),
.Y(n_93)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g91 ( 
.A(n_75),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_53),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_81),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_60),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_79),
.B(n_52),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_85),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_61),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_72),
.A2(n_63),
.B1(n_55),
.B2(n_56),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_86),
.A2(n_89),
.B1(n_75),
.B2(n_76),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_69),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_58),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_76),
.A2(n_68),
.B1(n_57),
.B2(n_65),
.Y(n_89)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

XNOR2x1_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_62),
.Y(n_96)
);

MAJx2_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_108),
.C(n_72),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_102),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_73),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_99),
.Y(n_130)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_71),
.Y(n_102)
);

BUFx4f_ASAP7_75t_SL g103 ( 
.A(n_88),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_103),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_89),
.B(n_59),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_104),
.B(n_112),
.Y(n_122)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_107),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_73),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_48),
.Y(n_108)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_110),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_70),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_111),
.A2(n_67),
.B1(n_65),
.B2(n_68),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_90),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_101),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_115),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_54),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_118),
.A2(n_123),
.B1(n_24),
.B2(n_46),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_111),
.A2(n_77),
.B1(n_90),
.B2(n_75),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_92),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_129),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_49),
.B(n_50),
.C(n_2),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_126),
.B(n_127),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_95),
.B(n_0),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_49),
.B(n_50),
.C(n_4),
.Y(n_128)
);

NOR3xp33_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_3),
.C(n_5),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_107),
.B(n_1),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_21),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_77),
.B1(n_92),
.B2(n_56),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_132),
.A2(n_47),
.B1(n_27),
.B2(n_29),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_125),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_135),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_67),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_133),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_144),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_130),
.A2(n_109),
.B(n_103),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_137),
.A2(n_148),
.B(n_154),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_138),
.A2(n_145),
.B1(n_140),
.B2(n_149),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_128),
.A2(n_3),
.B(n_5),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_140),
.A2(n_12),
.B(n_13),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_118),
.A2(n_123),
.B1(n_122),
.B2(n_124),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_11),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_9),
.Y(n_168)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_6),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_150),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_116),
.A2(n_6),
.B(n_7),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_120),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_8),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_152),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_131),
.A2(n_9),
.B(n_11),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_125),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_157),
.Y(n_174)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_121),
.Y(n_156)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_125),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_152),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_167),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_137),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_15),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_142),
.Y(n_169)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_169),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_170),
.A2(n_145),
.B1(n_148),
.B2(n_154),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_171),
.A2(n_138),
.B1(n_141),
.B2(n_16),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_172),
.A2(n_14),
.B(n_15),
.Y(n_182)
);

NOR3xp33_ASAP7_75t_SL g173 ( 
.A(n_139),
.B(n_32),
.C(n_40),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_173),
.B(n_175),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_143),
.B(n_44),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_17),
.C(n_19),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_180),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_178),
.A2(n_158),
.B1(n_165),
.B2(n_174),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_31),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_183),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_182),
.A2(n_184),
.B(n_172),
.Y(n_190)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_181),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_185),
.A2(n_191),
.B1(n_166),
.B2(n_159),
.Y(n_195)
);

XNOR2x2_ASAP7_75t_SL g186 ( 
.A(n_177),
.B(n_170),
.Y(n_186)
);

OAI21x1_ASAP7_75t_L g192 ( 
.A1(n_186),
.A2(n_164),
.B(n_162),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_189),
.B(n_161),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_190),
.A2(n_161),
.B(n_184),
.Y(n_194)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_179),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_193),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_188),
.Y(n_198)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_195),
.Y(n_196)
);

OAI221xp5_ASAP7_75t_L g199 ( 
.A1(n_198),
.A2(n_188),
.B1(n_173),
.B2(n_187),
.C(n_183),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_199),
.B(n_200),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_168),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_196),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_30),
.C(n_34),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_35),
.Y(n_204)
);


endmodule