module fake_jpeg_31744_n_49 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_49);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_49;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_5),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx6_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_4),
.B(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_0),
.B(n_2),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_13),
.B(n_0),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_19),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_10),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_1),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_20),
.A2(n_10),
.B1(n_14),
.B2(n_7),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_5),
.Y(n_21)
);

A2O1A1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_21),
.A2(n_8),
.B(n_12),
.C(n_6),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_22),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_28),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_15),
.A2(n_9),
.B1(n_8),
.B2(n_12),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_26),
.A2(n_19),
.B1(n_18),
.B2(n_9),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_18),
.A2(n_9),
.B1(n_2),
.B2(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_30),
.B(n_25),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_35),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_22),
.A2(n_17),
.B1(n_16),
.B2(n_20),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_36),
.B1(n_16),
.B2(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_SL g37 ( 
.A(n_32),
.B(n_29),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_1),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_38),
.A2(n_40),
.B1(n_36),
.B2(n_35),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_39),
.A2(n_34),
.B1(n_31),
.B2(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_43),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_43),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_44),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_37),
.C(n_44),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_48),
.A2(n_41),
.B(n_3),
.Y(n_49)
);


endmodule