module fake_jpeg_16225_n_301 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_301);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_301;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_259;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

INVx3_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx2_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_9),
.B(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_35),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_32),
.A2(n_15),
.B1(n_24),
.B2(n_17),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_40),
.A2(n_45),
.B1(n_50),
.B2(n_29),
.Y(n_76)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_41),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_20),
.C(n_17),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_49),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_33),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_32),
.A2(n_15),
.B1(n_24),
.B2(n_22),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_34),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_29),
.Y(n_82)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_36),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_72),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_47),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_60),
.B(n_61),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_51),
.Y(n_62)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_50),
.Y(n_63)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_15),
.B1(n_36),
.B2(n_24),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_64),
.A2(n_76),
.B1(n_80),
.B2(n_23),
.Y(n_103)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_24),
.B1(n_19),
.B2(n_28),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_66),
.A2(n_74),
.B1(n_22),
.B2(n_18),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_68),
.Y(n_100)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_45),
.A2(n_27),
.B(n_19),
.C(n_25),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_53),
.A2(n_21),
.B1(n_22),
.B2(n_16),
.Y(n_74)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_75),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_39),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_82),
.Y(n_95)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_48),
.A2(n_39),
.B1(n_29),
.B2(n_21),
.Y(n_80)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_79),
.A2(n_48),
.B1(n_18),
.B2(n_21),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_38),
.C(n_37),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_84),
.B(n_93),
.C(n_52),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_68),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_90),
.A2(n_70),
.B1(n_30),
.B2(n_23),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_38),
.C(n_37),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_70),
.Y(n_94)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_54),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_20),
.Y(n_133)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_103),
.B(n_89),
.Y(n_125)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_76),
.A2(n_25),
.B1(n_28),
.B2(n_41),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_110),
.A2(n_30),
.B1(n_27),
.B2(n_65),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_97),
.Y(n_111)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_107),
.A2(n_70),
.B1(n_81),
.B2(n_62),
.Y(n_112)
);

O2A1O1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_112),
.A2(n_114),
.B(n_122),
.C(n_67),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_113),
.A2(n_116),
.B1(n_125),
.B2(n_94),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_91),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_69),
.B1(n_55),
.B2(n_62),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_110),
.A2(n_72),
.B1(n_60),
.B2(n_56),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_SL g159 ( 
.A(n_118),
.B(n_123),
.C(n_133),
.Y(n_159)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_SL g121 ( 
.A1(n_89),
.A2(n_75),
.B(n_80),
.C(n_82),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_121),
.A2(n_20),
.B(n_1),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_88),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_67),
.Y(n_166)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_126),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_107),
.A2(n_61),
.B1(n_46),
.B2(n_43),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_127),
.A2(n_105),
.B1(n_67),
.B2(n_26),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_84),
.B(n_58),
.C(n_52),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_93),
.C(n_95),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_68),
.Y(n_129)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_86),
.A2(n_9),
.B1(n_10),
.B2(n_8),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_132),
.A2(n_134),
.B1(n_6),
.B2(n_14),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_86),
.A2(n_10),
.B1(n_7),
.B2(n_6),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_103),
.A2(n_17),
.B1(n_26),
.B2(n_14),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_135),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_85),
.Y(n_136)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_87),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_140),
.B(n_166),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_95),
.Y(n_141)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_141),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_142),
.B(n_148),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_83),
.Y(n_143)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_109),
.B(n_85),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_144),
.A2(n_145),
.B(n_146),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_109),
.Y(n_145)
);

OAI21x1_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_94),
.B(n_106),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_106),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_147),
.A2(n_149),
.B(n_155),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_130),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_104),
.B(n_98),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_88),
.Y(n_150)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_135),
.A2(n_105),
.B1(n_100),
.B2(n_96),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_112),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_154),
.B(n_162),
.Y(n_177)
);

OAI21xp33_ASAP7_75t_L g155 ( 
.A1(n_121),
.A2(n_26),
.B(n_98),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_112),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_108),
.Y(n_161)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_130),
.Y(n_162)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_164),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_165),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_119),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_168),
.B(n_169),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_112),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_126),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_170),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_122),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_171),
.B(n_179),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_174),
.A2(n_194),
.B(n_199),
.Y(n_210)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_176),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_114),
.Y(n_179)
);

OAI32xp33_ASAP7_75t_L g181 ( 
.A1(n_161),
.A2(n_121),
.A3(n_123),
.B1(n_115),
.B2(n_127),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_181),
.B(n_163),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_156),
.B(n_115),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_182),
.B(n_185),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_141),
.B(n_131),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_147),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_186),
.Y(n_207)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

INVx13_ASAP7_75t_L g209 ( 
.A(n_187),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_149),
.B(n_119),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_193),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_137),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_189),
.B(n_153),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_140),
.B(n_131),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_193),
.C(n_183),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_119),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_143),
.B(n_0),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_150),
.B(n_26),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_164),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_147),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_145),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_201),
.B(n_218),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_180),
.A2(n_160),
.B(n_144),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_203),
.A2(n_213),
.B(n_194),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_180),
.A2(n_169),
.B1(n_154),
.B2(n_138),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_204),
.A2(n_174),
.B1(n_198),
.B2(n_199),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_208),
.C(n_201),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_145),
.C(n_159),
.Y(n_208)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_188),
.A2(n_138),
.B(n_159),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_212),
.A2(n_194),
.B(n_178),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_192),
.A2(n_153),
.B(n_2),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_215),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_216),
.A2(n_198),
.B1(n_172),
.B2(n_178),
.Y(n_233)
);

MAJx2_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_14),
.C(n_13),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_173),
.B(n_1),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_219),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_173),
.B(n_1),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_219),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_175),
.B(n_177),
.Y(n_222)
);

OAI21xp33_ASAP7_75t_L g229 ( 
.A1(n_222),
.A2(n_172),
.B(n_190),
.Y(n_229)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_224),
.A2(n_238),
.B1(n_240),
.B2(n_213),
.Y(n_251)
);

XOR2x2_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_184),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_225),
.B(n_236),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_235),
.Y(n_246)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_228),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_200),
.C(n_196),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_231),
.Y(n_241)
);

FAx1_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_192),
.CI(n_181),
.CON(n_231),
.SN(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_176),
.Y(n_232)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_233),
.A2(n_205),
.B1(n_204),
.B2(n_218),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_212),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_202),
.A2(n_200),
.B1(n_197),
.B2(n_195),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_203),
.A2(n_195),
.B(n_197),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_234),
.A2(n_211),
.B1(n_207),
.B2(n_222),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_242),
.A2(n_243),
.B1(n_215),
.B2(n_237),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_225),
.A2(n_207),
.B1(n_216),
.B2(n_220),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_210),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_253),
.C(n_224),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_238),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_250),
.B(n_254),
.Y(n_264)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_251),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_239),
.B(n_217),
.Y(n_252)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_252),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_205),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_262),
.C(n_249),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_255),
.A2(n_226),
.B1(n_240),
.B2(n_231),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_258),
.A2(n_209),
.B1(n_187),
.B2(n_4),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_248),
.Y(n_259)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_259),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_242),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_261),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_226),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_241),
.A2(n_231),
.B(n_223),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_214),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_265),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_214),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_237),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_246),
.C(n_227),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_269),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_246),
.C(n_244),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_274),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_249),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_243),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_275),
.B(n_258),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_276),
.Y(n_281)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_277),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_284),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_271),
.A2(n_260),
.B1(n_264),
.B2(n_266),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_283),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_273),
.A2(n_259),
.B1(n_209),
.B2(n_10),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_269),
.A2(n_270),
.B1(n_276),
.B2(n_268),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_209),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_286),
.A2(n_290),
.B1(n_2),
.B2(n_3),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_11),
.C(n_13),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_287),
.A2(n_291),
.B(n_281),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_11),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_2),
.Y(n_291)
);

NOR2x1_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_278),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_292),
.A2(n_293),
.B1(n_294),
.B2(n_286),
.Y(n_295)
);

AOI21x1_ASAP7_75t_L g296 ( 
.A1(n_295),
.A2(n_289),
.B(n_3),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_296),
.B(n_2),
.Y(n_297)
);

OAI21xp33_ASAP7_75t_L g298 ( 
.A1(n_297),
.A2(n_4),
.B(n_5),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_4),
.C(n_5),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_4),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_300),
.B(n_5),
.Y(n_301)
);


endmodule