module fake_jpeg_4715_n_58 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_58);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_58;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

BUFx5_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_2),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

AND2x2_ASAP7_75t_L g13 ( 
.A(n_0),
.B(n_6),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

AND2x2_ASAP7_75t_SL g16 ( 
.A(n_5),
.B(n_1),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_18),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_16),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

AOI21xp33_ASAP7_75t_SL g20 ( 
.A1(n_16),
.A2(n_2),
.B(n_3),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_20),
.A2(n_11),
.B1(n_12),
.B2(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_26),
.B(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_21),
.C(n_20),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_31),
.C(n_11),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_32),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_28),
.C(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_34),
.B(n_35),
.Y(n_38)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_18),
.B(n_12),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_41),
.B(n_15),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_15),
.C(n_10),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_13),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_13),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_29),
.B(n_13),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_45),
.C(n_4),
.Y(n_49)
);

AOI221xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.C(n_14),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_44),
.A2(n_36),
.B1(n_5),
.B2(n_7),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_19),
.C(n_30),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx12f_ASAP7_75t_SL g50 ( 
.A(n_46),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_48),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_51),
.B(n_50),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_54),
.Y(n_55)
);

MAJx2_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_50),
.C(n_49),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_55),
.A2(n_52),
.B1(n_14),
.B2(n_30),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_8),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_14),
.Y(n_58)
);


endmodule