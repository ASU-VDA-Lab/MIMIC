module fake_ariane_2206_n_175 (n_8, n_24, n_7, n_22, n_43, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_41, n_38, n_2, n_18, n_32, n_28, n_37, n_9, n_11, n_34, n_26, n_3, n_14, n_0, n_36, n_33, n_19, n_30, n_39, n_40, n_31, n_42, n_16, n_5, n_12, n_15, n_21, n_23, n_35, n_10, n_25, n_175);

input n_8;
input n_24;
input n_7;
input n_22;
input n_43;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_41;
input n_38;
input n_2;
input n_18;
input n_32;
input n_28;
input n_37;
input n_9;
input n_11;
input n_34;
input n_26;
input n_3;
input n_14;
input n_0;
input n_36;
input n_33;
input n_19;
input n_30;
input n_39;
input n_40;
input n_31;
input n_42;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_35;
input n_10;
input n_25;

output n_175;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_160;
wire n_64;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_149;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_92;
wire n_143;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_91;
wire n_159;
wire n_107;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_82;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_48;
wire n_94;
wire n_101;
wire n_134;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_118;
wire n_93;
wire n_121;
wire n_61;
wire n_108;
wire n_102;
wire n_125;
wire n_168;
wire n_81;
wire n_87;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_63;
wire n_59;
wire n_99;
wire n_155;
wire n_127;
wire n_54;

OA21x2_ASAP7_75t_L g44 ( 
.A1(n_3),
.A2(n_15),
.B(n_36),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

AND2x4_ASAP7_75t_L g47 ( 
.A(n_19),
.B(n_34),
.Y(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_29),
.Y(n_48)
);

AND2x4_ASAP7_75t_L g49 ( 
.A(n_18),
.B(n_0),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_31),
.A2(n_41),
.B1(n_24),
.B2(n_30),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_0),
.B(n_43),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_13),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

AND2x4_ASAP7_75t_L g56 ( 
.A(n_25),
.B(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

OA21x2_ASAP7_75t_L g61 ( 
.A1(n_22),
.A2(n_14),
.B(n_1),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_4),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

OA21x2_ASAP7_75t_L g65 ( 
.A1(n_6),
.A2(n_38),
.B(n_8),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_20),
.B(n_28),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_27),
.Y(n_69)
);

CKINVDCx8_ASAP7_75t_R g70 ( 
.A(n_5),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_4),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_11),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_16),
.B(n_2),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_5),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_68),
.B1(n_74),
.B2(n_49),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_2),
.Y(n_77)
);

OR2x6_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_17),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_49),
.A2(n_59),
.B1(n_71),
.B2(n_61),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_33),
.Y(n_82)
);

CKINVDCx5p33_ASAP7_75t_R g83 ( 
.A(n_48),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

AND2x4_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_67),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_60),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_62),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_52),
.A2(n_67),
.B(n_50),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

AND2x6_ASAP7_75t_SL g95 ( 
.A(n_73),
.B(n_69),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_45),
.B(n_58),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_54),
.A2(n_51),
.B1(n_53),
.B2(n_47),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_45),
.B(n_58),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_56),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

NAND3xp33_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_56),
.C(n_61),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_103),
.Y(n_107)
);

AO32x2_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_61),
.A3(n_44),
.B1(n_65),
.B2(n_54),
.Y(n_108)
);

OAI21x1_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_102),
.B(n_82),
.Y(n_109)
);

AND3x2_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_69),
.C(n_66),
.Y(n_110)
);

AOI21x1_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_66),
.B(n_44),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_83),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_64),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_64),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_81),
.A2(n_44),
.B(n_65),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_81),
.A2(n_65),
.B(n_87),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_96),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_99),
.A2(n_85),
.B(n_103),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_95),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_76),
.A2(n_99),
.B(n_97),
.C(n_75),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_98),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_98),
.Y(n_126)
);

OA21x2_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_100),
.B(n_101),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

AO21x2_ASAP7_75t_L g131 ( 
.A1(n_116),
.A2(n_80),
.B(n_86),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_106),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

HB1xp67_ASAP7_75t_SL g137 ( 
.A(n_123),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

AOI33xp33_ASAP7_75t_L g139 ( 
.A1(n_126),
.A2(n_110),
.A3(n_133),
.B1(n_138),
.B2(n_124),
.B3(n_137),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_125),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_121),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_134),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

AND2x4_ASAP7_75t_SL g145 ( 
.A(n_133),
.B(n_78),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_143),
.B(n_135),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_146),
.Y(n_149)
);

AOI222xp33_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_134),
.B1(n_145),
.B2(n_105),
.C1(n_144),
.C2(n_140),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_146),
.B(n_130),
.Y(n_151)
);

NOR2x1_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_130),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_128),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_115),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_147),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_151),
.A2(n_124),
.B(n_117),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_151),
.B(n_150),
.Y(n_157)
);

AOI21xp33_ASAP7_75t_L g158 ( 
.A1(n_150),
.A2(n_78),
.B(n_128),
.Y(n_158)
);

OAI221xp5_ASAP7_75t_L g159 ( 
.A1(n_148),
.A2(n_78),
.B1(n_154),
.B2(n_152),
.C(n_128),
.Y(n_159)
);

OAI221xp5_ASAP7_75t_SL g160 ( 
.A1(n_153),
.A2(n_117),
.B1(n_108),
.B2(n_132),
.C(n_80),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_132),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_157),
.A2(n_132),
.B1(n_131),
.B2(n_104),
.Y(n_162)
);

NAND3xp33_ASAP7_75t_SL g163 ( 
.A(n_159),
.B(n_86),
.C(n_90),
.Y(n_163)
);

OAI211xp5_ASAP7_75t_SL g164 ( 
.A1(n_155),
.A2(n_104),
.B(n_90),
.C(n_129),
.Y(n_164)
);

NAND3xp33_ASAP7_75t_SL g165 ( 
.A(n_157),
.B(n_129),
.C(n_108),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_164),
.B(n_158),
.Y(n_166)
);

NAND4xp25_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_160),
.C(n_156),
.D(n_161),
.Y(n_167)
);

AND2x4_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_131),
.Y(n_168)
);

AND2x4_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_131),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_169),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_166),
.A2(n_127),
.B1(n_108),
.B2(n_111),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_127),
.Y(n_172)
);

AOI21xp33_ASAP7_75t_L g173 ( 
.A1(n_170),
.A2(n_168),
.B(n_127),
.Y(n_173)
);

OR2x6_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_127),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_171),
.B(n_173),
.Y(n_175)
);


endmodule