module fake_jpeg_27107_n_35 (n_3, n_2, n_1, n_0, n_4, n_5, n_35);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_35;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx5_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

INVx11_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_5),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

AO22x1_ASAP7_75t_SL g12 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_12),
.A2(n_16),
.B1(n_17),
.B2(n_11),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_9),
.B(n_0),
.Y(n_13)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_6),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_7),
.A2(n_10),
.B1(n_11),
.B2(n_8),
.Y(n_16)
);

OAI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_7),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_18),
.A2(n_20),
.B1(n_10),
.B2(n_7),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_13),
.A2(n_12),
.B1(n_7),
.B2(n_11),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_12),
.C(n_16),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_24),
.C(n_25),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_14),
.C(n_12),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_20),
.C(n_19),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_26),
.A2(n_18),
.B1(n_10),
.B2(n_15),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_9),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_31),
.C(n_14),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_14),
.C(n_8),
.Y(n_31)
);

OA21x2_ASAP7_75t_SL g33 ( 
.A1(n_32),
.A2(n_6),
.B(n_9),
.Y(n_33)
);

AOI221xp5_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_34),
.B1(n_31),
.B2(n_3),
.C(n_4),
.Y(n_35)
);


endmodule