module fake_netlist_1_11643_n_20 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_20);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_20;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_19;
NAND2xp5_ASAP7_75t_L g11 ( .A(n_4), .B(n_2), .Y(n_11) );
INVxp67_ASAP7_75t_SL g12 ( .A(n_8), .Y(n_12) );
BUFx3_ASAP7_75t_L g13 ( .A(n_7), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_10), .Y(n_14) );
OAI22xp5_ASAP7_75t_L g15 ( .A1(n_12), .A2(n_0), .B1(n_1), .B2(n_3), .Y(n_15) );
INVxp67_ASAP7_75t_L g16 ( .A(n_15), .Y(n_16) );
NOR2xp33_ASAP7_75t_L g17 ( .A(n_16), .B(n_14), .Y(n_17) );
AOI22xp5_ASAP7_75t_L g18 ( .A1(n_17), .A2(n_13), .B1(n_11), .B2(n_0), .Y(n_18) );
INVxp67_ASAP7_75t_L g19 ( .A(n_18), .Y(n_19) );
AOI22xp33_ASAP7_75t_SL g20 ( .A1(n_19), .A2(n_9), .B1(n_5), .B2(n_6), .Y(n_20) );
endmodule