module fake_netlist_1_3532_n_530 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_530);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_530;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g78 ( .A(n_36), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_7), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_33), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_41), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_63), .Y(n_82) );
INVxp67_ASAP7_75t_SL g83 ( .A(n_40), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_58), .Y(n_84) );
XOR2xp5_ASAP7_75t_L g85 ( .A(n_43), .B(n_22), .Y(n_85) );
CKINVDCx20_ASAP7_75t_R g86 ( .A(n_51), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_23), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_26), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_48), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_10), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_17), .Y(n_91) );
INVxp33_ASAP7_75t_SL g92 ( .A(n_56), .Y(n_92) );
CKINVDCx16_ASAP7_75t_R g93 ( .A(n_20), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_35), .Y(n_94) );
CKINVDCx16_ASAP7_75t_R g95 ( .A(n_65), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_62), .Y(n_96) );
BUFx3_ASAP7_75t_L g97 ( .A(n_54), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_10), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_16), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_32), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_12), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_31), .Y(n_102) );
INVxp33_ASAP7_75t_L g103 ( .A(n_8), .Y(n_103) );
INVxp33_ASAP7_75t_SL g104 ( .A(n_64), .Y(n_104) );
INVxp33_ASAP7_75t_SL g105 ( .A(n_6), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_44), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_13), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_73), .Y(n_108) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_6), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_2), .Y(n_110) );
CKINVDCx14_ASAP7_75t_R g111 ( .A(n_57), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_72), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_37), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_78), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_78), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_94), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_94), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_108), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_103), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_108), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_80), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_80), .Y(n_122) );
OAI22xp5_ASAP7_75t_L g123 ( .A1(n_93), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_81), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_81), .Y(n_125) );
INVx3_ASAP7_75t_L g126 ( .A(n_82), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_97), .Y(n_127) );
HB1xp67_ASAP7_75t_L g128 ( .A(n_109), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_82), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_96), .B(n_0), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_97), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g132 ( .A(n_105), .B(n_1), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_84), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_84), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_87), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_95), .B(n_3), .Y(n_136) );
INVx3_ASAP7_75t_L g137 ( .A(n_126), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_126), .Y(n_138) );
BUFx3_ASAP7_75t_L g139 ( .A(n_127), .Y(n_139) );
OAI22xp33_ASAP7_75t_SL g140 ( .A1(n_114), .A2(n_79), .B1(n_98), .B2(n_90), .Y(n_140) );
BUFx2_ASAP7_75t_L g141 ( .A(n_119), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_126), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_128), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_127), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_126), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_114), .B(n_113), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_120), .Y(n_147) );
BUFx10_ASAP7_75t_L g148 ( .A(n_115), .Y(n_148) );
BUFx2_ASAP7_75t_L g149 ( .A(n_136), .Y(n_149) );
INVx4_ASAP7_75t_L g150 ( .A(n_127), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_120), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_115), .B(n_87), .Y(n_152) );
AO22x2_ASAP7_75t_L g153 ( .A1(n_123), .A2(n_85), .B1(n_112), .B2(n_88), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_127), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_120), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_116), .Y(n_156) );
BUFx3_ASAP7_75t_L g157 ( .A(n_127), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g158 ( .A(n_136), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_122), .B(n_88), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_131), .Y(n_160) );
BUFx10_ASAP7_75t_L g161 ( .A(n_122), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_148), .B(n_125), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_137), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_137), .Y(n_164) );
INVxp67_ASAP7_75t_L g165 ( .A(n_141), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_141), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_148), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_148), .B(n_92), .Y(n_168) );
AOI211xp5_ASAP7_75t_L g169 ( .A1(n_140), .A2(n_132), .B(n_79), .C(n_90), .Y(n_169) );
AND2x4_ASAP7_75t_SL g170 ( .A(n_148), .B(n_86), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_148), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_137), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_143), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_161), .B(n_140), .Y(n_174) );
INVx2_ASAP7_75t_SL g175 ( .A(n_161), .Y(n_175) );
INVx2_ASAP7_75t_SL g176 ( .A(n_161), .Y(n_176) );
OR2x2_ASAP7_75t_L g177 ( .A(n_149), .B(n_85), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_158), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_149), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_137), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_137), .Y(n_181) );
INVx2_ASAP7_75t_SL g182 ( .A(n_161), .Y(n_182) );
BUFx3_ASAP7_75t_L g183 ( .A(n_161), .Y(n_183) );
INVx2_ASAP7_75t_SL g184 ( .A(n_146), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_138), .B(n_125), .Y(n_185) );
OAI221xp5_ASAP7_75t_L g186 ( .A1(n_146), .A2(n_129), .B1(n_133), .B2(n_135), .C(n_130), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_138), .Y(n_187) );
AND2x4_ASAP7_75t_L g188 ( .A(n_152), .B(n_129), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_142), .B(n_104), .Y(n_189) );
CKINVDCx8_ASAP7_75t_R g190 ( .A(n_159), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_142), .Y(n_191) );
INVx3_ASAP7_75t_L g192 ( .A(n_155), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_159), .B(n_133), .Y(n_193) );
INVx5_ASAP7_75t_L g194 ( .A(n_154), .Y(n_194) );
OR2x6_ASAP7_75t_L g195 ( .A(n_184), .B(n_153), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_184), .B(n_147), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_187), .Y(n_197) );
AOI221xp5_ASAP7_75t_L g198 ( .A1(n_165), .A2(n_153), .B1(n_135), .B2(n_107), .C(n_152), .Y(n_198) );
INVx1_ASAP7_75t_SL g199 ( .A(n_166), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_187), .Y(n_200) );
INVx3_ASAP7_75t_L g201 ( .A(n_183), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_187), .Y(n_202) );
INVxp67_ASAP7_75t_L g203 ( .A(n_177), .Y(n_203) );
AND2x2_ASAP7_75t_SL g204 ( .A(n_170), .B(n_89), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_191), .Y(n_205) );
BUFx2_ASAP7_75t_L g206 ( .A(n_183), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_193), .B(n_145), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_191), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_191), .Y(n_209) );
INVx2_ASAP7_75t_SL g210 ( .A(n_183), .Y(n_210) );
BUFx2_ASAP7_75t_SL g211 ( .A(n_167), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_163), .Y(n_212) );
AND3x1_ASAP7_75t_SL g213 ( .A(n_177), .B(n_153), .C(n_101), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_193), .B(n_145), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g215 ( .A1(n_169), .A2(n_153), .B1(n_151), .B2(n_147), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_162), .A2(n_151), .B(n_156), .Y(n_216) );
CKINVDCx11_ASAP7_75t_R g217 ( .A(n_190), .Y(n_217) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_167), .Y(n_218) );
AOI22xp5_ASAP7_75t_SL g219 ( .A1(n_178), .A2(n_153), .B1(n_99), .B2(n_111), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_162), .Y(n_220) );
AND3x2_ASAP7_75t_L g221 ( .A(n_169), .B(n_153), .C(n_83), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_174), .A2(n_156), .B1(n_155), .B2(n_121), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_179), .B(n_121), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_186), .A2(n_155), .B1(n_134), .B2(n_124), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_164), .Y(n_225) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_186), .A2(n_155), .B1(n_124), .B2(n_134), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_190), .B(n_155), .Y(n_227) );
BUFx4f_ASAP7_75t_SL g228 ( .A(n_199), .Y(n_228) );
BUFx2_ASAP7_75t_L g229 ( .A(n_206), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g230 ( .A1(n_195), .A2(n_170), .B1(n_173), .B2(n_188), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_205), .Y(n_231) );
AOI22xp33_ASAP7_75t_SL g232 ( .A1(n_219), .A2(n_170), .B1(n_91), .B2(n_98), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_220), .B(n_188), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_218), .Y(n_234) );
CKINVDCx9p33_ASAP7_75t_R g235 ( .A(n_204), .Y(n_235) );
INVx1_ASAP7_75t_SL g236 ( .A(n_211), .Y(n_236) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_195), .A2(n_185), .B1(n_188), .B2(n_117), .Y(n_237) );
NAND2x1p5_ASAP7_75t_L g238 ( .A(n_218), .B(n_167), .Y(n_238) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_218), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_195), .A2(n_188), .B1(n_192), .B2(n_189), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_195), .A2(n_192), .B1(n_172), .B2(n_181), .Y(n_241) );
BUFx2_ASAP7_75t_L g242 ( .A(n_206), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_217), .Y(n_243) );
OAI211xp5_ASAP7_75t_L g244 ( .A1(n_198), .A2(n_101), .B(n_110), .C(n_91), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_218), .Y(n_245) );
OAI22xp33_ASAP7_75t_L g246 ( .A1(n_215), .A2(n_185), .B1(n_167), .B2(n_171), .Y(n_246) );
NAND2x1_ASAP7_75t_L g247 ( .A(n_218), .B(n_163), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g248 ( .A(n_219), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_197), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g250 ( .A1(n_204), .A2(n_192), .B1(n_164), .B2(n_181), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_197), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_203), .B(n_168), .Y(n_252) );
AND2x4_ASAP7_75t_L g253 ( .A(n_220), .B(n_167), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_205), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_232), .A2(n_204), .B1(n_221), .B2(n_223), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_232), .A2(n_215), .B1(n_196), .B2(n_227), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_231), .Y(n_257) );
AO31x2_ASAP7_75t_L g258 ( .A1(n_237), .A2(n_208), .A3(n_200), .B(n_202), .Y(n_258) );
INVx5_ASAP7_75t_SL g259 ( .A(n_235), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_231), .Y(n_260) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_228), .Y(n_261) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_229), .Y(n_262) );
OAI22xp5_ASAP7_75t_L g263 ( .A1(n_237), .A2(n_226), .B1(n_208), .B2(n_196), .Y(n_263) );
OAI21x1_ASAP7_75t_L g264 ( .A1(n_247), .A2(n_222), .B(n_200), .Y(n_264) );
AO21x2_ASAP7_75t_L g265 ( .A1(n_246), .A2(n_222), .B(n_226), .Y(n_265) );
OAI21xp5_ASAP7_75t_L g266 ( .A1(n_233), .A2(n_216), .B(n_224), .Y(n_266) );
NOR2x1_ASAP7_75t_SL g267 ( .A(n_254), .B(n_211), .Y(n_267) );
A2O1A1Ixp33_ASAP7_75t_L g268 ( .A1(n_244), .A2(n_214), .B(n_207), .C(n_202), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_248), .A2(n_225), .B1(n_192), .B2(n_209), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_230), .A2(n_209), .B1(n_210), .B2(n_201), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_243), .Y(n_271) );
OAI221xp5_ASAP7_75t_L g272 ( .A1(n_252), .A2(n_244), .B1(n_240), .B2(n_250), .C(n_241), .Y(n_272) );
AOI221xp5_ASAP7_75t_L g273 ( .A1(n_233), .A2(n_110), .B1(n_225), .B2(n_117), .C(n_116), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_254), .B(n_201), .Y(n_274) );
CKINVDCx20_ASAP7_75t_R g275 ( .A(n_229), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_249), .Y(n_276) );
OAI31xp33_ASAP7_75t_L g277 ( .A1(n_263), .A2(n_242), .A3(n_253), .B(n_213), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_257), .B(n_249), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_276), .B(n_249), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g280 ( .A1(n_255), .A2(n_242), .B1(n_253), .B2(n_251), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_272), .A2(n_253), .B1(n_251), .B2(n_118), .Y(n_281) );
OAI222xp33_ASAP7_75t_L g282 ( .A1(n_263), .A2(n_236), .B1(n_251), .B2(n_253), .C1(n_238), .C2(n_89), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_276), .Y(n_283) );
AOI22xp33_ASAP7_75t_SL g284 ( .A1(n_259), .A2(n_236), .B1(n_239), .B2(n_238), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_257), .Y(n_285) );
OA21x2_ASAP7_75t_L g286 ( .A1(n_264), .A2(n_234), .B(n_245), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_260), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_260), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_258), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_258), .Y(n_290) );
BUFx2_ASAP7_75t_L g291 ( .A(n_258), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_256), .A2(n_118), .B1(n_201), .B2(n_210), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_274), .B(n_234), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_258), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g295 ( .A1(n_259), .A2(n_212), .B1(n_112), .B2(n_102), .Y(n_295) );
AOI222xp33_ASAP7_75t_L g296 ( .A1(n_259), .A2(n_100), .B1(n_102), .B2(n_212), .C1(n_172), .C2(n_180), .Y(n_296) );
OAI221xp5_ASAP7_75t_L g297 ( .A1(n_268), .A2(n_100), .B1(n_238), .B2(n_180), .C(n_150), .Y(n_297) );
AOI221xp5_ASAP7_75t_L g298 ( .A1(n_273), .A2(n_131), .B1(n_163), .B2(n_150), .C(n_106), .Y(n_298) );
INVxp67_ASAP7_75t_L g299 ( .A(n_279), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_285), .Y(n_300) );
OAI221xp5_ASAP7_75t_L g301 ( .A1(n_277), .A2(n_269), .B1(n_262), .B2(n_261), .C(n_266), .Y(n_301) );
AO21x2_ASAP7_75t_L g302 ( .A1(n_282), .A2(n_264), .B(n_265), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_290), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_285), .Y(n_304) );
INVx5_ASAP7_75t_SL g305 ( .A(n_283), .Y(n_305) );
BUFx2_ASAP7_75t_L g306 ( .A(n_291), .Y(n_306) );
NAND4xp25_ASAP7_75t_L g307 ( .A(n_277), .B(n_266), .C(n_150), .D(n_274), .Y(n_307) );
INVx4_ASAP7_75t_L g308 ( .A(n_279), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_288), .B(n_275), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_288), .B(n_274), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_285), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_287), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_283), .B(n_258), .Y(n_313) );
AOI21xp33_ASAP7_75t_L g314 ( .A1(n_296), .A2(n_270), .B(n_274), .Y(n_314) );
OAI31xp33_ASAP7_75t_L g315 ( .A1(n_282), .A2(n_259), .A3(n_245), .B(n_234), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_283), .B(n_258), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_290), .B(n_267), .Y(n_317) );
INVx3_ASAP7_75t_L g318 ( .A(n_286), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_287), .Y(n_319) );
INVxp67_ASAP7_75t_SL g320 ( .A(n_279), .Y(n_320) );
AOI322xp5_ASAP7_75t_L g321 ( .A1(n_280), .A2(n_287), .A3(n_281), .B1(n_278), .B2(n_291), .C1(n_289), .C2(n_290), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_294), .Y(n_322) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_278), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_289), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_294), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_292), .A2(n_259), .B1(n_265), .B2(n_245), .Y(n_326) );
INVx1_ASAP7_75t_SL g327 ( .A(n_293), .Y(n_327) );
AOI221xp5_ASAP7_75t_L g328 ( .A1(n_297), .A2(n_271), .B1(n_131), .B2(n_150), .C(n_265), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_313), .B(n_294), .Y(n_329) );
AND2x4_ASAP7_75t_L g330 ( .A(n_317), .B(n_293), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_313), .B(n_316), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_324), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_303), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_320), .B(n_296), .Y(n_334) );
NAND4xp25_ASAP7_75t_L g335 ( .A(n_309), .B(n_295), .C(n_297), .D(n_298), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_327), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_308), .A2(n_298), .B1(n_284), .B2(n_286), .Y(n_337) );
OR2x2_ASAP7_75t_L g338 ( .A(n_308), .B(n_286), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_317), .B(n_267), .Y(n_339) );
NOR2xp33_ASAP7_75t_SL g340 ( .A(n_315), .B(n_239), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_323), .B(n_286), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_324), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_303), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_303), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_300), .Y(n_345) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_308), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_300), .B(n_286), .Y(n_347) );
BUFx2_ASAP7_75t_L g348 ( .A(n_308), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_304), .Y(n_349) );
BUFx2_ASAP7_75t_L g350 ( .A(n_317), .Y(n_350) );
NOR3xp33_ASAP7_75t_SL g351 ( .A(n_301), .B(n_3), .C(n_4), .Y(n_351) );
INVxp67_ASAP7_75t_SL g352 ( .A(n_322), .Y(n_352) );
NAND2xp5_ASAP7_75t_SL g353 ( .A(n_315), .B(n_284), .Y(n_353) );
AND2x2_ASAP7_75t_SL g354 ( .A(n_306), .B(n_239), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_316), .B(n_325), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_322), .Y(n_356) );
BUFx3_ASAP7_75t_L g357 ( .A(n_317), .Y(n_357) );
NOR3xp33_ASAP7_75t_SL g358 ( .A(n_307), .B(n_4), .C(n_5), .Y(n_358) );
AND4x1_ASAP7_75t_L g359 ( .A(n_328), .B(n_5), .C(n_7), .D(n_8), .Y(n_359) );
OAI33xp33_ASAP7_75t_L g360 ( .A1(n_310), .A2(n_144), .A3(n_160), .B1(n_12), .B2(n_13), .B3(n_14), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_299), .B(n_9), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_325), .B(n_131), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_322), .Y(n_363) );
CKINVDCx16_ASAP7_75t_R g364 ( .A(n_306), .Y(n_364) );
BUFx2_ASAP7_75t_L g365 ( .A(n_318), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_304), .B(n_9), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_311), .B(n_131), .Y(n_367) );
AND2x4_ASAP7_75t_L g368 ( .A(n_318), .B(n_239), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_311), .B(n_150), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_312), .Y(n_370) );
NOR3xp33_ASAP7_75t_L g371 ( .A(n_314), .B(n_160), .C(n_144), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_312), .B(n_11), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_319), .B(n_144), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_331), .B(n_319), .Y(n_374) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_353), .A2(n_326), .B(n_302), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_331), .B(n_321), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_332), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_332), .Y(n_378) );
OAI211xp5_ASAP7_75t_L g379 ( .A1(n_348), .A2(n_321), .B(n_318), .C(n_160), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_336), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_329), .B(n_318), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_342), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_355), .B(n_305), .Y(n_383) );
NAND2xp5_ASAP7_75t_SL g384 ( .A(n_340), .B(n_305), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_345), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_345), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_329), .B(n_302), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_349), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_361), .B(n_11), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_349), .Y(n_390) );
NOR2x1_ASAP7_75t_L g391 ( .A(n_348), .B(n_302), .Y(n_391) );
AND2x4_ASAP7_75t_L g392 ( .A(n_357), .B(n_305), .Y(n_392) );
AOI21xp5_ASAP7_75t_L g393 ( .A1(n_340), .A2(n_247), .B(n_239), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_370), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_370), .Y(n_395) );
NAND2x1p5_ASAP7_75t_L g396 ( .A(n_339), .B(n_305), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_355), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_364), .B(n_305), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_364), .B(n_14), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_335), .A2(n_154), .B1(n_239), .B2(n_157), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_333), .Y(n_401) );
AOI21xp33_ASAP7_75t_L g402 ( .A1(n_372), .A2(n_15), .B(n_16), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_350), .B(n_154), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_346), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_350), .B(n_154), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_333), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_372), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_366), .Y(n_408) );
NOR3xp33_ASAP7_75t_L g409 ( .A(n_360), .B(n_335), .C(n_371), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_334), .B(n_15), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_330), .B(n_154), .Y(n_411) );
INVx1_ASAP7_75t_SL g412 ( .A(n_339), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_338), .B(n_17), .Y(n_413) );
NAND4xp25_ASAP7_75t_L g414 ( .A(n_337), .B(n_157), .C(n_139), .D(n_20), .Y(n_414) );
OAI21xp33_ASAP7_75t_L g415 ( .A1(n_351), .A2(n_154), .B(n_157), .Y(n_415) );
INVx1_ASAP7_75t_SL g416 ( .A(n_339), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_330), .B(n_154), .Y(n_417) );
NAND4xp25_ASAP7_75t_L g418 ( .A(n_338), .B(n_139), .C(n_18), .D(n_19), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_341), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_352), .B(n_18), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_330), .B(n_19), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_365), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_381), .B(n_365), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_374), .Y(n_424) );
OAI322xp33_ASAP7_75t_L g425 ( .A1(n_376), .A2(n_341), .A3(n_347), .B1(n_354), .B2(n_356), .C1(n_363), .C2(n_344), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_381), .B(n_357), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_374), .Y(n_427) );
NAND2xp5_ASAP7_75t_SL g428 ( .A(n_384), .B(n_354), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_397), .Y(n_429) );
NAND2xp5_ASAP7_75t_SL g430 ( .A(n_384), .B(n_354), .Y(n_430) );
INVx1_ASAP7_75t_SL g431 ( .A(n_380), .Y(n_431) );
OAI322xp33_ASAP7_75t_L g432 ( .A1(n_413), .A2(n_347), .A3(n_343), .B1(n_363), .B2(n_356), .C1(n_344), .C2(n_369), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_387), .B(n_357), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_377), .Y(n_434) );
NAND2xp5_ASAP7_75t_SL g435 ( .A(n_413), .B(n_339), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_419), .B(n_367), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_378), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_410), .B(n_359), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_387), .B(n_330), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_399), .B(n_359), .Y(n_440) );
OAI21xp5_ASAP7_75t_SL g441 ( .A1(n_418), .A2(n_358), .B(n_362), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_408), .B(n_367), .Y(n_442) );
AOI222xp33_ASAP7_75t_L g443 ( .A1(n_389), .A2(n_362), .B1(n_373), .B2(n_356), .C1(n_363), .C2(n_344), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_401), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_382), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_407), .B(n_343), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_412), .B(n_416), .Y(n_447) );
OAI32xp33_ASAP7_75t_L g448 ( .A1(n_396), .A2(n_369), .A3(n_373), .B1(n_368), .B2(n_139), .Y(n_448) );
XNOR2xp5_ASAP7_75t_L g449 ( .A(n_421), .B(n_368), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_404), .B(n_368), .Y(n_450) );
A2O1A1Ixp33_ASAP7_75t_L g451 ( .A1(n_414), .A2(n_21), .B(n_24), .C(n_25), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_385), .B(n_27), .Y(n_452) );
NAND2xp33_ASAP7_75t_L g453 ( .A(n_396), .B(n_171), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_386), .Y(n_454) );
XOR2x2_ASAP7_75t_L g455 ( .A(n_421), .B(n_28), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_388), .Y(n_456) );
INVx1_ASAP7_75t_SL g457 ( .A(n_398), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_389), .B(n_29), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_390), .Y(n_459) );
XOR2x2_ASAP7_75t_L g460 ( .A(n_396), .B(n_30), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_394), .B(n_34), .Y(n_461) );
BUFx2_ASAP7_75t_SL g462 ( .A(n_392), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_395), .B(n_38), .Y(n_463) );
AOI221xp5_ASAP7_75t_L g464 ( .A1(n_409), .A2(n_194), .B1(n_42), .B2(n_45), .C(n_46), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_420), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_379), .A2(n_194), .B1(n_47), .B2(n_49), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_375), .B(n_39), .Y(n_467) );
OAI221xp5_ASAP7_75t_L g468 ( .A1(n_400), .A2(n_402), .B1(n_415), .B2(n_391), .C(n_422), .Y(n_468) );
AOI221xp5_ASAP7_75t_L g469 ( .A1(n_400), .A2(n_194), .B1(n_52), .B2(n_53), .C(n_55), .Y(n_469) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_411), .A2(n_194), .B1(n_59), .B2(n_60), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_L g471 ( .A1(n_411), .A2(n_50), .B(n_61), .C(n_66), .Y(n_471) );
OAI321xp33_ASAP7_75t_L g472 ( .A1(n_383), .A2(n_67), .A3(n_68), .B1(n_69), .B2(n_70), .C(n_71), .Y(n_472) );
AOI211xp5_ASAP7_75t_L g473 ( .A1(n_392), .A2(n_74), .B(n_75), .C(n_76), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g474 ( .A1(n_417), .A2(n_194), .B1(n_77), .B2(n_175), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_406), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_403), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_417), .B(n_194), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_392), .B(n_167), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_405), .A2(n_403), .B1(n_393), .B2(n_176), .Y(n_479) );
XNOR2x1_ASAP7_75t_L g480 ( .A(n_405), .B(n_171), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_374), .Y(n_481) );
OAI221xp5_ASAP7_75t_L g482 ( .A1(n_409), .A2(n_175), .B1(n_176), .B2(n_182), .C(n_171), .Y(n_482) );
BUFx12f_ASAP7_75t_L g483 ( .A(n_421), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_374), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_376), .B(n_171), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g486 ( .A1(n_413), .A2(n_171), .B1(n_182), .B2(n_348), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_374), .Y(n_487) );
INVx2_ASAP7_75t_SL g488 ( .A(n_380), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_380), .B(n_410), .Y(n_489) );
NOR2xp67_ASAP7_75t_L g490 ( .A(n_380), .B(n_418), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_453), .A2(n_460), .B(n_430), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_465), .B(n_443), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_490), .A2(n_438), .B1(n_440), .B2(n_480), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_462), .A2(n_483), .B1(n_431), .B2(n_435), .Y(n_494) );
NOR2xp33_ASAP7_75t_SL g495 ( .A(n_488), .B(n_432), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_427), .B(n_424), .Y(n_496) );
AOI211xp5_ASAP7_75t_L g497 ( .A1(n_453), .A2(n_468), .B(n_425), .C(n_430), .Y(n_497) );
AOI22x1_ASAP7_75t_L g498 ( .A1(n_460), .A2(n_449), .B1(n_455), .B2(n_457), .Y(n_498) );
NOR4xp25_ASAP7_75t_L g499 ( .A(n_489), .B(n_441), .C(n_467), .D(n_451), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_446), .Y(n_500) );
OA22x2_ASAP7_75t_L g501 ( .A1(n_435), .A2(n_428), .B1(n_484), .B2(n_481), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_428), .A2(n_455), .B(n_451), .Y(n_502) );
NOR3xp33_ASAP7_75t_L g503 ( .A(n_464), .B(n_482), .C(n_472), .Y(n_503) );
NAND3xp33_ASAP7_75t_L g504 ( .A(n_485), .B(n_473), .C(n_466), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_487), .B(n_429), .Y(n_505) );
NAND4xp75_ASAP7_75t_L g506 ( .A(n_458), .B(n_442), .C(n_447), .D(n_479), .Y(n_506) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_423), .Y(n_507) );
AND2x4_ASAP7_75t_L g508 ( .A(n_491), .B(n_439), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_505), .Y(n_509) );
AOI211xp5_ASAP7_75t_L g510 ( .A1(n_491), .A2(n_448), .B(n_486), .C(n_466), .Y(n_510) );
AOI211xp5_ASAP7_75t_L g511 ( .A1(n_499), .A2(n_486), .B(n_472), .C(n_471), .Y(n_511) );
NAND3xp33_ASAP7_75t_SL g512 ( .A(n_497), .B(n_469), .C(n_470), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_492), .B(n_436), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_494), .B(n_439), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_506), .A2(n_447), .B1(n_433), .B2(n_423), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_496), .Y(n_516) );
NOR3xp33_ASAP7_75t_L g517 ( .A(n_512), .B(n_502), .C(n_503), .Y(n_517) );
NOR2x1_ASAP7_75t_L g518 ( .A(n_508), .B(n_504), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_L g519 ( .A1(n_511), .A2(n_495), .B(n_493), .C(n_507), .Y(n_519) );
NAND4xp25_ASAP7_75t_L g520 ( .A(n_510), .B(n_498), .C(n_474), .D(n_478), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_514), .A2(n_501), .B(n_500), .C(n_426), .Y(n_521) );
OAI222xp33_ASAP7_75t_L g522 ( .A1(n_518), .A2(n_501), .B1(n_513), .B2(n_515), .C1(n_509), .C2(n_516), .Y(n_522) );
AOI221xp5_ASAP7_75t_L g523 ( .A1(n_517), .A2(n_454), .B1(n_459), .B2(n_456), .C(n_434), .Y(n_523) );
OR3x1_ASAP7_75t_L g524 ( .A(n_520), .B(n_445), .C(n_437), .Y(n_524) );
AO22x2_ASAP7_75t_L g525 ( .A1(n_524), .A2(n_519), .B1(n_521), .B2(n_463), .Y(n_525) );
AND3x4_ASAP7_75t_L g526 ( .A(n_522), .B(n_476), .C(n_444), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_525), .B(n_523), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_527), .Y(n_528) );
OAI21xp5_ASAP7_75t_L g529 ( .A1(n_528), .A2(n_526), .B(n_461), .Y(n_529) );
AOI221xp5_ASAP7_75t_L g530 ( .A1(n_529), .A2(n_477), .B1(n_452), .B2(n_450), .C(n_475), .Y(n_530) );
endmodule