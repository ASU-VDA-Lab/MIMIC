module real_jpeg_31070_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_38;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_47;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_40;
wire n_36;
wire n_39;
wire n_41;
wire n_27;
wire n_32;
wire n_20;
wire n_19;
wire n_26;
wire n_48;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

INVx4_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_0),
.B(n_27),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_0),
.B(n_40),
.Y(n_42)
);

BUFx2_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

NAND2x1p5_ASAP7_75t_L g34 ( 
.A(n_1),
.B(n_13),
.Y(n_34)
);

AND2x4_ASAP7_75t_SL g7 ( 
.A(n_2),
.B(n_8),
.Y(n_7)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_2),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_2),
.B(n_27),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_2),
.B(n_37),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_3),
.B(n_21),
.Y(n_20)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

OA22x2_ASAP7_75t_L g11 ( 
.A1(n_4),
.A2(n_5),
.B1(n_12),
.B2(n_13),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

AO21x1_ASAP7_75t_L g37 ( 
.A1(n_4),
.A2(n_32),
.B(n_34),
.Y(n_37)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_5),
.B(n_33),
.Y(n_32)
);

O2A1O1Ixp33_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_16),
.B(n_19),
.C(n_22),
.Y(n_6)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_9),
.Y(n_8)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_9),
.B(n_18),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g9 ( 
.A1(n_10),
.A2(n_11),
.B1(n_14),
.B2(n_15),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_11),
.Y(n_10)
);

OA21x2_ASAP7_75t_L g31 ( 
.A1(n_12),
.A2(n_32),
.B(n_34),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_14),
.B(n_18),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_18),
.Y(n_23)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

INVx2_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_21),
.B(n_45),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B(n_26),
.C(n_28),
.Y(n_22)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

O2A1O1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_35),
.B(n_38),
.C(n_41),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B(n_44),
.C(n_47),
.Y(n_41)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);


endmodule