module fake_jpeg_11999_n_582 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_582);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_582;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_1),
.B(n_5),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_2),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_14),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_17),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_61),
.Y(n_163)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_62),
.Y(n_139)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

NOR2xp67_ASAP7_75t_L g64 ( 
.A(n_28),
.B(n_0),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_64),
.B(n_74),
.Y(n_129)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_65),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_67),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_68),
.Y(n_194)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_69),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_70),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_71),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_72),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_73),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_34),
.B(n_1),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_21),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_75),
.B(n_87),
.Y(n_133)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx5_ASAP7_75t_SL g148 ( 
.A(n_76),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_77),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_78),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_40),
.B(n_2),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_79),
.B(n_84),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_80),
.Y(n_204)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_82),
.Y(n_156)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_83),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_40),
.B(n_2),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_34),
.B(n_2),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_85),
.B(n_127),
.Y(n_162)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_86),
.Y(n_143)
);

BUFx16f_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_89),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_21),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_90),
.B(n_92),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_3),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_91),
.B(n_3),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_21),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_93),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_94),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_95),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_21),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_96),
.B(n_100),
.Y(n_164)
);

AND2x4_ASAP7_75t_SL g97 ( 
.A(n_33),
.B(n_47),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_97),
.B(n_99),
.Y(n_153)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_98),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_43),
.B(n_3),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_48),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_101),
.Y(n_152)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_22),
.Y(n_102)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_102),
.Y(n_176)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_23),
.Y(n_103)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_103),
.Y(n_192)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_23),
.Y(n_104)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_104),
.Y(n_197)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_44),
.Y(n_105)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_105),
.Y(n_178)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_35),
.Y(n_106)
);

INVx11_ASAP7_75t_L g206 ( 
.A(n_106),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_22),
.Y(n_107)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_108),
.Y(n_160)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_30),
.Y(n_109)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_109),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_22),
.Y(n_110)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

BUFx10_ASAP7_75t_L g111 ( 
.A(n_32),
.Y(n_111)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_32),
.Y(n_112)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

CKINVDCx9p33_ASAP7_75t_R g113 ( 
.A(n_19),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_113),
.B(n_121),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_41),
.Y(n_114)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_114),
.Y(n_183)
);

BUFx16f_ASAP7_75t_L g115 ( 
.A(n_41),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_115),
.B(n_120),
.Y(n_166)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_30),
.Y(n_116)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_116),
.Y(n_173)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_24),
.Y(n_117)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_117),
.Y(n_193)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_51),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_24),
.Y(n_119)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_119),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_41),
.B(n_3),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_27),
.Y(n_121)
);

INVx11_ASAP7_75t_SL g122 ( 
.A(n_41),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_122),
.B(n_124),
.Y(n_175)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_60),
.Y(n_123)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_123),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_51),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_51),
.Y(n_125)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_125),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_60),
.Y(n_126)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_126),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_60),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_89),
.A2(n_50),
.B1(n_52),
.B2(n_45),
.Y(n_128)
);

OAI22x1_ASAP7_75t_L g275 ( 
.A1(n_128),
.A2(n_130),
.B1(n_132),
.B2(n_189),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_70),
.A2(n_50),
.B1(n_52),
.B2(n_45),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_94),
.A2(n_50),
.B1(n_27),
.B2(n_46),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_83),
.A2(n_39),
.B1(n_42),
.B2(n_46),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_137),
.A2(n_151),
.B1(n_158),
.B2(n_190),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_93),
.A2(n_59),
.B1(n_26),
.B2(n_29),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_141),
.A2(n_161),
.B1(n_169),
.B2(n_171),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_95),
.A2(n_39),
.B1(n_42),
.B2(n_55),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_99),
.A2(n_25),
.B1(n_57),
.B2(n_55),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_66),
.A2(n_59),
.B1(n_19),
.B2(n_25),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_71),
.A2(n_57),
.B1(n_38),
.B2(n_37),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_73),
.A2(n_38),
.B1(n_37),
.B2(n_31),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_107),
.A2(n_31),
.B1(n_29),
.B2(n_26),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_172),
.A2(n_187),
.B1(n_209),
.B2(n_185),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_177),
.B(n_184),
.Y(n_211)
);

AND2x4_ASAP7_75t_SL g179 ( 
.A(n_97),
.B(n_50),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_179),
.B(n_61),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_87),
.B(n_5),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_115),
.B(n_120),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_186),
.B(n_191),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_110),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_94),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_112),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_124),
.B(n_10),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_82),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_198),
.A2(n_200),
.B1(n_201),
.B2(n_189),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_77),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_105),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_201)
);

OR2x4_ASAP7_75t_L g203 ( 
.A(n_97),
.B(n_16),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_203),
.B(n_205),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_124),
.B(n_16),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_72),
.B(n_88),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_208),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_114),
.B(n_81),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_78),
.A2(n_80),
.B1(n_126),
.B2(n_125),
.Y(n_209)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_199),
.Y(n_212)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_212),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_148),
.A2(n_62),
.B1(n_69),
.B2(n_65),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_213),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_162),
.B(n_118),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_214),
.B(n_225),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_131),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_215),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_131),
.Y(n_216)
);

INVx6_ASAP7_75t_L g318 ( 
.A(n_216),
.Y(n_318)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_143),
.Y(n_217)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_217),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_148),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_218),
.Y(n_301)
);

NAND2x1_ASAP7_75t_SL g219 ( 
.A(n_206),
.B(n_76),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_219),
.Y(n_298)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_202),
.Y(n_220)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_220),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_206),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_223),
.B(n_226),
.Y(n_297)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_224),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_153),
.B(n_102),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_164),
.B(n_123),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_188),
.Y(n_227)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_227),
.Y(n_305)
);

NOR2x1_ASAP7_75t_R g302 ( 
.A(n_228),
.B(n_233),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_153),
.B(n_127),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_229),
.B(n_258),
.Y(n_315)
);

INVx8_ASAP7_75t_L g230 ( 
.A(n_170),
.Y(n_230)
);

INVx5_ASAP7_75t_L g336 ( 
.A(n_230),
.Y(n_336)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_176),
.Y(n_231)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_231),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_138),
.B(n_111),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_232),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_179),
.B(n_68),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_233),
.B(n_245),
.C(n_251),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_147),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_234),
.B(n_235),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_157),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_158),
.B(n_111),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_236),
.B(n_242),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_210),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_238),
.Y(n_303)
);

BUFx4f_ASAP7_75t_SL g239 ( 
.A(n_174),
.Y(n_239)
);

INVx13_ASAP7_75t_L g323 ( 
.A(n_239),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_139),
.A2(n_67),
.B1(n_122),
.B2(n_106),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_240),
.Y(n_321)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_152),
.Y(n_241)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_241),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_175),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_192),
.Y(n_243)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_243),
.Y(n_309)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_174),
.Y(n_244)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_244),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_203),
.A2(n_196),
.B1(n_193),
.B2(n_136),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_151),
.A2(n_173),
.B1(n_167),
.B2(n_137),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_246),
.A2(n_253),
.B1(n_254),
.B2(n_263),
.Y(n_325)
);

BUFx12f_ASAP7_75t_L g247 ( 
.A(n_170),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_142),
.Y(n_248)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_248),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_129),
.B(n_133),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_250),
.B(n_256),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_179),
.A2(n_182),
.B(n_132),
.Y(n_251)
);

INVx8_ASAP7_75t_L g252 ( 
.A(n_181),
.Y(n_252)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_252),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_145),
.A2(n_163),
.B1(n_194),
.B2(n_149),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_160),
.Y(n_255)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_255),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_182),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_130),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_257),
.B(n_261),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_166),
.B(n_154),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_154),
.B(n_200),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_259),
.B(n_262),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_135),
.Y(n_260)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_260),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_146),
.B(n_159),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_134),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_163),
.A2(n_194),
.B1(n_155),
.B2(n_149),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_150),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_264),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_146),
.B(n_159),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_265),
.B(n_267),
.Y(n_311)
);

INVx8_ASAP7_75t_L g266 ( 
.A(n_181),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_266),
.Y(n_294)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_165),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_183),
.B(n_144),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_268),
.B(n_269),
.Y(n_327)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_165),
.Y(n_269)
);

INVx11_ASAP7_75t_L g270 ( 
.A(n_180),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_270),
.Y(n_300)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_185),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_271),
.B(n_276),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_273),
.A2(n_279),
.B1(n_280),
.B2(n_242),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_155),
.A2(n_150),
.B1(n_180),
.B2(n_183),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_274),
.A2(n_281),
.B1(n_218),
.B2(n_280),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_134),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_128),
.A2(n_197),
.B(n_144),
.Y(n_277)
);

FAx1_ASAP7_75t_SL g328 ( 
.A(n_277),
.B(n_219),
.CI(n_270),
.CON(n_328),
.SN(n_328)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_140),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_278),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_204),
.A2(n_135),
.B1(n_168),
.B2(n_140),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_204),
.A2(n_168),
.B1(n_178),
.B2(n_156),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_156),
.A2(n_70),
.B1(n_89),
.B2(n_56),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_197),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_282),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_283),
.A2(n_310),
.B(n_269),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_254),
.A2(n_259),
.B1(n_251),
.B2(n_237),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_287),
.A2(n_291),
.B1(n_313),
.B2(n_314),
.Y(n_344)
);

AOI32xp33_ASAP7_75t_L g289 ( 
.A1(n_229),
.A2(n_225),
.A3(n_214),
.B1(n_258),
.B2(n_256),
.Y(n_289)
);

NOR2x1_ASAP7_75t_L g348 ( 
.A(n_289),
.B(n_239),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_257),
.A2(n_237),
.B1(n_236),
.B2(n_245),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_302),
.B(n_308),
.Y(n_379)
);

NAND2xp33_ASAP7_75t_SL g310 ( 
.A(n_228),
.B(n_233),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_221),
.A2(n_275),
.B1(n_249),
.B2(n_222),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_221),
.A2(n_275),
.B1(n_272),
.B2(n_228),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_316),
.A2(n_317),
.B1(n_266),
.B2(n_252),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_217),
.A2(n_227),
.B1(n_277),
.B2(n_255),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_211),
.A2(n_243),
.B1(n_276),
.B2(n_234),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_326),
.A2(n_337),
.B1(n_239),
.B2(n_247),
.Y(n_362)
);

OR2x2_ASAP7_75t_L g378 ( 
.A(n_328),
.B(n_330),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_219),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_329),
.B(n_311),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_262),
.A2(n_212),
.B1(n_220),
.B2(n_241),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_320),
.B(n_248),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_338),
.B(n_343),
.C(n_351),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_293),
.B(n_224),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_339),
.B(n_346),
.Y(n_385)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_284),
.Y(n_340)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_340),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_301),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_341),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_334),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g390 ( 
.A(n_342),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_320),
.B(n_310),
.C(n_293),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_284),
.Y(n_345)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_345),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_315),
.B(n_235),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_295),
.B(n_231),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_347),
.B(n_359),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_348),
.A2(n_354),
.B(n_365),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_349),
.B(n_358),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_329),
.A2(n_282),
.B(n_264),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_350),
.A2(n_376),
.B(n_378),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_315),
.B(n_238),
.C(n_267),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_305),
.Y(n_352)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_352),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_290),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_353),
.B(n_367),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_291),
.A2(n_278),
.B1(n_271),
.B2(n_244),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_288),
.Y(n_355)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_355),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_356),
.A2(n_364),
.B1(n_370),
.B2(n_375),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_L g357 ( 
.A1(n_287),
.A2(n_230),
.B1(n_216),
.B2(n_215),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_SL g402 ( 
.A1(n_357),
.A2(n_288),
.B1(n_296),
.B2(n_333),
.Y(n_402)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_305),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_326),
.B(n_260),
.Y(n_359)
);

AND2x4_ASAP7_75t_L g360 ( 
.A(n_298),
.B(n_328),
.Y(n_360)
);

BUFx24_ASAP7_75t_L g389 ( 
.A(n_360),
.Y(n_389)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_309),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_361),
.B(n_362),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_312),
.B(n_247),
.Y(n_363)
);

CKINVDCx14_ASAP7_75t_R g411 ( 
.A(n_363),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_316),
.A2(n_247),
.B1(n_289),
.B2(n_332),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_307),
.A2(n_317),
.B(n_328),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_313),
.B(n_314),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_366),
.B(n_377),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_312),
.B(n_297),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_296),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_368),
.Y(n_404)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_309),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_369),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_332),
.A2(n_292),
.B1(n_283),
.B2(n_299),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_371),
.A2(n_378),
.B(n_285),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_337),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_372),
.B(n_374),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_302),
.B(n_327),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_373),
.B(n_286),
.C(n_304),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_306),
.B(n_319),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_299),
.A2(n_325),
.B1(n_321),
.B2(n_300),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_303),
.A2(n_330),
.B(n_319),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_286),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_379),
.B(n_380),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_308),
.B(n_322),
.Y(n_380)
);

MAJx2_ASAP7_75t_L g381 ( 
.A(n_343),
.B(n_335),
.C(n_322),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_381),
.B(n_391),
.C(n_395),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_344),
.A2(n_300),
.B1(n_294),
.B2(n_331),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_384),
.A2(n_397),
.B1(n_402),
.B2(n_403),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_394),
.A2(n_396),
.B(n_360),
.Y(n_417)
);

MAJx2_ASAP7_75t_L g395 ( 
.A(n_338),
.B(n_335),
.C(n_285),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_360),
.A2(n_304),
.B(n_294),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_344),
.A2(n_331),
.B1(n_324),
.B2(n_318),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_401),
.B(n_409),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_366),
.A2(n_378),
.B1(n_346),
.B2(n_364),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_363),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_405),
.B(n_412),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_379),
.B(n_333),
.C(n_324),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_339),
.B(n_336),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_377),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_413),
.B(n_340),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_360),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_416),
.B(n_360),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_417),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_398),
.A2(n_348),
.B1(n_354),
.B2(n_372),
.Y(n_419)
);

AOI22x1_ASAP7_75t_L g452 ( 
.A1(n_419),
.A2(n_442),
.B1(n_444),
.B2(n_446),
.Y(n_452)
);

NAND2xp33_ASAP7_75t_L g455 ( 
.A(n_420),
.B(n_408),
.Y(n_455)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_387),
.Y(n_421)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_421),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_389),
.A2(n_365),
.B(n_349),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_422),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_385),
.B(n_342),
.Y(n_423)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_423),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_385),
.B(n_380),
.Y(n_424)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_424),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_389),
.A2(n_362),
.B(n_370),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_425),
.B(n_439),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_393),
.B(n_353),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_426),
.B(n_427),
.Y(n_462)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_387),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_393),
.B(n_345),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_428),
.B(n_430),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_407),
.B(n_351),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_412),
.B(n_352),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_431),
.B(n_432),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_386),
.B(n_376),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_401),
.B(n_373),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_433),
.B(n_440),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_398),
.A2(n_356),
.B1(n_350),
.B2(n_375),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_435),
.A2(n_443),
.B1(n_410),
.B2(n_392),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_436),
.Y(n_450)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_388),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_438),
.Y(n_451)
);

INVx8_ASAP7_75t_L g439 ( 
.A(n_390),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_388),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_406),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_441),
.B(n_445),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_389),
.A2(n_369),
.B(n_361),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_396),
.A2(n_358),
.B1(n_318),
.B2(n_341),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_416),
.A2(n_355),
.B1(n_336),
.B2(n_288),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_406),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_389),
.A2(n_394),
.B(n_408),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_413),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_447),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_411),
.B(n_404),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_448),
.B(n_405),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_437),
.A2(n_403),
.B1(n_410),
.B2(n_409),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_449),
.A2(n_469),
.B1(n_419),
.B2(n_424),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_434),
.B(n_383),
.C(n_381),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_453),
.B(n_456),
.C(n_467),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_434),
.B(n_383),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_454),
.B(n_459),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_455),
.B(n_475),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_434),
.B(n_381),
.C(n_415),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_458),
.B(n_470),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_433),
.B(n_415),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_429),
.B(n_391),
.C(n_395),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_423),
.B(n_392),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_429),
.B(n_400),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_471),
.B(n_474),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_SL g474 ( 
.A(n_424),
.B(n_408),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_436),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_430),
.B(n_400),
.C(n_384),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_476),
.B(n_422),
.C(n_425),
.Y(n_499)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_462),
.Y(n_481)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_481),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_477),
.B(n_426),
.Y(n_482)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_482),
.Y(n_522)
);

MAJx2_ASAP7_75t_L g483 ( 
.A(n_456),
.B(n_453),
.C(n_459),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_483),
.B(n_499),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_476),
.A2(n_419),
.B1(n_435),
.B2(n_443),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_484),
.A2(n_490),
.B1(n_495),
.B2(n_496),
.Y(n_507)
);

FAx1_ASAP7_75t_L g485 ( 
.A(n_457),
.B(n_417),
.CI(n_446),
.CON(n_485),
.SN(n_485)
);

A2O1A1Ixp33_ASAP7_75t_SL g515 ( 
.A1(n_485),
.A2(n_452),
.B(n_417),
.C(n_425),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_477),
.B(n_428),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_486),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_465),
.B(n_439),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_488),
.B(n_491),
.Y(n_517)
);

BUFx24_ASAP7_75t_SL g491 ( 
.A(n_454),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_465),
.B(n_439),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_492),
.Y(n_521)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_462),
.Y(n_493)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_493),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_461),
.B(n_432),
.Y(n_494)
);

AO221x1_ASAP7_75t_L g518 ( 
.A1(n_494),
.A2(n_498),
.B1(n_468),
.B2(n_442),
.C(n_460),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_450),
.B(n_447),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_450),
.B(n_448),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_463),
.A2(n_437),
.B1(n_428),
.B2(n_418),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_497),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_449),
.B(n_404),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_471),
.B(n_422),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_500),
.B(n_467),
.Y(n_503)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_451),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_501),
.A2(n_502),
.B1(n_463),
.B2(n_466),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_475),
.B(n_382),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_503),
.B(n_509),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_480),
.A2(n_473),
.B(n_452),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_504),
.A2(n_518),
.B(n_466),
.Y(n_524)
);

INVxp33_ASAP7_75t_L g505 ( 
.A(n_482),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_505),
.B(n_510),
.Y(n_536)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_508),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_478),
.B(n_446),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_481),
.A2(n_493),
.B1(n_480),
.B2(n_486),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_478),
.B(n_457),
.C(n_472),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_513),
.B(n_514),
.C(n_519),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_489),
.B(n_472),
.C(n_452),
.Y(n_514)
);

AO21x1_ASAP7_75t_L g531 ( 
.A1(n_515),
.A2(n_485),
.B(n_420),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_489),
.B(n_468),
.C(n_442),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_524),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_506),
.B(n_483),
.C(n_499),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_525),
.B(n_529),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_519),
.B(n_484),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_526),
.B(n_531),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_507),
.A2(n_397),
.B1(n_501),
.B2(n_460),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_528),
.A2(n_538),
.B1(n_522),
.B2(n_511),
.Y(n_548)
);

OAI21x1_ASAP7_75t_L g529 ( 
.A1(n_517),
.A2(n_487),
.B(n_418),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_506),
.B(n_490),
.C(n_479),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_530),
.B(n_533),
.Y(n_547)
);

BUFx24_ASAP7_75t_SL g532 ( 
.A(n_504),
.Y(n_532)
);

BUFx24_ASAP7_75t_SL g539 ( 
.A(n_532),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_521),
.B(n_464),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_514),
.B(n_479),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_535),
.B(n_537),
.Y(n_543)
);

NOR2xp67_ASAP7_75t_L g537 ( 
.A(n_503),
.B(n_500),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_512),
.B(n_431),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_527),
.A2(n_513),
.B1(n_512),
.B2(n_505),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_540),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_523),
.B(n_509),
.C(n_515),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_542),
.B(n_545),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_523),
.B(n_515),
.C(n_516),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_536),
.A2(n_522),
.B1(n_511),
.B2(n_520),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g556 ( 
.A1(n_546),
.A2(n_550),
.B1(n_515),
.B2(n_438),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_548),
.A2(n_549),
.B1(n_414),
.B2(n_441),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_531),
.A2(n_510),
.B1(n_437),
.B2(n_516),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_530),
.A2(n_444),
.B1(n_414),
.B2(n_445),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_547),
.B(n_545),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_552),
.B(n_553),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_541),
.B(n_525),
.C(n_526),
.Y(n_553)
);

BUFx4f_ASAP7_75t_SL g554 ( 
.A(n_540),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_554),
.B(n_557),
.Y(n_567)
);

OAI21x1_ASAP7_75t_L g555 ( 
.A1(n_543),
.A2(n_535),
.B(n_534),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_L g568 ( 
.A1(n_555),
.A2(n_560),
.B(n_558),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_556),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_542),
.B(n_534),
.C(n_444),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_559),
.B(n_551),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_544),
.B(n_414),
.C(n_474),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_561),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_562),
.B(n_565),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_L g564 ( 
.A1(n_558),
.A2(n_544),
.B(n_551),
.Y(n_564)
);

AO21x1_ASAP7_75t_L g573 ( 
.A1(n_564),
.A2(n_567),
.B(n_563),
.Y(n_573)
);

OAI21xp33_ASAP7_75t_L g566 ( 
.A1(n_554),
.A2(n_539),
.B(n_485),
.Y(n_566)
);

NOR2xp67_ASAP7_75t_L g571 ( 
.A(n_566),
.B(n_554),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g570 ( 
.A(n_568),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_571),
.B(n_573),
.C(n_440),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g574 ( 
.A(n_567),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_574),
.B(n_569),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_SL g579 ( 
.A1(n_575),
.A2(n_576),
.B(n_399),
.Y(n_579)
);

BUFx24_ASAP7_75t_SL g576 ( 
.A(n_570),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_577),
.A2(n_572),
.B1(n_427),
.B2(n_421),
.Y(n_578)
);

AOI21x1_ASAP7_75t_L g580 ( 
.A1(n_578),
.A2(n_579),
.B(n_399),
.Y(n_580)
);

MAJx2_ASAP7_75t_L g581 ( 
.A(n_580),
.B(n_323),
.C(n_355),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_581),
.B(n_323),
.Y(n_582)
);


endmodule