module fake_aes_3407_n_36 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_36);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_36;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
OAI22x1_ASAP7_75t_R g11 ( .A1(n_7), .A2(n_6), .B1(n_8), .B2(n_5), .Y(n_11) );
OA21x2_ASAP7_75t_L g12 ( .A1(n_2), .A2(n_6), .B(n_0), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_9), .Y(n_13) );
INVxp67_ASAP7_75t_L g14 ( .A(n_0), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_5), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_15), .Y(n_16) );
BUFx3_ASAP7_75t_L g17 ( .A(n_12), .Y(n_17) );
INVx2_ASAP7_75t_SL g18 ( .A(n_15), .Y(n_18) );
OAI21x1_ASAP7_75t_L g19 ( .A1(n_16), .A2(n_12), .B(n_10), .Y(n_19) );
OAI21x1_ASAP7_75t_L g20 ( .A1(n_16), .A2(n_12), .B(n_14), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_19), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_19), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_21), .B(n_13), .Y(n_23) );
OR2x2_ASAP7_75t_L g24 ( .A(n_22), .B(n_13), .Y(n_24) );
INVxp67_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
NAND4xp25_ASAP7_75t_L g26 ( .A(n_23), .B(n_14), .C(n_11), .D(n_16), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
AOI221xp5_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_18), .B1(n_17), .B2(n_11), .C(n_12), .Y(n_28) );
OAI322xp33_ASAP7_75t_L g29 ( .A1(n_25), .A2(n_18), .A3(n_12), .B1(n_3), .B2(n_4), .C1(n_7), .C2(n_8), .Y(n_29) );
INVxp33_ASAP7_75t_SL g30 ( .A(n_28), .Y(n_30) );
NAND4xp25_ASAP7_75t_L g31 ( .A(n_27), .B(n_17), .C(n_2), .D(n_3), .Y(n_31) );
INVx2_ASAP7_75t_SL g32 ( .A(n_29), .Y(n_32) );
AOI21xp5_ASAP7_75t_L g33 ( .A1(n_31), .A2(n_20), .B(n_17), .Y(n_33) );
NOR2xp33_ASAP7_75t_L g34 ( .A(n_30), .B(n_12), .Y(n_34) );
AOI22xp33_ASAP7_75t_SL g35 ( .A1(n_34), .A2(n_32), .B1(n_20), .B2(n_9), .Y(n_35) );
AOI22x1_ASAP7_75t_L g36 ( .A1(n_35), .A2(n_33), .B1(n_1), .B2(n_4), .Y(n_36) );
endmodule