module real_jpeg_12766_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_0),
.Y(n_99)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_3),
.A2(n_58),
.B1(n_59),
.B2(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_62),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_3),
.A2(n_28),
.B1(n_31),
.B2(n_62),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_3),
.A2(n_42),
.B1(n_47),
.B2(n_62),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_4),
.A2(n_58),
.B1(n_59),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_4),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_67),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_4),
.A2(n_28),
.B1(n_31),
.B2(n_67),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_4),
.A2(n_42),
.B1(n_47),
.B2(n_67),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_5),
.A2(n_36),
.B1(n_58),
.B2(n_59),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_5),
.A2(n_28),
.B1(n_31),
.B2(n_36),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_5),
.A2(n_36),
.B1(n_42),
.B2(n_47),
.Y(n_135)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_7),
.A2(n_58),
.B1(n_59),
.B2(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_7),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_172),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_7),
.A2(n_28),
.B1(n_31),
.B2(n_172),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_7),
.A2(n_42),
.B1(n_47),
.B2(n_172),
.Y(n_277)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_9),
.Y(n_191)
);

AOI21xp33_ASAP7_75t_L g209 ( 
.A1(n_9),
.A2(n_58),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_9),
.B(n_82),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_9),
.B(n_33),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_L g262 ( 
.A1(n_9),
.A2(n_28),
.B1(n_31),
.B2(n_191),
.Y(n_262)
);

O2A1O1Ixp33_ASAP7_75t_L g264 ( 
.A1(n_9),
.A2(n_31),
.B(n_46),
.C(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_9),
.B(n_73),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_9),
.B(n_99),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_9),
.B(n_40),
.Y(n_289)
);

AOI21xp33_ASAP7_75t_L g298 ( 
.A1(n_9),
.A2(n_33),
.B(n_248),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_10),
.A2(n_58),
.B1(n_59),
.B2(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_10),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_199),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_10),
.A2(n_28),
.B1(n_31),
.B2(n_199),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_10),
.A2(n_42),
.B1(n_47),
.B2(n_199),
.Y(n_284)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_12),
.A2(n_58),
.B1(n_59),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_12),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_12),
.A2(n_33),
.B1(n_34),
.B2(n_107),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_12),
.A2(n_28),
.B1(n_31),
.B2(n_107),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_12),
.A2(n_42),
.B1(n_47),
.B2(n_107),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_13),
.A2(n_58),
.B1(n_59),
.B2(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_13),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_13),
.A2(n_33),
.B1(n_34),
.B2(n_144),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_13),
.A2(n_28),
.B1(n_31),
.B2(n_144),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_13),
.A2(n_42),
.B1(n_47),
.B2(n_144),
.Y(n_272)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_15),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_15),
.A2(n_28),
.B1(n_31),
.B2(n_38),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_15),
.A2(n_38),
.B1(n_42),
.B2(n_47),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_16),
.A2(n_58),
.B1(n_59),
.B2(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_16),
.A2(n_33),
.B1(n_34),
.B2(n_64),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_16),
.A2(n_28),
.B1(n_31),
.B2(n_64),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_16),
.A2(n_42),
.B1(n_47),
.B2(n_64),
.Y(n_163)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_88),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_86),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_74),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_21),
.B(n_74),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_65),
.C(n_68),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_22),
.A2(n_65),
.B1(n_115),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_22),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_52),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_39),
.B2(n_51),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_25),
.B(n_39),
.C(n_52),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_35),
.B2(n_37),
.Y(n_25)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_26),
.A2(n_27),
.B1(n_113),
.B2(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_26),
.A2(n_27),
.B1(n_141),
.B2(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_26),
.A2(n_27),
.B1(n_194),
.B2(n_213),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_26),
.A2(n_27),
.B1(n_223),
.B2(n_298),
.Y(n_297)
);

NAND2x1_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_32),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_27),
.Y(n_73)
);

OA22x2_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_27)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_28),
.A2(n_31),
.B1(n_45),
.B2(n_46),
.Y(n_49)
);

OAI32xp33_ASAP7_75t_L g246 ( 
.A1(n_28),
.A2(n_30),
.A3(n_33),
.B1(n_247),
.B2(n_249),
.Y(n_246)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_29),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_29),
.B(n_31),
.Y(n_249)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_33),
.A2(n_34),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_33),
.B(n_55),
.Y(n_189)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI32xp33_ASAP7_75t_L g188 ( 
.A1(n_34),
.A2(n_56),
.A3(n_58),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_35),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_37),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_39),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_65),
.C(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_39),
.A2(n_51),
.B1(n_69),
.B2(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_48),
.B(n_50),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_40),
.A2(n_48),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_40),
.A2(n_48),
.B1(n_50),
.B2(n_104),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_40),
.A2(n_48),
.B1(n_103),
.B2(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_40),
.A2(n_48),
.B1(n_166),
.B2(n_215),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_40),
.A2(n_48),
.B1(n_215),
.B2(n_241),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_40),
.A2(n_48),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_40),
.A2(n_48),
.B1(n_263),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_41),
.A2(n_139),
.B1(n_165),
.B2(n_167),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_41),
.A2(n_167),
.B1(n_242),
.B2(n_300),
.Y(n_299)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_41)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_42),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_42),
.B(n_286),
.Y(n_285)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp33_ASAP7_75t_L g265 ( 
.A1(n_45),
.A2(n_47),
.B(n_191),
.Y(n_265)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_48),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_61),
.B2(n_63),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_53),
.A2(n_54),
.B1(n_61),
.B2(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_53),
.A2(n_54),
.B1(n_66),
.B2(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_53),
.A2(n_54),
.B1(n_106),
.B2(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_53),
.A2(n_54),
.B1(n_143),
.B2(n_171),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_53),
.A2(n_54),
.B1(n_198),
.B2(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_54),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_59),
.B(n_191),
.Y(n_190)
);

BUFx16f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_63),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_65),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_68),
.B(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_70),
.A2(n_71),
.B1(n_73),
.B2(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_71),
.A2(n_73),
.B(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_71),
.A2(n_73),
.B1(n_193),
.B2(n_195),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_71),
.A2(n_73),
.B1(n_222),
.B2(n_224),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_85),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_78),
.B1(n_83),
.B2(n_84),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_76),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_80),
.A2(n_82),
.B1(n_197),
.B2(n_200),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AO21x1_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_150),
.B(n_320),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_145),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_121),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_91),
.B(n_121),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_108),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_92),
.B(n_114),
.C(n_119),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_96),
.B(n_105),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_93),
.A2(n_94),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_101),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_95),
.A2(n_96),
.B1(n_105),
.B2(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_95),
.A2(n_96),
.B1(n_101),
.B2(n_102),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_99),
.B(n_100),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_97),
.A2(n_99),
.B1(n_100),
.B2(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_97),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_97),
.A2(n_99),
.B1(n_163),
.B2(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_97),
.A2(n_99),
.B1(n_187),
.B2(n_227),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_97),
.A2(n_99),
.B1(n_227),
.B2(n_251),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_97),
.A2(n_99),
.B1(n_251),
.B2(n_272),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_97),
.A2(n_99),
.B1(n_191),
.B2(n_284),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_97),
.A2(n_99),
.B1(n_277),
.B2(n_284),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_98),
.A2(n_135),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_98),
.A2(n_161),
.B1(n_276),
.B2(n_278),
.Y(n_275)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_114),
.B1(n_119),
.B2(n_120),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_109),
.Y(n_119)
);

OAI21xp33_ASAP7_75t_L g128 ( 
.A1(n_109),
.A2(n_110),
.B(n_111),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_127),
.C(n_129),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_122),
.A2(n_123),
.B1(n_127),
.B2(n_128),
.Y(n_174)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_140),
.C(n_142),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_131),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_136),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_132),
.A2(n_133),
.B1(n_136),
.B2(n_137),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_142),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_145),
.A2(n_321),
.B(n_322),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_146),
.B(n_147),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_175),
.B(n_319),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_173),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_152),
.B(n_173),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.C(n_157),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_153),
.B(n_156),
.Y(n_202)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_157),
.B(n_202),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_168),
.C(n_170),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_158),
.A2(n_159),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_160),
.B(n_164),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_170),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_169),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_171),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_203),
.B(n_318),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_201),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_177),
.B(n_201),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_182),
.C(n_183),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_178),
.A2(n_179),
.B1(n_182),
.B2(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_182),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_183),
.B(n_315),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_192),
.C(n_196),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_184),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_188),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_185),
.A2(n_186),
.B1(n_188),
.B2(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_190),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_192),
.B(n_196),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

A2O1A1Ixp33_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_234),
.B(n_312),
.C(n_317),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_228),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_205),
.B(n_228),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_218),
.C(n_220),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_206),
.A2(n_207),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_212),
.C(n_217),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_214),
.B1(n_216),
.B2(n_217),
.Y(n_211)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_212),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_213),
.Y(n_224)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_214),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_218),
.B(n_220),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_225),
.C(n_226),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_221),
.B(n_239),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_226),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_232),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_230),
.B(n_231),
.C(n_232),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_311),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_255),
.B(n_310),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_252),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_237),
.B(n_252),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_240),
.C(n_243),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_238),
.B(n_307),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_240),
.A2(n_243),
.B1(n_244),
.B2(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_240),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_250),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_245),
.A2(n_246),
.B1(n_250),
.B2(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_250),
.Y(n_302)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_253),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_304),
.B(n_309),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_293),
.B(n_303),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_273),
.B(n_292),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_266),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_259),
.B(n_266),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_264),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_260),
.A2(n_261),
.B1(n_264),
.B2(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_264),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_271),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_268),
.B(n_269),
.C(n_271),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_270),
.Y(n_300)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_272),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_281),
.B(n_291),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_279),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_275),
.B(n_279),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_287),
.B(n_290),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_285),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_288),
.B(n_289),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_294),
.B(n_295),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_301),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_299),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_299),
.C(n_301),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_305),
.B(n_306),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_314),
.Y(n_317)
);


endmodule