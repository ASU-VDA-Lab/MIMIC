module real_aes_4835_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_919;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_918;
wire n_356;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_906;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_693;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_617;
wire n_602;
wire n_139;
wire n_402;
wire n_552;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_898;
wire n_115;
wire n_604;
wire n_110;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_288;
wire n_147;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_193;
wire n_397;
wire n_162;
wire n_293;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_899;
wire n_526;
wire n_637;
wire n_155;
wire n_653;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_103;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_237;
wire n_797;
wire n_862;
NAND2xp5_ASAP7_75t_L g637 ( .A(n_0), .B(n_202), .Y(n_637) );
CKINVDCx5p33_ASAP7_75t_R g651 ( .A(n_1), .Y(n_651) );
CKINVDCx5p33_ASAP7_75t_R g532 ( .A(n_2), .Y(n_532) );
INVx1_ASAP7_75t_L g300 ( .A(n_3), .Y(n_300) );
O2A1O1Ixp33_ASAP7_75t_SL g580 ( .A1(n_4), .A2(n_180), .B(n_581), .C(n_582), .Y(n_580) );
OAI22xp33_ASAP7_75t_L g642 ( .A1(n_5), .A2(n_80), .B1(n_144), .B2(n_172), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_6), .B(n_166), .Y(n_250) );
INVxp67_ASAP7_75t_L g108 ( .A(n_7), .Y(n_108) );
INVx1_ASAP7_75t_L g547 ( .A(n_7), .Y(n_547) );
INVx1_ASAP7_75t_L g898 ( .A(n_7), .Y(n_898) );
BUFx2_ASAP7_75t_L g920 ( .A(n_7), .Y(n_920) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_8), .B(n_252), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g216 ( .A1(n_9), .A2(n_36), .B1(n_165), .B2(n_217), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g127 ( .A1(n_10), .A2(n_41), .B1(n_128), .B2(n_132), .Y(n_127) );
AOI22xp5_ASAP7_75t_L g272 ( .A1(n_11), .A2(n_63), .B1(n_142), .B2(n_265), .Y(n_272) );
INVx1_ASAP7_75t_L g295 ( .A(n_12), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g670 ( .A(n_13), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_14), .A2(n_70), .B1(n_130), .B2(n_172), .Y(n_560) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_15), .Y(n_571) );
INVx1_ASAP7_75t_L g298 ( .A(n_16), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_17), .A2(n_59), .B1(n_144), .B2(n_176), .Y(n_559) );
OA21x2_ASAP7_75t_L g150 ( .A1(n_18), .A2(n_69), .B(n_151), .Y(n_150) );
OA21x2_ASAP7_75t_L g159 ( .A1(n_18), .A2(n_69), .B(n_151), .Y(n_159) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_19), .A2(n_66), .B1(n_142), .B2(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g292 ( .A(n_20), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g666 ( .A(n_21), .Y(n_666) );
BUFx3_ASAP7_75t_L g537 ( .A(n_22), .Y(n_537) );
BUFx8_ASAP7_75t_SL g911 ( .A(n_22), .Y(n_911) );
O2A1O1Ixp33_ASAP7_75t_L g586 ( .A1(n_23), .A2(n_271), .B(n_587), .C(n_588), .Y(n_586) );
OAI22xp33_ASAP7_75t_SL g640 ( .A1(n_24), .A2(n_45), .B1(n_134), .B2(n_144), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_25), .A2(n_34), .B1(n_134), .B2(n_248), .Y(n_630) );
AO22x1_ASAP7_75t_L g245 ( .A1(n_26), .A2(n_76), .B1(n_178), .B2(n_246), .Y(n_245) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_27), .Y(n_169) );
AND2x2_ASAP7_75t_L g188 ( .A(n_28), .B(n_132), .Y(n_188) );
OAI22xp5_ASAP7_75t_L g114 ( .A1(n_29), .A2(n_115), .B1(n_116), .B2(n_117), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_29), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_30), .B(n_178), .Y(n_177) );
O2A1O1Ixp5_ASAP7_75t_L g601 ( .A1(n_31), .A2(n_180), .B(n_602), .C(n_603), .Y(n_601) );
INVx1_ASAP7_75t_L g113 ( .A(n_32), .Y(n_113) );
AOI22x1_ASAP7_75t_L g139 ( .A1(n_33), .A2(n_94), .B1(n_140), .B2(n_142), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_35), .B(n_148), .Y(n_220) );
AND2x2_ASAP7_75t_L g918 ( .A(n_37), .B(n_919), .Y(n_918) );
CKINVDCx5p33_ASAP7_75t_R g604 ( .A(n_38), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_39), .B(n_617), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_40), .B(n_196), .Y(n_195) );
CKINVDCx5p33_ASAP7_75t_R g584 ( .A(n_42), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_43), .B(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_44), .B(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g151 ( .A(n_46), .Y(n_151) );
AND2x4_ASAP7_75t_L g153 ( .A(n_47), .B(n_154), .Y(n_153) );
AND2x4_ASAP7_75t_L g592 ( .A(n_47), .B(n_154), .Y(n_592) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_48), .Y(n_138) );
INVx2_ASAP7_75t_L g267 ( .A(n_49), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g649 ( .A(n_50), .Y(n_649) );
CKINVDCx5p33_ASAP7_75t_R g609 ( .A(n_51), .Y(n_609) );
INVx2_ASAP7_75t_L g575 ( .A(n_52), .Y(n_575) );
O2A1O1Ixp33_ASAP7_75t_L g667 ( .A1(n_53), .A2(n_180), .B(n_668), .C(n_669), .Y(n_667) );
CKINVDCx5p33_ASAP7_75t_R g648 ( .A(n_54), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_55), .A2(n_100), .B1(n_912), .B2(n_921), .Y(n_99) );
AOI22xp33_ASAP7_75t_L g213 ( .A1(n_56), .A2(n_72), .B1(n_140), .B2(n_165), .Y(n_213) );
CKINVDCx14_ASAP7_75t_R g254 ( .A(n_57), .Y(n_254) );
AND2x2_ASAP7_75t_L g193 ( .A(n_58), .B(n_178), .Y(n_193) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_60), .A2(n_78), .B1(n_129), .B2(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_61), .B(n_226), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_62), .B(n_236), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g652 ( .A(n_64), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_65), .B(n_226), .Y(n_225) );
NAND2xp33_ASAP7_75t_R g562 ( .A(n_67), .B(n_150), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_67), .A2(n_97), .B1(n_288), .B2(n_617), .Y(n_748) );
NAND2x1p5_ASAP7_75t_L g197 ( .A(n_68), .B(n_184), .Y(n_197) );
CKINVDCx14_ASAP7_75t_R g156 ( .A(n_71), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_73), .B(n_166), .Y(n_231) );
OR2x6_ASAP7_75t_L g110 ( .A(n_74), .B(n_111), .Y(n_110) );
AND3x1_ASAP7_75t_L g917 ( .A(n_74), .B(n_918), .C(n_920), .Y(n_917) );
CKINVDCx5p33_ASAP7_75t_R g574 ( .A(n_75), .Y(n_574) );
CKINVDCx5p33_ASAP7_75t_R g572 ( .A(n_77), .Y(n_572) );
INVx1_ASAP7_75t_L g112 ( .A(n_79), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g916 ( .A(n_79), .B(n_113), .Y(n_916) );
INVx1_ASAP7_75t_L g919 ( .A(n_81), .Y(n_919) );
INVx1_ASAP7_75t_L g131 ( .A(n_82), .Y(n_131) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_82), .Y(n_135) );
BUFx5_ASAP7_75t_L g144 ( .A(n_82), .Y(n_144) );
INVx2_ASAP7_75t_L g594 ( .A(n_83), .Y(n_594) );
INVx2_ASAP7_75t_L g302 ( .A(n_84), .Y(n_302) );
INVx2_ASAP7_75t_L g672 ( .A(n_85), .Y(n_672) );
CKINVDCx5p33_ASAP7_75t_R g589 ( .A(n_86), .Y(n_589) );
AOI221xp5_ASAP7_75t_L g540 ( .A1(n_87), .A2(n_541), .B1(n_542), .B2(n_899), .C(n_906), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_87), .Y(n_541) );
NAND2xp33_ASAP7_75t_L g190 ( .A(n_88), .B(n_141), .Y(n_190) );
CKINVDCx5p33_ASAP7_75t_R g907 ( .A(n_89), .Y(n_907) );
INVx2_ASAP7_75t_SL g154 ( .A(n_90), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_91), .B(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_92), .B(n_196), .Y(n_230) );
INVx1_ASAP7_75t_L g607 ( .A(n_93), .Y(n_607) );
INVx2_ASAP7_75t_L g612 ( .A(n_95), .Y(n_612) );
OAI21xp33_ASAP7_75t_SL g664 ( .A1(n_96), .A2(n_144), .B(n_665), .Y(n_664) );
INVxp67_ASAP7_75t_SL g577 ( .A(n_97), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_97), .B(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_98), .B(n_182), .Y(n_181) );
OR2x2_ASAP7_75t_L g100 ( .A(n_101), .B(n_538), .Y(n_100) );
NOR2xp33_ASAP7_75t_L g101 ( .A(n_102), .B(n_536), .Y(n_101) );
AOI21xp5_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_114), .B(n_531), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
BUFx8_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
BUFx12f_ASAP7_75t_L g535 ( .A(n_106), .Y(n_535) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
OR2x6_ASAP7_75t_L g897 ( .A(n_109), .B(n_898), .Y(n_897) );
INVx8_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_L g546 ( .A(n_110), .B(n_547), .Y(n_546) );
OR2x6_ASAP7_75t_L g909 ( .A(n_110), .B(n_547), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
BUFx3_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_118), .A2(n_543), .B1(n_548), .B2(n_897), .Y(n_542) );
INVx1_ASAP7_75t_L g904 ( .A(n_118), .Y(n_904) );
AND2x4_ASAP7_75t_L g118 ( .A(n_119), .B(n_420), .Y(n_118) );
NOR3xp33_ASAP7_75t_L g119 ( .A(n_120), .B(n_344), .C(n_390), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_310), .Y(n_120) );
AOI21xp33_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_221), .B(n_255), .Y(n_121) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_160), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_123), .B(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_124), .B(n_318), .Y(n_506) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND2x4_ASAP7_75t_L g277 ( .A(n_125), .B(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g386 ( .A(n_125), .B(n_186), .Y(n_386) );
AND2x2_ASAP7_75t_L g482 ( .A(n_125), .B(n_186), .Y(n_482) );
AO31x2_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_147), .A3(n_152), .B(n_155), .Y(n_125) );
AO31x2_ASAP7_75t_L g323 ( .A1(n_126), .A2(n_147), .A3(n_152), .B(n_155), .Y(n_323) );
OAI22x1_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_136), .B1(n_139), .B2(n_145), .Y(n_126) );
INVx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g581 ( .A(n_129), .Y(n_581) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g248 ( .A(n_131), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_132), .B(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g141 ( .A(n_134), .Y(n_141) );
INVx1_ASAP7_75t_L g196 ( .A(n_134), .Y(n_196) );
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_134), .A2(n_144), .B1(n_571), .B2(n_572), .Y(n_570) );
INVx2_ASAP7_75t_L g583 ( .A(n_134), .Y(n_583) );
INVx2_ASAP7_75t_SL g632 ( .A(n_134), .Y(n_632) );
AOI22xp33_ASAP7_75t_SL g647 ( .A1(n_134), .A2(n_144), .B1(n_648), .B2(n_649), .Y(n_647) );
INVx6_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g172 ( .A(n_135), .Y(n_172) );
INVx2_ASAP7_75t_L g176 ( .A(n_135), .Y(n_176) );
INVx3_ASAP7_75t_L g219 ( .A(n_135), .Y(n_219) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_137), .B(n_211), .Y(n_215) );
OA22x2_ASAP7_75t_L g629 ( .A1(n_137), .A2(n_146), .B1(n_630), .B2(n_631), .Y(n_629) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_138), .Y(n_146) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_138), .Y(n_180) );
INVxp67_ASAP7_75t_L g191 ( .A(n_138), .Y(n_191) );
INVx4_ASAP7_75t_L g262 ( .A(n_138), .Y(n_262) );
INVx3_ASAP7_75t_L g271 ( .A(n_138), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_138), .B(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_138), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_138), .B(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_SL g639 ( .A(n_138), .B(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g166 ( .A(n_144), .Y(n_166) );
INVx2_ASAP7_75t_L g178 ( .A(n_144), .Y(n_178) );
INVx2_ASAP7_75t_L g236 ( .A(n_144), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_144), .B(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_144), .B(n_609), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_144), .A2(n_176), .B1(n_651), .B2(n_652), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g665 ( .A(n_144), .B(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_145), .B(n_168), .Y(n_167) );
INVx4_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
OAI22xp5_ASAP7_75t_L g164 ( .A1(n_146), .A2(n_165), .B1(n_167), .B2(n_170), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_146), .B(n_211), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_146), .A2(n_230), .B(n_231), .Y(n_229) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_150), .B(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g263 ( .A(n_150), .Y(n_263) );
BUFx3_ASAP7_75t_L g568 ( .A(n_150), .Y(n_568) );
INVx1_ASAP7_75t_L g613 ( .A(n_150), .Y(n_613) );
INVx1_ASAP7_75t_L g662 ( .A(n_150), .Y(n_662) );
OAI21x1_ASAP7_75t_L g163 ( .A1(n_152), .A2(n_164), .B(n_173), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_152), .B(n_567), .Y(n_566) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx3_ASAP7_75t_L g204 ( .A(n_153), .Y(n_204) );
INVx3_ASAP7_75t_L g212 ( .A(n_153), .Y(n_212) );
INVx1_ASAP7_75t_L g242 ( .A(n_153), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_153), .B(n_185), .Y(n_643) );
OAI221xp5_ASAP7_75t_L g646 ( .A1(n_153), .A2(n_180), .B1(n_271), .B2(n_647), .C(n_650), .Y(n_646) );
NOR2xp67_ASAP7_75t_SL g155 ( .A(n_156), .B(n_157), .Y(n_155) );
OR2x2_ASAP7_75t_L g253 ( .A(n_157), .B(n_254), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g692 ( .A1(n_157), .A2(n_693), .B(n_694), .Y(n_692) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_158), .A2(n_163), .B(n_181), .Y(n_162) );
OA21x2_ASAP7_75t_L g282 ( .A1(n_158), .A2(n_163), .B(n_181), .Y(n_282) );
BUFx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx4_ASAP7_75t_L g185 ( .A(n_159), .Y(n_185) );
INVx2_ASAP7_75t_L g227 ( .A(n_159), .Y(n_227) );
AND2x2_ASAP7_75t_L g160 ( .A(n_161), .B(n_206), .Y(n_160) );
INVx2_ASAP7_75t_L g383 ( .A(n_161), .Y(n_383) );
AND2x2_ASAP7_75t_L g161 ( .A(n_162), .B(n_186), .Y(n_161) );
NAND2x1_ASAP7_75t_L g356 ( .A(n_162), .B(n_322), .Y(n_356) );
AND2x2_ASAP7_75t_L g397 ( .A(n_162), .B(n_208), .Y(n_397) );
AND2x2_ASAP7_75t_L g402 ( .A(n_162), .B(n_309), .Y(n_402) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_177), .B(n_179), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_175), .B(n_294), .Y(n_293) );
AOI22xp5_ASAP7_75t_L g296 ( .A1(n_175), .A2(n_178), .B1(n_297), .B2(n_299), .Y(n_296) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_176), .A2(n_248), .B1(n_574), .B2(n_575), .Y(n_573) );
INVx1_ASAP7_75t_L g587 ( .A(n_176), .Y(n_587) );
INVxp67_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_SL g199 ( .A(n_180), .Y(n_199) );
INVx1_ASAP7_75t_L g237 ( .A(n_180), .Y(n_237) );
INVx1_ASAP7_75t_L g244 ( .A(n_180), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_180), .A2(n_262), .B1(n_559), .B2(n_560), .Y(n_558) );
OAI22xp33_ASAP7_75t_L g569 ( .A1(n_180), .A2(n_262), .B1(n_570), .B2(n_573), .Y(n_569) );
OR2x2_ASAP7_75t_L g241 ( .A(n_182), .B(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
OR2x2_ASAP7_75t_L g266 ( .A(n_183), .B(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx3_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g202 ( .A(n_185), .Y(n_202) );
NOR2xp33_ASAP7_75t_SL g593 ( .A(n_185), .B(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g617 ( .A(n_185), .Y(n_617) );
AND2x4_ASAP7_75t_L g373 ( .A(n_186), .B(n_318), .Y(n_373) );
AO21x2_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_192), .B(n_200), .Y(n_186) );
AO21x2_ASAP7_75t_L g279 ( .A1(n_187), .A2(n_192), .B(n_200), .Y(n_279) );
OAI21x1_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_191), .Y(n_187) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
OAI21x1_ASAP7_75t_SL g192 ( .A1(n_193), .A2(n_194), .B(n_198), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_195), .B(n_197), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_197), .B(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g205 ( .A(n_197), .Y(n_205) );
AOI21x1_ASAP7_75t_L g249 ( .A1(n_199), .A2(n_250), .B(n_251), .Y(n_249) );
AOI21xp33_ASAP7_75t_SL g200 ( .A1(n_201), .A2(n_203), .B(n_205), .Y(n_200) );
OR2x2_ASAP7_75t_L g576 ( .A(n_201), .B(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g645 ( .A(n_201), .Y(n_645) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NOR2xp33_ASAP7_75t_SL g590 ( .A(n_202), .B(n_591), .Y(n_590) );
NAND3xp33_ASAP7_75t_SL g261 ( .A(n_203), .B(n_262), .C(n_263), .Y(n_261) );
NAND3xp33_ASAP7_75t_L g269 ( .A(n_203), .B(n_263), .C(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
NOR2x1_ASAP7_75t_L g238 ( .A(n_204), .B(n_226), .Y(n_238) );
INVx1_ASAP7_75t_L g478 ( .A(n_206), .Y(n_478) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g347 ( .A(n_207), .Y(n_347) );
OR2x2_ASAP7_75t_L g442 ( .A(n_207), .B(n_356), .Y(n_442) );
AND2x2_ASAP7_75t_L g450 ( .A(n_207), .B(n_321), .Y(n_450) );
INVx2_ASAP7_75t_SL g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_214), .Y(n_208) );
NAND2x1p5_ASAP7_75t_L g309 ( .A(n_209), .B(n_214), .Y(n_309) );
OR2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_213), .Y(n_209) );
OA21x2_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_216), .B(n_220), .Y(n_214) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g265 ( .A(n_218), .Y(n_265) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx2_ASAP7_75t_L g234 ( .A(n_219), .Y(n_234) );
INVx1_ASAP7_75t_L g252 ( .A(n_219), .Y(n_252) );
INVx1_ASAP7_75t_L g602 ( .A(n_219), .Y(n_602) );
INVx1_ASAP7_75t_L g668 ( .A(n_219), .Y(n_668) );
AOI32xp33_ASAP7_75t_L g446 ( .A1(n_221), .A2(n_443), .A3(n_447), .B1(n_449), .B2(n_450), .Y(n_446) );
AOI221x1_ASAP7_75t_L g464 ( .A1(n_221), .A2(n_465), .B1(n_468), .B2(n_470), .C(n_471), .Y(n_464) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
OR2x2_ASAP7_75t_L g332 ( .A(n_222), .B(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g475 ( .A(n_223), .B(n_363), .Y(n_475) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_239), .Y(n_223) );
INVx3_ASAP7_75t_L g275 ( .A(n_224), .Y(n_275) );
INVx2_ASAP7_75t_L g362 ( .A(n_224), .Y(n_362) );
AND2x2_ASAP7_75t_L g377 ( .A(n_224), .B(n_240), .Y(n_377) );
AND2x4_ASAP7_75t_L g224 ( .A(n_225), .B(n_228), .Y(n_224) );
NOR2xp67_ASAP7_75t_L g561 ( .A(n_226), .B(n_242), .Y(n_561) );
INVx3_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_227), .B(n_302), .Y(n_301) );
BUFx3_ASAP7_75t_L g610 ( .A(n_227), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_227), .B(n_672), .Y(n_671) );
OAI21x1_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_232), .B(n_238), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_235), .B(n_237), .Y(n_232) );
AOI221xp5_ASAP7_75t_L g619 ( .A1(n_237), .A2(n_591), .B1(n_620), .B2(n_621), .C(n_622), .Y(n_619) );
INVx1_ASAP7_75t_L g303 ( .A(n_239), .Y(n_303) );
INVx1_ASAP7_75t_L g330 ( .A(n_239), .Y(n_330) );
AND2x2_ASAP7_75t_L g438 ( .A(n_239), .B(n_286), .Y(n_438) );
INVx2_ASAP7_75t_SL g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g274 ( .A(n_240), .B(n_275), .Y(n_274) );
OAI21x1_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_243), .B(n_253), .Y(n_240) );
OAI21xp5_ASAP7_75t_L g343 ( .A1(n_241), .A2(n_243), .B(n_253), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_242), .B(n_288), .Y(n_287) );
AOI21x1_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_245), .B(n_249), .Y(n_243) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_248), .B(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g669 ( .A(n_248), .B(n_670), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_252), .A2(n_262), .B1(n_606), .B2(n_608), .Y(n_605) );
OAI22xp33_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_276), .B1(n_283), .B2(n_304), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_256), .A2(n_366), .B1(n_469), .B2(n_500), .Y(n_499) );
OR2x2_ASAP7_75t_SL g256 ( .A(n_257), .B(n_273), .Y(n_256) );
OR2x2_ASAP7_75t_L g350 ( .A(n_257), .B(n_328), .Y(n_350) );
INVx2_ASAP7_75t_L g448 ( .A(n_257), .Y(n_448) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g520 ( .A(n_258), .B(n_341), .Y(n_520) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NOR2x1_ASAP7_75t_L g314 ( .A(n_259), .B(n_315), .Y(n_314) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_259), .Y(n_340) );
AND2x2_ASAP7_75t_L g352 ( .A(n_259), .B(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g364 ( .A(n_259), .Y(n_364) );
AND2x2_ASAP7_75t_L g389 ( .A(n_259), .B(n_286), .Y(n_389) );
INVx1_ASAP7_75t_L g409 ( .A(n_259), .Y(n_409) );
INVx1_ASAP7_75t_L g436 ( .A(n_259), .Y(n_436) );
AND2x2_ASAP7_75t_L g512 ( .A(n_259), .B(n_275), .Y(n_512) );
OR2x6_ASAP7_75t_L g259 ( .A(n_260), .B(n_268), .Y(n_259) );
OAI21x1_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_264), .B(n_266), .Y(n_260) );
NOR2xp33_ASAP7_75t_SL g297 ( .A(n_262), .B(n_298), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_262), .B(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g620 ( .A(n_262), .Y(n_620) );
INVx1_ASAP7_75t_L g288 ( .A(n_263), .Y(n_288) );
NOR2xp67_ASAP7_75t_L g268 ( .A(n_269), .B(n_272), .Y(n_268) );
INVx3_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g641 ( .A1(n_271), .A2(n_642), .B(n_643), .Y(n_641) );
OR2x2_ASAP7_75t_L g469 ( .A(n_273), .B(n_436), .Y(n_469) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x4_ASAP7_75t_L g313 ( .A(n_274), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g351 ( .A(n_274), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g329 ( .A(n_275), .Y(n_329) );
OAI22xp33_ASAP7_75t_L g331 ( .A1(n_276), .A2(n_332), .B1(n_334), .B2(n_338), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_280), .Y(n_276) );
AND2x4_ASAP7_75t_L g460 ( .A(n_277), .B(n_397), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_277), .B(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g337 ( .A(n_278), .Y(n_337) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g306 ( .A(n_279), .Y(n_306) );
INVxp67_ASAP7_75t_L g348 ( .A(n_279), .Y(n_348) );
AND2x2_ASAP7_75t_L g399 ( .A(n_279), .B(n_322), .Y(n_399) );
AND3x2_ASAP7_75t_L g346 ( .A(n_280), .B(n_347), .C(n_348), .Y(n_346) );
OR2x2_ASAP7_75t_L g385 ( .A(n_280), .B(n_386), .Y(n_385) );
OR2x2_ASAP7_75t_L g466 ( .A(n_280), .B(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_281), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g326 ( .A(n_281), .B(n_309), .Y(n_326) );
AND2x2_ASAP7_75t_L g529 ( .A(n_281), .B(n_323), .Y(n_529) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g318 ( .A(n_282), .Y(n_318) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_282), .Y(n_336) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_303), .Y(n_284) );
NOR2xp67_ASAP7_75t_SL g327 ( .A(n_285), .B(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g370 ( .A(n_285), .Y(n_370) );
AND2x2_ASAP7_75t_L g457 ( .A(n_285), .B(n_361), .Y(n_457) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g315 ( .A(n_286), .Y(n_315) );
OR2x2_ASAP7_75t_L g342 ( .A(n_286), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g353 ( .A(n_286), .Y(n_353) );
INVxp67_ASAP7_75t_L g406 ( .A(n_286), .Y(n_406) );
AO21x2_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_289), .B(n_301), .Y(n_286) );
NAND3xp33_ASAP7_75t_SL g289 ( .A(n_290), .B(n_293), .C(n_296), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_303), .B(n_352), .Y(n_476) );
OR2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
INVx1_ASAP7_75t_L g358 ( .A(n_305), .Y(n_358) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_306), .B(n_309), .Y(n_467) );
INVxp67_ASAP7_75t_L g455 ( .A(n_307), .Y(n_455) );
AND2x2_ASAP7_75t_L g427 ( .A(n_308), .B(n_322), .Y(n_427) );
AND2x2_ASAP7_75t_L g473 ( .A(n_308), .B(n_373), .Y(n_473) );
INVx1_ASAP7_75t_L g510 ( .A(n_308), .Y(n_510) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g376 ( .A(n_309), .Y(n_376) );
INVx1_ASAP7_75t_L g486 ( .A(n_309), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_311), .B(n_331), .Y(n_310) );
OAI21xp5_ASAP7_75t_SL g311 ( .A1(n_312), .A2(n_316), .B(n_324), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g333 ( .A(n_314), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_319), .Y(n_316) );
INVxp67_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g381 ( .A(n_319), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g325 ( .A(n_320), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g372 ( .A(n_320), .B(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g430 ( .A(n_321), .Y(n_430) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g416 ( .A(n_322), .Y(n_416) );
INVx3_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2x1p5_ASAP7_75t_L g324 ( .A(n_325), .B(n_327), .Y(n_324) );
INVx1_ASAP7_75t_L g517 ( .A(n_325), .Y(n_517) );
INVx1_ASAP7_75t_L g431 ( .A(n_326), .Y(n_431) );
OR2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx1_ASAP7_75t_L g487 ( .A(n_329), .Y(n_487) );
INVxp67_ASAP7_75t_SL g496 ( .A(n_330), .Y(n_496) );
INVx1_ASAP7_75t_L g449 ( .A(n_332), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_332), .A2(n_476), .B(n_492), .Y(n_491) );
OR2x2_ASAP7_75t_L g498 ( .A(n_333), .B(n_361), .Y(n_498) );
INVxp33_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
INVx1_ASAP7_75t_L g528 ( .A(n_337), .Y(n_528) );
INVx2_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g392 ( .A(n_339), .Y(n_392) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_340), .Y(n_425) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g412 ( .A(n_342), .Y(n_412) );
OR2x2_ASAP7_75t_L g423 ( .A(n_342), .B(n_362), .Y(n_423) );
BUFx2_ASAP7_75t_L g408 ( .A(n_343), .Y(n_408) );
NAND3xp33_ASAP7_75t_L g344 ( .A(n_345), .B(n_368), .C(n_378), .Y(n_344) );
AOI222xp33_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_349), .B1(n_351), .B2(n_354), .C1(n_359), .C2(n_365), .Y(n_345) );
NAND2x1_ASAP7_75t_L g492 ( .A(n_347), .B(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_347), .B(n_399), .Y(n_500) );
AND2x2_ASAP7_75t_L g508 ( .A(n_347), .B(n_482), .Y(n_508) );
INVx1_ASAP7_75t_L g367 ( .A(n_348), .Y(n_367) );
AND2x2_ASAP7_75t_L g401 ( .A(n_348), .B(n_402), .Y(n_401) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_348), .Y(n_522) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_351), .B(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g363 ( .A(n_353), .B(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_SL g354 ( .A(n_355), .B(n_357), .Y(n_354) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g366 ( .A(n_356), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_363), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_362), .B(n_406), .Y(n_405) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_362), .Y(n_411) );
AND2x2_ASAP7_75t_L g435 ( .A(n_362), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NAND3xp33_ASAP7_75t_L g368 ( .A(n_369), .B(n_371), .C(n_374), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g480 ( .A1(n_369), .A2(n_481), .B1(n_483), .B2(n_488), .Y(n_480) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
O2A1O1Ixp5_ASAP7_75t_L g494 ( .A1(n_372), .A2(n_495), .B(n_497), .C(n_499), .Y(n_494) );
AND2x4_ASAP7_75t_SL g415 ( .A(n_373), .B(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_377), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g444 ( .A(n_376), .Y(n_444) );
INVx1_ASAP7_75t_L g490 ( .A(n_376), .Y(n_490) );
AND2x2_ASAP7_75t_L g388 ( .A(n_377), .B(n_389), .Y(n_388) );
OAI21xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_384), .B(n_387), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g445 ( .A(n_386), .Y(n_445) );
INVx2_ASAP7_75t_L g493 ( .A(n_386), .Y(n_493) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g495 ( .A(n_389), .B(n_496), .Y(n_495) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_389), .Y(n_516) );
OAI211xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_393), .B(n_403), .C(n_417), .Y(n_390) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_400), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_396), .B(n_398), .Y(n_395) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
BUFx3_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_399), .B(n_510), .Y(n_509) );
INVx2_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
O2A1O1Ixp5_ASAP7_75t_L g452 ( .A1(n_401), .A2(n_453), .B(n_456), .C(n_458), .Y(n_452) );
INVx1_ASAP7_75t_L g419 ( .A(n_402), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_402), .B(n_525), .Y(n_524) );
OAI21xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_410), .B(n_413), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_404), .A2(n_433), .B1(n_439), .B2(n_443), .Y(n_432) );
AND2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_407), .Y(n_404) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_406), .Y(n_463) );
AND2x2_ASAP7_75t_L g456 ( .A(n_407), .B(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_407), .B(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
AND2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g525 ( .A(n_416), .Y(n_525) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
NOR3xp33_ASAP7_75t_L g420 ( .A(n_421), .B(n_451), .C(n_501), .Y(n_420) );
OAI211xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_426), .B(n_432), .C(n_446), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_423), .Y(n_526) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AOI21x1_ASAP7_75t_L g458 ( .A1(n_429), .A2(n_459), .B(n_461), .Y(n_458) );
OR2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NAND2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_437), .Y(n_434) );
BUFx3_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AND2x4_ASAP7_75t_L g511 ( .A(n_438), .B(n_512), .Y(n_511) );
INVxp67_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_448), .A2(n_480), .B(n_491), .Y(n_479) );
NAND4xp25_ASAP7_75t_L g451 ( .A(n_452), .B(n_464), .C(n_479), .D(n_494), .Y(n_451) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g470 ( .A(n_467), .Y(n_470) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
OAI22x1_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_474), .B1(n_476), .B2(n_477), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g489 ( .A(n_482), .B(n_490), .Y(n_489) );
INVx2_ASAP7_75t_SL g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g519 ( .A(n_484), .B(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_487), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g530 ( .A(n_495), .Y(n_530) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_518), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_511), .B(n_513), .Y(n_502) );
NAND3xp33_ASAP7_75t_L g503 ( .A(n_504), .B(n_507), .C(n_509), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_SL g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g514 ( .A(n_512), .Y(n_514) );
AOI21xp33_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B(n_517), .Y(n_513) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AOI21xp33_ASAP7_75t_SL g518 ( .A1(n_519), .A2(n_521), .B(n_523), .Y(n_518) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_526), .B1(n_527), .B2(n_530), .Y(n_523) );
NAND2x1p5_ASAP7_75t_L g527 ( .A(n_528), .B(n_529), .Y(n_527) );
INVxp33_ASAP7_75t_L g539 ( .A(n_531), .Y(n_539) );
NOR2x1_ASAP7_75t_R g531 ( .A(n_532), .B(n_533), .Y(n_531) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
CKINVDCx5p33_ASAP7_75t_R g534 ( .A(n_535), .Y(n_534) );
BUFx3_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_540), .B(n_910), .Y(n_538) );
INVx4_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
BUFx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g905 ( .A(n_545), .Y(n_905) );
BUFx8_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g900 ( .A(n_548), .Y(n_900) );
AND2x4_ASAP7_75t_L g548 ( .A(n_549), .B(n_794), .Y(n_548) );
NOR3xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_707), .C(n_753), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_654), .Y(n_550) );
OAI21xp33_ASAP7_75t_SL g551 ( .A1(n_552), .A2(n_595), .B(n_623), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g864 ( .A1(n_552), .A2(n_865), .B(n_867), .Y(n_864) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_563), .Y(n_553) );
OR2x2_ASAP7_75t_L g792 ( .A(n_554), .B(n_793), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_554), .B(n_825), .Y(n_824) );
INVx2_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g677 ( .A(n_556), .Y(n_677) );
INVx2_ASAP7_75t_L g706 ( .A(n_556), .Y(n_706) );
AND2x2_ASAP7_75t_L g727 ( .A(n_556), .B(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g844 ( .A(n_556), .B(n_565), .Y(n_844) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_562), .Y(n_556) );
AND2x2_ASAP7_75t_L g747 ( .A(n_557), .B(n_748), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_561), .Y(n_557) );
INVx2_ASAP7_75t_SL g563 ( .A(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_564), .B(n_681), .Y(n_797) );
AND2x2_ASAP7_75t_L g884 ( .A(n_564), .B(n_828), .Y(n_884) );
AND2x4_ASAP7_75t_L g564 ( .A(n_565), .B(n_578), .Y(n_564) );
INVx1_ASAP7_75t_L g703 ( .A(n_565), .Y(n_703) );
OAI21x1_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_569), .B(n_576), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_567), .B(n_592), .Y(n_628) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g621 ( .A(n_570), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_573), .Y(n_622) );
OR2x2_ASAP7_75t_L g614 ( .A(n_578), .B(n_615), .Y(n_614) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_578), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_578), .B(n_599), .Y(n_686) );
INVx2_ASAP7_75t_L g705 ( .A(n_578), .Y(n_705) );
INVx1_ASAP7_75t_L g744 ( .A(n_578), .Y(n_744) );
INVx1_ASAP7_75t_L g783 ( .A(n_578), .Y(n_783) );
AND2x2_ASAP7_75t_L g818 ( .A(n_578), .B(n_615), .Y(n_818) );
HB1xp67_ASAP7_75t_L g873 ( .A(n_578), .Y(n_873) );
AO31x2_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_585), .A3(n_590), .B(n_593), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NOR3xp33_ASAP7_75t_L g600 ( .A(n_591), .B(n_601), .C(n_605), .Y(n_600) );
INVx4_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g661 ( .A(n_592), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_614), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g676 ( .A(n_599), .B(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g713 ( .A(n_599), .B(n_705), .Y(n_713) );
INVx2_ASAP7_75t_L g728 ( .A(n_599), .Y(n_728) );
INVx2_ASAP7_75t_L g752 ( .A(n_599), .Y(n_752) );
AO21x2_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_610), .B(n_611), .Y(n_599) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_610), .B(n_619), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_614), .Y(n_710) );
OR2x2_ASAP7_75t_L g725 ( .A(n_614), .B(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g800 ( .A(n_614), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_615), .B(n_752), .Y(n_751) );
HB1xp67_ASAP7_75t_L g804 ( .A(n_615), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g834 ( .A(n_615), .B(n_808), .Y(n_834) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_618), .Y(n_615) );
AND2x2_ASAP7_75t_L g746 ( .A(n_618), .B(n_747), .Y(n_746) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_620), .A2(n_664), .B(n_667), .Y(n_663) );
AOI322xp5_ASAP7_75t_L g826 ( .A1(n_623), .A2(n_766), .A3(n_804), .B1(n_827), .B2(n_829), .C1(n_830), .C2(n_831), .Y(n_826) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_634), .Y(n_623) );
AND2x2_ASAP7_75t_L g831 ( .A(n_624), .B(n_811), .Y(n_831) );
NOR2xp33_ASAP7_75t_L g846 ( .A(n_624), .B(n_847), .Y(n_846) );
AND2x2_ASAP7_75t_L g882 ( .A(n_624), .B(n_774), .Y(n_882) );
INVx3_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_625), .B(n_683), .Y(n_699) );
AND2x2_ASAP7_75t_L g758 ( .A(n_625), .B(n_759), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_625), .B(n_722), .Y(n_802) );
AND2x4_ASAP7_75t_L g839 ( .A(n_625), .B(n_634), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_625), .B(n_761), .Y(n_880) );
INVx3_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g673 ( .A(n_626), .B(n_644), .Y(n_673) );
INVx1_ASAP7_75t_L g720 ( .A(n_626), .Y(n_720) );
AND2x2_ASAP7_75t_L g862 ( .A(n_626), .B(n_697), .Y(n_862) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g684 ( .A(n_627), .Y(n_684) );
OAI21x1_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_629), .B(n_633), .Y(n_627) );
INVx1_ASAP7_75t_L g693 ( .A(n_629), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_633), .Y(n_694) );
INVx1_ASAP7_75t_SL g787 ( .A(n_634), .Y(n_787) );
AND2x4_ASAP7_75t_L g634 ( .A(n_635), .B(n_644), .Y(n_634) );
AND2x2_ASAP7_75t_L g683 ( .A(n_635), .B(n_659), .Y(n_683) );
INVx1_ASAP7_75t_L g722 ( .A(n_635), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_635), .B(n_658), .Y(n_896) );
INVx3_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g697 ( .A(n_636), .Y(n_697) );
INVx1_ASAP7_75t_L g739 ( .A(n_636), .Y(n_739) );
AND2x2_ASAP7_75t_L g761 ( .A(n_636), .B(n_644), .Y(n_761) );
AND2x2_ASAP7_75t_L g811 ( .A(n_636), .B(n_659), .Y(n_811) );
HB1xp67_ASAP7_75t_L g815 ( .A(n_636), .Y(n_815) );
AND2x4_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_639), .B(n_641), .Y(n_638) );
OR2x2_ASAP7_75t_L g691 ( .A(n_644), .B(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g719 ( .A(n_644), .B(n_720), .Y(n_719) );
OA21x2_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_646), .B(n_653), .Y(n_644) );
OA21x2_ASAP7_75t_L g734 ( .A1(n_645), .A2(n_646), .B(n_653), .Y(n_734) );
AOI221xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_674), .B1(n_681), .B2(n_685), .C(n_687), .Y(n_654) );
INVxp67_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_657), .B(n_673), .Y(n_656) );
AND2x2_ASAP7_75t_L g857 ( .A(n_657), .B(n_719), .Y(n_857) );
BUFx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
OR2x2_ASAP7_75t_L g871 ( .A(n_658), .B(n_752), .Y(n_871) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
OR2x2_ASAP7_75t_L g696 ( .A(n_659), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g717 ( .A(n_659), .Y(n_717) );
AND2x2_ASAP7_75t_L g740 ( .A(n_659), .B(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g760 ( .A(n_659), .Y(n_760) );
BUFx2_ASAP7_75t_L g848 ( .A(n_659), .Y(n_848) );
INVx3_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AOI21x1_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_663), .B(n_671), .Y(n_660) );
AOI21xp5_ASAP7_75t_L g736 ( .A1(n_673), .A2(n_695), .B(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g860 ( .A(n_673), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_674), .A2(n_709), .B1(n_714), .B2(n_721), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_675), .B(n_678), .Y(n_674) );
OR2x2_ASAP7_75t_L g768 ( .A(n_675), .B(n_769), .Y(n_768) );
INVx2_ASAP7_75t_SL g675 ( .A(n_676), .Y(n_675) );
AND2x4_ASAP7_75t_L g799 ( .A(n_676), .B(n_800), .Y(n_799) );
AND2x2_ASAP7_75t_L g817 ( .A(n_676), .B(n_818), .Y(n_817) );
INVxp67_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g891 ( .A(n_680), .B(n_807), .Y(n_891) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NOR2xp33_ASAP7_75t_SL g803 ( .A(n_682), .B(n_804), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
AND2x2_ASAP7_75t_L g779 ( .A(n_684), .B(n_760), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_684), .B(n_815), .Y(n_814) );
INVx2_ASAP7_75t_L g866 ( .A(n_684), .Y(n_866) );
OR2x2_ASAP7_75t_L g895 ( .A(n_684), .B(n_896), .Y(n_895) );
AND2x4_ASAP7_75t_L g863 ( .A(n_685), .B(n_844), .Y(n_863) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AOI21xp33_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_698), .B(n_700), .Y(n_687) );
INVx2_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_690), .B(n_695), .Y(n_689) );
AND2x2_ASAP7_75t_L g721 ( .A(n_690), .B(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g821 ( .A(n_690), .B(n_822), .Y(n_821) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AND2x4_ASAP7_75t_L g732 ( .A(n_692), .B(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AND2x4_ASAP7_75t_L g774 ( .A(n_697), .B(n_733), .Y(n_774) );
OAI21xp33_ASAP7_75t_L g892 ( .A1(n_698), .A2(n_781), .B(n_893), .Y(n_892) );
BUFx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_704), .Y(n_700) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
OR2x2_ASAP7_75t_L g874 ( .A(n_702), .B(n_875), .Y(n_874) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
AND2x2_ASAP7_75t_L g749 ( .A(n_704), .B(n_750), .Y(n_749) );
AND2x2_ASAP7_75t_L g833 ( .A(n_704), .B(n_834), .Y(n_833) );
AND2x2_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .Y(n_704) );
INVx1_ASAP7_75t_L g770 ( .A(n_705), .Y(n_770) );
INVx1_ASAP7_75t_L g809 ( .A(n_706), .Y(n_809) );
AND2x4_ASAP7_75t_L g828 ( .A(n_706), .B(n_752), .Y(n_828) );
INVx1_ASAP7_75t_SL g875 ( .A(n_706), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_708), .B(n_723), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .Y(n_709) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g843 ( .A(n_713), .B(n_844), .Y(n_843) );
NOR2x1_ASAP7_75t_L g714 ( .A(n_715), .B(n_718), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
OR2x2_ASAP7_75t_L g730 ( .A(n_716), .B(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g827 ( .A(n_716), .B(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_717), .B(n_741), .Y(n_889) );
INVx3_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_721), .B(n_742), .Y(n_775) );
AND2x2_ASAP7_75t_L g766 ( .A(n_722), .B(n_732), .Y(n_766) );
AOI222xp33_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_729), .B1(n_735), .B2(n_737), .C1(n_742), .C2(n_749), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
OAI21xp33_ASAP7_75t_L g772 ( .A1(n_725), .A2(n_773), .B(n_775), .Y(n_772) );
OAI221xp5_ASAP7_75t_L g840 ( .A1(n_725), .A2(n_841), .B1(n_842), .B2(n_845), .C(n_849), .Y(n_840) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
BUFx2_ASAP7_75t_L g755 ( .A(n_727), .Y(n_755) );
AND2x2_ASAP7_75t_L g784 ( .A(n_728), .B(n_746), .Y(n_784) );
INVx1_ASAP7_75t_L g808 ( .A(n_728), .Y(n_808) );
HB1xp67_ASAP7_75t_L g837 ( .A(n_728), .Y(n_837) );
OAI21xp5_ASAP7_75t_L g820 ( .A1(n_729), .A2(n_821), .B(n_823), .Y(n_820) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AND2x2_ASAP7_75t_L g851 ( .A(n_732), .B(n_822), .Y(n_851) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g741 ( .A(n_734), .Y(n_741) );
INVxp67_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
AND2x4_ASAP7_75t_L g737 ( .A(n_738), .B(n_740), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_740), .Y(n_765) );
INVx2_ASAP7_75t_L g816 ( .A(n_741), .Y(n_816) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
OR2x2_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .Y(n_743) );
OR2x2_ASAP7_75t_L g872 ( .A(n_745), .B(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g838 ( .A(n_746), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_749), .B(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
OR2x2_ASAP7_75t_L g793 ( .A(n_751), .B(n_770), .Y(n_793) );
NAND4xp25_ASAP7_75t_L g753 ( .A(n_754), .B(n_762), .C(n_771), .D(n_776), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .Y(n_754) );
A2O1A1Ixp33_ASAP7_75t_L g849 ( .A1(n_755), .A2(n_850), .B(n_851), .C(n_852), .Y(n_849) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
AND2x2_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
INVx1_ASAP7_75t_L g790 ( .A(n_760), .Y(n_790) );
INVx1_ASAP7_75t_L g822 ( .A(n_760), .Y(n_822) );
OAI21xp5_ASAP7_75t_SL g762 ( .A1(n_763), .A2(n_766), .B(n_767), .Y(n_762) );
INVxp67_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVxp33_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
NAND2x1p5_ASAP7_75t_L g853 ( .A(n_774), .B(n_848), .Y(n_853) );
AND2x4_ASAP7_75t_L g865 ( .A(n_774), .B(n_866), .Y(n_865) );
NAND2x1p5_ASAP7_75t_L g876 ( .A(n_774), .B(n_789), .Y(n_876) );
AOI22xp5_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_780), .B1(n_785), .B2(n_791), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
NAND2x1p5_ASAP7_75t_SL g781 ( .A(n_782), .B(n_784), .Y(n_781) );
INVx2_ASAP7_75t_SL g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g850 ( .A(n_783), .Y(n_850) );
HB1xp67_ASAP7_75t_L g830 ( .A(n_784), .Y(n_830) );
INVx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
OR2x2_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
OR2x2_ASAP7_75t_L g841 ( .A(n_788), .B(n_814), .Y(n_841) );
INVx2_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx2_ASAP7_75t_L g829 ( .A(n_793), .Y(n_829) );
AND2x2_ASAP7_75t_L g794 ( .A(n_795), .B(n_854), .Y(n_794) );
NOR3xp33_ASAP7_75t_L g795 ( .A(n_796), .B(n_819), .C(n_840), .Y(n_795) );
NAND3xp33_ASAP7_75t_L g796 ( .A(n_797), .B(n_798), .C(n_810), .Y(n_796) );
AOI22x1_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_801), .B1(n_803), .B2(n_805), .Y(n_798) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
BUFx2_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_808), .B(n_809), .Y(n_807) );
OAI21xp33_ASAP7_75t_SL g810 ( .A1(n_811), .A2(n_812), .B(n_817), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_813), .B(n_816), .Y(n_812) );
HB1xp67_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVxp67_ASAP7_75t_L g888 ( .A(n_815), .Y(n_888) );
INVx1_ASAP7_75t_L g868 ( .A(n_816), .Y(n_868) );
BUFx6f_ASAP7_75t_L g825 ( .A(n_818), .Y(n_825) );
NAND3xp33_ASAP7_75t_L g819 ( .A(n_820), .B(n_826), .C(n_832), .Y(n_819) );
INVx1_ASAP7_75t_L g861 ( .A(n_822), .Y(n_861) );
INVx2_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
OAI21xp5_ASAP7_75t_L g832 ( .A1(n_833), .A2(n_835), .B(n_839), .Y(n_832) );
AOI22xp5_ASAP7_75t_L g885 ( .A1(n_833), .A2(n_851), .B1(n_886), .B2(n_890), .Y(n_885) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
OR2x2_ASAP7_75t_L g836 ( .A(n_837), .B(n_838), .Y(n_836) );
INVx2_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVxp67_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
NOR3xp33_ASAP7_75t_L g854 ( .A(n_855), .B(n_877), .C(n_892), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_856), .B(n_864), .Y(n_855) );
OAI31xp33_ASAP7_75t_L g856 ( .A1(n_857), .A2(n_858), .A3(n_862), .B(n_863), .Y(n_856) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
OR2x2_ASAP7_75t_L g859 ( .A(n_860), .B(n_861), .Y(n_859) );
OAI22xp5_ASAP7_75t_L g867 ( .A1(n_868), .A2(n_869), .B1(n_874), .B2(n_876), .Y(n_867) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
NOR2x1_ASAP7_75t_L g870 ( .A(n_871), .B(n_872), .Y(n_870) );
A2O1A1Ixp33_ASAP7_75t_L g877 ( .A1(n_878), .A2(n_881), .B(n_883), .C(n_885), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
INVx2_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
OR2x2_ASAP7_75t_L g887 ( .A(n_888), .B(n_889), .Y(n_887) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
INVx2_ASAP7_75t_L g903 ( .A(n_897), .Y(n_903) );
OAI22x1_ASAP7_75t_L g899 ( .A1(n_900), .A2(n_901), .B1(n_904), .B2(n_905), .Y(n_899) );
BUFx12f_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
CKINVDCx11_ASAP7_75t_R g902 ( .A(n_903), .Y(n_902) );
NOR2xp33_ASAP7_75t_L g906 ( .A(n_907), .B(n_908), .Y(n_906) );
BUFx3_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
CKINVDCx20_ASAP7_75t_R g910 ( .A(n_911), .Y(n_910) );
BUFx3_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
BUFx3_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
CKINVDCx6p67_ASAP7_75t_R g921 ( .A(n_914), .Y(n_921) );
BUFx5_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
AND2x2_ASAP7_75t_L g915 ( .A(n_916), .B(n_917), .Y(n_915) );
endmodule