module real_jpeg_2431_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_173;
wire n_105;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_70;
wire n_41;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_167;
wire n_128;
wire n_244;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_1),
.B(n_48),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_1),
.B(n_34),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_1),
.B(n_42),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_1),
.B(n_39),
.Y(n_145)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_3),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_3),
.B(n_52),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_3),
.B(n_30),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_3),
.B(n_26),
.Y(n_146)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_3),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_3),
.B(n_34),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_3),
.B(n_42),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_4),
.B(n_26),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_4),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_4),
.B(n_30),
.Y(n_236)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_5),
.B(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_5),
.Y(n_62)
);

AND2x2_ASAP7_75t_SL g110 ( 
.A(n_5),
.B(n_39),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_5),
.B(n_52),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_6),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_6),
.B(n_52),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_6),
.B(n_39),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_6),
.Y(n_85)
);

AND2x2_ASAP7_75t_SL g123 ( 
.A(n_6),
.B(n_34),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_6),
.B(n_30),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_9),
.B(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_9),
.B(n_26),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_9),
.B(n_65),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_9),
.B(n_34),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_9),
.B(n_48),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_9),
.B(n_42),
.Y(n_200)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_13),
.B(n_34),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_13),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_13),
.B(n_48),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_14),
.B(n_52),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_14),
.B(n_42),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_14),
.B(n_48),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_14),
.B(n_39),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_152),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_150),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_116),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_19),
.B(n_116),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_79),
.C(n_102),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_20),
.B(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_53),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_21),
.B(n_54),
.C(n_70),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_36),
.C(n_44),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_22),
.B(n_171),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_28),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_23),
.B(n_32),
.C(n_35),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_24),
.B(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_24),
.B(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_24),
.B(n_61),
.Y(n_213)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_28)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_36),
.B(n_44),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_41),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_37),
.A2(n_38),
.B1(n_41),
.B2(n_124),
.Y(n_162)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_39),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_41),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_41),
.Y(n_124)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_47),
.C(n_49),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_45),
.B(n_49),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_47),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_47),
.Y(n_161)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_50),
.B(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_51),
.B(n_101),
.Y(n_197)
);

INVx3_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_69),
.B2(n_70),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_58),
.B2(n_68),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_57),
.B(n_60),
.C(n_63),
.Y(n_148)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_63),
.B2(n_67),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_59),
.A2(n_60),
.B1(n_83),
.B2(n_84),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_97),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_64),
.B(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_71),
.A2(n_72),
.B(n_73),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_71),
.B(n_75),
.C(n_78),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_77),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_79),
.B(n_102),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_91),
.C(n_93),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_80),
.A2(n_91),
.B1(n_92),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_80),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_87),
.C(n_89),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_81),
.A2(n_82),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_86),
.B(n_101),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_87),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_93),
.B(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_100),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_98),
.B2(n_99),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_99),
.C(n_100),
.Y(n_115)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_97),
.B(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_97),
.B(n_101),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_101),
.B(n_169),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_115),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_107),
.C(n_115),
.Y(n_139)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_113),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_108)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_109),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_110),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_112),
.C(n_113),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_149),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_138),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_127),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_125),
.B2(n_126),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_122),
.A2(n_123),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_123),
.B(n_204),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_125),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_134),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_135),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_148),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_146),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_177),
.B(n_258),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_175),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_154),
.B(n_175),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_170),
.C(n_172),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_155),
.A2(n_156),
.B1(n_170),
.B2(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_162),
.C(n_163),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_157),
.A2(n_158),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_162),
.B(n_163),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.C(n_168),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_166),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_168),
.B(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_170),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_172),
.B(n_255),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_252),
.B(n_257),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_240),
.B(n_251),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_226),
.B(n_239),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_207),
.B(n_225),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_190),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_182),
.B(n_190),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_187),
.C(n_189),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_183),
.A2(n_184),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_184),
.A2(n_185),
.B(n_186),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_189),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_198),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_199),
.C(n_203),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_197),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_193),
.B(n_196),
.C(n_197),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_195),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_202),
.B1(n_203),
.B2(n_206),
.Y(n_198)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_199),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_200),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_201),
.Y(n_218)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_206),
.A2(n_218),
.B(n_219),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_216),
.B(n_224),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_212),
.B(n_215),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_210),
.B(n_211),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_217),
.B(n_220),
.Y(n_224)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_227),
.B(n_228),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_234),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_233),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_233),
.C(n_234),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_238),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_237),
.C(n_238),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_241),
.B(n_242),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_246),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_247),
.C(n_248),
.Y(n_253)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_253),
.B(n_254),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);


endmodule