module real_jpeg_17665_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_553;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_556;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_487;
wire n_93;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_534;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_0),
.A2(n_97),
.B1(n_100),
.B2(n_101),
.Y(n_96)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_0),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_0),
.A2(n_100),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_0),
.A2(n_100),
.B1(n_427),
.B2(n_428),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_SL g486 ( 
.A1(n_0),
.A2(n_100),
.B1(n_487),
.B2(n_489),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_1),
.A2(n_149),
.B1(n_153),
.B2(n_157),
.Y(n_148)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_1),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_1),
.A2(n_157),
.B1(n_247),
.B2(n_250),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_1),
.A2(n_157),
.B1(n_341),
.B2(n_343),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g552 ( 
.A1(n_1),
.A2(n_37),
.B1(n_157),
.B2(n_553),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_2),
.A2(n_32),
.B1(n_36),
.B2(n_37),
.Y(n_31)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_2),
.A2(n_36),
.B1(n_308),
.B2(n_311),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_2),
.A2(n_36),
.B1(n_419),
.B2(n_423),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_2),
.A2(n_36),
.B1(n_459),
.B2(n_462),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_3),
.A2(n_19),
.B(n_569),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_3),
.B(n_570),
.Y(n_569)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_4),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_4),
.Y(n_87)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_5),
.Y(n_182)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_5),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_5),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_5),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g406 ( 
.A(n_5),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_6),
.A2(n_207),
.B1(n_208),
.B2(n_211),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_6),
.Y(n_207)
);

OAI22x1_ASAP7_75t_L g238 ( 
.A1(n_6),
.A2(n_207),
.B1(n_239),
.B2(n_242),
.Y(n_238)
);

OAI22x1_ASAP7_75t_SL g291 ( 
.A1(n_6),
.A2(n_207),
.B1(n_292),
.B2(n_294),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_6),
.A2(n_207),
.B1(n_379),
.B2(n_380),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_7),
.A2(n_109),
.B1(n_112),
.B2(n_113),
.Y(n_108)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_7),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_7),
.A2(n_112),
.B1(n_197),
.B2(n_201),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_7),
.A2(n_112),
.B1(n_266),
.B2(n_269),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_7),
.A2(n_37),
.B1(n_112),
.B2(n_347),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_8),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_8),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g237 ( 
.A(n_8),
.Y(n_237)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_8),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_9),
.Y(n_78)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_9),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g213 ( 
.A(n_9),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_9),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_9),
.Y(n_396)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_9),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_9),
.Y(n_417)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_9),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_10),
.Y(n_570)
);

OAI32xp33_ASAP7_75t_L g117 ( 
.A1(n_11),
.A2(n_118),
.A3(n_123),
.B1(n_125),
.B2(n_132),
.Y(n_117)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_11),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_11),
.A2(n_131),
.B1(n_216),
.B2(n_219),
.Y(n_215)
);

OAI32xp33_ASAP7_75t_L g304 ( 
.A1(n_11),
.A2(n_118),
.A3(n_123),
.B1(n_125),
.B2(n_132),
.Y(n_304)
);

NAND2xp33_ASAP7_75t_SL g315 ( 
.A(n_11),
.B(n_41),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_11),
.B(n_69),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_11),
.B(n_467),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_11),
.B(n_205),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_SL g495 ( 
.A1(n_11),
.A2(n_131),
.B1(n_312),
.B2(n_496),
.Y(n_495)
);

OAI32xp33_ASAP7_75t_L g499 ( 
.A1(n_11),
.A2(n_500),
.A3(n_503),
.B1(n_504),
.B2(n_507),
.Y(n_499)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_14),
.A2(n_55),
.B1(n_62),
.B2(n_65),
.Y(n_61)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_14),
.A2(n_65),
.B1(n_225),
.B2(n_229),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_14),
.A2(n_65),
.B1(n_435),
.B2(n_436),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_14),
.A2(n_65),
.B1(n_444),
.B2(n_445),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_15),
.Y(n_143)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_15),
.Y(n_152)
);

BUFx4f_ASAP7_75t_L g167 ( 
.A(n_15),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g193 ( 
.A(n_15),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_16),
.A2(n_163),
.B1(n_168),
.B2(n_172),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_16),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_16),
.A2(n_172),
.B1(n_276),
.B2(n_278),
.Y(n_275)
);

OAI22xp33_ASAP7_75t_L g365 ( 
.A1(n_16),
.A2(n_172),
.B1(n_366),
.B2(n_368),
.Y(n_365)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_542),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_536),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_386),
.Y(n_22)
);

NOR3xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_325),
.C(n_355),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_298),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_255),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_26),
.B(n_255),
.C(n_538),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_173),
.C(n_231),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_27),
.B(n_324),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_116),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_66),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_29),
.B(n_66),
.C(n_116),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_39),
.B1(n_41),
.B2(n_60),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_31),
.A2(n_40),
.B1(n_215),
.B2(n_222),
.Y(n_214)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_33),
.Y(n_124)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_34),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_37),
.Y(n_285)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_39),
.B(n_378),
.Y(n_554)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_L g283 ( 
.A1(n_40),
.A2(n_61),
.B1(n_222),
.B2(n_284),
.Y(n_283)
);

OAI21xp33_ASAP7_75t_L g344 ( 
.A1(n_40),
.A2(n_284),
.B(n_345),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_40),
.A2(n_376),
.B(n_377),
.Y(n_375)
);

OR2x6_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_50),
.Y(n_40)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_41),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_41),
.B(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_41),
.B(n_378),
.Y(n_377)
);

AO22x2_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_44),
.B1(n_46),
.B2(n_48),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_43),
.Y(n_52)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_44),
.Y(n_115)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_45),
.Y(n_293)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_46),
.Y(n_313)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_47),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_47),
.Y(n_130)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_49),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_53),
.B1(n_55),
.B2(n_57),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_54),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_55),
.Y(n_133)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_56),
.Y(n_381)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_64),
.Y(n_288)
);

BUFx12f_ASAP7_75t_L g348 ( 
.A(n_64),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_95),
.B(n_106),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_67),
.A2(n_69),
.B1(n_364),
.B2(n_365),
.Y(n_363)
);

AOI21x1_ASAP7_75t_L g558 ( 
.A1(n_67),
.A2(n_365),
.B(n_559),
.Y(n_558)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_68),
.A2(n_96),
.B1(n_107),
.B2(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_68),
.A2(n_108),
.B(n_290),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_68),
.A2(n_107),
.B1(n_224),
.B2(n_307),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_68),
.A2(n_107),
.B1(n_339),
.B2(n_340),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_68),
.A2(n_107),
.B1(n_307),
.B2(n_495),
.Y(n_494)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_83),
.Y(n_68)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_69),
.B(n_291),
.Y(n_290)
);

AO22x2_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_72),
.B1(n_76),
.B2(n_79),
.Y(n_69)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_70),
.Y(n_278)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_70),
.Y(n_506)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_71),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_71),
.Y(n_437)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_77),
.Y(n_178)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_77),
.Y(n_200)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_77),
.Y(n_253)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_77),
.Y(n_277)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_78),
.Y(n_210)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_88),
.B1(n_91),
.B2(n_92),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_87),
.Y(n_513)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_88),
.Y(n_368)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_90),
.Y(n_230)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_90),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_90),
.Y(n_497)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_94),
.Y(n_310)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_103),
.Y(n_343)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

NOR2xp67_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_111),
.Y(n_502)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_137),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_122),
.Y(n_367)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_131),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_129),
.Y(n_228)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_131),
.B(n_399),
.Y(n_398)
);

OAI21xp33_ASAP7_75t_SL g413 ( 
.A1(n_131),
.A2(n_398),
.B(n_414),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_131),
.A2(n_139),
.B1(n_455),
.B2(n_458),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g504 ( 
.A(n_131),
.B(n_505),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_137),
.B(n_304),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_148),
.B1(n_158),
.B2(n_162),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_138),
.A2(n_162),
.B(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_138),
.A2(n_442),
.B1(n_448),
.B2(n_449),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_138),
.A2(n_233),
.B(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_139),
.B(n_238),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_139),
.A2(n_265),
.B(n_332),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_139),
.A2(n_426),
.B(n_431),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_139),
.A2(n_443),
.B1(n_458),
.B2(n_474),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_144),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_142),
.Y(n_410)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_144),
.Y(n_332)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_147),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_148),
.A2(n_272),
.B(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_149),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_150),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_151),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_152),
.Y(n_156)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_156),
.Y(n_189)
);

BUFx5_ASAP7_75t_L g449 ( 
.A(n_158),
.Y(n_449)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_167),
.Y(n_241)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_167),
.Y(n_461)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_173),
.B(n_231),
.Y(n_324)
);

MAJx2_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_214),
.C(n_223),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_174),
.B(n_223),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_196),
.B(n_204),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_175),
.A2(n_188),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

OA21x2_ASAP7_75t_L g334 ( 
.A1(n_175),
.A2(n_204),
.B(n_275),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_175),
.A2(n_188),
.B1(n_485),
.B2(n_486),
.Y(n_484)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_176),
.B(n_206),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_176),
.A2(n_205),
.B1(n_413),
.B2(n_418),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_176),
.A2(n_205),
.B1(n_418),
.B2(n_434),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_176),
.A2(n_370),
.B(n_523),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g556 ( 
.A1(n_176),
.A2(n_205),
.B(n_557),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_188),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_183),
.B2(n_187),
.Y(n_177)
);

OAI32xp33_ASAP7_75t_L g392 ( 
.A1(n_179),
.A2(n_393),
.A3(n_397),
.B1(n_398),
.B2(n_403),
.Y(n_392)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_188),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_188),
.B(n_196),
.Y(n_370)
);

OA22x2_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_192),
.B2(n_194),
.Y(n_188)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_192),
.Y(n_243)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_192),
.Y(n_471)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_193),
.Y(n_271)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_193),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_196),
.Y(n_557)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_202),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_205),
.B(n_246),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_214),
.B(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_221),
.Y(n_379)
);

OAI21x1_ASAP7_75t_SL g551 ( 
.A1(n_222),
.A2(n_552),
.B(n_554),
.Y(n_551)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_230),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_244),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_232),
.B(n_244),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_238),
.Y(n_233)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx12f_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_254),
.Y(n_244)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_246),
.Y(n_274)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVxp33_ASAP7_75t_L g371 ( 
.A(n_254),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_256),
.B(n_279),
.C(n_297),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_279),
.B1(n_280),
.B2(n_297),
.Y(n_257)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_258),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_273),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_259),
.B(n_273),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_272),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_260),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_265),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVxp33_ASAP7_75t_SL g515 ( 
.A(n_265),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_269),
.Y(n_397)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_280),
.Y(n_279)
);

XOR2x2_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_281),
.B(n_352),
.C(n_353),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_289),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_283),
.Y(n_352)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_289),
.Y(n_353)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_290),
.Y(n_559)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_291),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_323),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_299),
.B(n_323),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_302),
.C(n_305),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_300),
.B(n_533),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_302),
.A2(n_303),
.B1(n_305),
.B2(n_534),
.Y(n_533)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_305),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_314),
.C(n_316),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_306),
.B(n_526),
.Y(n_525)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx3_ASAP7_75t_SL g311 ( 
.A(n_312),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_314),
.A2(n_315),
.B1(n_316),
.B2(n_527),
.Y(n_526)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_316),
.Y(n_527)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_319),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx4_ASAP7_75t_SL g468 ( 
.A(n_320),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_321),
.Y(n_457)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g536 ( 
.A1(n_326),
.A2(n_537),
.B(n_539),
.C(n_540),
.D(n_541),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_327),
.B(n_328),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_329),
.A2(n_350),
.B1(n_351),
.B2(n_354),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g354 ( 
.A(n_329),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_336),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_330),
.B(n_336),
.C(n_350),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_331),
.A2(n_333),
.B1(n_334),
.B2(n_335),
.Y(n_330)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_331),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_331),
.A2(n_335),
.B1(n_375),
.B2(n_382),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_331),
.B(n_334),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

AOI21xp33_ASAP7_75t_L g564 ( 
.A1(n_335),
.A2(n_382),
.B(n_565),
.Y(n_564)
);

XNOR2x1_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_349),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_344),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_338),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_340),
.Y(n_364)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_344),
.Y(n_359)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_346),
.Y(n_376)
);

INVx5_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_349),
.B(n_359),
.C(n_360),
.Y(n_358)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_355),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_357),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_356),
.B(n_357),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_361),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_358),
.B(n_385),
.C(n_567),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_362),
.A2(n_373),
.B1(n_384),
.B2(n_385),
.Y(n_361)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_362),
.Y(n_385)
);

OAI21xp33_ASAP7_75t_L g362 ( 
.A1(n_363),
.A2(n_369),
.B(n_372),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_363),
.B(n_369),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_367),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_372),
.Y(n_548)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_373),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g567 ( 
.A(n_373),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_383),
.Y(n_373)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_375),
.Y(n_382)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_379),
.Y(n_553)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVxp33_ASAP7_75t_L g565 ( 
.A(n_383),
.Y(n_565)
);

OAI21x1_ASAP7_75t_L g386 ( 
.A1(n_387),
.A2(n_530),
.B(n_535),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_388),
.A2(n_517),
.B(n_529),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_389),
.A2(n_480),
.B(n_516),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_390),
.A2(n_439),
.B(n_479),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_424),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_391),
.B(n_424),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_411),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_392),
.A2(n_411),
.B1(n_412),
.B2(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_392),
.Y(n_451)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_393),
.Y(n_503)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_402),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_407),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_410),
.Y(n_430)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_416),
.Y(n_488)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx5_ASAP7_75t_L g435 ( 
.A(n_423),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_432),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_425),
.B(n_433),
.C(n_438),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_426),
.Y(n_448)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_438),
.Y(n_432)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_434),
.Y(n_485)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_440),
.A2(n_452),
.B(n_478),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_450),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_441),
.B(n_450),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_453),
.A2(n_472),
.B(n_477),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_465),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_461),
.Y(n_464)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_466),
.B(n_469),
.Y(n_465)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_473),
.B(n_476),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_473),
.B(n_476),
.Y(n_477)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_482),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_481),
.B(n_482),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_498),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_494),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_484),
.B(n_494),
.C(n_498),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_486),
.Y(n_523)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_514),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_499),
.B(n_514),
.Y(n_521)
);

INVx8_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_511),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_518),
.B(n_519),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g529 ( 
.A(n_518),
.B(n_519),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_520),
.A2(n_524),
.B1(n_525),
.B2(n_528),
.Y(n_519)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_520),
.Y(n_528)
);

XOR2x1_ASAP7_75t_SL g520 ( 
.A(n_521),
.B(n_522),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_521),
.B(n_522),
.C(n_524),
.Y(n_531)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_531),
.B(n_532),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_531),
.B(n_532),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_543),
.B(n_568),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

NOR2xp67_ASAP7_75t_SL g544 ( 
.A(n_545),
.B(n_566),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_545),
.B(n_566),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_546),
.A2(n_547),
.B1(n_563),
.B2(n_564),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_548),
.A2(n_549),
.B1(n_561),
.B2(n_562),
.Y(n_547)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_548),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_549),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_550),
.A2(n_551),
.B1(n_555),
.B2(n_560),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_555),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_556),
.B(n_558),
.Y(n_555)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);


endmodule