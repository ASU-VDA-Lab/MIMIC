module fake_jpeg_3545_n_191 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_191);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_191;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_24),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_12),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_35),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_33),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_68),
.B(n_69),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_55),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_0),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_71),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_18),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_0),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_63),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_53),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_59),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_74),
.A2(n_58),
.B1(n_49),
.B2(n_48),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_80),
.B(n_54),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_78),
.B(n_1),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_64),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_71),
.A2(n_58),
.B1(n_48),
.B2(n_66),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_73),
.Y(n_81)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_60),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_53),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_74),
.A2(n_64),
.B1(n_53),
.B2(n_50),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_88),
.A2(n_64),
.B1(n_50),
.B2(n_66),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_91),
.B(n_93),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_56),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_100),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_65),
.Y(n_93)
);

OAI21xp33_ASAP7_75t_SL g116 ( 
.A1(n_94),
.A2(n_20),
.B(n_42),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_52),
.B(n_61),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_95),
.A2(n_85),
.B(n_61),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_101),
.Y(n_109)
);

INVx6_ASAP7_75t_SL g97 ( 
.A(n_81),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_97),
.Y(n_113)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_99),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_54),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_78),
.B(n_77),
.C(n_82),
.Y(n_102)
);

FAx1_ASAP7_75t_SL g119 ( 
.A(n_102),
.B(n_2),
.CI(n_3),
.CON(n_119),
.SN(n_119)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_86),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_105),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_82),
.B(n_1),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_116),
.Y(n_125)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_100),
.A2(n_84),
.B1(n_76),
.B2(n_82),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_108),
.A2(n_110),
.B1(n_117),
.B2(n_118),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_101),
.A2(n_76),
.B1(n_82),
.B2(n_4),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

AO21x2_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_17),
.B(n_41),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_119),
.Y(n_140)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_2),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_122),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_3),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_124),
.B(n_98),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_129),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_104),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_123),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_134),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_104),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_135),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_133),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_98),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_46),
.Y(n_136)
);

AOI322xp5_ASAP7_75t_SL g148 ( 
.A1(n_136),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_13),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_137),
.A2(n_26),
.B1(n_36),
.B2(n_34),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_4),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_145),
.C(n_8),
.Y(n_151)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_142),
.Y(n_150)
);

CKINVDCx10_ASAP7_75t_R g143 ( 
.A(n_117),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_143),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_111),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_144),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_21),
.C(n_37),
.Y(n_145)
);

A2O1A1Ixp33_ASAP7_75t_SL g146 ( 
.A1(n_128),
.A2(n_117),
.B(n_119),
.C(n_22),
.Y(n_146)
);

OA21x2_ASAP7_75t_L g171 ( 
.A1(n_146),
.A2(n_142),
.B(n_140),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_143),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_147),
.A2(n_159),
.B1(n_162),
.B2(n_125),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_151),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_149),
.A2(n_145),
.B1(n_136),
.B2(n_126),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_129),
.C(n_131),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_160),
.C(n_158),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_134),
.Y(n_157)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_157),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_138),
.A2(n_25),
.B1(n_31),
.B2(n_30),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_125),
.A2(n_16),
.B(n_28),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_164),
.B(n_169),
.Y(n_175)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_165),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_168),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_132),
.C(n_139),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_161),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_172),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_171),
.A2(n_152),
.B(n_150),
.Y(n_178)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_164),
.B(n_148),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_177),
.B(n_166),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_179),
.Y(n_182)
);

INVx13_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_180),
.A2(n_183),
.B1(n_173),
.B2(n_146),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_163),
.C(n_159),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_SL g184 ( 
.A1(n_181),
.A2(n_174),
.B(n_146),
.C(n_127),
.Y(n_184)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_176),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_184),
.A2(n_185),
.B1(n_156),
.B2(n_173),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_186),
.Y(n_187)
);

AOI221xp5_ASAP7_75t_L g188 ( 
.A1(n_187),
.A2(n_182),
.B1(n_179),
.B2(n_171),
.C(n_27),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_188),
.B(n_171),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_38),
.C(n_11),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_15),
.Y(n_191)
);


endmodule