module fake_jpeg_25987_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_32),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_0),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_32),
.A2(n_25),
.B1(n_13),
.B2(n_15),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_45),
.B1(n_15),
.B2(n_20),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_17),
.B1(n_24),
.B2(n_23),
.Y(n_45)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_29),
.Y(n_51)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_60),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_47),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_50),
.B(n_57),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_31),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_59),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_13),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_54),
.B(n_56),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_33),
.B1(n_28),
.B2(n_36),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_55),
.A2(n_66),
.B1(n_53),
.B2(n_58),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_22),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_20),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_30),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_30),
.Y(n_81)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_38),
.A2(n_22),
.B(n_27),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_23),
.C(n_19),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_45),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_64),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_45),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_19),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_40),
.A2(n_13),
.B1(n_27),
.B2(n_24),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_71),
.B(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_77),
.B(n_78),
.Y(n_90)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_82),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_64),
.Y(n_91)
);

OAI32xp33_ASAP7_75t_L g83 ( 
.A1(n_65),
.A2(n_17),
.A3(n_26),
.B1(n_21),
.B2(n_1),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_63),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_96),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_86),
.B(n_88),
.Y(n_104)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_91),
.Y(n_106)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_92),
.A2(n_67),
.B1(n_76),
.B2(n_57),
.Y(n_98)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

BUFx24_ASAP7_75t_SL g105 ( 
.A(n_93),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_62),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_71),
.C(n_52),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_96),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_90),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_69),
.C(n_82),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_95),
.C(n_88),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_84),
.A2(n_67),
.B(n_69),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_103),
.A2(n_107),
.B(n_68),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_91),
.A2(n_74),
.B(n_82),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_110),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_54),
.C(n_92),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_116),
.C(n_94),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_113),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_106),
.A2(n_50),
.B1(n_60),
.B2(n_49),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_114),
.B(n_115),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_101),
.A2(n_60),
.B1(n_49),
.B2(n_48),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_26),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_112),
.A2(n_100),
.B(n_101),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_117),
.A2(n_119),
.B(n_122),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_105),
.Y(n_121)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_122),
.B(n_108),
.Y(n_124)
);

AO21x1_ASAP7_75t_L g123 ( 
.A1(n_118),
.A2(n_108),
.B(n_21),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_124),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_126),
.A2(n_7),
.B(n_8),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_120),
.B(n_3),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_3),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_128),
.B(n_8),
.Y(n_132)
);

INVxp33_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

OAI21xp33_ASAP7_75t_L g134 ( 
.A1(n_129),
.A2(n_12),
.B(n_11),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_131),
.A2(n_125),
.B(n_11),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_133),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_130),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_134),
.Y(n_137)
);


endmodule