module real_jpeg_15844_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_493;
wire n_93;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_20),
.B(n_493),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_0),
.B(n_494),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_1),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_1),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_1),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_1),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_1),
.B(n_179),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_1),
.B(n_214),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_2),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_2),
.Y(n_249)
);

BUFx5_ASAP7_75t_L g354 ( 
.A(n_2),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_3),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_3),
.B(n_126),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_3),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_3),
.B(n_275),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_3),
.B(n_317),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_3),
.B(n_412),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_3),
.B(n_415),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_3),
.B(n_432),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_4),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_4),
.B(n_86),
.Y(n_85)
);

INVxp33_ASAP7_75t_L g112 ( 
.A(n_4),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_4),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_4),
.B(n_162),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_4),
.B(n_259),
.Y(n_258)
);

AND2x4_ASAP7_75t_SL g272 ( 
.A(n_4),
.B(n_273),
.Y(n_272)
);

AND2x2_ASAP7_75t_SL g309 ( 
.A(n_4),
.B(n_214),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_5),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_5),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_5),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_5),
.B(n_175),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_5),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_5),
.B(n_222),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_5),
.A2(n_12),
.B1(n_245),
.B2(n_250),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_5),
.Y(n_351)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_6),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_6),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_7),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_7),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_7),
.B(n_109),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_7),
.B(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_8),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_8),
.Y(n_273)
);

BUFx5_ASAP7_75t_L g315 ( 
.A(n_8),
.Y(n_315)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_8),
.Y(n_403)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_9),
.Y(n_262)
);

BUFx12f_ASAP7_75t_L g308 ( 
.A(n_9),
.Y(n_308)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_9),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_10),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_10),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_10),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_10),
.B(n_98),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_10),
.B(n_202),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_10),
.B(n_270),
.Y(n_269)
);

INVxp33_ASAP7_75t_L g306 ( 
.A(n_10),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_10),
.B(n_247),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_11),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_12),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_12),
.B(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_12),
.B(n_312),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_12),
.B(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_12),
.B(n_383),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_12),
.B(n_401),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_12),
.B(n_407),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_12),
.B(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

NAND2x1_ASAP7_75t_L g41 ( 
.A(n_13),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g205 ( 
.A(n_13),
.B(n_206),
.Y(n_205)
);

AND2x2_ASAP7_75t_SL g224 ( 
.A(n_13),
.B(n_225),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_13),
.B(n_266),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_13),
.B(n_315),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_13),
.B(n_358),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_13),
.B(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_14),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_14),
.Y(n_99)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_14),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_15),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_15),
.B(n_363),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_15),
.B(n_349),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_15),
.B(n_398),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_15),
.B(n_448),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_15),
.B(n_452),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_15),
.B(n_458),
.Y(n_457)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_16),
.Y(n_80)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_16),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_16),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_16),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_16),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_16),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_18),
.Y(n_127)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_18),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_184),
.Y(n_20)
);

NAND2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_183),
.Y(n_21)
);

INVxp33_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp67_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_150),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_24),
.B(n_150),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_105),
.C(n_119),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_25),
.A2(n_26),
.B1(n_105),
.B2(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_63),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_47),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_28),
.B(n_47),
.C(n_152),
.Y(n_151)
);

MAJx2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_41),
.C(n_43),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_29),
.A2(n_30),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

MAJx2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_35),
.C(n_37),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_31),
.A2(n_69),
.B1(n_70),
.B2(n_74),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_31),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_31),
.A2(n_35),
.B1(n_74),
.B2(n_134),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_32),
.B(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_33),
.Y(n_129)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_33),
.Y(n_458)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_34),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_35),
.B(n_125),
.C(n_128),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_35),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_35),
.A2(n_128),
.B1(n_134),
.B2(n_197),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_36),
.Y(n_412)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_36),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_37),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_37),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_37),
.A2(n_131),
.B1(n_258),
.B2(n_303),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_39),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_40),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_41),
.B(n_43),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_41),
.B(n_213),
.C(n_218),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_41),
.B(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_43),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_43),
.A2(n_145),
.B1(n_146),
.B2(n_230),
.Y(n_229)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_46),
.Y(n_181)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_46),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_48),
.B(n_57),
.C(n_62),
.Y(n_182)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_57),
.B1(n_58),
.B2(n_62),
.Y(n_51)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_55),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_56),
.Y(n_227)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_63),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_75),
.C(n_89),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_64),
.B(n_192),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_68),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_65),
.B(n_70),
.C(n_74),
.Y(n_117)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_69),
.A2(n_70),
.B1(n_108),
.B2(n_110),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_SL g159 ( 
.A(n_70),
.B(n_108),
.C(n_111),
.Y(n_159)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_75),
.B(n_89),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_81),
.C(n_85),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_76),
.B(n_85),
.Y(n_123)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_80),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_123),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_84),
.Y(n_222)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_88),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_94),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_95),
.C(n_100),
.Y(n_118)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_100),
.Y(n_94)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_99),
.Y(n_170)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_104),
.Y(n_266)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_105),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_116),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_106),
.B(n_117),
.C(n_118),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_111),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_108),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_108),
.A2(n_110),
.B1(n_167),
.B2(n_171),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_115),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_119),
.B(n_232),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_135),
.C(n_147),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_121),
.B(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_124),
.C(n_130),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_122),
.B(n_124),
.Y(n_287)
);

XNOR2x1_ASAP7_75t_L g195 ( 
.A(n_125),
.B(n_196),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_128),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_130),
.B(n_287),
.Y(n_286)
);

MAJx2_ASAP7_75t_L g254 ( 
.A(n_131),
.B(n_255),
.C(n_258),
.Y(n_254)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_135),
.B(n_147),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_145),
.C(n_146),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_136),
.B(n_229),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.C(n_144),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_137),
.B(n_144),
.Y(n_210)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_140),
.B(n_210),
.Y(n_209)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_145),
.Y(n_230)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_148),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_153),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_172),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

XOR2x1_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_166),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_164),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_167),
.Y(n_171)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_182),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_178),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_491),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_234),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_231),
.Y(n_187)
);

NOR2xp67_ASAP7_75t_SL g492 ( 
.A(n_188),
.B(n_231),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.C(n_193),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_189),
.B(n_191),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_193),
.B(n_327),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_211),
.C(n_228),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_194),
.B(n_285),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_198),
.C(n_209),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_195),
.B(n_198),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_201),
.C(n_204),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_199),
.A2(n_204),
.B1(n_205),
.B2(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_199),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_201),
.B(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVxp67_ASAP7_75t_SL g448 ( 
.A(n_203),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_204),
.B(n_381),
.C(n_382),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_204),
.A2(n_205),
.B1(n_381),
.B2(n_426),
.Y(n_425)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_207),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_208),
.Y(n_313)
);

XNOR2x1_ASAP7_75t_SL g295 ( 
.A(n_209),
.B(n_296),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_211),
.B(n_228),
.Y(n_285)
);

MAJx2_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_221),
.C(n_223),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_212),
.B(n_281),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_218),
.Y(n_242)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_217),
.Y(n_418)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_221),
.A2(n_223),
.B1(n_224),
.B2(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_221),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_223),
.A2(n_224),
.B1(n_361),
.B2(n_362),
.Y(n_474)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_224),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_224),
.B(n_356),
.C(n_361),
.Y(n_355)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

AO21x2_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_331),
.B(n_488),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_325),
.Y(n_235)
);

AND2x2_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_290),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g489 ( 
.A(n_237),
.B(n_290),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_283),
.Y(n_237)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_238),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_263),
.C(n_278),
.Y(n_238)
);

INVxp33_ASAP7_75t_SL g239 ( 
.A(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_240),
.B(n_293),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_243),
.C(n_254),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_241),
.B(n_366),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_243),
.A2(n_244),
.B1(n_254),
.B2(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_244),
.A2(n_347),
.B(n_350),
.Y(n_346)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_254),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_255),
.B(n_302),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_258),
.Y(n_303)
);

BUFx2_ASAP7_75t_SL g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_263),
.A2(n_279),
.B1(n_280),
.B2(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_263),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_271),
.C(n_274),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_264),
.B(n_320),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_267),
.C(n_269),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_265),
.A2(n_269),
.B1(n_344),
.B2(n_345),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_265),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_265),
.B(n_396),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_267),
.B(n_343),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_269),
.Y(n_345)
);

INVx6_ASAP7_75t_L g453 ( 
.A(n_270),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_271),
.A2(n_272),
.B1(n_274),
.B2(n_321),
.Y(n_320)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_274),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_277),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_286),
.B1(n_288),
.B2(n_289),
.Y(n_283)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_284),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_286),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_286),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_288),
.B(n_329),
.C(n_330),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_295),
.C(n_297),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_291),
.A2(n_292),
.B1(n_295),
.B2(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_295),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g297 ( 
.A(n_298),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_298),
.B(n_335),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_319),
.C(n_322),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_299),
.B(n_340),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_304),
.C(n_310),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

XNOR2x1_ASAP7_75t_L g386 ( 
.A(n_301),
.B(n_387),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_304),
.B(n_310),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_309),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_305),
.B(n_309),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx5_ASAP7_75t_L g359 ( 
.A(n_308),
.Y(n_359)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_308),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_314),
.C(n_316),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_311),
.A2(n_314),
.B1(n_377),
.B2(n_378),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_311),
.Y(n_377)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_314),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_314),
.A2(n_378),
.B1(n_446),
.B2(n_447),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_314),
.B(n_442),
.C(n_446),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_315),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_316),
.B(n_376),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_319),
.B(n_322),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_325),
.A2(n_489),
.B(n_490),
.Y(n_488)
);

AND2x2_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_328),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g490 ( 
.A(n_326),
.B(n_328),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_388),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_337),
.C(n_368),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_334),
.B(n_338),
.Y(n_487)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_341),
.C(n_364),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_339),
.B(n_370),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_341),
.B(n_365),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_346),
.C(n_355),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_342),
.B(n_346),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_344),
.B(n_397),
.C(n_400),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

INVx6_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

BUFx12f_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_355),
.B(n_373),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_SL g473 ( 
.A(n_356),
.B(n_474),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_360),
.Y(n_356)
);

XNOR2x1_ASAP7_75t_SL g430 ( 
.A(n_357),
.B(n_360),
.Y(n_430)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_357),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_357),
.A2(n_437),
.B1(n_438),
.B2(n_455),
.Y(n_454)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

NOR2xp67_ASAP7_75t_SL g368 ( 
.A(n_369),
.B(n_371),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_369),
.B(n_371),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_374),
.C(n_386),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_372),
.B(n_484),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_374),
.B(n_386),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_379),
.C(n_384),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_375),
.B(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_380),
.B(n_385),
.Y(n_479)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_381),
.Y(n_426)
);

XOR2x1_ASAP7_75t_L g424 ( 
.A(n_382),
.B(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

NAND3xp33_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_390),
.C(n_487),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_391),
.A2(n_482),
.B(n_486),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_392),
.A2(n_468),
.B(n_481),
.Y(n_391)
);

OAI21x1_ASAP7_75t_L g392 ( 
.A1(n_393),
.A2(n_433),
.B(n_467),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_421),
.Y(n_393)
);

OR2x2_ASAP7_75t_L g467 ( 
.A(n_394),
.B(n_421),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_404),
.C(n_413),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_395),
.B(n_463),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_400),
.Y(n_396)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_404),
.A2(n_405),
.B1(n_413),
.B2(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_411),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_SL g443 ( 
.A(n_406),
.B(n_411),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx4_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_413),
.Y(n_464)
);

AO22x1_ASAP7_75t_SL g413 ( 
.A1(n_414),
.A2(n_417),
.B1(n_419),
.B2(n_420),
.Y(n_413)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_414),
.Y(n_419)
);

INVx4_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_417),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_417),
.B(n_419),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_420),
.B(n_457),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_427),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_423),
.B(n_424),
.C(n_427),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_429),
.Y(n_427)
);

MAJx2_ASAP7_75t_L g476 ( 
.A(n_428),
.B(n_430),
.C(n_431),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_431),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_434),
.A2(n_461),
.B(n_466),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_435),
.A2(n_449),
.B(n_460),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_441),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_436),
.B(n_441),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_437),
.B(n_438),
.Y(n_436)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_438),
.Y(n_455)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_442),
.A2(n_443),
.B1(n_444),
.B2(n_445),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_450),
.A2(n_456),
.B(n_459),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_454),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_451),
.B(n_454),
.Y(n_459)
);

INVx4_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_462),
.B(n_465),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_462),
.B(n_465),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_469),
.B(n_480),
.Y(n_468)
);

NOR2xp67_ASAP7_75t_SL g481 ( 
.A(n_469),
.B(n_480),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_470),
.A2(n_471),
.B1(n_477),
.B2(n_478),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_472),
.A2(n_473),
.B1(n_475),
.B2(n_476),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_472),
.B(n_476),
.C(n_477),
.Y(n_485)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_485),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_483),
.B(n_485),
.Y(n_486)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);


endmodule