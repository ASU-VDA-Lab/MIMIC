module fake_netlist_5_582_n_1667 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1667);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1667;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_254;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_368;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_139),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_80),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_136),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_9),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_117),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_40),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_41),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_7),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_74),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_51),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_50),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_97),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_110),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_96),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_68),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_19),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_129),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_69),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_75),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_91),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_21),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_128),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_90),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_130),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_79),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_141),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_84),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_71),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_34),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_12),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_104),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_142),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_124),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_102),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_52),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_10),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_111),
.Y(n_191)
);

BUFx5_ASAP7_75t_L g192 ( 
.A(n_78),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_29),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_7),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_22),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_26),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_95),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_1),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_59),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_92),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_39),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_70),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_25),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_12),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_8),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_148),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_18),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_46),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_98),
.Y(n_209)
);

BUFx10_ASAP7_75t_L g210 ( 
.A(n_8),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_17),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_145),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_43),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_131),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_149),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_3),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_61),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_87),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_55),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_119),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_82),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_99),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_135),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_140),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_138),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_133),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_103),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_45),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_89),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_16),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_4),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_16),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_32),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_112),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_9),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_21),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_29),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_5),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_34),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_35),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_83),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_127),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_37),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_25),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_26),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_38),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_35),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_54),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_101),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_4),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_146),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_122),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_137),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_94),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_3),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_41),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_2),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_27),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_150),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_126),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_17),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_13),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_114),
.Y(n_263)
);

BUFx10_ASAP7_75t_L g264 ( 
.A(n_63),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_125),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_123),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_152),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_5),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_118),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_62),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_18),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_11),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_6),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_42),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_49),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_132),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_47),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_20),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_0),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_121),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_1),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_76),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_6),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_113),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_65),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_109),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_31),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_116),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_100),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_33),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_23),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_77),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_147),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_38),
.Y(n_294)
);

BUFx8_ASAP7_75t_SL g295 ( 
.A(n_57),
.Y(n_295)
);

INVx4_ASAP7_75t_R g296 ( 
.A(n_120),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_30),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_107),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_13),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_32),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_144),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_53),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_14),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_67),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_43),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_40),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_260),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_211),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_211),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_257),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_192),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_257),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_279),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_210),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_163),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_279),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_210),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_287),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_287),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_192),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_159),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_159),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_179),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_200),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_265),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_160),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_160),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_193),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_295),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_193),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_239),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_239),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_181),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_170),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_188),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_169),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_200),
.Y(n_337)
);

INVxp67_ASAP7_75t_SL g338 ( 
.A(n_284),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_183),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_189),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_184),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_201),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_286),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_168),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_249),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_157),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_187),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_203),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_263),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_205),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_293),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_206),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_231),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_208),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_233),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_245),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_209),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_235),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_237),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_264),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_215),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_240),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_247),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_256),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_220),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_192),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_268),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_297),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_192),
.Y(n_369)
);

BUFx6f_ASAP7_75t_SL g370 ( 
.A(n_264),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_221),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_223),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_299),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_224),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_300),
.Y(n_375)
);

AND2x4_ASAP7_75t_L g376 ( 
.A(n_349),
.B(n_263),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_334),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_338),
.A2(n_198),
.B1(n_294),
.B2(n_281),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_336),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_334),
.Y(n_380)
);

NOR2x1_ASAP7_75t_L g381 ( 
.A(n_344),
.B(n_263),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_324),
.B(n_264),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_336),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_341),
.Y(n_384)
);

OA21x2_ASAP7_75t_L g385 ( 
.A1(n_311),
.A2(n_303),
.B(n_186),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_344),
.B(n_180),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_324),
.B(n_337),
.Y(n_387)
);

OAI21x1_ASAP7_75t_L g388 ( 
.A1(n_311),
.A2(n_186),
.B(n_168),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_333),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_344),
.B(n_180),
.Y(n_390)
);

NOR2x1_ASAP7_75t_L g391 ( 
.A(n_360),
.B(n_248),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_341),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_336),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_337),
.B(n_217),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_342),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_336),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_336),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_342),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_321),
.B(n_217),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_320),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_321),
.B(n_222),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_320),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_366),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_335),
.B(n_340),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_366),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_369),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_369),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_356),
.B(n_210),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_348),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_322),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_348),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_322),
.B(n_222),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_307),
.B(n_305),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_308),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_326),
.B(n_327),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_308),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_350),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_326),
.B(n_248),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_315),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_350),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_309),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_323),
.A2(n_232),
.B1(n_204),
.B2(n_216),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_345),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_327),
.B(n_154),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_309),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_328),
.B(n_154),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_346),
.Y(n_427)
);

AND2x6_ASAP7_75t_L g428 ( 
.A(n_360),
.B(n_169),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_353),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_314),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_310),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_328),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_325),
.B(n_157),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_310),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_330),
.B(n_155),
.Y(n_435)
);

AND2x6_ASAP7_75t_L g436 ( 
.A(n_312),
.B(n_169),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_317),
.A2(n_306),
.B1(n_175),
.B2(n_161),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_312),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_376),
.B(n_352),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_400),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_400),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_385),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_376),
.B(n_354),
.Y(n_443)
);

NAND3xp33_ASAP7_75t_L g444 ( 
.A(n_424),
.B(n_347),
.C(n_357),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_400),
.Y(n_445)
);

INVx2_ASAP7_75t_SL g446 ( 
.A(n_387),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_396),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_376),
.B(n_361),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_376),
.B(n_269),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_404),
.B(n_371),
.Y(n_450)
);

INVxp33_ASAP7_75t_L g451 ( 
.A(n_430),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_387),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_410),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_406),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_412),
.B(n_330),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_396),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_427),
.A2(n_343),
.B1(n_365),
.B2(n_372),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_430),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_402),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_433),
.B(n_374),
.Y(n_460)
);

INVx2_ASAP7_75t_SL g461 ( 
.A(n_382),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_402),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_396),
.Y(n_463)
);

NAND2xp33_ASAP7_75t_SL g464 ( 
.A(n_382),
.B(n_370),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_402),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_385),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_403),
.Y(n_467)
);

INVx2_ASAP7_75t_SL g468 ( 
.A(n_394),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_394),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_410),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_412),
.B(n_331),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_385),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_385),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_385),
.Y(n_474)
);

NAND2xp33_ASAP7_75t_R g475 ( 
.A(n_389),
.B(n_329),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_403),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_396),
.Y(n_477)
);

INVx4_ASAP7_75t_L g478 ( 
.A(n_406),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_403),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_433),
.A2(n_370),
.B1(n_351),
.B2(n_172),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_396),
.Y(n_481)
);

NAND2xp33_ASAP7_75t_L g482 ( 
.A(n_428),
.B(n_169),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_405),
.Y(n_483)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_424),
.B(n_331),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_419),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_413),
.B(n_155),
.Y(n_486)
);

INVx2_ASAP7_75t_SL g487 ( 
.A(n_394),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_405),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_405),
.Y(n_489)
);

INVx2_ASAP7_75t_SL g490 ( 
.A(n_394),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_423),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_427),
.B(n_370),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_413),
.B(n_156),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_L g494 ( 
.A1(n_418),
.A2(n_302),
.B1(n_269),
.B2(n_285),
.Y(n_494)
);

BUFx4f_ASAP7_75t_L g495 ( 
.A(n_428),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_425),
.Y(n_496)
);

INVxp33_ASAP7_75t_L g497 ( 
.A(n_422),
.Y(n_497)
);

INVxp33_ASAP7_75t_SL g498 ( 
.A(n_408),
.Y(n_498)
);

AND2x6_ASAP7_75t_L g499 ( 
.A(n_381),
.B(n_285),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_422),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_396),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_425),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_418),
.A2(n_302),
.B1(n_339),
.B2(n_292),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_425),
.Y(n_504)
);

INVxp33_ASAP7_75t_L g505 ( 
.A(n_437),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_426),
.B(n_332),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_L g507 ( 
.A1(n_418),
.A2(n_169),
.B1(n_182),
.B2(n_292),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_426),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_408),
.B(n_156),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_410),
.B(n_332),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_406),
.B(n_158),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_407),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_432),
.B(n_375),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_425),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g515 ( 
.A(n_435),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_435),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_391),
.B(n_166),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_407),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_432),
.B(n_254),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_406),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_406),
.Y(n_521)
);

AO22x2_ASAP7_75t_L g522 ( 
.A1(n_437),
.A2(n_212),
.B1(n_276),
.B2(n_266),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_432),
.B(n_313),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_428),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g525 ( 
.A1(n_418),
.A2(n_182),
.B1(n_292),
.B2(n_375),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_391),
.B(n_259),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_377),
.B(n_313),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_407),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_407),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_428),
.B(n_226),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_388),
.Y(n_531)
);

BUFx2_ASAP7_75t_L g532 ( 
.A(n_378),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_425),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_399),
.B(n_166),
.Y(n_534)
);

INVx2_ASAP7_75t_SL g535 ( 
.A(n_381),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_388),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_388),
.Y(n_537)
);

NAND2xp33_ASAP7_75t_L g538 ( 
.A(n_428),
.B(n_182),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_378),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_377),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_380),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_386),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_425),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_380),
.Y(n_544)
);

INVx5_ASAP7_75t_L g545 ( 
.A(n_436),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_434),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_384),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_386),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_384),
.A2(n_182),
.B1(n_292),
.B2(n_367),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_434),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_434),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_434),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_434),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_399),
.B(n_171),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_434),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_392),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_428),
.B(n_227),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_392),
.Y(n_558)
);

INVxp67_ASAP7_75t_SL g559 ( 
.A(n_397),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_395),
.B(n_316),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_395),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_397),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_397),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_428),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_401),
.B(n_171),
.Y(n_565)
);

OAI22xp33_ASAP7_75t_L g566 ( 
.A1(n_415),
.A2(n_236),
.B1(n_195),
.B2(n_190),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_L g567 ( 
.A1(n_398),
.A2(n_182),
.B1(n_292),
.B2(n_373),
.Y(n_567)
);

OR2x6_ASAP7_75t_L g568 ( 
.A(n_415),
.B(n_401),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_398),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_409),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_428),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_397),
.Y(n_572)
);

INVx8_ASAP7_75t_L g573 ( 
.A(n_428),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_379),
.B(n_229),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_421),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_409),
.B(n_316),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_411),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_411),
.B(n_172),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_417),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_417),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_420),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_420),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_429),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_429),
.B(n_318),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_508),
.A2(n_234),
.B1(n_241),
.B2(n_251),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_508),
.A2(n_275),
.B1(n_252),
.B2(n_267),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_516),
.B(n_173),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_440),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_451),
.B(n_353),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_579),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_579),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_540),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_540),
.Y(n_593)
);

A2O1A1Ixp33_ASAP7_75t_L g594 ( 
.A1(n_515),
.A2(n_202),
.B(n_162),
.C(n_253),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_461),
.B(n_173),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_475),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_541),
.Y(n_597)
);

BUFx6f_ASAP7_75t_SL g598 ( 
.A(n_515),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_544),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_461),
.B(n_174),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_544),
.Y(n_601)
);

NAND3xp33_ASAP7_75t_L g602 ( 
.A(n_534),
.B(n_207),
.C(n_213),
.Y(n_602)
);

INVxp67_ASAP7_75t_SL g603 ( 
.A(n_442),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_542),
.B(n_548),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_547),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_440),
.Y(n_606)
);

O2A1O1Ixp33_ASAP7_75t_L g607 ( 
.A1(n_484),
.A2(n_390),
.B(n_355),
.C(n_364),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_542),
.B(n_421),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_452),
.B(n_355),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_505),
.A2(n_291),
.B1(n_278),
.B2(n_283),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_548),
.B(n_468),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_526),
.B(n_174),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_491),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_468),
.B(n_176),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_469),
.A2(n_270),
.B1(n_177),
.B2(n_178),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_469),
.B(n_421),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_487),
.B(n_421),
.Y(n_617)
);

OR2x6_ASAP7_75t_L g618 ( 
.A(n_532),
.B(n_358),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_487),
.B(n_431),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_490),
.B(n_431),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_547),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_556),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_454),
.A2(n_390),
.B(n_379),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_490),
.A2(n_176),
.B1(n_177),
.B2(n_304),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_452),
.B(n_358),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_556),
.Y(n_626)
);

NAND2x1p5_ASAP7_75t_L g627 ( 
.A(n_495),
.B(n_164),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_558),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_558),
.Y(n_629)
);

INVx8_ASAP7_75t_L g630 ( 
.A(n_568),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_561),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_561),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_449),
.A2(n_199),
.B1(n_165),
.B2(n_242),
.Y(n_633)
);

INVx6_ASAP7_75t_L g634 ( 
.A(n_513),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_446),
.B(n_359),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_450),
.B(n_178),
.Y(n_636)
);

AO22x1_ASAP7_75t_L g637 ( 
.A1(n_497),
.A2(n_291),
.B1(n_278),
.B2(n_283),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_446),
.B(n_359),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_506),
.B(n_362),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_441),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_442),
.B(n_431),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_466),
.B(n_431),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_439),
.B(n_277),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_455),
.B(n_362),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_455),
.B(n_363),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_510),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_466),
.B(n_438),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_443),
.B(n_277),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_448),
.B(n_444),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_457),
.B(n_280),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_472),
.B(n_438),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_486),
.B(n_280),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_472),
.B(n_438),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_519),
.B(n_282),
.Y(n_654)
);

INVx1_ASAP7_75t_SL g655 ( 
.A(n_458),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_473),
.B(n_383),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_441),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_453),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_569),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_445),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_569),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_473),
.B(n_383),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_554),
.B(n_282),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_565),
.B(n_288),
.Y(n_664)
);

AOI22x1_ASAP7_75t_L g665 ( 
.A1(n_474),
.A2(n_185),
.B1(n_225),
.B2(n_219),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_471),
.B(n_363),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_570),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_449),
.A2(n_288),
.B1(n_304),
.B2(n_301),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_535),
.B(n_383),
.Y(n_669)
);

A2O1A1Ixp33_ASAP7_75t_L g670 ( 
.A1(n_449),
.A2(n_167),
.B(n_218),
.C(n_214),
.Y(n_670)
);

BUFx4f_ASAP7_75t_L g671 ( 
.A(n_568),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_570),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_492),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_445),
.Y(n_674)
);

NAND2xp33_ASAP7_75t_L g675 ( 
.A(n_564),
.B(n_192),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_493),
.B(n_289),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_577),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_459),
.Y(n_678)
);

AND2x6_ASAP7_75t_SL g679 ( 
.A(n_500),
.B(n_364),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_453),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_474),
.B(n_393),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_484),
.B(n_535),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_470),
.B(n_289),
.Y(n_683)
);

OAI21xp33_ASAP7_75t_L g684 ( 
.A1(n_471),
.A2(n_373),
.B(n_368),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_510),
.B(n_568),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_449),
.B(n_393),
.Y(n_686)
);

NAND2xp33_ASAP7_75t_L g687 ( 
.A(n_564),
.B(n_192),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_470),
.B(n_298),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_460),
.B(n_298),
.Y(n_689)
);

HB1xp67_ASAP7_75t_L g690 ( 
.A(n_568),
.Y(n_690)
);

INVxp67_ASAP7_75t_L g691 ( 
.A(n_509),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_491),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_566),
.B(n_301),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_485),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_SL g695 ( 
.A(n_498),
.B(n_161),
.Y(n_695)
);

NAND2xp33_ASAP7_75t_L g696 ( 
.A(n_573),
.B(n_499),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_513),
.A2(n_228),
.B1(n_197),
.B2(n_191),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_577),
.B(n_414),
.Y(n_698)
);

NOR2xp67_ASAP7_75t_L g699 ( 
.A(n_480),
.B(n_414),
.Y(n_699)
);

NAND3xp33_ASAP7_75t_L g700 ( 
.A(n_578),
.B(n_243),
.C(n_238),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_580),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_580),
.B(n_414),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_513),
.B(n_194),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_581),
.B(n_582),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_581),
.Y(n_705)
);

BUFx5_ASAP7_75t_L g706 ( 
.A(n_531),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_498),
.B(n_196),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_582),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_583),
.B(n_511),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_517),
.B(n_230),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_523),
.B(n_527),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_583),
.B(n_271),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_559),
.B(n_416),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_532),
.B(n_262),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_459),
.Y(n_715)
);

NAND2x1p5_ASAP7_75t_L g716 ( 
.A(n_495),
.B(n_416),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_499),
.A2(n_192),
.B1(n_436),
.B2(n_416),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_575),
.B(n_192),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_495),
.B(n_273),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_524),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_523),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_527),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_464),
.B(n_274),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_539),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_539),
.B(n_261),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_575),
.B(n_436),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_574),
.B(n_258),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_560),
.B(n_272),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_562),
.B(n_563),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_560),
.B(n_576),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_576),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_584),
.B(n_244),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_476),
.B(n_436),
.Y(n_733)
);

INVx2_ASAP7_75t_SL g734 ( 
.A(n_584),
.Y(n_734)
);

NAND3xp33_ASAP7_75t_L g735 ( 
.A(n_494),
.B(n_246),
.C(n_250),
.Y(n_735)
);

AND2x2_ASAP7_75t_SL g736 ( 
.A(n_507),
.B(n_368),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_512),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_524),
.Y(n_738)
);

INVx4_ASAP7_75t_L g739 ( 
.A(n_573),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_512),
.Y(n_740)
);

NAND3xp33_ASAP7_75t_L g741 ( 
.A(n_503),
.B(n_255),
.C(n_175),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_525),
.B(n_290),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_462),
.Y(n_743)
);

NAND2x1p5_ASAP7_75t_L g744 ( 
.A(n_571),
.B(n_367),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_571),
.B(n_318),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_562),
.B(n_290),
.Y(n_746)
);

BUFx2_ASAP7_75t_L g747 ( 
.A(n_522),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_573),
.A2(n_319),
.B(n_296),
.Y(n_748)
);

OR2x2_ASAP7_75t_L g749 ( 
.A(n_531),
.B(n_306),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_476),
.B(n_436),
.Y(n_750)
);

OR2x2_ASAP7_75t_L g751 ( 
.A(n_536),
.B(n_319),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_530),
.B(n_0),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_462),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_720),
.Y(n_754)
);

NOR2x1p5_ASAP7_75t_L g755 ( 
.A(n_596),
.B(n_694),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_636),
.B(n_518),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_639),
.B(n_518),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_737),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_589),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_740),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_587),
.B(n_562),
.Y(n_761)
);

HB1xp67_ASAP7_75t_L g762 ( 
.A(n_655),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_603),
.B(n_528),
.Y(n_763)
);

INVx4_ASAP7_75t_L g764 ( 
.A(n_720),
.Y(n_764)
);

OR2x6_ASAP7_75t_L g765 ( 
.A(n_630),
.B(n_522),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_720),
.Y(n_766)
);

OR2x6_ASAP7_75t_L g767 ( 
.A(n_630),
.B(n_522),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_711),
.B(n_528),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_592),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_709),
.B(n_529),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_588),
.Y(n_771)
);

NOR2xp67_ASAP7_75t_L g772 ( 
.A(n_673),
.B(n_557),
.Y(n_772)
);

AND2x4_ASAP7_75t_SL g773 ( 
.A(n_680),
.B(n_563),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_685),
.A2(n_522),
.B1(n_499),
.B2(n_529),
.Y(n_774)
);

AND3x2_ASAP7_75t_SL g775 ( 
.A(n_679),
.B(n_2),
.C(n_10),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_722),
.A2(n_499),
.B1(n_537),
.B2(n_536),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_738),
.Y(n_777)
);

INVx5_ASAP7_75t_L g778 ( 
.A(n_618),
.Y(n_778)
);

OR2x6_ASAP7_75t_L g779 ( 
.A(n_630),
.B(n_573),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_734),
.B(n_537),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_593),
.Y(n_781)
);

AND2x4_ASAP7_75t_L g782 ( 
.A(n_646),
.B(n_563),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_SL g783 ( 
.A1(n_695),
.A2(n_499),
.B1(n_573),
.B2(n_538),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_655),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_649),
.B(n_521),
.Y(n_785)
);

HB1xp67_ASAP7_75t_L g786 ( 
.A(n_618),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_682),
.A2(n_499),
.B1(n_483),
.B2(n_467),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_597),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_604),
.B(n_572),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_725),
.B(n_572),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_599),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_680),
.B(n_521),
.Y(n_792)
);

INVx3_ASAP7_75t_L g793 ( 
.A(n_738),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_695),
.B(n_572),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_747),
.A2(n_499),
.B1(n_483),
.B2(n_479),
.Y(n_795)
);

OR2x2_ASAP7_75t_L g796 ( 
.A(n_724),
.B(n_465),
.Y(n_796)
);

NOR3xp33_ASAP7_75t_L g797 ( 
.A(n_650),
.B(n_482),
.C(n_520),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_730),
.A2(n_489),
.B1(n_488),
.B2(n_479),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_704),
.B(n_465),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_738),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_680),
.B(n_611),
.Y(n_801)
);

INVx2_ASAP7_75t_SL g802 ( 
.A(n_618),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_SL g803 ( 
.A1(n_714),
.A2(n_520),
.B1(n_533),
.B2(n_496),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_601),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_691),
.B(n_478),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_606),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_721),
.B(n_521),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_605),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_621),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_622),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_613),
.Y(n_811)
);

CKINVDCx20_ASAP7_75t_R g812 ( 
.A(n_692),
.Y(n_812)
);

BUFx4f_ASAP7_75t_L g813 ( 
.A(n_634),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_609),
.B(n_496),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_635),
.B(n_521),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_739),
.A2(n_478),
.B(n_521),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_640),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_626),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_R g819 ( 
.A(n_598),
.B(n_447),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_657),
.Y(n_820)
);

INVxp33_ASAP7_75t_L g821 ( 
.A(n_707),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_644),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_608),
.B(n_488),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_628),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_731),
.A2(n_489),
.B1(n_555),
.B2(n_553),
.Y(n_825)
);

INVx4_ASAP7_75t_L g826 ( 
.A(n_634),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_629),
.Y(n_827)
);

AOI21x1_ASAP7_75t_L g828 ( 
.A1(n_656),
.A2(n_514),
.B(n_555),
.Y(n_828)
);

NOR2x1_ASAP7_75t_R g829 ( 
.A(n_723),
.B(n_545),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_609),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_706),
.B(n_514),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_625),
.B(n_533),
.Y(n_832)
);

HB1xp67_ASAP7_75t_L g833 ( 
.A(n_690),
.Y(n_833)
);

BUFx12f_ASAP7_75t_L g834 ( 
.A(n_635),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_693),
.A2(n_504),
.B1(n_553),
.B2(n_552),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_625),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_638),
.B(n_545),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_752),
.A2(n_502),
.B1(n_552),
.B2(n_551),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_638),
.B(n_545),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_631),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_598),
.B(n_478),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_632),
.Y(n_842)
);

INVxp67_ASAP7_75t_L g843 ( 
.A(n_728),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_659),
.B(n_477),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_661),
.B(n_477),
.Y(n_845)
);

NOR2x2_ASAP7_75t_L g846 ( 
.A(n_637),
.B(n_502),
.Y(n_846)
);

OR2x6_ASAP7_75t_L g847 ( 
.A(n_699),
.B(n_645),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_706),
.B(n_504),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_666),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_590),
.B(n_543),
.Y(n_850)
);

BUFx2_ASAP7_75t_L g851 ( 
.A(n_591),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_658),
.B(n_543),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_667),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_706),
.B(n_546),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_672),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_706),
.B(n_677),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_706),
.B(n_546),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_701),
.B(n_551),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_658),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_705),
.B(n_447),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_736),
.A2(n_550),
.B1(n_567),
.B2(n_549),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_708),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_665),
.A2(n_550),
.B1(n_477),
.B2(n_501),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_689),
.B(n_447),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_643),
.B(n_648),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_727),
.B(n_501),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_712),
.B(n_501),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_698),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_746),
.B(n_481),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_660),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_674),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_678),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_745),
.B(n_481),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_671),
.B(n_545),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_745),
.B(n_481),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_671),
.A2(n_436),
.B1(n_481),
.B2(n_463),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_607),
.B(n_481),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_744),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_698),
.Y(n_879)
);

INVxp67_ASAP7_75t_L g880 ( 
.A(n_732),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_652),
.A2(n_436),
.B1(n_463),
.B2(n_456),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_702),
.Y(n_882)
);

AND2x6_ASAP7_75t_L g883 ( 
.A(n_641),
.B(n_463),
.Y(n_883)
);

INVxp33_ASAP7_75t_SL g884 ( 
.A(n_676),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_702),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_749),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_710),
.B(n_545),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_715),
.Y(n_888)
);

AOI22xp5_ASAP7_75t_L g889 ( 
.A1(n_686),
.A2(n_436),
.B1(n_463),
.B2(n_456),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_654),
.B(n_456),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_751),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_612),
.B(n_463),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_663),
.B(n_456),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_664),
.B(n_456),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_686),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_743),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_753),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_669),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_675),
.A2(n_436),
.B1(n_545),
.B2(n_58),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_641),
.B(n_11),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_L g901 ( 
.A1(n_687),
.A2(n_56),
.B1(n_143),
.B2(n_134),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_616),
.Y(n_902)
);

NOR2x1p5_ASAP7_75t_L g903 ( 
.A(n_700),
.B(n_14),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_617),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_744),
.Y(n_905)
);

OR2x2_ASAP7_75t_L g906 ( 
.A(n_610),
.B(n_15),
.Y(n_906)
);

AND2x4_ASAP7_75t_L g907 ( 
.A(n_703),
.B(n_48),
.Y(n_907)
);

BUFx3_ASAP7_75t_L g908 ( 
.A(n_718),
.Y(n_908)
);

BUFx3_ASAP7_75t_L g909 ( 
.A(n_718),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_619),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_595),
.B(n_15),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_600),
.B(n_19),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_602),
.B(n_20),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_620),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_713),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_684),
.A2(n_633),
.B1(n_653),
.B2(n_651),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_642),
.B(n_22),
.Y(n_917)
);

BUFx4f_ASAP7_75t_L g918 ( 
.A(n_627),
.Y(n_918)
);

AND2x6_ASAP7_75t_L g919 ( 
.A(n_642),
.B(n_64),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_683),
.B(n_66),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_656),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_586),
.B(n_60),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_662),
.Y(n_923)
);

NAND3xp33_ASAP7_75t_SL g924 ( 
.A(n_585),
.B(n_23),
.C(n_24),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_610),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_662),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_688),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_681),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_615),
.Y(n_929)
);

AO22x1_ASAP7_75t_L g930 ( 
.A1(n_729),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_614),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_681),
.Y(n_932)
);

INVxp67_ASAP7_75t_L g933 ( 
.A(n_735),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_647),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_647),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_651),
.B(n_28),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_653),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_716),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_726),
.Y(n_939)
);

BUFx12f_ASAP7_75t_L g940 ( 
.A(n_784),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_771),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_884),
.B(n_865),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_769),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_754),
.Y(n_944)
);

AOI21x1_ASAP7_75t_L g945 ( 
.A1(n_785),
.A2(n_623),
.B(n_748),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_762),
.Y(n_946)
);

NOR2xp67_ASAP7_75t_SL g947 ( 
.A(n_778),
.B(n_741),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_790),
.A2(n_668),
.B1(n_719),
.B2(n_624),
.Y(n_948)
);

OAI22xp5_ASAP7_75t_L g949 ( 
.A1(n_923),
.A2(n_627),
.B1(n_716),
.B2(n_697),
.Y(n_949)
);

AOI221xp5_ASAP7_75t_L g950 ( 
.A1(n_925),
.A2(n_742),
.B1(n_594),
.B2(n_670),
.C(n_717),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_915),
.B(n_750),
.Y(n_951)
);

NAND3xp33_ASAP7_75t_SL g952 ( 
.A(n_911),
.B(n_912),
.C(n_913),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_843),
.A2(n_750),
.B1(n_733),
.B2(n_85),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_868),
.B(n_733),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_822),
.B(n_73),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_806),
.Y(n_956)
);

INVx1_ASAP7_75t_SL g957 ( 
.A(n_796),
.Y(n_957)
);

INVx2_ASAP7_75t_SL g958 ( 
.A(n_786),
.Y(n_958)
);

OAI21xp33_ASAP7_75t_L g959 ( 
.A1(n_759),
.A2(n_849),
.B(n_906),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_886),
.B(n_30),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_817),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_781),
.Y(n_962)
);

INVx3_ASAP7_75t_L g963 ( 
.A(n_754),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_799),
.A2(n_81),
.B(n_115),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_788),
.Y(n_965)
);

BUFx2_ASAP7_75t_L g966 ( 
.A(n_812),
.Y(n_966)
);

BUFx2_ASAP7_75t_L g967 ( 
.A(n_834),
.Y(n_967)
);

A2O1A1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_794),
.A2(n_31),
.B(n_33),
.C(n_36),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_791),
.Y(n_969)
);

NAND2x1p5_ASAP7_75t_L g970 ( 
.A(n_764),
.B(n_86),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_804),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_866),
.A2(n_88),
.B(n_108),
.Y(n_972)
);

INVxp67_ASAP7_75t_SL g973 ( 
.A(n_754),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_808),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_809),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_811),
.Y(n_976)
);

INVx3_ASAP7_75t_SL g977 ( 
.A(n_846),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_830),
.B(n_36),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_R g979 ( 
.A(n_813),
.B(n_72),
.Y(n_979)
);

BUFx10_ASAP7_75t_L g980 ( 
.A(n_755),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_820),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_833),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_932),
.A2(n_37),
.B1(n_39),
.B2(n_42),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_813),
.B(n_93),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_831),
.A2(n_105),
.B(n_106),
.Y(n_985)
);

AOI22xp33_ASAP7_75t_L g986 ( 
.A1(n_907),
.A2(n_44),
.B1(n_153),
.B2(n_920),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_921),
.A2(n_44),
.B1(n_928),
.B2(n_926),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_821),
.B(n_929),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_848),
.A2(n_857),
.B(n_854),
.Y(n_989)
);

AOI22xp5_ASAP7_75t_L g990 ( 
.A1(n_880),
.A2(n_931),
.B1(n_933),
.B2(n_927),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_836),
.B(n_891),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_766),
.B(n_777),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_851),
.B(n_761),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_766),
.B(n_777),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_870),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_826),
.B(n_847),
.Y(n_996)
);

NAND2x1_ASAP7_75t_L g997 ( 
.A(n_764),
.B(n_766),
.Y(n_997)
);

NOR2x1_ASAP7_75t_L g998 ( 
.A(n_826),
.B(n_793),
.Y(n_998)
);

NOR2x1_ASAP7_75t_SL g999 ( 
.A(n_779),
.B(n_938),
.Y(n_999)
);

NOR2x1_ASAP7_75t_L g1000 ( 
.A(n_793),
.B(n_924),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_879),
.B(n_882),
.Y(n_1001)
);

OR2x2_ASAP7_75t_SL g1002 ( 
.A(n_775),
.B(n_810),
.Y(n_1002)
);

INVx3_ASAP7_75t_L g1003 ( 
.A(n_777),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_885),
.A2(n_774),
.B1(n_916),
.B2(n_934),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_778),
.B(n_818),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_802),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_816),
.A2(n_875),
.B(n_873),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_871),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_895),
.A2(n_856),
.B(n_770),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_778),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_898),
.B(n_935),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_856),
.A2(n_770),
.B(n_867),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_800),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_937),
.B(n_757),
.Y(n_1014)
);

OAI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_916),
.A2(n_939),
.B(n_936),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_887),
.A2(n_864),
.B(n_763),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_824),
.B(n_827),
.Y(n_1017)
);

AND2x4_ASAP7_75t_SL g1018 ( 
.A(n_847),
.B(n_878),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_840),
.B(n_842),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_763),
.A2(n_756),
.B(n_823),
.Y(n_1020)
);

AOI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_847),
.A2(n_772),
.B1(n_832),
.B2(n_814),
.Y(n_1021)
);

NOR3xp33_ASAP7_75t_SL g1022 ( 
.A(n_841),
.B(n_862),
.C(n_853),
.Y(n_1022)
);

O2A1O1Ixp5_ASAP7_75t_SL g1023 ( 
.A1(n_922),
.A2(n_801),
.B(n_917),
.C(n_900),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_R g1024 ( 
.A(n_918),
.B(n_905),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_872),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_888),
.Y(n_1026)
);

INVx5_ASAP7_75t_L g1027 ( 
.A(n_779),
.Y(n_1027)
);

OAI22x1_ASAP7_75t_L g1028 ( 
.A1(n_903),
.A2(n_855),
.B1(n_795),
.B2(n_760),
.Y(n_1028)
);

AOI222xp33_ASAP7_75t_L g1029 ( 
.A1(n_930),
.A2(n_758),
.B1(n_768),
.B2(n_904),
.C1(n_902),
.C2(n_914),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_768),
.A2(n_910),
.B(n_877),
.C(n_815),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_789),
.A2(n_893),
.B(n_894),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_776),
.A2(n_861),
.B1(n_795),
.B2(n_918),
.Y(n_1032)
);

OR2x6_ASAP7_75t_L g1033 ( 
.A(n_779),
.B(n_765),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_765),
.A2(n_767),
.B1(n_783),
.B2(n_901),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_859),
.B(n_814),
.Y(n_1035)
);

NAND3xp33_ASAP7_75t_SL g1036 ( 
.A(n_901),
.B(n_797),
.C(n_805),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_890),
.A2(n_837),
.B(n_839),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_908),
.B(n_909),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_782),
.B(n_765),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_782),
.B(n_767),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_874),
.A2(n_892),
.B(n_792),
.Y(n_1041)
);

INVx1_ASAP7_75t_SL g1042 ( 
.A(n_780),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_R g1043 ( 
.A(n_905),
.B(n_878),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_859),
.B(n_832),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_859),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_787),
.A2(n_896),
.B(n_897),
.C(n_858),
.Y(n_1046)
);

NOR3xp33_ASAP7_75t_L g1047 ( 
.A(n_807),
.B(n_829),
.C(n_803),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_852),
.A2(n_773),
.B(n_860),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_767),
.A2(n_850),
.B1(n_852),
.B2(n_878),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_850),
.B(n_938),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_919),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_819),
.B(n_825),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_844),
.B(n_845),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_SL g1054 ( 
.A1(n_835),
.A2(n_881),
.B(n_863),
.C(n_876),
.Y(n_1054)
);

AOI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_883),
.A2(n_919),
.B1(n_825),
.B2(n_838),
.Y(n_1055)
);

INVx6_ASAP7_75t_L g1056 ( 
.A(n_919),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_798),
.A2(n_889),
.B(n_876),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_798),
.B(n_889),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_919),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_899),
.B(n_883),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_SL g1061 ( 
.A1(n_899),
.A2(n_500),
.B1(n_724),
.B2(n_422),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_R g1062 ( 
.A(n_811),
.B(n_485),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_759),
.B(n_516),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_865),
.B(n_508),
.Y(n_1064)
);

INVx1_ASAP7_75t_SL g1065 ( 
.A(n_762),
.Y(n_1065)
);

O2A1O1Ixp33_ASAP7_75t_SL g1066 ( 
.A1(n_922),
.A2(n_932),
.B(n_923),
.C(n_934),
.Y(n_1066)
);

NOR2x1_ASAP7_75t_SL g1067 ( 
.A(n_779),
.B(n_938),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_769),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_865),
.A2(n_636),
.B(n_649),
.C(n_911),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_865),
.B(n_508),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_869),
.A2(n_739),
.B(n_696),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_869),
.A2(n_739),
.B(n_696),
.Y(n_1072)
);

NOR2x1_ASAP7_75t_SL g1073 ( 
.A(n_779),
.B(n_938),
.Y(n_1073)
);

OAI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_923),
.A2(n_932),
.B1(n_921),
.B2(n_928),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_884),
.B(n_498),
.Y(n_1075)
);

NAND2x1p5_ASAP7_75t_L g1076 ( 
.A(n_764),
.B(n_754),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_762),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_1071),
.A2(n_1072),
.B(n_989),
.Y(n_1078)
);

INVx4_ASAP7_75t_L g1079 ( 
.A(n_944),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_1063),
.B(n_957),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_1069),
.A2(n_986),
.B1(n_1001),
.B2(n_1014),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_1027),
.Y(n_1082)
);

A2O1A1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_952),
.A2(n_948),
.B(n_1030),
.C(n_1058),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1011),
.B(n_1074),
.Y(n_1084)
);

OR2x6_ASAP7_75t_L g1085 ( 
.A(n_1033),
.B(n_996),
.Y(n_1085)
);

AO22x2_ASAP7_75t_L g1086 ( 
.A1(n_1034),
.A2(n_1032),
.B1(n_987),
.B2(n_983),
.Y(n_1086)
);

AO31x2_ASAP7_75t_L g1087 ( 
.A1(n_1004),
.A2(n_1031),
.A3(n_1032),
.B(n_1046),
.Y(n_1087)
);

INVxp67_ASAP7_75t_SL g1088 ( 
.A(n_1077),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_1012),
.A2(n_1020),
.B(n_1009),
.Y(n_1089)
);

OAI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_1015),
.A2(n_1023),
.B(n_1016),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_1057),
.A2(n_1041),
.B(n_1037),
.Y(n_1091)
);

CKINVDCx14_ASAP7_75t_R g1092 ( 
.A(n_1062),
.Y(n_1092)
);

BUFx3_ASAP7_75t_L g1093 ( 
.A(n_940),
.Y(n_1093)
);

OAI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_1015),
.A2(n_1036),
.B(n_1004),
.Y(n_1094)
);

INVxp67_ASAP7_75t_SL g1095 ( 
.A(n_1038),
.Y(n_1095)
);

AO21x1_ASAP7_75t_L g1096 ( 
.A1(n_1034),
.A2(n_949),
.B(n_1047),
.Y(n_1096)
);

OAI22x1_ASAP7_75t_L g1097 ( 
.A1(n_993),
.A2(n_977),
.B1(n_1021),
.B2(n_942),
.Y(n_1097)
);

NAND2x1_ASAP7_75t_L g1098 ( 
.A(n_1045),
.B(n_963),
.Y(n_1098)
);

AOI21xp33_ASAP7_75t_L g1099 ( 
.A1(n_1029),
.A2(n_1028),
.B(n_987),
.Y(n_1099)
);

O2A1O1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_968),
.A2(n_959),
.B(n_1064),
.C(n_1070),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_1048),
.A2(n_1051),
.B(n_1053),
.Y(n_1101)
);

NOR2x1_ASAP7_75t_L g1102 ( 
.A(n_982),
.B(n_1050),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_1027),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1066),
.A2(n_949),
.B(n_1054),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_957),
.B(n_1075),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1055),
.A2(n_954),
.B(n_953),
.Y(n_1106)
);

BUFx2_ASAP7_75t_L g1107 ( 
.A(n_946),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_SL g1108 ( 
.A1(n_999),
.A2(n_1073),
.B(n_1067),
.Y(n_1108)
);

OAI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_951),
.A2(n_1074),
.B(n_1060),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_962),
.Y(n_1110)
);

AND2x4_ASAP7_75t_L g1111 ( 
.A(n_996),
.B(n_1018),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_950),
.A2(n_1000),
.B(n_1022),
.C(n_1017),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1035),
.A2(n_1044),
.B(n_972),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_1051),
.A2(n_964),
.B(n_985),
.Y(n_1114)
);

AOI221xp5_ASAP7_75t_L g1115 ( 
.A1(n_1061),
.A2(n_983),
.B1(n_1019),
.B2(n_988),
.C(n_969),
.Y(n_1115)
);

AO21x2_ASAP7_75t_L g1116 ( 
.A1(n_992),
.A2(n_994),
.B(n_1049),
.Y(n_1116)
);

AO31x2_ASAP7_75t_L g1117 ( 
.A1(n_1005),
.A2(n_1068),
.A3(n_975),
.B(n_974),
.Y(n_1117)
);

NOR4xp25_ASAP7_75t_L g1118 ( 
.A(n_1042),
.B(n_1052),
.C(n_955),
.D(n_984),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_970),
.A2(n_998),
.B(n_1076),
.Y(n_1119)
);

INVx2_ASAP7_75t_SL g1120 ( 
.A(n_946),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1042),
.B(n_971),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1027),
.A2(n_1059),
.B(n_973),
.Y(n_1122)
);

INVx2_ASAP7_75t_SL g1123 ( 
.A(n_1065),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_970),
.A2(n_1076),
.B(n_997),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_991),
.B(n_1065),
.Y(n_1125)
);

HB1xp67_ASAP7_75t_L g1126 ( 
.A(n_958),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_965),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_941),
.A2(n_1026),
.B(n_981),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1029),
.B(n_961),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_990),
.A2(n_947),
.B(n_1039),
.C(n_1040),
.Y(n_1130)
);

OR2x2_ASAP7_75t_L g1131 ( 
.A(n_966),
.B(n_956),
.Y(n_1131)
);

CKINVDCx11_ASAP7_75t_R g1132 ( 
.A(n_980),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_995),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_1033),
.B(n_1027),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1008),
.B(n_1025),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_963),
.A2(n_1003),
.B(n_1010),
.Y(n_1136)
);

AOI221x1_ASAP7_75t_L g1137 ( 
.A1(n_978),
.A2(n_960),
.B1(n_1003),
.B2(n_1013),
.C(n_1045),
.Y(n_1137)
);

NOR2xp67_ASAP7_75t_L g1138 ( 
.A(n_976),
.B(n_1006),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1013),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_1033),
.B(n_1045),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1043),
.Y(n_1141)
);

OR2x6_ASAP7_75t_L g1142 ( 
.A(n_967),
.B(n_1056),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1024),
.B(n_980),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1056),
.Y(n_1144)
);

INVx2_ASAP7_75t_SL g1145 ( 
.A(n_979),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1002),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_1069),
.A2(n_865),
.B(n_952),
.C(n_636),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_SL g1148 ( 
.A(n_976),
.B(n_884),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_952),
.A2(n_1069),
.B(n_884),
.C(n_636),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_1075),
.B(n_884),
.Y(n_1150)
);

INVx3_ASAP7_75t_L g1151 ( 
.A(n_1027),
.Y(n_1151)
);

NOR2x1_ASAP7_75t_SL g1152 ( 
.A(n_1027),
.B(n_1033),
.Y(n_1152)
);

BUFx2_ASAP7_75t_L g1153 ( 
.A(n_940),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1001),
.B(n_1014),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_976),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_943),
.Y(n_1156)
);

OR2x2_ASAP7_75t_L g1157 ( 
.A(n_957),
.B(n_516),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1007),
.A2(n_828),
.B(n_945),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_1007),
.A2(n_828),
.B(n_945),
.Y(n_1159)
);

AO21x2_ASAP7_75t_L g1160 ( 
.A1(n_1036),
.A2(n_1015),
.B(n_1031),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_1007),
.A2(n_828),
.B(n_945),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1007),
.A2(n_828),
.B(n_945),
.Y(n_1162)
);

AO21x2_ASAP7_75t_L g1163 ( 
.A1(n_1036),
.A2(n_1015),
.B(n_1031),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_943),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_957),
.B(n_884),
.Y(n_1165)
);

AOI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_952),
.A2(n_884),
.B1(n_636),
.B2(n_724),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_943),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_976),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1063),
.B(n_516),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1001),
.B(n_1014),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_943),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1069),
.A2(n_865),
.B(n_952),
.C(n_636),
.Y(n_1172)
);

O2A1O1Ixp33_ASAP7_75t_SL g1173 ( 
.A1(n_1069),
.A2(n_1054),
.B(n_922),
.C(n_952),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_943),
.Y(n_1174)
);

INVx3_ASAP7_75t_SL g1175 ( 
.A(n_976),
.Y(n_1175)
);

BUFx2_ASAP7_75t_L g1176 ( 
.A(n_940),
.Y(n_1176)
);

OA21x2_ASAP7_75t_L g1177 ( 
.A1(n_1015),
.A2(n_1031),
.B(n_1016),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_943),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1001),
.B(n_1014),
.Y(n_1179)
);

INVx4_ASAP7_75t_L g1180 ( 
.A(n_944),
.Y(n_1180)
);

INVx3_ASAP7_75t_SL g1181 ( 
.A(n_976),
.Y(n_1181)
);

AOI21x1_ASAP7_75t_SL g1182 ( 
.A1(n_1064),
.A2(n_865),
.B(n_1070),
.Y(n_1182)
);

AND2x2_ASAP7_75t_SL g1183 ( 
.A(n_986),
.B(n_865),
.Y(n_1183)
);

NOR2xp67_ASAP7_75t_SL g1184 ( 
.A(n_976),
.B(n_811),
.Y(n_1184)
);

AOI221x1_ASAP7_75t_L g1185 ( 
.A1(n_952),
.A2(n_1069),
.B1(n_1036),
.B2(n_1028),
.C(n_1034),
.Y(n_1185)
);

NAND3xp33_ASAP7_75t_SL g1186 ( 
.A(n_1069),
.B(n_408),
.C(n_636),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_957),
.B(n_884),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_940),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_1075),
.B(n_884),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_944),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1007),
.A2(n_828),
.B(n_945),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1001),
.B(n_1014),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1069),
.A2(n_986),
.B1(n_1001),
.B2(n_884),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_1075),
.B(n_884),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1069),
.A2(n_1015),
.B(n_1012),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1069),
.A2(n_986),
.B1(n_1001),
.B2(n_884),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_957),
.B(n_884),
.Y(n_1197)
);

BUFx2_ASAP7_75t_R g1198 ( 
.A(n_976),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_943),
.Y(n_1199)
);

OA21x2_ASAP7_75t_L g1200 ( 
.A1(n_1015),
.A2(n_1031),
.B(n_1016),
.Y(n_1200)
);

OAI22x1_ASAP7_75t_L g1201 ( 
.A1(n_993),
.A2(n_925),
.B1(n_977),
.B2(n_539),
.Y(n_1201)
);

AO31x2_ASAP7_75t_L g1202 ( 
.A1(n_1004),
.A2(n_1031),
.A3(n_1032),
.B(n_1058),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1012),
.A2(n_1020),
.B(n_1031),
.Y(n_1203)
);

OAI22x1_ASAP7_75t_L g1204 ( 
.A1(n_993),
.A2(n_925),
.B1(n_977),
.B2(n_539),
.Y(n_1204)
);

OAI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_952),
.A2(n_413),
.B1(n_695),
.B2(n_408),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1001),
.B(n_1014),
.Y(n_1206)
);

NAND3x1_ASAP7_75t_L g1207 ( 
.A(n_1075),
.B(n_650),
.C(n_378),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1105),
.B(n_1205),
.Y(n_1208)
);

OAI221xp5_ASAP7_75t_L g1209 ( 
.A1(n_1166),
.A2(n_1149),
.B1(n_1147),
.B2(n_1172),
.C(n_1083),
.Y(n_1209)
);

AOI21xp33_ASAP7_75t_L g1210 ( 
.A1(n_1183),
.A2(n_1196),
.B(n_1193),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_SL g1211 ( 
.A1(n_1152),
.A2(n_1100),
.B(n_1096),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1174),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1169),
.B(n_1154),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_1107),
.Y(n_1214)
);

AO21x2_ASAP7_75t_L g1215 ( 
.A1(n_1090),
.A2(n_1104),
.B(n_1203),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1178),
.Y(n_1216)
);

CKINVDCx6p67_ASAP7_75t_R g1217 ( 
.A(n_1175),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1154),
.B(n_1170),
.Y(n_1218)
);

OR2x2_ASAP7_75t_L g1219 ( 
.A(n_1157),
.B(n_1080),
.Y(n_1219)
);

AO21x1_ASAP7_75t_L g1220 ( 
.A1(n_1081),
.A2(n_1196),
.B(n_1193),
.Y(n_1220)
);

OAI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1186),
.A2(n_1112),
.B(n_1207),
.Y(n_1221)
);

HB1xp67_ASAP7_75t_L g1222 ( 
.A(n_1125),
.Y(n_1222)
);

NOR2xp67_ASAP7_75t_L g1223 ( 
.A(n_1155),
.B(n_1168),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1081),
.A2(n_1094),
.B(n_1185),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1127),
.Y(n_1225)
);

INVx4_ASAP7_75t_L g1226 ( 
.A(n_1134),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1156),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1094),
.A2(n_1115),
.B1(n_1099),
.B2(n_1106),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1115),
.A2(n_1099),
.B1(n_1106),
.B2(n_1195),
.Y(n_1229)
);

OR2x2_ASAP7_75t_L g1230 ( 
.A(n_1121),
.B(n_1131),
.Y(n_1230)
);

OR2x2_ASAP7_75t_L g1231 ( 
.A(n_1121),
.B(n_1165),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1170),
.B(n_1179),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1179),
.B(n_1192),
.Y(n_1233)
);

CKINVDCx6p67_ASAP7_75t_R g1234 ( 
.A(n_1181),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_SL g1235 ( 
.A(n_1198),
.B(n_1184),
.Y(n_1235)
);

INVx1_ASAP7_75t_SL g1236 ( 
.A(n_1187),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1198),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1164),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1167),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1161),
.A2(n_1162),
.B(n_1191),
.Y(n_1240)
);

O2A1O1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1173),
.A2(n_1130),
.B(n_1146),
.C(n_1197),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1171),
.Y(n_1242)
);

BUFx2_ASAP7_75t_L g1243 ( 
.A(n_1120),
.Y(n_1243)
);

OA21x2_ASAP7_75t_L g1244 ( 
.A1(n_1078),
.A2(n_1091),
.B(n_1114),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1199),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1192),
.A2(n_1206),
.B1(n_1150),
.B2(n_1189),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1206),
.B(n_1202),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_SL g1248 ( 
.A1(n_1084),
.A2(n_1129),
.B(n_1113),
.Y(n_1248)
);

BUFx10_ASAP7_75t_L g1249 ( 
.A(n_1111),
.Y(n_1249)
);

AO21x2_ASAP7_75t_L g1250 ( 
.A1(n_1160),
.A2(n_1163),
.B(n_1118),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_SL g1251 ( 
.A1(n_1084),
.A2(n_1129),
.B(n_1122),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1101),
.A2(n_1182),
.B(n_1119),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1202),
.B(n_1095),
.Y(n_1253)
);

O2A1O1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1194),
.A2(n_1141),
.B(n_1118),
.C(n_1123),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1177),
.A2(n_1200),
.B(n_1124),
.Y(n_1255)
);

AO21x2_ASAP7_75t_L g1256 ( 
.A1(n_1116),
.A2(n_1136),
.B(n_1128),
.Y(n_1256)
);

OA21x2_ASAP7_75t_L g1257 ( 
.A1(n_1137),
.A2(n_1135),
.B(n_1133),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1135),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1177),
.A2(n_1200),
.B(n_1082),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1082),
.A2(n_1103),
.B(n_1151),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1103),
.A2(n_1151),
.B(n_1108),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1102),
.A2(n_1145),
.B(n_1148),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1087),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1098),
.A2(n_1144),
.B(n_1139),
.Y(n_1264)
);

CKINVDCx11_ASAP7_75t_R g1265 ( 
.A(n_1132),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1087),
.A2(n_1202),
.B(n_1143),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1117),
.Y(n_1267)
);

INVx2_ASAP7_75t_SL g1268 ( 
.A(n_1111),
.Y(n_1268)
);

NOR2x1_ASAP7_75t_SL g1269 ( 
.A(n_1116),
.B(n_1085),
.Y(n_1269)
);

CKINVDCx11_ASAP7_75t_R g1270 ( 
.A(n_1153),
.Y(n_1270)
);

OAI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1148),
.A2(n_1088),
.B(n_1126),
.Y(n_1271)
);

INVx1_ASAP7_75t_SL g1272 ( 
.A(n_1201),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1204),
.B(n_1097),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1117),
.Y(n_1274)
);

OR2x2_ASAP7_75t_L g1275 ( 
.A(n_1085),
.B(n_1142),
.Y(n_1275)
);

BUFx3_ASAP7_75t_L g1276 ( 
.A(n_1142),
.Y(n_1276)
);

OR2x6_ASAP7_75t_L g1277 ( 
.A(n_1085),
.B(n_1142),
.Y(n_1277)
);

NAND2x1p5_ASAP7_75t_L g1278 ( 
.A(n_1140),
.B(n_1138),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1079),
.A2(n_1180),
.B(n_1190),
.Y(n_1279)
);

AO21x2_ASAP7_75t_L g1280 ( 
.A1(n_1092),
.A2(n_1176),
.B(n_1188),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1093),
.A2(n_952),
.B1(n_1183),
.B2(n_1205),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1183),
.A2(n_952),
.B1(n_1205),
.B2(n_1186),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_SL g1283 ( 
.A1(n_1183),
.A2(n_498),
.B1(n_408),
.B2(n_884),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1134),
.B(n_1085),
.Y(n_1284)
);

BUFx2_ASAP7_75t_L g1285 ( 
.A(n_1107),
.Y(n_1285)
);

NAND2x1p5_ASAP7_75t_L g1286 ( 
.A(n_1134),
.B(n_1027),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_SL g1287 ( 
.A1(n_1152),
.A2(n_1100),
.B(n_1096),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1169),
.B(n_1154),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1110),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1107),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1110),
.Y(n_1291)
);

NAND2xp33_ASAP7_75t_SL g1292 ( 
.A(n_1154),
.B(n_1024),
.Y(n_1292)
);

OAI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1147),
.A2(n_1069),
.B(n_636),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1158),
.A2(n_1161),
.B(n_1159),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_SL g1295 ( 
.A1(n_1183),
.A2(n_498),
.B1(n_408),
.B2(n_884),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1158),
.A2(n_1161),
.B(n_1159),
.Y(n_1296)
);

INVx2_ASAP7_75t_SL g1297 ( 
.A(n_1120),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1110),
.Y(n_1298)
);

AND2x4_ASAP7_75t_L g1299 ( 
.A(n_1134),
.B(n_1085),
.Y(n_1299)
);

BUFx3_ASAP7_75t_L g1300 ( 
.A(n_1107),
.Y(n_1300)
);

NAND2x1p5_ASAP7_75t_L g1301 ( 
.A(n_1134),
.B(n_1027),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1110),
.Y(n_1302)
);

OAI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1147),
.A2(n_1069),
.B(n_636),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1198),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1109),
.B(n_1086),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1110),
.Y(n_1306)
);

NOR2xp67_ASAP7_75t_L g1307 ( 
.A(n_1155),
.B(n_976),
.Y(n_1307)
);

AOI21xp33_ASAP7_75t_L g1308 ( 
.A1(n_1149),
.A2(n_865),
.B(n_636),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1169),
.B(n_1154),
.Y(n_1309)
);

OAI222xp33_ASAP7_75t_L g1310 ( 
.A1(n_1205),
.A2(n_986),
.B1(n_925),
.B2(n_906),
.C1(n_1196),
.C2(n_1193),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1183),
.A2(n_952),
.B1(n_1205),
.B2(n_1186),
.Y(n_1311)
);

OAI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1147),
.A2(n_1069),
.B(n_636),
.Y(n_1312)
);

OA21x2_ASAP7_75t_L g1313 ( 
.A1(n_1090),
.A2(n_1104),
.B(n_1089),
.Y(n_1313)
);

BUFx4f_ASAP7_75t_L g1314 ( 
.A(n_1085),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1169),
.B(n_1154),
.Y(n_1315)
);

NAND2x1p5_ASAP7_75t_L g1316 ( 
.A(n_1134),
.B(n_1027),
.Y(n_1316)
);

AOI21x1_ASAP7_75t_SL g1317 ( 
.A1(n_1273),
.A2(n_1233),
.B(n_1218),
.Y(n_1317)
);

CKINVDCx20_ASAP7_75t_R g1318 ( 
.A(n_1265),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1232),
.B(n_1247),
.Y(n_1319)
);

BUFx6f_ASAP7_75t_L g1320 ( 
.A(n_1276),
.Y(n_1320)
);

OA21x2_ASAP7_75t_L g1321 ( 
.A1(n_1224),
.A2(n_1255),
.B(n_1259),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1232),
.B(n_1247),
.Y(n_1322)
);

OA21x2_ASAP7_75t_L g1323 ( 
.A1(n_1255),
.A2(n_1259),
.B(n_1240),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1228),
.B(n_1229),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1208),
.B(n_1222),
.Y(n_1325)
);

INVx1_ASAP7_75t_SL g1326 ( 
.A(n_1231),
.Y(n_1326)
);

A2O1A1Ixp33_ASAP7_75t_L g1327 ( 
.A1(n_1221),
.A2(n_1308),
.B(n_1312),
.C(n_1303),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1208),
.B(n_1219),
.Y(n_1328)
);

O2A1O1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1310),
.A2(n_1293),
.B(n_1209),
.C(n_1246),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1228),
.A2(n_1229),
.B1(n_1295),
.B2(n_1283),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1282),
.A2(n_1311),
.B1(n_1281),
.B2(n_1315),
.Y(n_1331)
);

O2A1O1Ixp5_ASAP7_75t_L g1332 ( 
.A1(n_1220),
.A2(n_1210),
.B(n_1292),
.C(n_1271),
.Y(n_1332)
);

INVxp67_ASAP7_75t_L g1333 ( 
.A(n_1290),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1213),
.B(n_1288),
.Y(n_1334)
);

AOI221x1_ASAP7_75t_SL g1335 ( 
.A1(n_1309),
.A2(n_1238),
.B1(n_1242),
.B2(n_1245),
.C(n_1227),
.Y(n_1335)
);

O2A1O1Ixp5_ASAP7_75t_L g1336 ( 
.A1(n_1292),
.A2(n_1263),
.B(n_1267),
.C(n_1274),
.Y(n_1336)
);

O2A1O1Ixp33_ASAP7_75t_L g1337 ( 
.A1(n_1241),
.A2(n_1254),
.B(n_1311),
.C(n_1282),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1281),
.A2(n_1314),
.B1(n_1230),
.B2(n_1277),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1253),
.B(n_1305),
.Y(n_1339)
);

INVx1_ASAP7_75t_SL g1340 ( 
.A(n_1285),
.Y(n_1340)
);

AND2x4_ASAP7_75t_L g1341 ( 
.A(n_1284),
.B(n_1299),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_SL g1342 ( 
.A1(n_1262),
.A2(n_1277),
.B(n_1286),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1314),
.A2(n_1277),
.B1(n_1236),
.B2(n_1272),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1314),
.A2(n_1277),
.B1(n_1239),
.B2(n_1305),
.Y(n_1344)
);

AND2x4_ASAP7_75t_L g1345 ( 
.A(n_1284),
.B(n_1299),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1212),
.A2(n_1289),
.B1(n_1306),
.B2(n_1298),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1216),
.A2(n_1278),
.B1(n_1276),
.B2(n_1275),
.Y(n_1347)
);

NOR2xp67_ASAP7_75t_L g1348 ( 
.A(n_1307),
.B(n_1297),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1214),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1258),
.B(n_1248),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1300),
.B(n_1291),
.Y(n_1351)
);

O2A1O1Ixp33_ASAP7_75t_L g1352 ( 
.A1(n_1251),
.A2(n_1211),
.B(n_1287),
.C(n_1278),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1266),
.B(n_1263),
.Y(n_1353)
);

NOR2xp67_ASAP7_75t_L g1354 ( 
.A(n_1223),
.B(n_1226),
.Y(n_1354)
);

CKINVDCx6p67_ASAP7_75t_R g1355 ( 
.A(n_1265),
.Y(n_1355)
);

AOI21x1_ASAP7_75t_SL g1356 ( 
.A1(n_1217),
.A2(n_1234),
.B(n_1269),
.Y(n_1356)
);

OAI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1237),
.A2(n_1304),
.B1(n_1302),
.B2(n_1243),
.Y(n_1357)
);

AND2x4_ASAP7_75t_L g1358 ( 
.A(n_1268),
.B(n_1280),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_SL g1359 ( 
.A1(n_1286),
.A2(n_1316),
.B(n_1301),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1257),
.B(n_1215),
.Y(n_1360)
);

OR2x2_ASAP7_75t_L g1361 ( 
.A(n_1280),
.B(n_1257),
.Y(n_1361)
);

INVx1_ASAP7_75t_SL g1362 ( 
.A(n_1280),
.Y(n_1362)
);

AOI21x1_ASAP7_75t_SL g1363 ( 
.A1(n_1217),
.A2(n_1234),
.B(n_1235),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1264),
.Y(n_1364)
);

AOI21x1_ASAP7_75t_SL g1365 ( 
.A1(n_1270),
.A2(n_1304),
.B(n_1237),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1260),
.Y(n_1366)
);

INVx3_ASAP7_75t_SL g1367 ( 
.A(n_1249),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1250),
.B(n_1316),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1249),
.B(n_1301),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1260),
.Y(n_1370)
);

CKINVDCx8_ASAP7_75t_R g1371 ( 
.A(n_1270),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1250),
.B(n_1313),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1256),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1250),
.B(n_1313),
.Y(n_1374)
);

OR2x6_ASAP7_75t_L g1375 ( 
.A(n_1261),
.B(n_1252),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1244),
.A2(n_1279),
.B1(n_1294),
.B2(n_1296),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1225),
.Y(n_1377)
);

NOR2x1_ASAP7_75t_L g1378 ( 
.A(n_1246),
.B(n_1262),
.Y(n_1378)
);

CKINVDCx20_ASAP7_75t_R g1379 ( 
.A(n_1265),
.Y(n_1379)
);

OA21x2_ASAP7_75t_L g1380 ( 
.A1(n_1224),
.A2(n_1090),
.B(n_1104),
.Y(n_1380)
);

NOR2x1_ASAP7_75t_SL g1381 ( 
.A(n_1344),
.B(n_1368),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1366),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1370),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1339),
.B(n_1360),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1339),
.B(n_1360),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_SL g1386 ( 
.A1(n_1329),
.A2(n_1327),
.B(n_1337),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1323),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_1358),
.Y(n_1388)
);

HB1xp67_ASAP7_75t_L g1389 ( 
.A(n_1353),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1361),
.B(n_1374),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1372),
.B(n_1362),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_1362),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1380),
.B(n_1319),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1380),
.B(n_1319),
.Y(n_1394)
);

NOR2x1_ASAP7_75t_SL g1395 ( 
.A(n_1344),
.B(n_1350),
.Y(n_1395)
);

CKINVDCx11_ASAP7_75t_R g1396 ( 
.A(n_1379),
.Y(n_1396)
);

BUFx6f_ASAP7_75t_L g1397 ( 
.A(n_1321),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1322),
.B(n_1335),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1322),
.B(n_1321),
.Y(n_1399)
);

INVx3_ASAP7_75t_L g1400 ( 
.A(n_1375),
.Y(n_1400)
);

AND4x1_ASAP7_75t_L g1401 ( 
.A(n_1378),
.B(n_1332),
.C(n_1342),
.D(n_1352),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1330),
.A2(n_1331),
.B1(n_1324),
.B2(n_1328),
.Y(n_1402)
);

BUFx8_ASAP7_75t_SL g1403 ( 
.A(n_1318),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1373),
.B(n_1326),
.Y(n_1404)
);

AND2x4_ASAP7_75t_L g1405 ( 
.A(n_1375),
.B(n_1364),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1377),
.Y(n_1406)
);

BUFx2_ASAP7_75t_L g1407 ( 
.A(n_1375),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1350),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1335),
.B(n_1326),
.Y(n_1409)
);

INVx5_ASAP7_75t_L g1410 ( 
.A(n_1358),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1376),
.A2(n_1336),
.B(n_1356),
.Y(n_1411)
);

OR2x2_ASAP7_75t_L g1412 ( 
.A(n_1325),
.B(n_1351),
.Y(n_1412)
);

INVx2_ASAP7_75t_SL g1413 ( 
.A(n_1341),
.Y(n_1413)
);

BUFx2_ASAP7_75t_SL g1414 ( 
.A(n_1347),
.Y(n_1414)
);

OA21x2_ASAP7_75t_L g1415 ( 
.A1(n_1346),
.A2(n_1330),
.B(n_1338),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1334),
.B(n_1331),
.Y(n_1416)
);

BUFx3_ASAP7_75t_L g1417 ( 
.A(n_1341),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1392),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1393),
.B(n_1394),
.Y(n_1419)
);

NOR2x1_ASAP7_75t_L g1420 ( 
.A(n_1408),
.B(n_1346),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1393),
.B(n_1340),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1392),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1389),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1382),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1394),
.B(n_1340),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1384),
.B(n_1333),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1384),
.B(n_1347),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_1403),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1389),
.Y(n_1429)
);

NAND2x1_ASAP7_75t_L g1430 ( 
.A(n_1405),
.B(n_1359),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1399),
.B(n_1345),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1399),
.B(n_1338),
.Y(n_1432)
);

OR2x6_ASAP7_75t_L g1433 ( 
.A(n_1414),
.B(n_1343),
.Y(n_1433)
);

AOI221xp5_ASAP7_75t_L g1434 ( 
.A1(n_1386),
.A2(n_1402),
.B1(n_1398),
.B2(n_1416),
.C(n_1409),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1384),
.B(n_1349),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1383),
.Y(n_1436)
);

OAI221xp5_ASAP7_75t_L g1437 ( 
.A1(n_1402),
.A2(n_1371),
.B1(n_1357),
.B2(n_1348),
.C(n_1354),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1385),
.B(n_1357),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_SL g1439 ( 
.A(n_1401),
.B(n_1320),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1436),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1424),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1436),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1418),
.Y(n_1443)
);

OAI31xp33_ASAP7_75t_L g1444 ( 
.A1(n_1437),
.A2(n_1416),
.A3(n_1409),
.B(n_1401),
.Y(n_1444)
);

NAND3xp33_ASAP7_75t_SL g1445 ( 
.A(n_1434),
.B(n_1398),
.C(n_1408),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1419),
.B(n_1410),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1422),
.Y(n_1447)
);

HB1xp67_ASAP7_75t_L g1448 ( 
.A(n_1422),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1419),
.B(n_1410),
.Y(n_1449)
);

AOI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1434),
.A2(n_1415),
.B1(n_1414),
.B2(n_1355),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1423),
.B(n_1385),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1437),
.A2(n_1415),
.B1(n_1414),
.B2(n_1413),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_1430),
.Y(n_1453)
);

NAND3xp33_ASAP7_75t_L g1454 ( 
.A(n_1420),
.B(n_1415),
.C(n_1404),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_SL g1455 ( 
.A1(n_1433),
.A2(n_1415),
.B1(n_1413),
.B2(n_1395),
.Y(n_1455)
);

OA21x2_ASAP7_75t_L g1456 ( 
.A1(n_1424),
.A2(n_1411),
.B(n_1387),
.Y(n_1456)
);

NAND4xp25_ASAP7_75t_L g1457 ( 
.A(n_1420),
.B(n_1404),
.C(n_1390),
.D(n_1391),
.Y(n_1457)
);

INVxp67_ASAP7_75t_L g1458 ( 
.A(n_1435),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1433),
.A2(n_1415),
.B1(n_1413),
.B2(n_1417),
.Y(n_1459)
);

INVx2_ASAP7_75t_SL g1460 ( 
.A(n_1431),
.Y(n_1460)
);

NOR2x1_ASAP7_75t_SL g1461 ( 
.A(n_1433),
.B(n_1439),
.Y(n_1461)
);

BUFx2_ASAP7_75t_L g1462 ( 
.A(n_1423),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1419),
.B(n_1410),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1439),
.A2(n_1415),
.B1(n_1433),
.B2(n_1438),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_1428),
.Y(n_1465)
);

OAI31xp33_ASAP7_75t_SL g1466 ( 
.A1(n_1432),
.A2(n_1395),
.A3(n_1411),
.B(n_1369),
.Y(n_1466)
);

OAI221xp5_ASAP7_75t_L g1467 ( 
.A1(n_1438),
.A2(n_1407),
.B1(n_1390),
.B2(n_1400),
.C(n_1412),
.Y(n_1467)
);

NOR4xp25_ASAP7_75t_SL g1468 ( 
.A(n_1428),
.B(n_1407),
.C(n_1381),
.D(n_1406),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_SL g1469 ( 
.A1(n_1433),
.A2(n_1381),
.B1(n_1410),
.B2(n_1388),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1433),
.A2(n_1417),
.B1(n_1388),
.B2(n_1412),
.Y(n_1470)
);

AOI211xp5_ASAP7_75t_L g1471 ( 
.A1(n_1432),
.A2(n_1367),
.B(n_1397),
.C(n_1317),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1440),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1457),
.B(n_1429),
.Y(n_1473)
);

NOR2x1_ASAP7_75t_L g1474 ( 
.A(n_1454),
.B(n_1433),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1456),
.Y(n_1475)
);

BUFx3_ASAP7_75t_L g1476 ( 
.A(n_1453),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1446),
.B(n_1421),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1456),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1453),
.Y(n_1479)
);

INVxp67_ASAP7_75t_L g1480 ( 
.A(n_1443),
.Y(n_1480)
);

INVx3_ASAP7_75t_L g1481 ( 
.A(n_1453),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1462),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1442),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1462),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1447),
.Y(n_1485)
);

NOR2x1p5_ASAP7_75t_L g1486 ( 
.A(n_1445),
.B(n_1454),
.Y(n_1486)
);

INVx4_ASAP7_75t_SL g1487 ( 
.A(n_1455),
.Y(n_1487)
);

INVxp67_ASAP7_75t_L g1488 ( 
.A(n_1448),
.Y(n_1488)
);

OR2x6_ASAP7_75t_L g1489 ( 
.A(n_1455),
.B(n_1400),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1446),
.B(n_1421),
.Y(n_1490)
);

NAND3xp33_ASAP7_75t_L g1491 ( 
.A(n_1444),
.B(n_1426),
.C(n_1396),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1457),
.B(n_1429),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1449),
.B(n_1421),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1486),
.B(n_1458),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1474),
.B(n_1449),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1472),
.Y(n_1496)
);

INVxp67_ASAP7_75t_SL g1497 ( 
.A(n_1486),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1474),
.B(n_1463),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1479),
.B(n_1463),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1475),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1479),
.B(n_1461),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1491),
.A2(n_1464),
.B1(n_1444),
.B2(n_1450),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_SL g1503 ( 
.A(n_1491),
.B(n_1471),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1472),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1479),
.B(n_1461),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1472),
.Y(n_1506)
);

NAND4xp25_ASAP7_75t_L g1507 ( 
.A(n_1473),
.B(n_1450),
.C(n_1452),
.D(n_1471),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1475),
.Y(n_1508)
);

AND2x4_ASAP7_75t_L g1509 ( 
.A(n_1487),
.B(n_1441),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1475),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1484),
.Y(n_1511)
);

AOI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1487),
.A2(n_1464),
.B1(n_1459),
.B2(n_1432),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1487),
.B(n_1477),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1480),
.B(n_1451),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1487),
.B(n_1466),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1480),
.B(n_1451),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1483),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1488),
.B(n_1425),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1487),
.B(n_1477),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1475),
.Y(n_1520)
);

INVx1_ASAP7_75t_SL g1521 ( 
.A(n_1482),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1487),
.B(n_1466),
.Y(n_1522)
);

OAI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1473),
.A2(n_1469),
.B(n_1467),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1487),
.B(n_1460),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1477),
.B(n_1490),
.Y(n_1525)
);

INVx2_ASAP7_75t_SL g1526 ( 
.A(n_1482),
.Y(n_1526)
);

OR2x6_ASAP7_75t_L g1527 ( 
.A(n_1489),
.B(n_1476),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1473),
.B(n_1427),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1490),
.B(n_1460),
.Y(n_1529)
);

BUFx2_ASAP7_75t_L g1530 ( 
.A(n_1484),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1490),
.B(n_1468),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1478),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1488),
.B(n_1425),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1513),
.B(n_1476),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1511),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1511),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1528),
.B(n_1492),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1513),
.B(n_1476),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1526),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1513),
.B(n_1519),
.Y(n_1540)
);

INVx2_ASAP7_75t_SL g1541 ( 
.A(n_1526),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1519),
.B(n_1476),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_SL g1543 ( 
.A(n_1497),
.B(n_1465),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1497),
.B(n_1494),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1496),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1519),
.B(n_1481),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1496),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1504),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1528),
.B(n_1492),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1514),
.B(n_1492),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1514),
.B(n_1485),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1515),
.B(n_1522),
.Y(n_1552)
);

INVx2_ASAP7_75t_SL g1553 ( 
.A(n_1526),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1530),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1516),
.B(n_1485),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1515),
.B(n_1481),
.Y(n_1556)
);

OAI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1502),
.A2(n_1489),
.B1(n_1470),
.B2(n_1468),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1530),
.Y(n_1558)
);

HB1xp67_ASAP7_75t_L g1559 ( 
.A(n_1521),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1504),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1525),
.Y(n_1561)
);

INVxp67_ASAP7_75t_L g1562 ( 
.A(n_1494),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1506),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1506),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1503),
.B(n_1493),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1517),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1516),
.B(n_1499),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1517),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1544),
.B(n_1507),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1540),
.B(n_1499),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1565),
.B(n_1507),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1567),
.B(n_1518),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1543),
.B(n_1403),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1562),
.B(n_1518),
.Y(n_1574)
);

CKINVDCx16_ASAP7_75t_R g1575 ( 
.A(n_1540),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1534),
.B(n_1499),
.Y(n_1576)
);

AND2x4_ASAP7_75t_SL g1577 ( 
.A(n_1538),
.B(n_1524),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1535),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_1559),
.Y(n_1579)
);

INVx1_ASAP7_75t_SL g1580 ( 
.A(n_1534),
.Y(n_1580)
);

NAND3xp33_ASAP7_75t_L g1581 ( 
.A(n_1557),
.B(n_1523),
.C(n_1512),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1558),
.B(n_1396),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1552),
.A2(n_1523),
.B1(n_1512),
.B2(n_1515),
.Y(n_1583)
);

NAND2x1_ASAP7_75t_L g1584 ( 
.A(n_1538),
.B(n_1501),
.Y(n_1584)
);

INVx1_ASAP7_75t_SL g1585 ( 
.A(n_1542),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1545),
.Y(n_1586)
);

INVx1_ASAP7_75t_SL g1587 ( 
.A(n_1542),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1554),
.B(n_1525),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1541),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1545),
.Y(n_1590)
);

INVxp33_ASAP7_75t_L g1591 ( 
.A(n_1552),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1554),
.B(n_1525),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1550),
.B(n_1533),
.Y(n_1593)
);

AOI21xp33_ASAP7_75t_L g1594 ( 
.A1(n_1591),
.A2(n_1553),
.B(n_1541),
.Y(n_1594)
);

OAI221xp5_ASAP7_75t_L g1595 ( 
.A1(n_1581),
.A2(n_1550),
.B1(n_1522),
.B2(n_1527),
.C(n_1537),
.Y(n_1595)
);

OAI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1569),
.A2(n_1527),
.B1(n_1549),
.B2(n_1537),
.Y(n_1596)
);

AOI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1583),
.A2(n_1522),
.B1(n_1538),
.B2(n_1527),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1573),
.B(n_1582),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1586),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1580),
.B(n_1536),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1575),
.B(n_1551),
.Y(n_1601)
);

INVx1_ASAP7_75t_SL g1602 ( 
.A(n_1577),
.Y(n_1602)
);

OAI31xp33_ASAP7_75t_L g1603 ( 
.A1(n_1583),
.A2(n_1501),
.A3(n_1505),
.B(n_1521),
.Y(n_1603)
);

XNOR2x1_ASAP7_75t_L g1604 ( 
.A(n_1571),
.B(n_1527),
.Y(n_1604)
);

NAND2x1_ASAP7_75t_L g1605 ( 
.A(n_1570),
.B(n_1553),
.Y(n_1605)
);

AOI221xp5_ASAP7_75t_SL g1606 ( 
.A1(n_1585),
.A2(n_1546),
.B1(n_1556),
.B2(n_1531),
.C(n_1501),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1576),
.B(n_1546),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1587),
.B(n_1536),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1579),
.B(n_1561),
.Y(n_1609)
);

OAI21xp33_ASAP7_75t_L g1610 ( 
.A1(n_1591),
.A2(n_1549),
.B(n_1551),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1582),
.A2(n_1527),
.B1(n_1561),
.B2(n_1531),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1578),
.A2(n_1527),
.B1(n_1531),
.B2(n_1555),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1602),
.B(n_1589),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1601),
.B(n_1589),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1605),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_L g1616 ( 
.A(n_1598),
.B(n_1573),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1600),
.B(n_1588),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1607),
.B(n_1577),
.Y(n_1618)
);

INVx1_ASAP7_75t_SL g1619 ( 
.A(n_1604),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1608),
.Y(n_1620)
);

AOI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1597),
.A2(n_1592),
.B1(n_1590),
.B2(n_1584),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1610),
.B(n_1574),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1611),
.B(n_1556),
.Y(n_1623)
);

AOI222xp33_ASAP7_75t_L g1624 ( 
.A1(n_1622),
.A2(n_1595),
.B1(n_1612),
.B2(n_1596),
.C1(n_1609),
.C2(n_1599),
.Y(n_1624)
);

AOI211xp5_ASAP7_75t_L g1625 ( 
.A1(n_1616),
.A2(n_1596),
.B(n_1594),
.C(n_1603),
.Y(n_1625)
);

AOI221xp5_ASAP7_75t_L g1626 ( 
.A1(n_1620),
.A2(n_1612),
.B1(n_1606),
.B2(n_1539),
.C(n_1593),
.Y(n_1626)
);

O2A1O1Ixp33_ASAP7_75t_L g1627 ( 
.A1(n_1614),
.A2(n_1539),
.B(n_1555),
.C(n_1572),
.Y(n_1627)
);

AOI31xp33_ASAP7_75t_L g1628 ( 
.A1(n_1619),
.A2(n_1505),
.A3(n_1495),
.B(n_1498),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1613),
.Y(n_1629)
);

AOI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1623),
.A2(n_1505),
.B1(n_1524),
.B2(n_1495),
.Y(n_1630)
);

NOR3x1_ASAP7_75t_L g1631 ( 
.A(n_1617),
.B(n_1564),
.C(n_1563),
.Y(n_1631)
);

NAND2xp33_ASAP7_75t_R g1632 ( 
.A(n_1615),
.B(n_1524),
.Y(n_1632)
);

AOI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1621),
.A2(n_1568),
.B(n_1548),
.Y(n_1633)
);

AOI221xp5_ASAP7_75t_L g1634 ( 
.A1(n_1621),
.A2(n_1568),
.B1(n_1566),
.B2(n_1560),
.C(n_1548),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1629),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1627),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_1632),
.Y(n_1637)
);

OAI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1624),
.A2(n_1618),
.B(n_1498),
.Y(n_1638)
);

OAI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1625),
.A2(n_1509),
.B1(n_1495),
.B2(n_1498),
.Y(n_1639)
);

INVxp67_ASAP7_75t_SL g1640 ( 
.A(n_1638),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1635),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1637),
.B(n_1626),
.Y(n_1642)
);

INVx1_ASAP7_75t_SL g1643 ( 
.A(n_1636),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1639),
.B(n_1628),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1637),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1641),
.Y(n_1646)
);

INVx1_ASAP7_75t_SL g1647 ( 
.A(n_1643),
.Y(n_1647)
);

OAI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1640),
.A2(n_1633),
.B(n_1634),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1645),
.Y(n_1649)
);

NOR2x1p5_ASAP7_75t_L g1650 ( 
.A(n_1642),
.B(n_1631),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1647),
.B(n_1644),
.Y(n_1651)
);

NOR3xp33_ASAP7_75t_L g1652 ( 
.A(n_1649),
.B(n_1630),
.C(n_1566),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1650),
.B(n_1529),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1653),
.B(n_1646),
.Y(n_1654)
);

OAI211xp5_ASAP7_75t_SL g1655 ( 
.A1(n_1654),
.A2(n_1651),
.B(n_1648),
.C(n_1652),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1655),
.B(n_1547),
.Y(n_1656)
);

AOI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1656),
.A2(n_1560),
.B(n_1547),
.Y(n_1657)
);

AOI22x1_ASAP7_75t_L g1658 ( 
.A1(n_1657),
.A2(n_1500),
.B1(n_1520),
.B2(n_1508),
.Y(n_1658)
);

XNOR2xp5_ASAP7_75t_L g1659 ( 
.A(n_1658),
.B(n_1365),
.Y(n_1659)
);

XOR2xp5_ASAP7_75t_L g1660 ( 
.A(n_1658),
.B(n_1363),
.Y(n_1660)
);

AOI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1659),
.A2(n_1510),
.B(n_1500),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1660),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1662),
.Y(n_1663)
);

NAND3xp33_ASAP7_75t_L g1664 ( 
.A(n_1661),
.B(n_1520),
.C(n_1508),
.Y(n_1664)
);

AOI21xp5_ASAP7_75t_SL g1665 ( 
.A1(n_1663),
.A2(n_1664),
.B(n_1509),
.Y(n_1665)
);

AOI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1665),
.A2(n_1508),
.B1(n_1510),
.B2(n_1532),
.Y(n_1666)
);

AOI211xp5_ASAP7_75t_L g1667 ( 
.A1(n_1666),
.A2(n_1510),
.B(n_1500),
.C(n_1532),
.Y(n_1667)
);


endmodule