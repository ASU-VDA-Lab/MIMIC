module fake_jpeg_9471_n_110 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_110);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_110;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_9),
.B(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_15),
.A2(n_23),
.B1(n_18),
.B2(n_14),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_25),
.A2(n_18),
.B1(n_16),
.B2(n_19),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_29),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_12),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_31),
.Y(n_35)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_19),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_31),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_41),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_20),
.B1(n_17),
.B2(n_13),
.Y(n_54)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_33),
.A2(n_25),
.B1(n_30),
.B2(n_13),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_44),
.A2(n_48),
.B1(n_55),
.B2(n_42),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_42),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_27),
.B1(n_16),
.B2(n_11),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_24),
.C(n_20),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_53),
.Y(n_56)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_50),
.B(n_51),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_21),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_54),
.A2(n_40),
.B1(n_42),
.B2(n_32),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_11),
.B1(n_17),
.B2(n_21),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_37),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_58),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_38),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_34),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_59),
.B(n_62),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_60),
.Y(n_72)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_61),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_47),
.B(n_10),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_22),
.B(n_2),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_65),
.B1(n_66),
.B2(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_47),
.B(n_8),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_67),
.B(n_1),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_SL g78 ( 
.A1(n_68),
.A2(n_73),
.B(n_63),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_56),
.A2(n_44),
.B1(n_55),
.B2(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_57),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_56),
.A2(n_54),
.B1(n_43),
.B2(n_52),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_58),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_75),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_76),
.B(n_64),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_78),
.A2(n_75),
.B1(n_74),
.B2(n_72),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_73),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_79),
.B(n_83),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_81),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_70),
.A2(n_22),
.B(n_21),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_86),
.Y(n_90)
);

BUFx24_ASAP7_75t_SL g83 ( 
.A(n_77),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_77),
.Y(n_84)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_45),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_52),
.B1(n_34),
.B2(n_24),
.Y(n_96)
);

MAJx2_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_69),
.C(n_32),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_92),
.A2(n_93),
.B(n_88),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_71),
.C(n_45),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_89),
.B(n_43),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_96),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_92),
.A2(n_52),
.B1(n_43),
.B2(n_61),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_97),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_90),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_87),
.C(n_3),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_97),
.A2(n_24),
.B1(n_3),
.B2(n_4),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_101),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_105),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_2),
.C(n_5),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_104),
.B(n_6),
.Y(n_107)
);

AO21x1_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_99),
.B(n_101),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_106),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_7),
.Y(n_110)
);


endmodule