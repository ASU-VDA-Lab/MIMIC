module fake_jpeg_22624_n_206 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_206);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_35),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_27),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_34),
.B(n_27),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_24),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVxp33_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_26),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_53),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_32),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_52),
.Y(n_63)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_23),
.B1(n_30),
.B2(n_24),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_54),
.A2(n_55),
.B1(n_56),
.B2(n_26),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_26),
.B1(n_25),
.B2(n_21),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_30),
.B1(n_26),
.B2(n_19),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_60),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_61),
.B(n_75),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_34),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_73),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_64),
.A2(n_17),
.B1(n_60),
.B2(n_42),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_41),
.B1(n_35),
.B2(n_22),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_66),
.A2(n_78),
.B1(n_48),
.B2(n_55),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_44),
.A2(n_15),
.B1(n_19),
.B2(n_40),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_69),
.B1(n_74),
.B2(n_43),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_53),
.A2(n_39),
.B1(n_20),
.B2(n_28),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_51),
.B(n_50),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_44),
.A2(n_15),
.B1(n_18),
.B2(n_22),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_29),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_79),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_43),
.A2(n_18),
.B1(n_28),
.B2(n_22),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_28),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_82),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_69),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_90),
.B1(n_99),
.B2(n_65),
.Y(n_105)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_84),
.B(n_86),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_63),
.A2(n_58),
.B(n_49),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_95),
.C(n_68),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_63),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_77),
.Y(n_89)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_62),
.A2(n_48),
.B1(n_18),
.B2(n_17),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_59),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_67),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_66),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_93),
.B(n_100),
.Y(n_109)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_0),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_71),
.B1(n_3),
.B2(n_4),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_64),
.A2(n_17),
.B1(n_42),
.B2(n_59),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_72),
.B(n_13),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_86),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_102),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_116),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_105),
.A2(n_108),
.B1(n_111),
.B2(n_118),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_72),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_95),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_99),
.A2(n_83),
.B1(n_92),
.B2(n_84),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_85),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_110),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_98),
.A2(n_74),
.B1(n_76),
.B2(n_73),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_87),
.B(n_68),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_112),
.B(n_87),
.Y(n_121)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_119),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_81),
.B(n_71),
.C(n_13),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_100),
.C(n_95),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_130),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_88),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_120),
.C(n_111),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_126),
.B(n_133),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_110),
.Y(n_127)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_132),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_113),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_102),
.B(n_91),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_109),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_137),
.Y(n_151)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_103),
.A2(n_89),
.B1(n_97),
.B2(n_94),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_138),
.A2(n_89),
.B1(n_114),
.B2(n_117),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_104),
.Y(n_140)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_129),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_141),
.Y(n_167)
);

AOI21x1_ASAP7_75t_SL g146 ( 
.A1(n_127),
.A2(n_103),
.B(n_116),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_146),
.A2(n_128),
.B1(n_136),
.B2(n_123),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_149),
.C(n_122),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_105),
.C(n_117),
.Y(n_149)
);

AOI21xp33_ASAP7_75t_L g150 ( 
.A1(n_125),
.A2(n_12),
.B(n_11),
.Y(n_150)
);

AOI321xp33_ASAP7_75t_L g158 ( 
.A1(n_150),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_154),
.Y(n_166)
);

AOI322xp5_ASAP7_75t_L g153 ( 
.A1(n_128),
.A2(n_114),
.A3(n_96),
.B1(n_101),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_153)
);

MAJx2_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_4),
.C(n_8),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_149),
.A2(n_137),
.B1(n_136),
.B2(n_131),
.Y(n_156)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_160),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_158),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_146),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_148),
.A2(n_122),
.B1(n_130),
.B2(n_101),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_139),
.B(n_126),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_163),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_147),
.C(n_145),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_164),
.A2(n_143),
.B1(n_154),
.B2(n_148),
.Y(n_170)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_165),
.A2(n_142),
.B(n_152),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_167),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_172),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_170),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_L g171 ( 
.A1(n_166),
.A2(n_141),
.B1(n_140),
.B2(n_143),
.Y(n_171)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_140),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_173),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_172),
.Y(n_184)
);

NOR2xp67_ASAP7_75t_SL g179 ( 
.A(n_174),
.B(n_162),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_179),
.A2(n_184),
.B(n_185),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_156),
.Y(n_181)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_181),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_159),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_177),
.C(n_160),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_171),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_188),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_180),
.A2(n_184),
.B(n_175),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_189),
.A2(n_164),
.B(n_158),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_180),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_190),
.A2(n_96),
.B1(n_9),
.B2(n_10),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_170),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_193),
.B(n_192),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_194),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_195),
.A2(n_191),
.B(n_9),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_196),
.A2(n_198),
.B1(n_197),
.B2(n_8),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_8),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_200),
.B(n_198),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_202),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_201),
.C(n_203),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_10),
.Y(n_206)
);


endmodule