module fake_jpeg_32078_n_151 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_151);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_151;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_33),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_27),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_13),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_38),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_40),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_13),
.B(n_0),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_15),
.B(n_5),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_22),
.B1(n_17),
.B2(n_20),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_43),
.A2(n_50),
.B1(n_51),
.B2(n_35),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_38),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_44),
.B(n_45),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_34),
.B(n_15),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_20),
.B1(n_14),
.B2(n_17),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_14),
.B1(n_26),
.B2(n_21),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_29),
.B(n_25),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_36),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_24),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_24),
.Y(n_66)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_53),
.A2(n_28),
.B1(n_26),
.B2(n_39),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_65),
.B1(n_35),
.B2(n_49),
.Y(n_82)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_30),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_0),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_46),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_68),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_70),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx24_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_18),
.Y(n_70)
);

INVxp67_ASAP7_75t_SL g71 ( 
.A(n_52),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_71),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_18),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_73),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_21),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_43),
.B(n_19),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_74),
.B(n_77),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_28),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_78),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_52),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_16),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_80),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_41),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_82),
.A2(n_86),
.B1(n_97),
.B2(n_67),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_68),
.A2(n_39),
.B1(n_47),
.B2(n_16),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_16),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_75),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_63),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_91),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_106),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_99),
.A2(n_74),
.B(n_80),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_101),
.A2(n_110),
.B(n_113),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_103),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_77),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_79),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_88),
.B(n_64),
.Y(n_109)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_90),
.A2(n_58),
.B(n_60),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_57),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_111),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_112),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_84),
.B(n_62),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_103),
.A2(n_82),
.B1(n_86),
.B2(n_89),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_101),
.B1(n_108),
.B2(n_111),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_124),
.A2(n_128),
.B1(n_114),
.B2(n_118),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_107),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_126),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_115),
.A2(n_108),
.B1(n_102),
.B2(n_106),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_127),
.A2(n_129),
.B(n_130),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_115),
.A2(n_110),
.B1(n_87),
.B2(n_83),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

INVxp67_ASAP7_75t_SL g130 ( 
.A(n_116),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_85),
.Y(n_131)
);

NOR3xp33_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_96),
.C(n_121),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_132),
.B(n_133),
.Y(n_140)
);

FAx1_ASAP7_75t_SL g134 ( 
.A(n_124),
.B(n_117),
.CI(n_118),
.CON(n_134),
.SN(n_134)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_134),
.B(n_135),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_117),
.C(n_114),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_135),
.A2(n_129),
.B1(n_127),
.B2(n_87),
.Y(n_138)
);

AOI322xp5_ASAP7_75t_L g144 ( 
.A1(n_138),
.A2(n_83),
.A3(n_93),
.B1(n_59),
.B2(n_2),
.C1(n_10),
.C2(n_11),
.Y(n_144)
);

NOR3xp33_ASAP7_75t_L g139 ( 
.A(n_136),
.B(n_93),
.C(n_5),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_139),
.B(n_12),
.Y(n_142)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_142),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_SL g143 ( 
.A1(n_140),
.A2(n_132),
.B(n_134),
.C(n_137),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_143),
.B(n_144),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_145),
.A2(n_141),
.B(n_138),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_147),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_146),
.A2(n_93),
.B(n_8),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_148),
.C(n_11),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_2),
.Y(n_151)
);


endmodule