module real_jpeg_30143_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_0),
.B(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_0),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_SL g82 ( 
.A1(n_0),
.A2(n_26),
.B(n_43),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_0),
.A2(n_71),
.B1(n_83),
.B2(n_105),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_0),
.A2(n_34),
.B(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_0),
.B(n_34),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_0),
.B(n_39),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_0),
.A2(n_74),
.B1(n_76),
.B2(n_146),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_0),
.A2(n_25),
.B(n_162),
.Y(n_161)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_2),
.A2(n_34),
.B1(n_35),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_2),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_64),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_2),
.A2(n_47),
.B1(n_52),
.B2(n_64),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_3),
.A2(n_47),
.B1(n_52),
.B2(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_3),
.Y(n_87)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_5),
.A2(n_34),
.B1(n_35),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_5),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_5),
.A2(n_47),
.B1(n_52),
.B2(n_66),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_7),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_8),
.A2(n_47),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_8),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g101 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_53),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_L g37 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_38),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_9),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_9),
.A2(n_38),
.B1(n_47),
.B2(n_52),
.Y(n_139)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_11),
.A2(n_27),
.B1(n_83),
.B2(n_105),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_11),
.A2(n_27),
.B1(n_34),
.B2(n_35),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_11),
.A2(n_27),
.B1(n_47),
.B2(n_52),
.Y(n_146)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_13),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g48 ( 
.A(n_14),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_15),
.A2(n_47),
.B1(n_52),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_15),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_112),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_110),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_78),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_19),
.B(n_78),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_56),
.C(n_67),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_20),
.A2(n_21),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_40),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_22),
.B(n_41),
.C(n_45),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_37),
.B2(n_39),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_24),
.A2(n_29),
.B1(n_33),
.B2(n_161),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_30),
.B(n_32),
.C(n_33),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_30),
.Y(n_32)
);

AO22x1_ASAP7_75t_L g42 ( 
.A1(n_25),
.A2(n_26),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

OAI32xp33_ASAP7_75t_L g69 ( 
.A1(n_25),
.A2(n_30),
.A3(n_35),
.B1(n_70),
.B2(n_72),
.Y(n_69)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_26),
.B(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_29),
.A2(n_33),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_34),
.A2(n_35),
.B1(n_59),
.B2(n_60),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_34),
.B(n_36),
.Y(n_72)
);

OAI32xp33_ASAP7_75t_L g123 ( 
.A1(n_34),
.A2(n_52),
.A3(n_59),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_37),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_45),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_42),
.A2(n_104),
.B1(n_107),
.B2(n_108),
.Y(n_103)
);

O2A1O1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_42),
.A2(n_43),
.B(n_105),
.C(n_106),
.Y(n_104)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

NAND2xp33_ASAP7_75t_SL g106 ( 
.A(n_43),
.B(n_105),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_44),
.A2(n_71),
.B(n_82),
.C(n_83),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_49),
.B1(n_51),
.B2(n_54),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_46),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_46),
.A2(n_49),
.B1(n_54),
.B2(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_46),
.A2(n_138),
.B1(n_140),
.B2(n_141),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_49),
.Y(n_46)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_52),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_47),
.B(n_60),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_47),
.B(n_152),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx5_ASAP7_75t_SL g147 ( 
.A(n_49),
.Y(n_147)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_51),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_56),
.A2(n_67),
.B1(n_68),
.B2(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_56),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_62),
.B2(n_65),
.Y(n_56)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_57),
.A2(n_58),
.B1(n_119),
.B2(n_121),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_57),
.A2(n_58),
.B1(n_121),
.B2(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_58),
.B(n_71),
.Y(n_148)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_63),
.A2(n_100),
.B1(n_102),
.B2(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_65),
.Y(n_99)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_73),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_69),
.B(n_73),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_70),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_71),
.B(n_76),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_74),
.A2(n_139),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_91),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_80),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_85),
.Y(n_80)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_103),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_97),
.B2(n_98),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_171),
.B(n_177),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_156),
.B(n_170),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_135),
.B(n_155),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_126),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_116),
.B(n_126),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_122),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_117),
.A2(n_118),
.B1(n_122),
.B2(n_123),
.Y(n_142)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_120),
.Y(n_124)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_133),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_131),
.C(n_133),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_132),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_134),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_143),
.B(n_154),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_142),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_137),
.B(n_142),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_149),
.B(n_153),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_148),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_145),
.B(n_148),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_157),
.B(n_158),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_158)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_159),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_163),
.B1(n_165),
.B2(n_166),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_160),
.Y(n_166)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_163),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_166),
.C(n_169),
.Y(n_172)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_167),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_172),
.B(n_173),
.Y(n_177)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);


endmodule