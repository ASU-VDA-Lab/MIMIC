module fake_ariane_3350_n_160 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_17, n_4, n_2, n_18, n_28, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_160);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_17;
input n_4;
input n_2;
input n_18;
input n_28;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_160;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_124;
wire n_119;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_149;
wire n_34;
wire n_158;
wire n_69;
wire n_95;
wire n_92;
wire n_143;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_152;
wire n_120;
wire n_106;
wire n_53;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_100;
wire n_50;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_30;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_85;
wire n_130;
wire n_144;
wire n_48;
wire n_101;
wire n_94;
wire n_134;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_52;
wire n_157;
wire n_135;
wire n_73;
wire n_77;
wire n_118;
wire n_93;
wire n_121;
wire n_61;
wire n_108;
wire n_102;
wire n_125;
wire n_43;
wire n_81;
wire n_87;
wire n_29;
wire n_41;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_88;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_39;
wire n_63;
wire n_59;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_25),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVxp33_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_22),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_3),
.B(n_10),
.Y(n_38)
);

CKINVDCx5p33_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_11),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVxp67_ASAP7_75t_SL g48 ( 
.A(n_17),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_0),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_41),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_30),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_5),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_35),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NAND2xp33_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_6),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_31),
.B(n_8),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_50),
.B(n_12),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_16),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_42),
.B(n_23),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_70),
.B(n_52),
.Y(n_72)
);

NAND2xp33_ASAP7_75t_SL g73 ( 
.A(n_71),
.B(n_45),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_69),
.B(n_45),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_69),
.B(n_68),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_69),
.B(n_30),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_68),
.B(n_34),
.Y(n_77)
);

NAND2xp33_ASAP7_75t_SL g78 ( 
.A(n_56),
.B(n_34),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_68),
.B(n_33),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_58),
.B(n_42),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_62),
.B(n_66),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_61),
.B(n_24),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_61),
.B(n_64),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_64),
.B(n_26),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_60),
.B(n_27),
.Y(n_85)
);

NAND2xp33_ASAP7_75t_SL g86 ( 
.A(n_56),
.B(n_55),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_54),
.B(n_63),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_54),
.B(n_63),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_57),
.B(n_53),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_59),
.Y(n_90)
);

OAI21x1_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_65),
.B(n_53),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_89),
.B(n_53),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

BUFx10_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

BUFx8_ASAP7_75t_SL g95 ( 
.A(n_78),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

AOI221x1_ASAP7_75t_SL g97 ( 
.A1(n_86),
.A2(n_72),
.B1(n_60),
.B2(n_67),
.C(n_73),
.Y(n_97)
);

OAI22x1_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_59),
.B1(n_67),
.B2(n_74),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_85),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_59),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_59),
.B1(n_67),
.B2(n_87),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_81),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

OAI21x1_ASAP7_75t_L g106 ( 
.A1(n_81),
.A2(n_75),
.B(n_66),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_95),
.Y(n_107)
);

AND2x4_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_96),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

AND2x4_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_93),
.Y(n_110)
);

AND2x4_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_101),
.Y(n_111)
);

OR2x6_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_98),
.Y(n_112)
);

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_98),
.Y(n_113)
);

NAND2xp33_ASAP7_75t_R g114 ( 
.A(n_104),
.B(n_90),
.Y(n_114)
);

NAND2xp33_ASAP7_75t_R g115 ( 
.A(n_104),
.B(n_90),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_94),
.Y(n_116)
);

AND2x4_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_105),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_R g120 ( 
.A(n_94),
.B(n_102),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

OR2x6_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_91),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

NOR3xp33_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_106),
.C(n_102),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

AO21x2_ASAP7_75t_L g127 ( 
.A1(n_124),
.A2(n_97),
.B(n_94),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_118),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g129 ( 
.A(n_116),
.B(n_97),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_103),
.Y(n_130)
);

OAI222xp33_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_103),
.B1(n_113),
.B2(n_111),
.C1(n_108),
.C2(n_117),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_111),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_112),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_121),
.Y(n_136)
);

NAND3xp33_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_115),
.C(n_122),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

NOR2x1_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_122),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_129),
.A2(n_114),
.B1(n_115),
.B2(n_133),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_120),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

AO221x2_ASAP7_75t_L g143 ( 
.A1(n_131),
.A2(n_119),
.B1(n_123),
.B2(n_129),
.C(n_130),
.Y(n_143)
);

NOR2x1_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_119),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_135),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_142),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_L g148 ( 
.A1(n_140),
.A2(n_134),
.B1(n_135),
.B2(n_132),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_147),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_147),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_148),
.Y(n_151)
);

NAND3xp33_ASAP7_75t_L g152 ( 
.A(n_150),
.B(n_125),
.C(n_146),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_149),
.Y(n_153)
);

NAND2xp33_ASAP7_75t_SL g154 ( 
.A(n_153),
.B(n_141),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_R g155 ( 
.A(n_152),
.B(n_151),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_154),
.A2(n_143),
.B1(n_151),
.B2(n_139),
.Y(n_156)
);

OAI21x1_ASAP7_75t_L g157 ( 
.A1(n_155),
.A2(n_138),
.B(n_137),
.Y(n_157)
);

AOI31xp33_ASAP7_75t_L g158 ( 
.A1(n_156),
.A2(n_137),
.A3(n_144),
.B(n_138),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_157),
.B1(n_134),
.B2(n_136),
.Y(n_159)
);

AOI221xp5_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_127),
.B1(n_136),
.B2(n_128),
.C(n_132),
.Y(n_160)
);


endmodule