module fake_netlist_6_4466_n_1097 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_256, n_18, n_21, n_193, n_147, n_258, n_154, n_191, n_88, n_3, n_209, n_98, n_260, n_265, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_252, n_266, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_247, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_245, n_0, n_87, n_195, n_261, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_257, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_254, n_142, n_20, n_143, n_207, n_2, n_242, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_263, n_122, n_264, n_45, n_255, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_251, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_246, n_38, n_110, n_151, n_61, n_112, n_172, n_237, n_81, n_59, n_244, n_181, n_76, n_36, n_182, n_26, n_124, n_238, n_239, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_240, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_259, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_243, n_9, n_248, n_107, n_10, n_71, n_74, n_229, n_253, n_6, n_190, n_14, n_123, n_262, n_136, n_72, n_187, n_89, n_249, n_173, n_201, n_250, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_241, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_1097);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_256;
input n_18;
input n_21;
input n_193;
input n_147;
input n_258;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_260;
input n_265;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_252;
input n_266;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_247;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_245;
input n_0;
input n_87;
input n_195;
input n_261;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_257;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_254;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_242;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_263;
input n_122;
input n_264;
input n_45;
input n_255;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_251;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_246;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_244;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_238;
input n_239;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_240;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_259;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_243;
input n_9;
input n_248;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_253;
input n_6;
input n_190;
input n_14;
input n_123;
input n_262;
input n_136;
input n_72;
input n_187;
input n_89;
input n_249;
input n_173;
input n_201;
input n_250;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_241;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1097;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_278;
wire n_1079;
wire n_341;
wire n_362;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_988;
wire n_969;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_898;
wire n_617;
wire n_698;
wire n_1074;
wire n_1032;
wire n_845;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1095;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_1057;
wire n_360;
wire n_977;
wire n_945;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1017;
wire n_1004;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_638;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_653;
wire n_887;
wire n_1087;
wire n_908;
wire n_752;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_1043;
wire n_1011;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_1084;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_870;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_1085;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_757;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_1078;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_543;
wire n_889;
wire n_357;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_584;
wire n_399;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_322;
wire n_707;
wire n_993;
wire n_345;
wire n_409;
wire n_689;
wire n_354;
wire n_799;
wire n_505;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_1092;
wire n_441;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_582;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_518;
wire n_299;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_834;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_401;
wire n_324;
wire n_743;
wire n_816;
wire n_766;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_228),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_189),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_94),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_112),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_6),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_185),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_226),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_21),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_150),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_248),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_133),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_18),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_214),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_11),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_79),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_264),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_159),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_83),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_181),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_241),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_148),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_216),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_165),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_160),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_128),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_186),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_108),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_12),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_145),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_184),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_170),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_15),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_180),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_78),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_253),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_105),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_53),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_249),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_175),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_256),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_35),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_121),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_209),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_106),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_201),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_125),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_153),
.Y(n_313)
);

INVx2_ASAP7_75t_SL g314 ( 
.A(n_87),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_42),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_88),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_254),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_237),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_203),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_250),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_163),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_174),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_122),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_119),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_16),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_130),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_84),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_57),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_103),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_23),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_314),
.B(n_297),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_267),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_280),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_268),
.Y(n_334)
);

NOR2xp67_ASAP7_75t_L g335 ( 
.A(n_294),
.B(n_0),
.Y(n_335)
);

NOR2xp67_ASAP7_75t_L g336 ( 
.A(n_309),
.B(n_0),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_286),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_286),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_271),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_269),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_310),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_310),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_276),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_274),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_272),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_282),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_284),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_288),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_277),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_279),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_281),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_273),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_283),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_287),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_289),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_291),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_292),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_295),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_278),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_298),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_296),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_325),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_309),
.B(n_1),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_315),
.B(n_1),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_330),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_285),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_290),
.Y(n_367)
);

INVxp33_ASAP7_75t_SL g368 ( 
.A(n_299),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_275),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_316),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_303),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_301),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_302),
.Y(n_373)
);

NOR2xp67_ASAP7_75t_L g374 ( 
.A(n_319),
.B(n_2),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_352),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_343),
.Y(n_376)
);

INVxp33_ASAP7_75t_SL g377 ( 
.A(n_332),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_369),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_346),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_347),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_352),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_354),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_355),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_356),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_344),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_365),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_357),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_358),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_361),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_370),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_333),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_337),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_338),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_342),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_341),
.B(n_328),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_364),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_334),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_331),
.B(n_270),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_363),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_339),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_348),
.B(n_323),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_374),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_340),
.B(n_304),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_345),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_349),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_336),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_335),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_350),
.B(n_273),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_351),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_353),
.B(n_329),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_366),
.B(n_305),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_367),
.B(n_273),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_372),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_373),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_365),
.Y(n_415)
);

OA21x2_ASAP7_75t_L g416 ( 
.A1(n_368),
.A2(n_308),
.B(n_306),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_368),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_359),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_359),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_360),
.A2(n_307),
.B1(n_312),
.B2(n_311),
.Y(n_420)
);

NAND2xp33_ASAP7_75t_L g421 ( 
.A(n_360),
.B(n_273),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_362),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_362),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_399),
.B(n_313),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_390),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_390),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_395),
.B(n_317),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_390),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_397),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_381),
.Y(n_430)
);

INVx4_ASAP7_75t_L g431 ( 
.A(n_408),
.Y(n_431)
);

INVxp33_ASAP7_75t_L g432 ( 
.A(n_419),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_395),
.B(n_318),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_400),
.B(n_398),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_381),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_376),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_381),
.Y(n_437)
);

INVx5_ASAP7_75t_L g438 ( 
.A(n_399),
.Y(n_438)
);

NAND2x1p5_ASAP7_75t_L g439 ( 
.A(n_397),
.B(n_293),
.Y(n_439)
);

NAND2xp33_ASAP7_75t_L g440 ( 
.A(n_399),
.B(n_293),
.Y(n_440)
);

INVx5_ASAP7_75t_L g441 ( 
.A(n_399),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_378),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_381),
.Y(n_443)
);

INVx4_ASAP7_75t_L g444 ( 
.A(n_408),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_399),
.B(n_320),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_381),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_379),
.Y(n_447)
);

NAND2xp33_ASAP7_75t_L g448 ( 
.A(n_396),
.B(n_293),
.Y(n_448)
);

AND2x2_ASAP7_75t_SL g449 ( 
.A(n_401),
.B(n_293),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_392),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_380),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_414),
.Y(n_452)
);

OR2x6_ASAP7_75t_L g453 ( 
.A(n_419),
.B(n_300),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_414),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_392),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g456 ( 
.A(n_395),
.B(n_321),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_382),
.Y(n_457)
);

BUFx10_ASAP7_75t_L g458 ( 
.A(n_405),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_382),
.Y(n_459)
);

AND2x4_ASAP7_75t_L g460 ( 
.A(n_408),
.B(n_322),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_383),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_383),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_384),
.Y(n_463)
);

AO21x2_ASAP7_75t_L g464 ( 
.A1(n_403),
.A2(n_326),
.B(n_324),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_375),
.Y(n_465)
);

INVx4_ASAP7_75t_L g466 ( 
.A(n_412),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_387),
.Y(n_467)
);

INVx6_ASAP7_75t_L g468 ( 
.A(n_412),
.Y(n_468)
);

BUFx4f_ASAP7_75t_L g469 ( 
.A(n_416),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_375),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_404),
.B(n_369),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_400),
.B(n_327),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_412),
.B(n_300),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_388),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_398),
.B(n_300),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_391),
.Y(n_476)
);

AND2x6_ASAP7_75t_L g477 ( 
.A(n_404),
.B(n_300),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_413),
.B(n_371),
.Y(n_478)
);

AND2x6_ASAP7_75t_L g479 ( 
.A(n_413),
.B(n_402),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_389),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_391),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_393),
.B(n_36),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_394),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_416),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_407),
.Y(n_485)
);

BUFx4f_ASAP7_75t_L g486 ( 
.A(n_416),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_385),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_410),
.B(n_371),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_406),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_434),
.B(n_417),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_474),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_474),
.Y(n_492)
);

AO22x2_ASAP7_75t_L g493 ( 
.A1(n_485),
.A2(n_423),
.B1(n_418),
.B2(n_422),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_425),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_487),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_480),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g497 ( 
.A(n_453),
.Y(n_497)
);

AO22x2_ASAP7_75t_L g498 ( 
.A1(n_485),
.A2(n_423),
.B1(n_418),
.B2(n_415),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_480),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_468),
.A2(n_421),
.B1(n_386),
.B2(n_377),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_438),
.B(n_411),
.Y(n_501)
);

OAI22xp33_ASAP7_75t_L g502 ( 
.A1(n_475),
.A2(n_420),
.B1(n_405),
.B2(n_409),
.Y(n_502)
);

BUFx8_ASAP7_75t_L g503 ( 
.A(n_442),
.Y(n_503)
);

CKINVDCx16_ASAP7_75t_R g504 ( 
.A(n_458),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_483),
.Y(n_505)
);

BUFx8_ASAP7_75t_L g506 ( 
.A(n_429),
.Y(n_506)
);

AO22x2_ASAP7_75t_L g507 ( 
.A1(n_449),
.A2(n_421),
.B1(n_4),
.B2(n_2),
.Y(n_507)
);

OR2x2_ASAP7_75t_SL g508 ( 
.A(n_489),
.B(n_419),
.Y(n_508)
);

AO22x2_ASAP7_75t_L g509 ( 
.A1(n_452),
.A2(n_454),
.B1(n_433),
.B2(n_427),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_483),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_453),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_425),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_468),
.A2(n_377),
.B1(n_409),
.B2(n_419),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_450),
.Y(n_514)
);

INVx1_ASAP7_75t_SL g515 ( 
.A(n_458),
.Y(n_515)
);

OR2x6_ASAP7_75t_L g516 ( 
.A(n_439),
.B(n_419),
.Y(n_516)
);

AO21x1_ASAP7_75t_L g517 ( 
.A1(n_440),
.A2(n_445),
.B(n_424),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_436),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_427),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_432),
.B(n_378),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_447),
.Y(n_521)
);

AO22x2_ASAP7_75t_L g522 ( 
.A1(n_433),
.A2(n_456),
.B1(n_473),
.B2(n_460),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_451),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_455),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_476),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_489),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_426),
.Y(n_527)
);

AO22x2_ASAP7_75t_L g528 ( 
.A1(n_456),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_481),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_426),
.Y(n_530)
);

NAND2x1p5_ASAP7_75t_L g531 ( 
.A(n_431),
.B(n_37),
.Y(n_531)
);

AO22x2_ASAP7_75t_L g532 ( 
.A1(n_473),
.A2(n_460),
.B1(n_472),
.B2(n_428),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_471),
.B(n_3),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_428),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_438),
.B(n_38),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_465),
.Y(n_536)
);

INVxp67_ASAP7_75t_SL g537 ( 
.A(n_430),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_489),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_457),
.Y(n_539)
);

AO22x2_ASAP7_75t_L g540 ( 
.A1(n_431),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_540)
);

OAI221xp5_ASAP7_75t_L g541 ( 
.A1(n_457),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_541)
);

AO22x2_ASAP7_75t_L g542 ( 
.A1(n_444),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_542)
);

OAI221xp5_ASAP7_75t_L g543 ( 
.A1(n_461),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.C(n_14),
.Y(n_543)
);

AO22x2_ASAP7_75t_L g544 ( 
.A1(n_444),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_544)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_478),
.Y(n_545)
);

OAI221xp5_ASAP7_75t_L g546 ( 
.A1(n_461),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.C(n_19),
.Y(n_546)
);

AO22x2_ASAP7_75t_L g547 ( 
.A1(n_466),
.A2(n_20),
.B1(n_17),
.B2(n_19),
.Y(n_547)
);

NAND2x1p5_ASAP7_75t_L g548 ( 
.A(n_466),
.B(n_39),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_438),
.B(n_40),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_470),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_488),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_479),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_482),
.Y(n_553)
);

AO22x2_ASAP7_75t_L g554 ( 
.A1(n_482),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_463),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_462),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_462),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_441),
.B(n_41),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_441),
.B(n_43),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_459),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_459),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_463),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_555),
.B(n_545),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_555),
.B(n_441),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_555),
.B(n_463),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_490),
.B(n_467),
.Y(n_566)
);

AND2x4_ASAP7_75t_SL g567 ( 
.A(n_519),
.B(n_467),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_513),
.B(n_467),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_500),
.B(n_459),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_553),
.B(n_479),
.Y(n_570)
);

NAND2xp33_ASAP7_75t_SL g571 ( 
.A(n_533),
.B(n_464),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_502),
.B(n_469),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_551),
.B(n_469),
.Y(n_573)
);

NAND2xp33_ASAP7_75t_SL g574 ( 
.A(n_497),
.B(n_464),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_538),
.B(n_486),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_495),
.B(n_484),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_526),
.B(n_486),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_491),
.B(n_484),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_492),
.B(n_496),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_499),
.B(n_484),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_505),
.B(n_430),
.Y(n_581)
);

NAND2xp33_ASAP7_75t_SL g582 ( 
.A(n_511),
.B(n_437),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_510),
.B(n_562),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_518),
.B(n_430),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_521),
.B(n_435),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_539),
.B(n_479),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_520),
.B(n_479),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_523),
.B(n_536),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_516),
.B(n_443),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_550),
.B(n_435),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_514),
.B(n_524),
.Y(n_591)
);

NAND2xp33_ASAP7_75t_SL g592 ( 
.A(n_501),
.B(n_435),
.Y(n_592)
);

NAND2xp33_ASAP7_75t_SL g593 ( 
.A(n_508),
.B(n_446),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_556),
.B(n_446),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_525),
.B(n_529),
.Y(n_595)
);

NAND2xp33_ASAP7_75t_SL g596 ( 
.A(n_494),
.B(n_448),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_557),
.B(n_504),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_515),
.B(n_477),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_516),
.B(n_44),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_560),
.B(n_477),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_561),
.B(n_477),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_517),
.B(n_477),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_494),
.B(n_45),
.Y(n_603)
);

AND2x2_ASAP7_75t_SL g604 ( 
.A(n_507),
.B(n_46),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_512),
.B(n_47),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_512),
.B(n_48),
.Y(n_606)
);

NAND2xp33_ASAP7_75t_SL g607 ( 
.A(n_527),
.B(n_530),
.Y(n_607)
);

NAND2xp33_ASAP7_75t_SL g608 ( 
.A(n_534),
.B(n_24),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_532),
.B(n_25),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_531),
.B(n_49),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_532),
.B(n_25),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_SL g612 ( 
.A(n_535),
.B(n_26),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_548),
.B(n_50),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_552),
.B(n_506),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_506),
.B(n_51),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_537),
.B(n_26),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_549),
.B(n_52),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_558),
.B(n_54),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_559),
.B(n_55),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_SL g620 ( 
.A(n_522),
.B(n_27),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_503),
.B(n_56),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_522),
.B(n_27),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_503),
.B(n_58),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_509),
.B(n_59),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_509),
.B(n_60),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_507),
.B(n_61),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_498),
.B(n_28),
.Y(n_627)
);

AND2x2_ASAP7_75t_SL g628 ( 
.A(n_554),
.B(n_62),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_SL g629 ( 
.A(n_628),
.B(n_541),
.Y(n_629)
);

NOR2xp67_ASAP7_75t_L g630 ( 
.A(n_597),
.B(n_543),
.Y(n_630)
);

AO31x2_ASAP7_75t_L g631 ( 
.A1(n_609),
.A2(n_498),
.A3(n_493),
.B(n_542),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_566),
.B(n_493),
.Y(n_632)
);

OAI21x1_ASAP7_75t_L g633 ( 
.A1(n_586),
.A2(n_64),
.B(n_63),
.Y(n_633)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_576),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_567),
.B(n_528),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_579),
.B(n_554),
.Y(n_636)
);

OAI21xp5_ASAP7_75t_SL g637 ( 
.A1(n_614),
.A2(n_546),
.B(n_528),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_589),
.Y(n_638)
);

OAI21x1_ASAP7_75t_SL g639 ( 
.A1(n_611),
.A2(n_542),
.B(n_540),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_577),
.A2(n_547),
.B(n_544),
.Y(n_640)
);

NAND3x1_ASAP7_75t_L g641 ( 
.A(n_622),
.B(n_544),
.C(n_540),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_594),
.Y(n_642)
);

OAI21x1_ASAP7_75t_L g643 ( 
.A1(n_575),
.A2(n_66),
.B(n_65),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_568),
.A2(n_547),
.B(n_68),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_589),
.Y(n_645)
);

OA21x2_ASAP7_75t_L g646 ( 
.A1(n_602),
.A2(n_69),
.B(n_67),
.Y(n_646)
);

OAI22x1_ASAP7_75t_L g647 ( 
.A1(n_626),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_647)
);

INVx2_ASAP7_75t_SL g648 ( 
.A(n_563),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_574),
.Y(n_649)
);

OAI22xp5_ASAP7_75t_L g650 ( 
.A1(n_572),
.A2(n_172),
.B1(n_265),
.B2(n_263),
.Y(n_650)
);

BUFx5_ASAP7_75t_L g651 ( 
.A(n_587),
.Y(n_651)
);

AO21x2_ASAP7_75t_L g652 ( 
.A1(n_569),
.A2(n_71),
.B(n_70),
.Y(n_652)
);

INVx1_ASAP7_75t_SL g653 ( 
.A(n_627),
.Y(n_653)
);

OAI21x1_ASAP7_75t_L g654 ( 
.A1(n_578),
.A2(n_73),
.B(n_72),
.Y(n_654)
);

OAI21x1_ASAP7_75t_L g655 ( 
.A1(n_580),
.A2(n_75),
.B(n_74),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_588),
.B(n_573),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_628),
.B(n_29),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_L g658 ( 
.A1(n_604),
.A2(n_570),
.B1(n_583),
.B2(n_599),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_571),
.A2(n_177),
.B1(n_262),
.B2(n_261),
.Y(n_659)
);

OAI21x1_ASAP7_75t_L g660 ( 
.A1(n_565),
.A2(n_77),
.B(n_76),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_591),
.Y(n_661)
);

AOI21x1_ASAP7_75t_SL g662 ( 
.A1(n_616),
.A2(n_30),
.B(n_31),
.Y(n_662)
);

BUFx2_ASAP7_75t_L g663 ( 
.A(n_599),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_595),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_590),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_604),
.B(n_31),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_607),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_624),
.B(n_32),
.Y(n_668)
);

INVxp67_ASAP7_75t_SL g669 ( 
.A(n_564),
.Y(n_669)
);

AOI21x1_ASAP7_75t_SL g670 ( 
.A1(n_620),
.A2(n_32),
.B(n_33),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_581),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_R g672 ( 
.A(n_593),
.B(n_80),
.Y(n_672)
);

INVx5_ASAP7_75t_L g673 ( 
.A(n_608),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_621),
.B(n_33),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_592),
.A2(n_596),
.B(n_610),
.Y(n_675)
);

OAI21x1_ASAP7_75t_SL g676 ( 
.A1(n_625),
.A2(n_82),
.B(n_81),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_584),
.B(n_34),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_585),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_613),
.A2(n_86),
.B(n_85),
.Y(n_679)
);

NAND2xp33_ASAP7_75t_R g680 ( 
.A(n_582),
.B(n_89),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_612),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_623),
.B(n_34),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_603),
.Y(n_683)
);

NAND3x1_ASAP7_75t_L g684 ( 
.A(n_615),
.B(n_90),
.C(n_91),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_598),
.B(n_92),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_605),
.B(n_93),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_606),
.B(n_95),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_617),
.B(n_618),
.Y(n_688)
);

INVx5_ASAP7_75t_L g689 ( 
.A(n_619),
.Y(n_689)
);

OAI21x1_ASAP7_75t_L g690 ( 
.A1(n_600),
.A2(n_96),
.B(n_97),
.Y(n_690)
);

INVx1_ASAP7_75t_SL g691 ( 
.A(n_634),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_661),
.Y(n_692)
);

OR2x2_ASAP7_75t_L g693 ( 
.A(n_653),
.B(n_601),
.Y(n_693)
);

A2O1A1Ixp33_ASAP7_75t_L g694 ( 
.A1(n_629),
.A2(n_98),
.B(n_99),
.C(n_100),
.Y(n_694)
);

BUFx2_ASAP7_75t_SL g695 ( 
.A(n_638),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_642),
.B(n_651),
.Y(n_696)
);

AO21x2_ASAP7_75t_L g697 ( 
.A1(n_675),
.A2(n_101),
.B(n_102),
.Y(n_697)
);

OAI21x1_ASAP7_75t_L g698 ( 
.A1(n_654),
.A2(n_104),
.B(n_107),
.Y(n_698)
);

AOI22x1_ASAP7_75t_L g699 ( 
.A1(n_667),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_699)
);

CKINVDCx11_ASAP7_75t_R g700 ( 
.A(n_649),
.Y(n_700)
);

OAI21x1_ASAP7_75t_L g701 ( 
.A1(n_655),
.A2(n_113),
.B(n_114),
.Y(n_701)
);

OAI21x1_ASAP7_75t_L g702 ( 
.A1(n_643),
.A2(n_115),
.B(n_116),
.Y(n_702)
);

AOI221xp5_ASAP7_75t_L g703 ( 
.A1(n_666),
.A2(n_117),
.B1(n_118),
.B2(n_120),
.C(n_123),
.Y(n_703)
);

NOR2xp67_ASAP7_75t_L g704 ( 
.A(n_689),
.B(n_124),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_661),
.Y(n_705)
);

OAI21x1_ASAP7_75t_L g706 ( 
.A1(n_633),
.A2(n_126),
.B(n_127),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_664),
.Y(n_707)
);

AO31x2_ASAP7_75t_L g708 ( 
.A1(n_667),
.A2(n_129),
.A3(n_131),
.B(n_132),
.Y(n_708)
);

O2A1O1Ixp5_ASAP7_75t_L g709 ( 
.A1(n_644),
.A2(n_658),
.B(n_681),
.C(n_688),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_632),
.Y(n_710)
);

AO21x2_ASAP7_75t_L g711 ( 
.A1(n_640),
.A2(n_134),
.B(n_135),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_665),
.Y(n_712)
);

OAI21x1_ASAP7_75t_L g713 ( 
.A1(n_660),
.A2(n_136),
.B(n_137),
.Y(n_713)
);

OA21x2_ASAP7_75t_L g714 ( 
.A1(n_683),
.A2(n_138),
.B(n_139),
.Y(n_714)
);

AOI21x1_ASAP7_75t_L g715 ( 
.A1(n_656),
.A2(n_683),
.B(n_642),
.Y(n_715)
);

OAI21x1_ASAP7_75t_SL g716 ( 
.A1(n_676),
.A2(n_140),
.B(n_141),
.Y(n_716)
);

OAI21xp5_ASAP7_75t_L g717 ( 
.A1(n_630),
.A2(n_266),
.B(n_143),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_638),
.Y(n_718)
);

AO31x2_ASAP7_75t_L g719 ( 
.A1(n_647),
.A2(n_650),
.A3(n_668),
.B(n_687),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_671),
.Y(n_720)
);

INVx4_ASAP7_75t_L g721 ( 
.A(n_645),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_663),
.B(n_142),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_645),
.Y(n_723)
);

INVx1_ASAP7_75t_SL g724 ( 
.A(n_636),
.Y(n_724)
);

AND2x4_ASAP7_75t_L g725 ( 
.A(n_648),
.B(n_144),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_669),
.Y(n_726)
);

BUFx8_ASAP7_75t_L g727 ( 
.A(n_674),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_651),
.B(n_673),
.Y(n_728)
);

OA21x2_ASAP7_75t_L g729 ( 
.A1(n_690),
.A2(n_685),
.B(n_659),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_678),
.Y(n_730)
);

BUFx12f_ASAP7_75t_L g731 ( 
.A(n_682),
.Y(n_731)
);

AND2x4_ASAP7_75t_L g732 ( 
.A(n_673),
.B(n_260),
.Y(n_732)
);

OAI21x1_ASAP7_75t_L g733 ( 
.A1(n_646),
.A2(n_679),
.B(n_670),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_SL g734 ( 
.A1(n_657),
.A2(n_146),
.B1(n_147),
.B2(n_149),
.Y(n_734)
);

OAI22xp33_ASAP7_75t_L g735 ( 
.A1(n_637),
.A2(n_673),
.B1(n_680),
.B2(n_677),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_641),
.A2(n_151),
.B1(n_152),
.B2(n_154),
.Y(n_736)
);

OAI21xp5_ASAP7_75t_L g737 ( 
.A1(n_686),
.A2(n_155),
.B(n_156),
.Y(n_737)
);

OAI21x1_ASAP7_75t_L g738 ( 
.A1(n_646),
.A2(n_157),
.B(n_158),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_631),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_635),
.B(n_161),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_678),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_SL g742 ( 
.A(n_639),
.B(n_162),
.Y(n_742)
);

OR2x6_ASAP7_75t_L g743 ( 
.A(n_678),
.B(n_164),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_651),
.Y(n_744)
);

A2O1A1Ixp33_ASAP7_75t_L g745 ( 
.A1(n_689),
.A2(n_166),
.B(n_167),
.C(n_168),
.Y(n_745)
);

NAND2x1p5_ASAP7_75t_L g746 ( 
.A(n_689),
.B(n_169),
.Y(n_746)
);

INVxp67_ASAP7_75t_SL g747 ( 
.A(n_696),
.Y(n_747)
);

BUFx3_ASAP7_75t_L g748 ( 
.A(n_741),
.Y(n_748)
);

INVx4_ASAP7_75t_L g749 ( 
.A(n_744),
.Y(n_749)
);

HB1xp67_ASAP7_75t_L g750 ( 
.A(n_691),
.Y(n_750)
);

OAI22xp33_ASAP7_75t_L g751 ( 
.A1(n_736),
.A2(n_684),
.B1(n_672),
.B2(n_662),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_698),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_710),
.B(n_631),
.Y(n_753)
);

INVxp67_ASAP7_75t_L g754 ( 
.A(n_691),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_739),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_715),
.Y(n_756)
);

AOI21x1_ASAP7_75t_L g757 ( 
.A1(n_733),
.A2(n_652),
.B(n_651),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_696),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_692),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_705),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_720),
.Y(n_761)
);

OAI21x1_ASAP7_75t_L g762 ( 
.A1(n_706),
.A2(n_652),
.B(n_651),
.Y(n_762)
);

INVx3_ASAP7_75t_L g763 ( 
.A(n_701),
.Y(n_763)
);

NAND2xp33_ASAP7_75t_L g764 ( 
.A(n_728),
.B(n_631),
.Y(n_764)
);

AO21x2_ASAP7_75t_L g765 ( 
.A1(n_717),
.A2(n_171),
.B(n_173),
.Y(n_765)
);

NOR2x1_ASAP7_75t_R g766 ( 
.A(n_700),
.B(n_176),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_730),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_714),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_724),
.B(n_178),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_707),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_714),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_724),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_712),
.B(n_259),
.Y(n_773)
);

INVx1_ASAP7_75t_SL g774 ( 
.A(n_731),
.Y(n_774)
);

INVx1_ASAP7_75t_SL g775 ( 
.A(n_693),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_738),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_713),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_736),
.B(n_179),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_711),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_709),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_737),
.B(n_258),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_728),
.B(n_182),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_711),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_708),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_697),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_737),
.B(n_257),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_735),
.B(n_183),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_708),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_697),
.Y(n_789)
);

INVx3_ASAP7_75t_L g790 ( 
.A(n_702),
.Y(n_790)
);

INVx3_ASAP7_75t_L g791 ( 
.A(n_729),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_726),
.B(n_725),
.Y(n_792)
);

NAND2xp33_ASAP7_75t_R g793 ( 
.A(n_732),
.B(n_187),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_708),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_699),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_729),
.Y(n_796)
);

OAI21x1_ASAP7_75t_L g797 ( 
.A1(n_716),
.A2(n_188),
.B(n_190),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_719),
.Y(n_798)
);

O2A1O1Ixp33_ASAP7_75t_SL g799 ( 
.A1(n_694),
.A2(n_745),
.B(n_717),
.C(n_703),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_719),
.Y(n_800)
);

HB1xp67_ASAP7_75t_L g801 ( 
.A(n_730),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_742),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_719),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_718),
.Y(n_804)
);

OAI21x1_ASAP7_75t_L g805 ( 
.A1(n_746),
.A2(n_194),
.B(n_195),
.Y(n_805)
);

HB1xp67_ASAP7_75t_L g806 ( 
.A(n_723),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_746),
.Y(n_807)
);

BUFx12f_ASAP7_75t_L g808 ( 
.A(n_727),
.Y(n_808)
);

OR2x4_ASAP7_75t_L g809 ( 
.A(n_782),
.B(n_727),
.Y(n_809)
);

AND2x4_ASAP7_75t_L g810 ( 
.A(n_748),
.B(n_743),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_748),
.Y(n_811)
);

AND2x4_ASAP7_75t_L g812 ( 
.A(n_748),
.B(n_743),
.Y(n_812)
);

BUFx10_ASAP7_75t_L g813 ( 
.A(n_750),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_808),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_749),
.B(n_743),
.Y(n_815)
);

XOR2xp5_ASAP7_75t_L g816 ( 
.A(n_774),
.B(n_734),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_R g817 ( 
.A(n_793),
.B(n_740),
.Y(n_817)
);

AND2x4_ASAP7_75t_L g818 ( 
.A(n_749),
.B(n_732),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_R g819 ( 
.A(n_808),
.B(n_722),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_749),
.B(n_725),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_R g821 ( 
.A(n_808),
.B(n_742),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_749),
.B(n_721),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_775),
.B(n_695),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_772),
.B(n_721),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_759),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_R g826 ( 
.A(n_792),
.B(n_767),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_806),
.B(n_704),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_755),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_769),
.B(n_754),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_755),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_759),
.B(n_704),
.Y(n_831)
);

XNOR2xp5_ASAP7_75t_L g832 ( 
.A(n_801),
.B(n_255),
.Y(n_832)
);

NAND2xp33_ASAP7_75t_R g833 ( 
.A(n_778),
.B(n_196),
.Y(n_833)
);

OR2x6_ASAP7_75t_L g834 ( 
.A(n_805),
.B(n_197),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_747),
.B(n_198),
.Y(n_835)
);

NAND2xp33_ASAP7_75t_R g836 ( 
.A(n_778),
.B(n_199),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_R g837 ( 
.A(n_767),
.B(n_200),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_759),
.B(n_202),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_760),
.Y(n_839)
);

BUFx3_ASAP7_75t_L g840 ( 
.A(n_761),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_769),
.B(n_204),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_R g842 ( 
.A(n_764),
.B(n_252),
.Y(n_842)
);

AND2x4_ASAP7_75t_L g843 ( 
.A(n_760),
.B(n_205),
.Y(n_843)
);

BUFx3_ASAP7_75t_L g844 ( 
.A(n_761),
.Y(n_844)
);

INVxp67_ASAP7_75t_L g845 ( 
.A(n_770),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_770),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_R g847 ( 
.A(n_782),
.B(n_251),
.Y(n_847)
);

INVxp67_ASAP7_75t_L g848 ( 
.A(n_753),
.Y(n_848)
);

XNOR2xp5_ASAP7_75t_L g849 ( 
.A(n_781),
.B(n_206),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_760),
.B(n_207),
.Y(n_850)
);

NAND2xp33_ASAP7_75t_R g851 ( 
.A(n_781),
.B(n_208),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_804),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_804),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_758),
.B(n_210),
.Y(n_854)
);

BUFx3_ASAP7_75t_L g855 ( 
.A(n_804),
.Y(n_855)
);

INVxp67_ASAP7_75t_L g856 ( 
.A(n_753),
.Y(n_856)
);

INVxp67_ASAP7_75t_L g857 ( 
.A(n_773),
.Y(n_857)
);

BUFx3_ASAP7_75t_L g858 ( 
.A(n_807),
.Y(n_858)
);

NAND2xp33_ASAP7_75t_R g859 ( 
.A(n_786),
.B(n_211),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_755),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_758),
.Y(n_861)
);

OR2x2_ASAP7_75t_L g862 ( 
.A(n_848),
.B(n_856),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_828),
.B(n_800),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_828),
.B(n_800),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_830),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_830),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_860),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_816),
.A2(n_802),
.B1(n_751),
.B2(n_786),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_860),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_825),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_817),
.A2(n_765),
.B1(n_787),
.B2(n_795),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_845),
.Y(n_872)
);

NOR2x1p5_ASAP7_75t_L g873 ( 
.A(n_814),
.B(n_807),
.Y(n_873)
);

OR2x2_ASAP7_75t_L g874 ( 
.A(n_840),
.B(n_798),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_858),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_L g876 ( 
.A1(n_849),
.A2(n_765),
.B1(n_795),
.B2(n_780),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_829),
.B(n_758),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_844),
.B(n_800),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_811),
.Y(n_879)
);

INVxp67_ASAP7_75t_SL g880 ( 
.A(n_852),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_839),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_846),
.Y(n_882)
);

BUFx2_ASAP7_75t_L g883 ( 
.A(n_826),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_861),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_824),
.B(n_798),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_853),
.B(n_803),
.Y(n_886)
);

OR2x2_ASAP7_75t_L g887 ( 
.A(n_855),
.B(n_803),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_823),
.B(n_807),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_857),
.B(n_784),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_819),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_827),
.B(n_813),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_813),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_831),
.Y(n_893)
);

NAND2x1p5_ASAP7_75t_L g894 ( 
.A(n_815),
.B(n_756),
.Y(n_894)
);

INVxp67_ASAP7_75t_SL g895 ( 
.A(n_831),
.Y(n_895)
);

BUFx2_ASAP7_75t_L g896 ( 
.A(n_809),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_810),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_810),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_838),
.B(n_784),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_854),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_838),
.B(n_788),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_815),
.B(n_788),
.Y(n_902)
);

OAI22xp33_ASAP7_75t_L g903 ( 
.A1(n_833),
.A2(n_780),
.B1(n_779),
.B2(n_799),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_812),
.B(n_794),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_843),
.B(n_794),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_812),
.B(n_780),
.Y(n_906)
);

INVx1_ASAP7_75t_SL g907 ( 
.A(n_847),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_820),
.B(n_756),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_835),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_843),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_818),
.B(n_756),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_850),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_818),
.B(n_773),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_850),
.B(n_796),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_820),
.B(n_796),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_834),
.A2(n_765),
.B(n_779),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_834),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_841),
.B(n_796),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_866),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_903),
.A2(n_832),
.B1(n_836),
.B2(n_859),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_866),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_865),
.Y(n_922)
);

NAND4xp25_ASAP7_75t_L g923 ( 
.A(n_876),
.B(n_851),
.C(n_785),
.D(n_789),
.Y(n_923)
);

INVx5_ASAP7_75t_SL g924 ( 
.A(n_902),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_893),
.B(n_902),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_878),
.B(n_791),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_869),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_885),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_878),
.B(n_791),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_867),
.Y(n_930)
);

OAI31xp33_ASAP7_75t_L g931 ( 
.A1(n_903),
.A2(n_821),
.A3(n_842),
.B(n_822),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_867),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_886),
.B(n_791),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_886),
.B(n_791),
.Y(n_934)
);

INVxp67_ASAP7_75t_L g935 ( 
.A(n_891),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_883),
.B(n_822),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_904),
.B(n_789),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_870),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_888),
.B(n_789),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_872),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_881),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_918),
.B(n_785),
.Y(n_942)
);

NAND2xp33_ASAP7_75t_SL g943 ( 
.A(n_890),
.B(n_837),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_863),
.Y(n_944)
);

OAI33xp33_ASAP7_75t_L g945 ( 
.A1(n_909),
.A2(n_868),
.A3(n_862),
.B1(n_892),
.B2(n_882),
.B3(n_877),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_918),
.B(n_785),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_917),
.A2(n_765),
.B1(n_797),
.B2(n_805),
.Y(n_947)
);

AOI31xp33_ASAP7_75t_L g948 ( 
.A1(n_890),
.A2(n_766),
.A3(n_783),
.B(n_768),
.Y(n_948)
);

OR2x2_ASAP7_75t_L g949 ( 
.A(n_874),
.B(n_783),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_879),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_863),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_864),
.Y(n_952)
);

INVxp67_ASAP7_75t_L g953 ( 
.A(n_880),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_889),
.B(n_783),
.Y(n_954)
);

AO21x2_ASAP7_75t_L g955 ( 
.A1(n_916),
.A2(n_768),
.B(n_771),
.Y(n_955)
);

INVxp67_ASAP7_75t_L g956 ( 
.A(n_928),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_938),
.Y(n_957)
);

NOR2xp67_ASAP7_75t_L g958 ( 
.A(n_935),
.B(n_897),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_920),
.A2(n_876),
.B1(n_871),
.B2(n_917),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_925),
.B(n_902),
.Y(n_960)
);

INVxp67_ASAP7_75t_SL g961 ( 
.A(n_953),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_925),
.B(n_895),
.Y(n_962)
);

AOI211xp5_ASAP7_75t_L g963 ( 
.A1(n_923),
.A2(n_907),
.B(n_766),
.C(n_906),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_940),
.B(n_911),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_925),
.B(n_897),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_936),
.B(n_896),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_938),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_941),
.B(n_908),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_941),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_919),
.Y(n_970)
);

NOR2x1p5_ASAP7_75t_L g971 ( 
.A(n_950),
.B(n_898),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_919),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_922),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_950),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_951),
.B(n_952),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_951),
.B(n_887),
.Y(n_976)
);

HB1xp67_ASAP7_75t_SL g977 ( 
.A(n_943),
.Y(n_977)
);

HB1xp67_ASAP7_75t_L g978 ( 
.A(n_944),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_952),
.B(n_894),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_926),
.B(n_894),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_921),
.Y(n_981)
);

OR2x2_ASAP7_75t_L g982 ( 
.A(n_944),
.B(n_915),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_921),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_R g984 ( 
.A(n_977),
.B(n_943),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_963),
.A2(n_871),
.B1(n_948),
.B2(n_924),
.Y(n_985)
);

OAI22xp33_ASAP7_75t_L g986 ( 
.A1(n_959),
.A2(n_947),
.B1(n_910),
.B2(n_912),
.Y(n_986)
);

AO221x2_ASAP7_75t_L g987 ( 
.A1(n_964),
.A2(n_945),
.B1(n_931),
.B2(n_927),
.C(n_913),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_961),
.B(n_937),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_956),
.B(n_937),
.Y(n_989)
);

NOR4xp25_ASAP7_75t_SL g990 ( 
.A(n_971),
.B(n_924),
.C(n_884),
.D(n_955),
.Y(n_990)
);

OAI22xp33_ASAP7_75t_L g991 ( 
.A1(n_958),
.A2(n_898),
.B1(n_900),
.B2(n_879),
.Y(n_991)
);

AO221x2_ASAP7_75t_L g992 ( 
.A1(n_973),
.A2(n_930),
.B1(n_932),
.B2(n_900),
.C(n_924),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_974),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_SL g994 ( 
.A(n_966),
.B(n_908),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_968),
.B(n_939),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_960),
.B(n_924),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_962),
.B(n_939),
.Y(n_997)
);

OAI22xp33_ASAP7_75t_L g998 ( 
.A1(n_974),
.A2(n_949),
.B1(n_875),
.B2(n_901),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_962),
.B(n_942),
.Y(n_999)
);

NAND2xp33_ASAP7_75t_SL g1000 ( 
.A(n_965),
.B(n_873),
.Y(n_1000)
);

OR2x2_ASAP7_75t_L g1001 ( 
.A(n_997),
.B(n_982),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_984),
.Y(n_1002)
);

OR2x2_ASAP7_75t_L g1003 ( 
.A(n_999),
.B(n_982),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_989),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_993),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_988),
.Y(n_1006)
);

INVx1_ASAP7_75t_SL g1007 ( 
.A(n_1000),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_995),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_987),
.Y(n_1009)
);

BUFx2_ASAP7_75t_L g1010 ( 
.A(n_996),
.Y(n_1010)
);

CKINVDCx16_ASAP7_75t_R g1011 ( 
.A(n_994),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_992),
.Y(n_1012)
);

NOR2x1_ASAP7_75t_L g1013 ( 
.A(n_991),
.B(n_983),
.Y(n_1013)
);

OAI221xp5_ASAP7_75t_L g1014 ( 
.A1(n_1009),
.A2(n_985),
.B1(n_987),
.B2(n_969),
.C(n_957),
.Y(n_1014)
);

O2A1O1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_1007),
.A2(n_986),
.B(n_998),
.C(n_955),
.Y(n_1015)
);

OAI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_1011),
.A2(n_992),
.B1(n_976),
.B2(n_978),
.Y(n_1016)
);

XNOR2xp5_ASAP7_75t_L g1017 ( 
.A(n_1002),
.B(n_965),
.Y(n_1017)
);

AO22x1_ASAP7_75t_L g1018 ( 
.A1(n_1007),
.A2(n_990),
.B1(n_960),
.B2(n_980),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_1006),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_1012),
.A2(n_979),
.B(n_980),
.C(n_797),
.Y(n_1020)
);

OAI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_1012),
.A2(n_976),
.B1(n_875),
.B2(n_967),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_1014),
.A2(n_1013),
.B(n_1005),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_1017),
.B(n_1004),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_1019),
.Y(n_1024)
);

AOI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_1016),
.A2(n_1010),
.B1(n_1008),
.B2(n_1003),
.Y(n_1025)
);

NAND2x1_ASAP7_75t_SL g1026 ( 
.A(n_1018),
.B(n_979),
.Y(n_1026)
);

BUFx4_ASAP7_75t_SL g1027 ( 
.A(n_1023),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1024),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1025),
.Y(n_1029)
);

INVxp33_ASAP7_75t_SL g1030 ( 
.A(n_1022),
.Y(n_1030)
);

INVx2_ASAP7_75t_SL g1031 ( 
.A(n_1026),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_1030),
.B(n_1015),
.Y(n_1032)
);

NAND3xp33_ASAP7_75t_L g1033 ( 
.A(n_1029),
.B(n_1020),
.C(n_1021),
.Y(n_1033)
);

NAND4xp25_ASAP7_75t_L g1034 ( 
.A(n_1030),
.B(n_1003),
.C(n_1001),
.D(n_875),
.Y(n_1034)
);

AOI211xp5_ASAP7_75t_L g1035 ( 
.A1(n_1031),
.A2(n_983),
.B(n_901),
.C(n_905),
.Y(n_1035)
);

INVxp33_ASAP7_75t_L g1036 ( 
.A(n_1028),
.Y(n_1036)
);

NAND4xp25_ASAP7_75t_L g1037 ( 
.A(n_1027),
.B(n_908),
.C(n_899),
.D(n_905),
.Y(n_1037)
);

NAND4xp75_ASAP7_75t_L g1038 ( 
.A(n_1031),
.B(n_899),
.C(n_933),
.D(n_934),
.Y(n_1038)
);

OAI221xp5_ASAP7_75t_SL g1039 ( 
.A1(n_1033),
.A2(n_981),
.B1(n_972),
.B2(n_970),
.C(n_949),
.Y(n_1039)
);

AOI222xp33_ASAP7_75t_L g1040 ( 
.A1(n_1032),
.A2(n_975),
.B1(n_981),
.B2(n_972),
.C1(n_970),
.C2(n_930),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1036),
.Y(n_1041)
);

AOI21xp33_ASAP7_75t_SL g1042 ( 
.A1(n_1034),
.A2(n_212),
.B(n_213),
.Y(n_1042)
);

NAND3xp33_ASAP7_75t_L g1043 ( 
.A(n_1035),
.B(n_932),
.C(n_934),
.Y(n_1043)
);

AOI21xp33_ASAP7_75t_L g1044 ( 
.A1(n_1038),
.A2(n_1037),
.B(n_955),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_1041),
.B(n_975),
.Y(n_1045)
);

NOR2x1_ASAP7_75t_L g1046 ( 
.A(n_1043),
.B(n_790),
.Y(n_1046)
);

XOR2x2_ASAP7_75t_L g1047 ( 
.A(n_1039),
.B(n_215),
.Y(n_1047)
);

NOR3xp33_ASAP7_75t_L g1048 ( 
.A(n_1042),
.B(n_790),
.C(n_763),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_1040),
.B(n_933),
.Y(n_1049)
);

INVxp33_ASAP7_75t_SL g1050 ( 
.A(n_1044),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_1041),
.B(n_929),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_1050),
.B(n_946),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_1048),
.B(n_946),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1047),
.B(n_929),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_R g1055 ( 
.A(n_1045),
.B(n_217),
.Y(n_1055)
);

NAND2xp33_ASAP7_75t_SL g1056 ( 
.A(n_1051),
.B(n_954),
.Y(n_1056)
);

NAND3xp33_ASAP7_75t_SL g1057 ( 
.A(n_1046),
.B(n_942),
.C(n_914),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_R g1058 ( 
.A(n_1049),
.B(n_218),
.Y(n_1058)
);

XNOR2xp5_ASAP7_75t_L g1059 ( 
.A(n_1047),
.B(n_219),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_1050),
.B(n_954),
.Y(n_1060)
);

OAI222xp33_ASAP7_75t_L g1061 ( 
.A1(n_1052),
.A2(n_926),
.B1(n_757),
.B2(n_776),
.C1(n_914),
.C2(n_777),
.Y(n_1061)
);

CKINVDCx20_ASAP7_75t_R g1062 ( 
.A(n_1059),
.Y(n_1062)
);

AOI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_1060),
.A2(n_752),
.B1(n_790),
.B2(n_777),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1054),
.Y(n_1064)
);

INVxp33_ASAP7_75t_SL g1065 ( 
.A(n_1055),
.Y(n_1065)
);

BUFx2_ASAP7_75t_L g1066 ( 
.A(n_1058),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_1053),
.B(n_864),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1056),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_SL g1069 ( 
.A1(n_1057),
.A2(n_771),
.B1(n_768),
.B2(n_776),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_1054),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_1059),
.B(n_220),
.Y(n_1071)
);

NAND2xp33_ASAP7_75t_SL g1072 ( 
.A(n_1055),
.B(n_771),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1054),
.Y(n_1073)
);

XOR2x1_ASAP7_75t_L g1074 ( 
.A(n_1070),
.B(n_221),
.Y(n_1074)
);

OAI221xp5_ASAP7_75t_R g1075 ( 
.A1(n_1062),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.C(n_225),
.Y(n_1075)
);

AOI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_1065),
.A2(n_790),
.B1(n_777),
.B2(n_763),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1066),
.Y(n_1077)
);

AND3x1_ASAP7_75t_L g1078 ( 
.A(n_1068),
.B(n_227),
.C(n_229),
.Y(n_1078)
);

OA22x2_ASAP7_75t_L g1079 ( 
.A1(n_1064),
.A2(n_776),
.B1(n_777),
.B2(n_763),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_SL g1080 ( 
.A1(n_1073),
.A2(n_763),
.B1(n_752),
.B2(n_232),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1071),
.Y(n_1081)
);

AND2x2_ASAP7_75t_SL g1082 ( 
.A(n_1078),
.B(n_1071),
.Y(n_1082)
);

AO22x2_ASAP7_75t_L g1083 ( 
.A1(n_1077),
.A2(n_1067),
.B1(n_1072),
.B2(n_1069),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1074),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1081),
.Y(n_1085)
);

NAND2x1_ASAP7_75t_SL g1086 ( 
.A(n_1075),
.B(n_1063),
.Y(n_1086)
);

AOI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_1084),
.A2(n_1080),
.B1(n_1079),
.B2(n_1076),
.Y(n_1087)
);

AOI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_1082),
.A2(n_1061),
.B1(n_752),
.B2(n_762),
.Y(n_1088)
);

AOI31xp33_ASAP7_75t_L g1089 ( 
.A1(n_1085),
.A2(n_230),
.A3(n_231),
.B(n_233),
.Y(n_1089)
);

AOI31xp33_ASAP7_75t_L g1090 ( 
.A1(n_1086),
.A2(n_1083),
.A3(n_235),
.B(n_236),
.Y(n_1090)
);

XNOR2xp5_ASAP7_75t_L g1091 ( 
.A(n_1087),
.B(n_234),
.Y(n_1091)
);

AOI222xp33_ASAP7_75t_L g1092 ( 
.A1(n_1091),
.A2(n_1088),
.B1(n_1090),
.B2(n_1089),
.C1(n_752),
.C2(n_242),
.Y(n_1092)
);

AOI22xp33_ASAP7_75t_SL g1093 ( 
.A1(n_1091),
.A2(n_762),
.B1(n_239),
.B2(n_240),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_1092),
.Y(n_1094)
);

AND2x4_ASAP7_75t_L g1095 ( 
.A(n_1093),
.B(n_238),
.Y(n_1095)
);

OAI221xp5_ASAP7_75t_L g1096 ( 
.A1(n_1094),
.A2(n_1095),
.B1(n_243),
.B2(n_244),
.C(n_245),
.Y(n_1096)
);

AOI211xp5_ASAP7_75t_L g1097 ( 
.A1(n_1096),
.A2(n_1095),
.B(n_246),
.C(n_247),
.Y(n_1097)
);


endmodule