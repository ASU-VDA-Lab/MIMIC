module fake_netlist_5_1022_n_37 (n_8, n_10, n_4, n_5, n_7, n_0, n_12, n_9, n_14, n_2, n_13, n_3, n_11, n_6, n_1, n_37);

input n_8;
input n_10;
input n_4;
input n_5;
input n_7;
input n_0;
input n_12;
input n_9;
input n_14;
input n_2;
input n_13;
input n_3;
input n_11;
input n_6;
input n_1;

output n_37;

wire n_29;
wire n_16;
wire n_36;
wire n_25;
wire n_18;
wire n_27;
wire n_22;
wire n_28;
wire n_24;
wire n_21;
wire n_34;
wire n_32;
wire n_35;
wire n_17;
wire n_19;
wire n_15;
wire n_26;
wire n_30;
wire n_33;
wire n_31;
wire n_23;
wire n_20;

CKINVDCx5p33_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_2),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_6),
.B(n_13),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_17),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_7),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

NAND3xp33_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_22),
.C(n_20),
.Y(n_27)
);

OAI21x1_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_18),
.B(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_29),
.B(n_24),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_30),
.A2(n_27),
.B1(n_15),
.B2(n_19),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_8),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_26),
.B(n_12),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_0),
.Y(n_34)
);

NAND2x1p5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_26),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_33),
.Y(n_37)
);


endmodule