module fake_jpeg_9917_n_330 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx5_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_37),
.Y(n_52)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_26),
.Y(n_38)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_22),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_0),
.Y(n_42)
);

AOI21xp33_ASAP7_75t_L g71 ( 
.A1(n_42),
.A2(n_43),
.B(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_22),
.B(n_1),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_22),
.B(n_1),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_19),
.B1(n_29),
.B2(n_17),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_46),
.A2(n_62),
.B1(n_34),
.B2(n_28),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_47),
.Y(n_83)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_49),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_40),
.B(n_21),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_17),
.B1(n_19),
.B2(n_29),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_51),
.A2(n_70),
.B1(n_30),
.B2(n_38),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_40),
.B(n_21),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_59),
.B(n_63),
.Y(n_95)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_44),
.A2(n_26),
.B1(n_19),
.B2(n_29),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_23),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_68),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_36),
.A2(n_17),
.B1(n_30),
.B2(n_26),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_66),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_76),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_45),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_36),
.B1(n_30),
.B2(n_42),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_78),
.A2(n_87),
.B1(n_88),
.B2(n_20),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_55),
.A2(n_30),
.B1(n_25),
.B2(n_23),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_69),
.A2(n_34),
.B1(n_28),
.B2(n_23),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_86),
.A2(n_90),
.B1(n_91),
.B2(n_38),
.Y(n_102)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_48),
.A2(n_38),
.B1(n_25),
.B2(n_22),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_69),
.A2(n_34),
.B1(n_28),
.B2(n_25),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_55),
.A2(n_33),
.B1(n_38),
.B2(n_20),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_45),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_32),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_43),
.C(n_42),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_32),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_47),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_97),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_47),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_75),
.A2(n_43),
.B(n_50),
.C(n_33),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_103),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_101),
.B(n_83),
.C(n_88),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_102),
.A2(n_110),
.B1(n_120),
.B2(n_73),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_76),
.B(n_67),
.Y(n_103)
);

INVxp33_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_121),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_73),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_105),
.B(n_109),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_67),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_113),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_74),
.B(n_33),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_93),
.A2(n_50),
.B1(n_60),
.B2(n_63),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_111),
.B(n_125),
.Y(n_151)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_112),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_95),
.B(n_57),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_58),
.Y(n_115)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_64),
.Y(n_116)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_77),
.B(n_47),
.Y(n_117)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_77),
.B(n_32),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_118),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_95),
.B(n_31),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_61),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_82),
.A2(n_54),
.B1(n_53),
.B2(n_65),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_86),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_123),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_73),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_124),
.A2(n_126),
.B1(n_90),
.B2(n_91),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_87),
.A2(n_65),
.B1(n_61),
.B2(n_20),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_129),
.A2(n_136),
.B1(n_137),
.B2(n_145),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_140),
.Y(n_175)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_105),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_110),
.A2(n_75),
.B1(n_78),
.B2(n_98),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_101),
.B(n_75),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_149),
.C(n_157),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_98),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_79),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_119),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_122),
.A2(n_106),
.B(n_114),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_144),
.A2(n_148),
.B(n_120),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_124),
.A2(n_85),
.B1(n_79),
.B2(n_88),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_97),
.Y(n_146)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_94),
.Y(n_147)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_101),
.B(n_88),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_81),
.Y(n_150)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_150),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_81),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_152),
.B(n_116),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_96),
.B1(n_72),
.B2(n_80),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_153),
.A2(n_154),
.B1(n_129),
.B2(n_145),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_126),
.A2(n_100),
.B1(n_111),
.B2(n_102),
.Y(n_154)
);

BUFx24_ASAP7_75t_L g155 ( 
.A(n_99),
.Y(n_155)
);

INVx5_ASAP7_75t_SL g163 ( 
.A(n_155),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_110),
.B(n_88),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_144),
.A2(n_102),
.B1(n_100),
.B2(n_120),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_159),
.A2(n_179),
.B(n_183),
.Y(n_190)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_160),
.Y(n_215)
);

AND2x6_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_99),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_164),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_123),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_165),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_131),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_166),
.B(n_169),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_128),
.B(n_125),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_167),
.B(n_32),
.Y(n_207)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_170),
.Y(n_203)
);

AND2x6_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_103),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_171),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_133),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_172),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_127),
.B(n_109),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_173),
.Y(n_216)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_176),
.Y(n_200)
);

AND2x6_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_108),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_141),
.B(n_117),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_181),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_113),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_188),
.C(n_130),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_139),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_151),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_140),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_128),
.B(n_118),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_143),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_189),
.A2(n_132),
.B1(n_154),
.B2(n_151),
.Y(n_191)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_183),
.A2(n_155),
.B(n_132),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_194),
.A2(n_201),
.B(n_202),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_195),
.B(n_196),
.C(n_197),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_137),
.C(n_157),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_136),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_130),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_199),
.B(n_204),
.C(n_210),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_159),
.A2(n_142),
.B(n_127),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_179),
.A2(n_155),
.B(n_142),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_167),
.B(n_141),
.C(n_155),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_161),
.A2(n_126),
.B1(n_83),
.B2(n_96),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_206),
.A2(n_169),
.B1(n_186),
.B2(n_158),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_207),
.B(n_181),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_174),
.A2(n_72),
.B1(n_83),
.B2(n_31),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_208),
.A2(n_213),
.B1(n_168),
.B2(n_170),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_189),
.C(n_188),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_161),
.A2(n_31),
.B1(n_27),
.B2(n_20),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_175),
.B(n_171),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_163),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_164),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_238),
.C(n_201),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_214),
.B(n_177),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_223),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_220),
.A2(n_213),
.B1(n_191),
.B2(n_204),
.Y(n_250)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_221),
.B(n_235),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_202),
.A2(n_163),
.B1(n_178),
.B2(n_175),
.Y(n_222)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_222),
.Y(n_253)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_205),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_224),
.B(n_230),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_190),
.Y(n_248)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_231),
.Y(n_247)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_228),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_31),
.Y(n_229)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_229),
.Y(n_260)
);

XNOR2x1_ASAP7_75t_L g230 ( 
.A(n_190),
.B(n_32),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_27),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_198),
.B(n_18),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_232),
.B(n_234),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_192),
.B(n_18),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_200),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_240),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_196),
.B(n_32),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_194),
.Y(n_239)
);

INVxp33_ASAP7_75t_SL g244 ( 
.A(n_239),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_203),
.B(n_10),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_208),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_243),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_10),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_245),
.B(n_248),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_230),
.A2(n_209),
.B1(n_193),
.B2(n_217),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_249),
.A2(n_265),
.B1(n_9),
.B2(n_15),
.Y(n_275)
);

O2A1O1Ixp33_ASAP7_75t_L g270 ( 
.A1(n_250),
.A2(n_228),
.B(n_224),
.C(n_238),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_225),
.A2(n_215),
.B(n_210),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_251),
.A2(n_233),
.B(n_231),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_195),
.C(n_199),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_236),
.C(n_241),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_218),
.B(n_207),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_8),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_221),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_2),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_225),
.A2(n_206),
.B1(n_215),
.B2(n_27),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_261),
.A2(n_264),
.B1(n_11),
.B2(n_15),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_227),
.A2(n_27),
.B1(n_18),
.B2(n_9),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_220),
.A2(n_233),
.B1(n_242),
.B2(n_226),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_279),
.C(n_280),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_267),
.A2(n_251),
.B(n_256),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_229),
.Y(n_268)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_268),
.Y(n_286)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_247),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_281),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_270),
.A2(n_255),
.B1(n_258),
.B2(n_248),
.Y(n_290)
);

O2A1O1Ixp33_ASAP7_75t_L g271 ( 
.A1(n_244),
.A2(n_241),
.B(n_2),
.C(n_3),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_271),
.A2(n_249),
.B1(n_255),
.B2(n_262),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_280),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_257),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_273),
.A2(n_275),
.B1(n_256),
.B2(n_254),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_274),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_246),
.B(n_11),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_276),
.B(n_277),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_252),
.B(n_8),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_245),
.B(n_16),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_16),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_261),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_289),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_267),
.A2(n_253),
.B1(n_260),
.B2(n_265),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_283),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_302)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_284),
.Y(n_297)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_287),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_271),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_13),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_293),
.B(n_278),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_294),
.A2(n_270),
.B(n_272),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_266),
.B(n_247),
.C(n_254),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_278),
.C(n_14),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_296),
.A2(n_283),
.B(n_292),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_279),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_303),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_300),
.A2(n_302),
.B1(n_287),
.B2(n_291),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_305),
.C(n_288),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_12),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_12),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_304),
.B(n_306),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_14),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_308),
.A2(n_307),
.B(n_296),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_6),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_286),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_314),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_313),
.B(n_7),
.Y(n_323)
);

AOI31xp67_ASAP7_75t_L g314 ( 
.A1(n_302),
.A2(n_284),
.A3(n_288),
.B(n_6),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_4),
.C(n_5),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_316),
.C(n_7),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_4),
.C(n_5),
.Y(n_316)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_317),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_311),
.B(n_305),
.Y(n_318)
);

NOR3xp33_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_319),
.C(n_320),
.Y(n_325)
);

MAJx2_ASAP7_75t_L g319 ( 
.A(n_316),
.B(n_5),
.C(n_6),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_322),
.A2(n_323),
.B(n_312),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_318),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_327),
.B(n_321),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_324),
.B(n_309),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_325),
.Y(n_330)
);


endmodule