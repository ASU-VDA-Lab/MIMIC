module real_jpeg_23220_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_213;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_1),
.A2(n_35),
.B1(n_36),
.B2(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_1),
.A2(n_60),
.B1(n_69),
.B2(n_70),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_1),
.A2(n_53),
.B1(n_54),
.B2(n_60),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

INVx8_ASAP7_75t_SL g34 ( 
.A(n_4),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_5),
.A2(n_69),
.B1(n_70),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_5),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_5),
.A2(n_53),
.B1(n_54),
.B2(n_84),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_6),
.A2(n_69),
.B1(n_70),
.B2(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_6),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_7),
.A2(n_53),
.B1(n_54),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_7),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_7),
.A2(n_35),
.B1(n_36),
.B2(n_73),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_7),
.A2(n_69),
.B1(n_70),
.B2(n_73),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_8),
.B(n_41),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_8),
.B(n_65),
.C(n_69),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_8),
.A2(n_28),
.B1(n_53),
.B2(n_54),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_8),
.B(n_58),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_8),
.A2(n_85),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_12),
.A2(n_35),
.B1(n_36),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_12),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_12),
.A2(n_27),
.B1(n_40),
.B2(n_49),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_12),
.A2(n_49),
.B1(n_53),
.B2(n_54),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_12),
.A2(n_49),
.B1(n_69),
.B2(n_70),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_13),
.A2(n_53),
.B1(n_54),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_13),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_13),
.A2(n_69),
.B1(n_70),
.B2(n_76),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_14),
.A2(n_24),
.B1(n_39),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_14),
.A2(n_35),
.B1(n_36),
.B2(n_44),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_14),
.A2(n_44),
.B1(n_53),
.B2(n_54),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_14),
.A2(n_44),
.B1(n_69),
.B2(n_70),
.Y(n_169)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_15),
.Y(n_86)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_15),
.Y(n_89)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_15),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_133),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_131),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_103),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_20),
.B(n_103),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_78),
.C(n_90),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_21),
.B(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_45),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_22),
.B(n_47),
.C(n_61),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_31),
.B1(n_41),
.B2(n_42),
.Y(n_22)
);

OAI21xp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B(n_29),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_28),
.B(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_28),
.B(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_28),
.B(n_68),
.Y(n_178)
);

HAxp5_ASAP7_75t_SL g187 ( 
.A(n_28),
.B(n_36),
.CON(n_187),
.SN(n_187)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_29),
.A2(n_33),
.B(n_36),
.C(n_80),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_33),
.B1(n_34),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_31),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_38),
.Y(n_31)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_32),
.A2(n_43),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND3xp33_ASAP7_75t_L g80 ( 
.A(n_34),
.B(n_35),
.C(n_40),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_36),
.B1(n_52),
.B2(n_56),
.Y(n_57)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND3xp33_ASAP7_75t_L g188 ( 
.A(n_36),
.B(n_53),
.C(n_56),
.Y(n_188)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_47),
.B1(n_61),
.B2(n_62),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_50),
.B1(n_58),
.B2(n_59),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_48),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_50),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_50),
.A2(n_58),
.B1(n_93),
.B2(n_187),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_57),
.Y(n_50)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_51),
.A2(n_92),
.B1(n_94),
.B2(n_95),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_51)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_52),
.A2(n_54),
.B(n_187),
.C(n_188),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_53),
.A2(n_54),
.B1(n_65),
.B2(n_67),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_54),
.B(n_140),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_58),
.B(n_128),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_59),
.Y(n_126)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_71),
.B(n_74),
.Y(n_62)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_63),
.A2(n_68),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_63),
.A2(n_68),
.B1(n_144),
.B2(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_63),
.A2(n_209),
.B(n_210),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_68),
.Y(n_63)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_67),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

BUFx24_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_68),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_68),
.A2(n_113),
.B(n_114),
.Y(n_112)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_70),
.B(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_72),
.B(n_77),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_77),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_75),
.B(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_77),
.A2(n_115),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_78),
.B(n_90),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_79),
.B(n_81),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_85),
.B1(n_87),
.B2(n_89),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_85),
.A2(n_87),
.B(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_85),
.A2(n_153),
.B(n_154),
.Y(n_152)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_85),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_85),
.A2(n_162),
.B1(n_169),
.B2(n_175),
.Y(n_179)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_86),
.Y(n_100)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_86),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_96),
.C(n_98),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_91),
.B(n_204),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_126),
.B(n_127),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_204)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_100),
.A2(n_160),
.B1(n_161),
.B2(n_163),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_110),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_118),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_116),
.B2(n_117),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_112),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_109),
.A2(n_156),
.B(n_160),
.Y(n_189)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_110),
.Y(n_155)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_129),
.B2(n_130),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_125),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_129),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_214),
.B(n_218),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_199),
.B(n_213),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_183),
.B(n_198),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_157),
.B(n_182),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_145),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_145),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_139),
.A2(n_141),
.B1(n_142),
.B2(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_139),
.Y(n_165)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_152),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_147),
.B(n_150),
.C(n_152),
.Y(n_197)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_151),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_153),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_166),
.B(n_181),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_164),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_164),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_177),
.B(n_180),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_173),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_178),
.B(n_179),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_197),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_197),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_192),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_193),
.C(n_196),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_186),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_191),
.Y(n_207)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_189),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_196),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_195),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_200),
.B(n_201),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_205),
.B2(n_206),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_208),
.C(n_211),
.Y(n_217)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_211),
.B2(n_212),
.Y(n_206)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_208),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_217),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_217),
.Y(n_218)
);


endmodule