module fake_jpeg_1906_n_541 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_541);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_541;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_13),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_57),
.Y(n_136)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_58),
.Y(n_185)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_62),
.Y(n_184)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_63),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_28),
.C(n_20),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_64),
.B(n_24),
.C(n_51),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_65),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_20),
.B(n_28),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_66),
.B(n_110),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_67),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_68),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_69),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_72),
.Y(n_186)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_73),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_74),
.Y(n_164)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_76),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_77),
.Y(n_177)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_78),
.Y(n_153)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_79),
.Y(n_133)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g171 ( 
.A(n_80),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_82),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_83),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_84),
.Y(n_183)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_85),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_54),
.B(n_0),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_86),
.B(n_118),
.Y(n_199)
);

BUFx8_ASAP7_75t_L g87 ( 
.A(n_18),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g205 ( 
.A(n_87),
.Y(n_205)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_89),
.Y(n_190)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_90),
.Y(n_162)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_91),
.Y(n_150)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_92),
.Y(n_176)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_93),
.Y(n_151)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g182 ( 
.A(n_94),
.Y(n_182)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_95),
.Y(n_154)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_96),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_27),
.B(n_16),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_97),
.B(n_114),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_98),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_99),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_101),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_18),
.Y(n_102)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_102),
.Y(n_172)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_103),
.Y(n_192)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_19),
.Y(n_104)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_104),
.Y(n_193)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_105),
.Y(n_194)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_106),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_18),
.Y(n_107)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_107),
.Y(n_197)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_21),
.Y(n_108)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_25),
.Y(n_109)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_109),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_56),
.B(n_15),
.Y(n_110)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_111),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_19),
.Y(n_112)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_112),
.Y(n_173)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_21),
.Y(n_113)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_113),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_27),
.B(n_0),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_41),
.Y(n_115)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_115),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_41),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_116),
.Y(n_137)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_49),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_49),
.Y(n_126)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_25),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_25),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_119),
.B(n_39),
.Y(n_200)
);

AOI21xp33_ASAP7_75t_L g120 ( 
.A1(n_22),
.A2(n_0),
.B(n_1),
.Y(n_120)
);

OR2x2_ASAP7_75t_SL g148 ( 
.A(n_120),
.B(n_121),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_25),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_25),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_47),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_86),
.A2(n_41),
.B1(n_47),
.B2(n_49),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_124),
.A2(n_204),
.B1(n_185),
.B2(n_190),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_126),
.B(n_200),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_127),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_97),
.A2(n_41),
.B1(n_47),
.B2(n_52),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_128),
.A2(n_134),
.B1(n_149),
.B2(n_170),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_56),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_130),
.B(n_132),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_70),
.B(n_53),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_62),
.A2(n_47),
.B1(n_31),
.B2(n_30),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_81),
.B(n_52),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_135),
.B(n_143),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_138),
.B(n_15),
.C(n_9),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_43),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_62),
.A2(n_87),
.B1(n_57),
.B2(n_39),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_68),
.B(n_24),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_158),
.B(n_160),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_90),
.B(n_50),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_61),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_166),
.B(n_181),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_74),
.B(n_22),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_168),
.B(n_169),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_92),
.B(n_29),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_77),
.A2(n_29),
.B1(n_50),
.B2(n_32),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_106),
.A2(n_30),
.B1(n_31),
.B2(n_39),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_174),
.A2(n_188),
.B1(n_202),
.B2(n_8),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_83),
.A2(n_32),
.B1(n_51),
.B2(n_34),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_46),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_111),
.B(n_53),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_84),
.A2(n_38),
.B1(n_43),
.B2(n_40),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_89),
.B(n_40),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_189),
.B(n_11),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_99),
.A2(n_38),
.B1(n_34),
.B2(n_31),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_101),
.A2(n_116),
.B1(n_115),
.B2(n_112),
.Y(n_204)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_193),
.Y(n_206)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_206),
.Y(n_288)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_192),
.Y(n_207)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_207),
.Y(n_293)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_142),
.Y(n_208)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_208),
.Y(n_289)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_152),
.Y(n_210)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_210),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_147),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_211),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_199),
.A2(n_30),
.B1(n_46),
.B2(n_33),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_212),
.A2(n_155),
.B(n_176),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_184),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_213),
.Y(n_281)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_180),
.Y(n_214)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_214),
.Y(n_309)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_125),
.Y(n_215)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_215),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_216),
.B(n_247),
.Y(n_283)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_142),
.Y(n_217)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_217),
.Y(n_319)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_184),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_218),
.Y(n_313)
);

AOI21xp33_ASAP7_75t_L g219 ( 
.A1(n_148),
.A2(n_46),
.B(n_2),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_219),
.A2(n_187),
.B(n_203),
.Y(n_299)
);

FAx1_ASAP7_75t_SL g220 ( 
.A(n_148),
.B(n_123),
.CI(n_165),
.CON(n_220),
.SN(n_220)
);

OAI32xp33_ASAP7_75t_L g276 ( 
.A1(n_220),
.A2(n_198),
.A3(n_171),
.B1(n_175),
.B2(n_191),
.Y(n_276)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_140),
.Y(n_222)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_222),
.Y(n_311)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_147),
.Y(n_223)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_223),
.Y(n_320)
);

OAI22xp33_ASAP7_75t_L g224 ( 
.A1(n_137),
.A2(n_104),
.B1(n_73),
.B2(n_3),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_224),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_310)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_145),
.Y(n_225)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_225),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_165),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_L g227 ( 
.A1(n_134),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_204),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_228)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_162),
.Y(n_230)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_230),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_144),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_231),
.Y(n_277)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_146),
.Y(n_232)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_232),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_163),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_233),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_157),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_234),
.Y(n_317)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_150),
.Y(n_235)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_235),
.Y(n_326)
);

INVx8_ASAP7_75t_L g237 ( 
.A(n_196),
.Y(n_237)
);

INVx5_ASAP7_75t_L g301 ( 
.A(n_237),
.Y(n_301)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_151),
.Y(n_238)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_238),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_131),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_239),
.A2(n_241),
.B1(n_253),
.B2(n_258),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_161),
.Y(n_240)
);

INVxp33_ASAP7_75t_L g300 ( 
.A(n_240),
.Y(n_300)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_133),
.Y(n_242)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_242),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_243),
.B(n_182),
.Y(n_324)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_173),
.Y(n_244)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_244),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_167),
.Y(n_245)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_245),
.Y(n_298)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_201),
.Y(n_246)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_246),
.Y(n_316)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_156),
.Y(n_247)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_195),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_250),
.B(n_254),
.Y(n_307)
);

OAI22xp33_ASAP7_75t_L g251 ( 
.A1(n_174),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_251),
.A2(n_267),
.B1(n_273),
.B2(n_185),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_129),
.B(n_9),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_252),
.B(n_255),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_139),
.A2(n_159),
.B1(n_194),
.B2(n_154),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_129),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_141),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_197),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_257),
.Y(n_275)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_153),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_172),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_262),
.Y(n_286)
);

INVx8_ASAP7_75t_L g260 ( 
.A(n_196),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_260),
.A2(n_261),
.B1(n_268),
.B2(n_191),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_141),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_153),
.B(n_12),
.Y(n_262)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_136),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_263),
.Y(n_322)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_139),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_264),
.B(n_265),
.Y(n_302)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_186),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_159),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_266),
.B(n_269),
.Y(n_306)
);

OAI22xp33_ASAP7_75t_L g267 ( 
.A1(n_149),
.A2(n_14),
.B1(n_15),
.B2(n_178),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_157),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_186),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_162),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_270),
.B(n_272),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_205),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_276),
.B(n_212),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_279),
.A2(n_182),
.B1(n_268),
.B2(n_297),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_229),
.A2(n_178),
.B1(n_190),
.B2(n_164),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_282),
.A2(n_323),
.B1(n_261),
.B2(n_216),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_285),
.A2(n_299),
.B(n_283),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_287),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_243),
.B(n_136),
.C(n_175),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_291),
.B(n_324),
.Y(n_340)
);

OAI32xp33_ASAP7_75t_L g295 ( 
.A1(n_271),
.A2(n_220),
.A3(n_209),
.B1(n_248),
.B2(n_274),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_295),
.B(n_220),
.Y(n_332)
);

O2A1O1Ixp33_ASAP7_75t_L g296 ( 
.A1(n_219),
.A2(n_198),
.B(n_155),
.C(n_176),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_296),
.A2(n_227),
.B(n_230),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_273),
.A2(n_164),
.B1(n_177),
.B2(n_183),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_297),
.A2(n_224),
.B1(n_253),
.B2(n_304),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_271),
.B(n_177),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_304),
.B(n_314),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_249),
.B(n_183),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_236),
.B(n_171),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_315),
.B(n_263),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_L g323 ( 
.A1(n_228),
.A2(n_187),
.B1(n_203),
.B2(n_171),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_327),
.Y(n_367)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_302),
.Y(n_328)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_328),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_286),
.B(n_221),
.Y(n_329)
);

NAND3xp33_ASAP7_75t_L g370 ( 
.A(n_329),
.B(n_332),
.C(n_344),
.Y(n_370)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_294),
.Y(n_330)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_330),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_SL g388 ( 
.A1(n_331),
.A2(n_355),
.B1(n_358),
.B2(n_359),
.Y(n_388)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_306),
.Y(n_334)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_334),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_335),
.A2(n_345),
.B1(n_356),
.B2(n_362),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_296),
.A2(n_226),
.B(n_258),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_337),
.A2(n_342),
.B(n_307),
.Y(n_371)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_278),
.Y(n_338)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_338),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_308),
.B(n_315),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_339),
.B(n_343),
.Y(n_381)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_313),
.Y(n_341)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_341),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_299),
.A2(n_239),
.B(n_251),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_311),
.B(n_217),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_314),
.B(n_208),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_284),
.A2(n_260),
.B1(n_237),
.B2(n_267),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_318),
.B(n_298),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_346),
.Y(n_394)
);

INVx5_ASAP7_75t_L g347 ( 
.A(n_301),
.Y(n_347)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_347),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_348),
.B(n_352),
.Y(n_390)
);

OAI21xp33_ASAP7_75t_SL g373 ( 
.A1(n_349),
.A2(n_353),
.B(n_360),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_324),
.B(n_206),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_350),
.B(n_351),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_291),
.B(n_213),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_295),
.B(n_234),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_303),
.B(n_218),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_275),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_354),
.Y(n_377)
);

BUFx12f_ASAP7_75t_L g355 ( 
.A(n_289),
.Y(n_355)
);

AO22x2_ASAP7_75t_L g357 ( 
.A1(n_310),
.A2(n_182),
.B1(n_276),
.B2(n_285),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_357),
.B(n_361),
.Y(n_391)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_288),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_313),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_283),
.B(n_322),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_283),
.A2(n_310),
.B1(n_298),
.B2(n_325),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_325),
.B(n_290),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_363),
.B(n_305),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_280),
.A2(n_313),
.B(n_277),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_364),
.A2(n_280),
.B(n_319),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_290),
.A2(n_292),
.B1(n_301),
.B2(n_326),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_365),
.A2(n_316),
.B1(n_294),
.B2(n_277),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_292),
.B(n_312),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_366),
.B(n_307),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_368),
.A2(n_371),
.B(n_379),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_372),
.B(n_357),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_L g410 ( 
.A1(n_374),
.A2(n_361),
.B1(n_330),
.B2(n_348),
.Y(n_410)
);

OAI32xp33_ASAP7_75t_L g375 ( 
.A1(n_352),
.A2(n_316),
.A3(n_307),
.B1(n_288),
.B2(n_303),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_375),
.B(n_392),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_360),
.A2(n_300),
.B(n_320),
.Y(n_379)
);

MAJx2_ASAP7_75t_L g380 ( 
.A(n_332),
.B(n_300),
.C(n_321),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_380),
.B(n_395),
.C(n_351),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_363),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_383),
.B(n_389),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_349),
.A2(n_289),
.B(n_319),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_386),
.A2(n_393),
.B(n_398),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_365),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_342),
.A2(n_317),
.B1(n_293),
.B2(n_320),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_337),
.A2(n_305),
.B(n_309),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_340),
.B(n_293),
.Y(n_395)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_396),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_336),
.B(n_281),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_397),
.B(n_366),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_333),
.A2(n_309),
.B(n_321),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_369),
.B(n_340),
.C(n_350),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_400),
.B(n_426),
.C(n_382),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_397),
.Y(n_402)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_402),
.Y(n_439)
);

OA21x2_ASAP7_75t_L g403 ( 
.A1(n_391),
.A2(n_362),
.B(n_357),
.Y(n_403)
);

INVx1_ASAP7_75t_SL g452 ( 
.A(n_403),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_396),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_L g453 ( 
.A1(n_406),
.A2(n_419),
.B1(n_420),
.B2(n_423),
.Y(n_453)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_407),
.Y(n_441)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_378),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_408),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_410),
.A2(n_421),
.B1(n_398),
.B2(n_384),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_371),
.A2(n_333),
.B(n_364),
.Y(n_411)
);

AOI21x1_ASAP7_75t_SL g436 ( 
.A1(n_411),
.A2(n_412),
.B(n_414),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_379),
.B(n_357),
.Y(n_412)
);

XNOR2x1_ASAP7_75t_L g429 ( 
.A(n_413),
.B(n_382),
.Y(n_429)
);

A2O1A1O1Ixp25_ASAP7_75t_L g414 ( 
.A1(n_391),
.A2(n_332),
.B(n_336),
.C(n_327),
.D(n_357),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_381),
.B(n_354),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_416),
.B(n_418),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g437 ( 
.A(n_417),
.B(n_370),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_367),
.A2(n_347),
.B(n_335),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_394),
.B(n_359),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_377),
.B(n_341),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_383),
.A2(n_317),
.B1(n_355),
.B2(n_281),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_380),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_422),
.B(n_424),
.Y(n_445)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_378),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_394),
.B(n_355),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_390),
.A2(n_355),
.B1(n_367),
.B2(n_389),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_425),
.A2(n_392),
.B1(n_373),
.B2(n_368),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_395),
.B(n_369),
.C(n_372),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_374),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g438 ( 
.A(n_427),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_429),
.B(n_437),
.Y(n_460)
);

INVx4_ASAP7_75t_L g430 ( 
.A(n_412),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_430),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_415),
.A2(n_390),
.B1(n_386),
.B2(n_388),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_432),
.B(n_433),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_415),
.A2(n_393),
.B1(n_377),
.B2(n_375),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_434),
.A2(n_442),
.B1(n_448),
.B2(n_405),
.Y(n_458)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_435),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_440),
.B(n_444),
.C(n_446),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_427),
.A2(n_376),
.B1(n_399),
.B2(n_387),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_416),
.A2(n_401),
.B1(n_376),
.B2(n_410),
.Y(n_443)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_443),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_400),
.B(n_387),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_400),
.B(n_399),
.C(n_385),
.Y(n_446)
);

XOR2x2_ASAP7_75t_L g447 ( 
.A(n_413),
.B(n_417),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_447),
.B(n_403),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_412),
.A2(n_385),
.B1(n_401),
.B2(n_425),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_426),
.B(n_407),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_449),
.B(n_451),
.C(n_412),
.Y(n_463)
);

FAx1_ASAP7_75t_SL g450 ( 
.A(n_414),
.B(n_406),
.CI(n_403),
.CON(n_450),
.SN(n_450)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_450),
.B(n_408),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_414),
.B(n_403),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_433),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_454),
.B(n_467),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_456),
.B(n_451),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_458),
.A2(n_452),
.B1(n_445),
.B2(n_450),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_439),
.B(n_424),
.Y(n_459)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_459),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_441),
.B(n_419),
.Y(n_461)
);

CKINVDCx14_ASAP7_75t_R g477 ( 
.A(n_461),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_428),
.A2(n_409),
.B(n_418),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_462),
.A2(n_466),
.B(n_472),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_463),
.B(n_444),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_452),
.A2(n_405),
.B1(n_404),
.B2(n_411),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_464),
.A2(n_473),
.B1(n_474),
.B2(n_432),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_430),
.A2(n_409),
.B(n_420),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_431),
.B(n_404),
.Y(n_467)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_431),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_469),
.B(n_470),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_442),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_453),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_438),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_475),
.B(n_484),
.Y(n_492)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_478),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_479),
.B(n_482),
.Y(n_494)
);

XNOR2x1_ASAP7_75t_L g482 ( 
.A(n_463),
.B(n_437),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_455),
.B(n_446),
.C(n_440),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_483),
.B(n_488),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_455),
.B(n_449),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_485),
.A2(n_436),
.B(n_465),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_456),
.B(n_429),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_487),
.B(n_489),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_462),
.A2(n_436),
.B(n_448),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_460),
.B(n_447),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_460),
.B(n_441),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_490),
.B(n_461),
.Y(n_498)
);

BUFx24_ASAP7_75t_SL g491 ( 
.A(n_476),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_491),
.B(n_499),
.Y(n_511)
);

INVx11_ASAP7_75t_L g496 ( 
.A(n_477),
.Y(n_496)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_496),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_498),
.B(n_501),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_486),
.B(n_454),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_480),
.A2(n_457),
.B1(n_468),
.B2(n_473),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_500),
.A2(n_478),
.B1(n_465),
.B2(n_485),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_483),
.B(n_468),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_502),
.B(n_503),
.Y(n_513)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_481),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_492),
.B(n_484),
.C(n_479),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_504),
.B(n_505),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_494),
.B(n_490),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_496),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_508),
.B(n_510),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_509),
.A2(n_514),
.B1(n_464),
.B2(n_500),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_492),
.B(n_487),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_494),
.B(n_489),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_512),
.B(n_482),
.C(n_497),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_495),
.A2(n_457),
.B1(n_472),
.B2(n_458),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_515),
.B(n_516),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_513),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_518),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_504),
.B(n_493),
.C(n_498),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_520),
.B(n_522),
.Y(n_524)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_506),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_521),
.B(n_469),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_514),
.A2(n_501),
.B(n_470),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_511),
.A2(n_471),
.B1(n_450),
.B2(n_475),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_523),
.B(n_507),
.C(n_510),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_526),
.B(n_528),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_520),
.B(n_507),
.C(n_505),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_529),
.B(n_530),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_517),
.B(n_512),
.C(n_474),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_SL g531 ( 
.A1(n_524),
.A2(n_519),
.B(n_522),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_531),
.A2(n_527),
.B(n_523),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_525),
.B(n_459),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_532),
.A2(n_518),
.B(n_497),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_535),
.A2(n_536),
.B(n_534),
.Y(n_537)
);

O2A1O1Ixp33_ASAP7_75t_SL g538 ( 
.A1(n_537),
.A2(n_533),
.B(n_467),
.C(n_423),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_538),
.B(n_421),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_539),
.B(n_434),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_540),
.B(n_466),
.Y(n_541)
);


endmodule