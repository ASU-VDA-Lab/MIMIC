module real_jpeg_6900_n_19 (n_17, n_123, n_8, n_116, n_0, n_2, n_125, n_10, n_9, n_12, n_124, n_6, n_121, n_11, n_14, n_7, n_117, n_18, n_3, n_119, n_5, n_4, n_122, n_1, n_118, n_16, n_15, n_13, n_120, n_19);

input n_17;
input n_123;
input n_8;
input n_116;
input n_0;
input n_2;
input n_125;
input n_10;
input n_9;
input n_12;
input n_124;
input n_6;
input n_121;
input n_11;
input n_14;
input n_7;
input n_117;
input n_18;
input n_3;
input n_119;
input n_5;
input n_4;
input n_122;
input n_1;
input n_118;
input n_16;
input n_15;
input n_13;
input n_120;

output n_19;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

INVx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_0),
.B(n_80),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_1),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_1),
.B(n_112),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_3),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_3),
.B(n_33),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_4),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_4),
.B(n_45),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_5),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_5),
.B(n_48),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_6),
.B(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_9),
.B(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_9),
.B(n_23),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_10),
.B(n_39),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_10),
.B(n_39),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_11),
.Y(n_81)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_12),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_13),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_13),
.B(n_97),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_14),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_15),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_16),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_16),
.B(n_84),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_17),
.B(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_17),
.B(n_57),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_18),
.B(n_60),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_18),
.B(n_60),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_29),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_28),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_25),
.B(n_70),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_25),
.B(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_25),
.B(n_113),
.Y(n_112)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_26),
.B(n_85),
.Y(n_84)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_114),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_52),
.B(n_102),
.C(n_111),
.Y(n_30)
);

NOR4xp25_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_38),
.C(n_44),
.D(n_47),
.Y(n_31)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_32),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_37),
.B(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_38),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_44),
.A2(n_106),
.B(n_107),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI21x1_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_96),
.B(n_101),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_91),
.B(n_95),
.Y(n_53)
);

AO221x1_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_66),
.B1(n_88),
.B2(n_89),
.C(n_90),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AO21x1_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_72),
.B(n_87),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_71),
.Y(n_87)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_83),
.B(n_86),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_77),
.B(n_82),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_81),
.Y(n_82)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_94),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_94),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

A2O1A1O1Ixp25_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B(n_108),
.C(n_109),
.D(n_110),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_116),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_117),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_118),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_119),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_120),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_121),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_122),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_123),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_124),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_125),
.Y(n_98)
);


endmodule