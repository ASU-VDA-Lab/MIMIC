module fake_jpeg_16113_n_168 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_168);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_5),
.B(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_34),
.B(n_22),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_36),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_24),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_19),
.B(n_1),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_20),
.B(n_19),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_26),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_43),
.A2(n_40),
.B(n_18),
.Y(n_59)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

AOI21xp33_ASAP7_75t_L g51 ( 
.A1(n_34),
.A2(n_40),
.B(n_26),
.Y(n_51)
);

AOI21xp33_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_23),
.B(n_17),
.Y(n_77)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_55),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_40),
.B(n_20),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_46),
.A2(n_36),
.B1(n_37),
.B2(n_22),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

XOR2x1_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_71),
.Y(n_90)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_46),
.A2(n_28),
.B1(n_21),
.B2(n_25),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_39),
.B1(n_33),
.B2(n_31),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_25),
.B1(n_32),
.B2(n_16),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_69),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_29),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_29),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_72),
.Y(n_99)
);

AO22x1_ASAP7_75t_L g71 ( 
.A1(n_43),
.A2(n_39),
.B1(n_33),
.B2(n_31),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_27),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_15),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_76),
.C(n_80),
.Y(n_91)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_15),
.Y(n_76)
);

FAx1_ASAP7_75t_SL g97 ( 
.A(n_77),
.B(n_79),
.CI(n_25),
.CON(n_97),
.SN(n_97)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_23),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_15),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_59),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_95),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_67),
.Y(n_101)
);

NOR3xp33_ASAP7_75t_SL g84 ( 
.A(n_68),
.B(n_25),
.C(n_17),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_16),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_100),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_57),
.B(n_2),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_101),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_90),
.A2(n_81),
.B(n_97),
.C(n_66),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_107),
.Y(n_130)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_74),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_58),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_108),
.A2(n_111),
.B(n_86),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_85),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_112),
.C(n_116),
.Y(n_118)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_65),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_56),
.C(n_73),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_115),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_61),
.Y(n_114)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_56),
.C(n_78),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_117),
.A2(n_108),
.B(n_111),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_107),
.C(n_112),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_126),
.C(n_132),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_105),
.B(n_84),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_102),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_99),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_110),
.A2(n_82),
.B1(n_86),
.B2(n_93),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_127),
.A2(n_101),
.B(n_3),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_108),
.A2(n_82),
.B1(n_95),
.B2(n_89),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_128),
.A2(n_122),
.B1(n_117),
.B2(n_132),
.Y(n_141)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_129),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_87),
.C(n_89),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_134),
.A2(n_137),
.B(n_142),
.Y(n_150)
);

AOI321xp33_ASAP7_75t_L g151 ( 
.A1(n_135),
.A2(n_121),
.A3(n_120),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_151)
);

OAI321xp33_ASAP7_75t_L g136 ( 
.A1(n_130),
.A2(n_101),
.A3(n_111),
.B1(n_62),
.B2(n_13),
.C(n_6),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_139),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_2),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_118),
.C(n_125),
.Y(n_146)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_126),
.B(n_10),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_143),
.B(n_118),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_151),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_148),
.C(n_149),
.Y(n_157)
);

XNOR2x1_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_130),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_143),
.B(n_131),
.C(n_128),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_131),
.C(n_121),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_144),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_147),
.A2(n_139),
.B1(n_133),
.B2(n_140),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_154),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_150),
.A2(n_135),
.B(n_133),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

OAI321xp33_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_146),
.A3(n_145),
.B1(n_124),
.B2(n_8),
.C(n_4),
.Y(n_160)
);

OAI211xp5_ASAP7_75t_L g163 ( 
.A1(n_160),
.A2(n_4),
.B(n_7),
.C(n_9),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_158),
.A2(n_156),
.B1(n_157),
.B2(n_153),
.Y(n_161)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_161),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_4),
.C(n_5),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_162),
.B(n_163),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_165),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_164),
.B(n_161),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_7),
.Y(n_168)
);


endmodule