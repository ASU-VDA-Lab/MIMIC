module real_jpeg_4944_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_1),
.A2(n_60),
.B1(n_61),
.B2(n_63),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_1),
.A2(n_176),
.B1(n_178),
.B2(n_179),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_1),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_2),
.A2(n_22),
.B1(n_26),
.B2(n_27),
.Y(n_21)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_2),
.A2(n_26),
.B1(n_75),
.B2(n_77),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_2),
.A2(n_26),
.B1(n_82),
.B2(n_86),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_2),
.A2(n_26),
.B1(n_116),
.B2(n_119),
.Y(n_115)
);

O2A1O1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_2),
.A2(n_201),
.B(n_204),
.C(n_207),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_2),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_2),
.B(n_41),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_2),
.B(n_246),
.C(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_2),
.B(n_255),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_2),
.B(n_107),
.C(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_2),
.B(n_121),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_3),
.A2(n_156),
.B1(n_160),
.B2(n_161),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_3),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_4),
.A2(n_40),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_4),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_4),
.A2(n_51),
.B1(n_119),
.B2(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_4),
.A2(n_51),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_4),
.A2(n_51),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_5),
.Y(n_159)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_6),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_7),
.Y(n_72)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_7),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_7),
.Y(n_217)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_8),
.Y(n_124)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_8),
.Y(n_130)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_8),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_8),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g206 ( 
.A(n_8),
.Y(n_206)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_9),
.Y(n_85)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_10),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_10),
.Y(n_119)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_10),
.Y(n_129)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_10),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_10),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_11),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_220),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_218),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_189),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_15),
.B(n_189),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_138),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_79),
.C(n_114),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_18),
.B(n_192),
.Y(n_191)
);

NOR2xp67_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_55),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_19),
.A2(n_240),
.B1(n_241),
.B2(n_248),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_19),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_19),
.A2(n_142),
.B1(n_143),
.B2(n_240),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_19),
.A2(n_55),
.B1(n_240),
.B2(n_312),
.Y(n_311)
);

AND2x2_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_49),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_20),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_30),
.Y(n_20)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_21),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_21),
.B(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_22),
.Y(n_177)
);

INVx4_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_24),
.Y(n_107)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_25),
.Y(n_111)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_25),
.Y(n_181)
);

OAI21xp33_ASAP7_75t_L g204 ( 
.A1(n_26),
.A2(n_82),
.B(n_205),
.Y(n_204)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_30),
.Y(n_169)
);

NOR2x1_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_41),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_34),
.B1(n_37),
.B2(n_39),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AO22x1_ASAP7_75t_SL g41 ( 
.A1(n_37),
.A2(n_42),
.B1(n_44),
.B2(n_47),
.Y(n_41)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_41),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_41),
.A2(n_175),
.B(n_182),
.Y(n_174)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_43),
.Y(n_214)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_50),
.Y(n_168)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_55),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_59),
.B(n_64),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_57),
.A2(n_66),
.B1(n_74),
.B2(n_210),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_59),
.Y(n_153)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_63),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_73),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_65),
.A2(n_153),
.B1(n_154),
.B2(n_163),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_65),
.B(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_66),
.A2(n_74),
.B1(n_210),
.B2(n_215),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_72),
.Y(n_187)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_72),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_74),
.B(n_184),
.Y(n_270)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_76),
.Y(n_162)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_76),
.Y(n_211)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_79),
.A2(n_114),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_79),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_90),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_81),
.A2(n_91),
.B1(n_105),
.B2(n_144),
.Y(n_143)
);

OA22x2_ASAP7_75t_L g198 ( 
.A1(n_81),
.A2(n_91),
.B1(n_105),
.B2(n_144),
.Y(n_198)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_105),
.Y(n_90)
);

NAND2x1_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_105),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_98),
.B1(n_100),
.B2(n_103),
.Y(n_92)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx6_ASAP7_75t_L g269 ( 
.A(n_102),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_105),
.Y(n_255)
);

AOI22x1_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_108),
.B1(n_110),
.B2(n_112),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_114),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_114),
.A2(n_193),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_114),
.B(n_143),
.C(n_295),
.Y(n_313)
);

OA22x2_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_120),
.B1(n_134),
.B2(n_137),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_120),
.B1(n_134),
.B2(n_137),
.Y(n_141)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_119),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_127),
.Y(n_120)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_121)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_172),
.Y(n_138)
);

XNOR2x1_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_151),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_150),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_141),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_141),
.B(n_198),
.C(n_199),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_141),
.A2(n_150),
.B1(n_198),
.B2(n_285),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_142),
.B(n_240),
.C(n_262),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_142),
.A2(n_143),
.B1(n_295),
.B2(n_297),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_149),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_166),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_152),
.A2(n_166),
.B1(n_167),
.B2(n_196),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_184),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_161),
.Y(n_247)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_166),
.A2(n_167),
.B1(n_254),
.B2(n_256),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_166),
.A2(n_167),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_167),
.B(n_209),
.C(n_254),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_167),
.B(n_277),
.C(n_279),
.Y(n_290)
);

OA22x2_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_169),
.B(n_170),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_183),
.B2(n_188),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_181),
.Y(n_244)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_195),
.C(n_197),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_190),
.A2(n_191),
.B1(n_195),
.B2(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_195),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_197),
.B(n_319),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_198),
.A2(n_281),
.B1(n_282),
.B2(n_285),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_198),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_199),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_208),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_200),
.A2(n_208),
.B1(n_209),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_200),
.Y(n_303)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_SL g205 ( 
.A(n_206),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_208),
.A2(n_209),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_235),
.Y(n_236)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_305),
.B(n_321),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_289),
.B(n_304),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_274),
.B(n_288),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_259),
.B(n_273),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_250),
.B(n_258),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_237),
.B(n_249),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_234),
.B(n_236),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_233),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_233),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_233),
.A2(n_238),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_239),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_238),
.B(n_283),
.C(n_285),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_248),
.Y(n_257)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_241),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_257),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_257),
.Y(n_258)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_254),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_261),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_272),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_270),
.B2(n_271),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_271),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_268),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_270),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_287),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_287),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_279),
.B1(n_280),
.B2(n_286),
.Y(n_275)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_276),
.Y(n_286)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_277),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_291),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_298),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_292),
.B(n_300),
.C(n_301),
.Y(n_314)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_295),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_301),
.B2(n_302),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NOR2x1_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_315),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_314),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_307),
.B(n_314),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_310),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_308),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_313),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_313),
.C(n_317),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_315),
.A2(n_322),
.B(n_323),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_318),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_318),
.Y(n_323)
);


endmodule