module fake_jpeg_11301_n_144 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_144);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_7),
.B(n_12),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_25),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_32),
.Y(n_46)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_8),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

NAND2x1p5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_0),
.Y(n_34)
);

HAxp5_ASAP7_75t_SL g59 ( 
.A(n_34),
.B(n_1),
.CON(n_59),
.SN(n_59)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_3),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_41),
.Y(n_48)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_13),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_42),
.B(n_20),
.Y(n_44)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_17),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_44),
.B(n_51),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_27),
.B1(n_17),
.B2(n_22),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_45),
.A2(n_28),
.B1(n_21),
.B2(n_19),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_27),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_20),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_22),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_30),
.B(n_28),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_55),
.B(n_52),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_59),
.A2(n_33),
.B1(n_39),
.B2(n_36),
.Y(n_67)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_68),
.Y(n_88)
);

BUFx24_ASAP7_75t_SL g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_63),
.B(n_69),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVxp33_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_54),
.A2(n_31),
.B1(n_41),
.B2(n_40),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_66),
.A2(n_83),
.B1(n_60),
.B2(n_61),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_80),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_16),
.Y(n_69)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_74),
.Y(n_96)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_21),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_76),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_33),
.C(n_37),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_81),
.C(n_67),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_78),
.A2(n_82),
.B1(n_61),
.B2(n_60),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_19),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_70),
.Y(n_84)
);

MAJx2_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_16),
.C(n_2),
.Y(n_81)
);

INVx3_ASAP7_75t_SL g82 ( 
.A(n_56),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_58),
.A2(n_3),
.B1(n_9),
.B2(n_10),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_87),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g85 ( 
.A(n_77),
.B(n_9),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_90),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_86),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_78),
.A2(n_60),
.B1(n_61),
.B2(n_56),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_91),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_11),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_64),
.A2(n_11),
.B1(n_67),
.B2(n_73),
.Y(n_91)
);

O2A1O1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_67),
.A2(n_64),
.B(n_65),
.C(n_68),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_95),
.A2(n_94),
.B(n_86),
.C(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_99),
.Y(n_108)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_104),
.Y(n_117)
);

AO22x1_ASAP7_75t_L g104 ( 
.A1(n_94),
.A2(n_71),
.B1(n_82),
.B2(n_76),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_109),
.Y(n_115)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_111),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_99),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_114),
.C(n_116),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_85),
.C(n_90),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_84),
.C(n_92),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_121),
.B(n_123),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_95),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_122),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_105),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_117),
.A2(n_107),
.B1(n_103),
.B2(n_106),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_124),
.A2(n_127),
.B1(n_106),
.B2(n_100),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_100),
.Y(n_126)
);

OA21x2_ASAP7_75t_SL g132 ( 
.A1(n_126),
.A2(n_128),
.B(n_103),
.Y(n_132)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_118),
.Y(n_128)
);

AOI31xp67_ASAP7_75t_L g135 ( 
.A1(n_129),
.A2(n_132),
.A3(n_104),
.B(n_133),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_125),
.B(n_112),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_125),
.C(n_116),
.Y(n_134)
);

NOR2x1_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_135),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_114),
.C(n_101),
.Y(n_136)
);

NOR2xp67_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_124),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_138),
.B(n_122),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_121),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_139),
.A2(n_140),
.B(n_129),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_92),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_93),
.Y(n_144)
);


endmodule