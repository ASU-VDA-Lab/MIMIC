module fake_netlist_1_6365_n_1265 (n_117, n_219, n_44, n_133, n_149, n_289, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_292, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_291, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_283, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_145, n_270, n_246, n_153, n_61, n_259, n_290, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1265);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_289;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_292;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_291;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_283;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1265;
wire n_963;
wire n_1034;
wire n_949;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_830;
wire n_1112;
wire n_517;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_673;
wire n_1071;
wire n_1079;
wire n_409;
wire n_315;
wire n_295;
wire n_677;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_1246;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_293;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_867;
wire n_1070;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_366;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_427;
wire n_703;
wire n_415;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1043;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_385;
wire n_1127;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_303;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_948;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_639;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_335;
wire n_700;
wire n_534;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
INVx1_ASAP7_75t_L g293 ( .A(n_202), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_215), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_85), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_44), .Y(n_296) );
AND2x4_ASAP7_75t_L g297 ( .A(n_87), .B(n_237), .Y(n_297) );
INVxp67_ASAP7_75t_SL g298 ( .A(n_94), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_7), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_26), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_52), .Y(n_301) );
INVxp33_ASAP7_75t_SL g302 ( .A(n_96), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_122), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_72), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_275), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_274), .Y(n_306) );
INVxp67_ASAP7_75t_SL g307 ( .A(n_253), .Y(n_307) );
INVxp67_ASAP7_75t_L g308 ( .A(n_19), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_286), .Y(n_309) );
CKINVDCx16_ASAP7_75t_R g310 ( .A(n_153), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_164), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_71), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_70), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_58), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_2), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_238), .Y(n_316) );
INVxp67_ASAP7_75t_SL g317 ( .A(n_133), .Y(n_317) );
INVxp67_ASAP7_75t_L g318 ( .A(n_211), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_262), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_292), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_278), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_170), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_201), .Y(n_323) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_219), .Y(n_324) );
CKINVDCx20_ASAP7_75t_R g325 ( .A(n_176), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_214), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_146), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_142), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_12), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_150), .Y(n_330) );
INVxp67_ASAP7_75t_SL g331 ( .A(n_224), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_79), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_216), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_130), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_198), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_177), .Y(n_336) );
NOR2xp67_ASAP7_75t_L g337 ( .A(n_149), .B(n_37), .Y(n_337) );
INVxp33_ASAP7_75t_SL g338 ( .A(n_279), .Y(n_338) );
CKINVDCx20_ASAP7_75t_R g339 ( .A(n_99), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_4), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_131), .Y(n_341) );
CKINVDCx16_ASAP7_75t_R g342 ( .A(n_123), .Y(n_342) );
BUFx3_ASAP7_75t_L g343 ( .A(n_20), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_30), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_108), .Y(n_345) );
INVxp67_ASAP7_75t_SL g346 ( .A(n_50), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_55), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_183), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_140), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_111), .Y(n_350) );
INVxp33_ASAP7_75t_L g351 ( .A(n_228), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_241), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_47), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_163), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_250), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_185), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_103), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_234), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_247), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_34), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_48), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_19), .Y(n_362) );
NOR2xp67_ASAP7_75t_L g363 ( .A(n_13), .B(n_263), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_1), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_116), .Y(n_365) );
CKINVDCx5p33_ASAP7_75t_R g366 ( .A(n_287), .Y(n_366) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_191), .Y(n_367) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_268), .Y(n_368) );
INVxp33_ASAP7_75t_L g369 ( .A(n_252), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_233), .Y(n_370) );
INVx1_ASAP7_75t_SL g371 ( .A(n_217), .Y(n_371) );
INVxp33_ASAP7_75t_L g372 ( .A(n_244), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_239), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_132), .Y(n_374) );
BUFx6f_ASAP7_75t_L g375 ( .A(n_281), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_88), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_209), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_161), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_222), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_193), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_169), .Y(n_381) );
INVx3_ASAP7_75t_L g382 ( .A(n_102), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_76), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_256), .Y(n_384) );
INVxp33_ASAP7_75t_SL g385 ( .A(n_226), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_255), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_89), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_83), .Y(n_388) );
BUFx2_ASAP7_75t_L g389 ( .A(n_151), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_49), .Y(n_390) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_156), .Y(n_391) );
BUFx3_ASAP7_75t_L g392 ( .A(n_288), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_115), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g394 ( .A(n_2), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_54), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_186), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_276), .Y(n_397) );
INVxp33_ASAP7_75t_L g398 ( .A(n_27), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_189), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_97), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_10), .Y(n_401) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_157), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_20), .Y(n_403) );
CKINVDCx20_ASAP7_75t_R g404 ( .A(n_154), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_40), .Y(n_405) );
INVxp33_ASAP7_75t_SL g406 ( .A(n_37), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_155), .Y(n_407) );
XOR2x2_ASAP7_75t_L g408 ( .A(n_68), .B(n_44), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_1), .Y(n_409) );
CKINVDCx16_ASAP7_75t_R g410 ( .A(n_28), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_178), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_46), .Y(n_412) );
INVxp67_ASAP7_75t_L g413 ( .A(n_175), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_28), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_134), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_167), .Y(n_416) );
CKINVDCx14_ASAP7_75t_R g417 ( .A(n_264), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_70), .Y(n_418) );
CKINVDCx16_ASAP7_75t_R g419 ( .A(n_14), .Y(n_419) );
INVxp67_ASAP7_75t_L g420 ( .A(n_197), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_42), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_194), .Y(n_422) );
INVxp67_ASAP7_75t_SL g423 ( .A(n_15), .Y(n_423) );
INVxp67_ASAP7_75t_L g424 ( .A(n_81), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_114), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_66), .Y(n_426) );
CKINVDCx5p33_ASAP7_75t_R g427 ( .A(n_61), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_229), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_98), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_128), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_173), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_259), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_195), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_93), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_204), .Y(n_435) );
BUFx3_ASAP7_75t_L g436 ( .A(n_242), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_138), .Y(n_437) );
INVxp33_ASAP7_75t_L g438 ( .A(n_230), .Y(n_438) );
BUFx3_ASAP7_75t_L g439 ( .A(n_152), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_323), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_382), .Y(n_441) );
OA21x2_ASAP7_75t_L g442 ( .A1(n_323), .A2(n_78), .B(n_77), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_382), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_389), .B(n_0), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_382), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_375), .Y(n_446) );
AND2x4_ASAP7_75t_L g447 ( .A(n_389), .B(n_0), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_324), .B(n_3), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_375), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_367), .B(n_3), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_327), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_375), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_327), .Y(n_453) );
OAI22xp5_ASAP7_75t_SL g454 ( .A1(n_410), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_375), .B(n_5), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_375), .Y(n_456) );
CKINVDCx5p33_ASAP7_75t_R g457 ( .A(n_310), .Y(n_457) );
OA21x2_ASAP7_75t_L g458 ( .A1(n_328), .A2(n_82), .B(n_80), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_419), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_368), .B(n_8), .Y(n_460) );
CKINVDCx5p33_ASAP7_75t_R g461 ( .A(n_342), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_398), .B(n_9), .Y(n_462) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_402), .Y(n_463) );
OAI22xp33_ASAP7_75t_R g464 ( .A1(n_346), .A2(n_423), .B1(n_408), .B2(n_329), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_328), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_398), .B(n_9), .Y(n_466) );
CKINVDCx16_ASAP7_75t_R g467 ( .A(n_417), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_330), .Y(n_468) );
NOR2x1_ASAP7_75t_L g469 ( .A(n_343), .B(n_10), .Y(n_469) );
CKINVDCx5p33_ASAP7_75t_R g470 ( .A(n_325), .Y(n_470) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_343), .Y(n_471) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_402), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_330), .Y(n_473) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_402), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_402), .Y(n_475) );
BUFx10_ASAP7_75t_L g476 ( .A(n_447), .Y(n_476) );
INVx4_ASAP7_75t_L g477 ( .A(n_447), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_467), .B(n_351), .Y(n_478) );
INVx2_ASAP7_75t_SL g479 ( .A(n_471), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_466), .A2(n_329), .B1(n_299), .B2(n_300), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_441), .Y(n_481) );
BUFx3_ASAP7_75t_L g482 ( .A(n_441), .Y(n_482) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_474), .Y(n_483) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_474), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_467), .B(n_297), .Y(n_485) );
INVx4_ASAP7_75t_SL g486 ( .A(n_447), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_463), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_447), .B(n_297), .Y(n_488) );
CKINVDCx16_ASAP7_75t_R g489 ( .A(n_466), .Y(n_489) );
CKINVDCx5p33_ASAP7_75t_R g490 ( .A(n_470), .Y(n_490) );
INVxp67_ASAP7_75t_SL g491 ( .A(n_471), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_441), .Y(n_492) );
BUFx6f_ASAP7_75t_L g493 ( .A(n_474), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_463), .Y(n_494) );
BUFx6f_ASAP7_75t_L g495 ( .A(n_474), .Y(n_495) );
NAND3x1_ASAP7_75t_L g496 ( .A(n_444), .B(n_408), .C(n_301), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_444), .B(n_351), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_444), .B(n_369), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_443), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_443), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_440), .B(n_369), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_440), .B(n_372), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_463), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_451), .B(n_297), .Y(n_504) );
INVx4_ASAP7_75t_L g505 ( .A(n_442), .Y(n_505) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_466), .Y(n_506) );
INVx4_ASAP7_75t_L g507 ( .A(n_442), .Y(n_507) );
INVx4_ASAP7_75t_L g508 ( .A(n_442), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_463), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_462), .B(n_340), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_443), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_462), .A2(n_304), .B1(n_312), .B2(n_296), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_451), .B(n_372), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_463), .Y(n_514) );
OAI221xp5_ASAP7_75t_L g515 ( .A1(n_453), .A2(n_308), .B1(n_347), .B2(n_353), .C(n_313), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_445), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_453), .B(n_438), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_465), .B(n_295), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_463), .Y(n_519) );
BUFx10_ASAP7_75t_L g520 ( .A(n_457), .Y(n_520) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_474), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_472), .Y(n_522) );
INVx3_ASAP7_75t_L g523 ( .A(n_445), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_489), .A2(n_464), .B1(n_461), .B2(n_448), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_477), .A2(n_473), .B1(n_468), .B2(n_445), .Y(n_525) );
BUFx4f_ASAP7_75t_L g526 ( .A(n_479), .Y(n_526) );
CKINVDCx8_ASAP7_75t_R g527 ( .A(n_490), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_486), .B(n_476), .Y(n_528) );
NOR2x2_ASAP7_75t_L g529 ( .A(n_496), .B(n_464), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_477), .A2(n_473), .B1(n_468), .B2(n_454), .Y(n_530) );
INVx1_ASAP7_75t_SL g531 ( .A(n_510), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_498), .B(n_450), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_506), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_482), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_501), .B(n_460), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_489), .A2(n_406), .B1(n_454), .B2(n_339), .Y(n_536) );
INVx4_ASAP7_75t_L g537 ( .A(n_486), .Y(n_537) );
INVx3_ASAP7_75t_L g538 ( .A(n_477), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_481), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_502), .B(n_295), .Y(n_540) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_486), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_481), .Y(n_542) );
INVxp67_ASAP7_75t_SL g543 ( .A(n_497), .Y(n_543) );
INVxp67_ASAP7_75t_L g544 ( .A(n_510), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_482), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_477), .A2(n_406), .B1(n_469), .B2(n_364), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_492), .Y(n_547) );
NOR2xp67_ASAP7_75t_L g548 ( .A(n_515), .B(n_459), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_488), .A2(n_458), .B(n_442), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_497), .B(n_340), .Y(n_550) );
NOR2xp33_ASAP7_75t_R g551 ( .A(n_520), .B(n_325), .Y(n_551) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_486), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_486), .B(n_320), .Y(n_553) );
INVx5_ASAP7_75t_L g554 ( .A(n_476), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_492), .A2(n_469), .B1(n_383), .B2(n_395), .Y(n_555) );
INVx5_ASAP7_75t_L g556 ( .A(n_476), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_485), .B(n_302), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_491), .B(n_361), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_476), .B(n_320), .Y(n_559) );
INVx3_ASAP7_75t_L g560 ( .A(n_523), .Y(n_560) );
OAI22xp5_ASAP7_75t_SL g561 ( .A1(n_496), .A2(n_459), .B1(n_404), .B2(n_339), .Y(n_561) );
AND2x6_ASAP7_75t_SL g562 ( .A(n_478), .B(n_362), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_523), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_513), .B(n_302), .Y(n_564) );
INVxp67_ASAP7_75t_L g565 ( .A(n_518), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_499), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_523), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_523), .Y(n_568) );
INVx5_ASAP7_75t_L g569 ( .A(n_483), .Y(n_569) );
INVx4_ASAP7_75t_L g570 ( .A(n_520), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_499), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_480), .B(n_345), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_500), .A2(n_403), .B1(n_405), .B2(n_401), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_500), .Y(n_574) );
XOR2xp5_ASAP7_75t_L g575 ( .A(n_512), .B(n_404), .Y(n_575) );
NOR2xp67_ASAP7_75t_L g576 ( .A(n_504), .B(n_345), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_511), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_517), .B(n_352), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_520), .B(n_352), .Y(n_579) );
INVxp67_ASAP7_75t_L g580 ( .A(n_511), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_516), .B(n_338), .Y(n_581) );
INVx4_ASAP7_75t_L g582 ( .A(n_516), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_505), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_505), .A2(n_361), .B1(n_394), .B2(n_390), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_505), .A2(n_394), .B1(n_409), .B2(n_390), .Y(n_585) );
INVxp67_ASAP7_75t_L g586 ( .A(n_487), .Y(n_586) );
BUFx2_ASAP7_75t_L g587 ( .A(n_505), .Y(n_587) );
NAND2x1p5_ASAP7_75t_L g588 ( .A(n_507), .B(n_412), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_507), .Y(n_589) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_507), .A2(n_421), .B1(n_427), .B2(n_409), .Y(n_590) );
INVx2_ASAP7_75t_SL g591 ( .A(n_507), .Y(n_591) );
INVx2_ASAP7_75t_SL g592 ( .A(n_508), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_508), .B(n_366), .Y(n_593) );
AND2x2_ASAP7_75t_SL g594 ( .A(n_508), .B(n_442), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_487), .B(n_366), .Y(n_595) );
INVx1_ASAP7_75t_SL g596 ( .A(n_487), .Y(n_596) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_483), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_522), .B(n_338), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g599 ( .A1(n_494), .A2(n_458), .B(n_455), .Y(n_599) );
AND2x6_ASAP7_75t_SL g600 ( .A(n_494), .B(n_414), .Y(n_600) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_483), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_503), .B(n_418), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_503), .B(n_381), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_509), .B(n_381), .Y(n_604) );
OAI21xp5_ASAP7_75t_L g605 ( .A1(n_509), .A2(n_458), .B(n_434), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_509), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_514), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_514), .Y(n_608) );
BUFx12f_ASAP7_75t_L g609 ( .A(n_483), .Y(n_609) );
BUFx6f_ASAP7_75t_L g610 ( .A(n_483), .Y(n_610) );
OR2x2_ASAP7_75t_SL g611 ( .A(n_514), .B(n_458), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_519), .B(n_426), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_519), .B(n_391), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_519), .B(n_314), .Y(n_614) );
NAND2xp5_ASAP7_75t_SL g615 ( .A(n_483), .B(n_391), .Y(n_615) );
NOR3xp33_ASAP7_75t_L g616 ( .A(n_561), .B(n_413), .C(n_318), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_531), .B(n_314), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_582), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_544), .B(n_315), .Y(n_619) );
INVx2_ASAP7_75t_SL g620 ( .A(n_526), .Y(n_620) );
BUFx6f_ASAP7_75t_L g621 ( .A(n_554), .Y(n_621) );
INVx2_ASAP7_75t_SL g622 ( .A(n_526), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_582), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_589), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_583), .Y(n_625) );
O2A1O1Ixp33_ASAP7_75t_L g626 ( .A1(n_543), .A2(n_344), .B(n_360), .C(n_315), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_591), .A2(n_307), .B(n_298), .Y(n_627) );
AND2x4_ASAP7_75t_SL g628 ( .A(n_570), .B(n_344), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_543), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_548), .A2(n_385), .B1(n_360), .B2(n_434), .Y(n_630) );
AND2x4_ASAP7_75t_L g631 ( .A(n_565), .B(n_337), .Y(n_631) );
NOR2xp33_ASAP7_75t_SL g632 ( .A(n_537), .B(n_385), .Y(n_632) );
AOI21xp5_ASAP7_75t_L g633 ( .A1(n_549), .A2(n_594), .B(n_593), .Y(n_633) );
AOI21xp5_ASAP7_75t_SL g634 ( .A1(n_537), .A2(n_331), .B(n_317), .Y(n_634) );
BUFx3_ASAP7_75t_L g635 ( .A(n_527), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_580), .B(n_433), .Y(n_636) );
BUFx2_ASAP7_75t_L g637 ( .A(n_551), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_550), .B(n_433), .Y(n_638) );
A2O1A1Ixp33_ASAP7_75t_L g639 ( .A1(n_581), .A2(n_363), .B(n_294), .C(n_303), .Y(n_639) );
BUFx6f_ASAP7_75t_L g640 ( .A(n_554), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_538), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_533), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_525), .B(n_293), .Y(n_643) );
AOI21xp5_ASAP7_75t_L g644 ( .A1(n_549), .A2(n_306), .B(n_305), .Y(n_644) );
INVx3_ASAP7_75t_L g645 ( .A(n_554), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_530), .A2(n_311), .B1(n_316), .B2(n_309), .Y(n_646) );
INVx3_ASAP7_75t_L g647 ( .A(n_554), .Y(n_647) );
A2O1A1Ixp33_ASAP7_75t_L g648 ( .A1(n_581), .A2(n_321), .B(n_332), .C(n_319), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_530), .A2(n_334), .B1(n_336), .B2(n_333), .Y(n_649) );
INVx1_ASAP7_75t_SL g650 ( .A(n_556), .Y(n_650) );
O2A1O1Ixp33_ASAP7_75t_L g651 ( .A1(n_532), .A2(n_424), .B(n_420), .C(n_348), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_538), .Y(n_652) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_558), .Y(n_653) );
OAI22xp33_ASAP7_75t_L g654 ( .A1(n_536), .A2(n_349), .B1(n_350), .B2(n_341), .Y(n_654) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_594), .A2(n_355), .B(n_354), .Y(n_655) );
O2A1O1Ixp33_ASAP7_75t_SL g656 ( .A1(n_592), .A2(n_357), .B(n_359), .C(n_356), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_539), .Y(n_657) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_587), .A2(n_370), .B(n_365), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_535), .B(n_11), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_525), .B(n_373), .Y(n_660) );
O2A1O1Ixp33_ASAP7_75t_L g661 ( .A1(n_572), .A2(n_377), .B(n_378), .C(n_374), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_546), .B(n_379), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_534), .Y(n_663) );
NAND2xp33_ASAP7_75t_L g664 ( .A(n_556), .B(n_402), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_542), .Y(n_665) );
BUFx6f_ASAP7_75t_L g666 ( .A(n_556), .Y(n_666) );
AOI21xp5_ASAP7_75t_L g667 ( .A1(n_528), .A2(n_522), .B(n_384), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_546), .A2(n_386), .B1(n_387), .B2(n_380), .Y(n_668) );
INVxp67_ASAP7_75t_SL g669 ( .A(n_588), .Y(n_669) );
O2A1O1Ixp33_ASAP7_75t_L g670 ( .A1(n_540), .A2(n_393), .B(n_396), .C(n_388), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_547), .Y(n_671) );
NOR2x1_ASAP7_75t_L g672 ( .A(n_579), .B(n_397), .Y(n_672) );
AOI222xp33_ASAP7_75t_L g673 ( .A1(n_529), .A2(n_425), .B1(n_429), .B2(n_437), .C1(n_428), .C2(n_431), .Y(n_673) );
BUFx12f_ASAP7_75t_L g674 ( .A(n_562), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_566), .Y(n_675) );
INVx4_ASAP7_75t_L g676 ( .A(n_556), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_557), .B(n_371), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_571), .Y(n_678) );
INVx4_ASAP7_75t_L g679 ( .A(n_609), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_577), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_574), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_545), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_602), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_573), .A2(n_400), .B1(n_407), .B2(n_399), .Y(n_684) );
BUFx2_ASAP7_75t_L g685 ( .A(n_600), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_612), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_588), .Y(n_687) );
NAND2xp5_ASAP7_75t_SL g688 ( .A(n_541), .B(n_552), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_560), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_560), .Y(n_690) );
AOI22xp33_ASAP7_75t_SL g691 ( .A1(n_557), .A2(n_436), .B1(n_439), .B2(n_392), .Y(n_691) );
BUFx12f_ASAP7_75t_L g692 ( .A(n_614), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_563), .Y(n_693) );
AOI21xp5_ASAP7_75t_L g694 ( .A1(n_605), .A2(n_416), .B(n_411), .Y(n_694) );
BUFx3_ASAP7_75t_L g695 ( .A(n_567), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_568), .Y(n_696) );
AOI21x1_ASAP7_75t_L g697 ( .A1(n_599), .A2(n_522), .B(n_432), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_565), .B(n_524), .Y(n_698) );
BUFx4f_ASAP7_75t_SL g699 ( .A(n_578), .Y(n_699) );
BUFx6f_ASAP7_75t_L g700 ( .A(n_569), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_564), .A2(n_435), .B1(n_422), .B2(n_326), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_584), .Y(n_702) );
BUFx3_ASAP7_75t_L g703 ( .A(n_585), .Y(n_703) );
BUFx8_ASAP7_75t_L g704 ( .A(n_606), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_590), .B(n_11), .Y(n_705) );
NAND2x1p5_ASAP7_75t_L g706 ( .A(n_559), .B(n_439), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_541), .Y(n_707) );
CKINVDCx5p33_ASAP7_75t_R g708 ( .A(n_573), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_576), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_598), .Y(n_710) );
A2O1A1Ixp33_ASAP7_75t_L g711 ( .A1(n_598), .A2(n_326), .B(n_335), .C(n_322), .Y(n_711) );
AND3x1_ASAP7_75t_L g712 ( .A(n_555), .B(n_335), .C(n_322), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_555), .A2(n_358), .B1(n_376), .B2(n_415), .Y(n_713) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_552), .Y(n_714) );
INVx4_ASAP7_75t_L g715 ( .A(n_569), .Y(n_715) );
NOR3xp33_ASAP7_75t_L g716 ( .A(n_553), .B(n_376), .C(n_358), .Y(n_716) );
OAI22xp5_ASAP7_75t_SL g717 ( .A1(n_611), .A2(n_430), .B1(n_415), .B2(n_595), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_615), .A2(n_430), .B1(n_446), .B2(n_449), .Y(n_718) );
A2O1A1Ixp33_ASAP7_75t_L g719 ( .A1(n_599), .A2(n_446), .B(n_449), .C(n_452), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_603), .B(n_12), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_604), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_613), .Y(n_722) );
OR2x6_ASAP7_75t_L g723 ( .A(n_586), .B(n_446), .Y(n_723) );
BUFx2_ASAP7_75t_SL g724 ( .A(n_569), .Y(n_724) );
INVx2_ASAP7_75t_L g725 ( .A(n_607), .Y(n_725) );
BUFx6f_ASAP7_75t_L g726 ( .A(n_569), .Y(n_726) );
BUFx6f_ASAP7_75t_L g727 ( .A(n_597), .Y(n_727) );
INVx2_ASAP7_75t_SL g728 ( .A(n_608), .Y(n_728) );
OAI21xp33_ASAP7_75t_L g729 ( .A1(n_586), .A2(n_452), .B(n_449), .Y(n_729) );
AND2x2_ASAP7_75t_L g730 ( .A(n_596), .B(n_13), .Y(n_730) );
INVx3_ASAP7_75t_L g731 ( .A(n_597), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_601), .B(n_452), .Y(n_732) );
INVx4_ASAP7_75t_L g733 ( .A(n_601), .Y(n_733) );
OR2x2_ASAP7_75t_L g734 ( .A(n_601), .B(n_14), .Y(n_734) );
BUFx6f_ASAP7_75t_L g735 ( .A(n_610), .Y(n_735) );
O2A1O1Ixp33_ASAP7_75t_L g736 ( .A1(n_610), .A2(n_456), .B(n_475), .C(n_17), .Y(n_736) );
NAND2xp33_ASAP7_75t_L g737 ( .A(n_554), .B(n_472), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_582), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_531), .A2(n_475), .B1(n_456), .B2(n_472), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_544), .B(n_456), .Y(n_740) );
AOI221xp5_ASAP7_75t_L g741 ( .A1(n_543), .A2(n_475), .B1(n_472), .B2(n_474), .C(n_484), .Y(n_741) );
OR2x6_ASAP7_75t_SL g742 ( .A(n_551), .B(n_15), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_544), .B(n_16), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_544), .B(n_16), .Y(n_744) );
AND2x2_ASAP7_75t_L g745 ( .A(n_531), .B(n_17), .Y(n_745) );
INVx2_ASAP7_75t_SL g746 ( .A(n_526), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_582), .Y(n_747) );
NAND2x2_ASAP7_75t_L g748 ( .A(n_529), .B(n_18), .Y(n_748) );
INVx2_ASAP7_75t_L g749 ( .A(n_582), .Y(n_749) );
CKINVDCx14_ASAP7_75t_R g750 ( .A(n_742), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_642), .Y(n_751) );
OAI22xp33_ASAP7_75t_L g752 ( .A1(n_708), .A2(n_472), .B1(n_474), .B2(n_22), .Y(n_752) );
HB1xp67_ASAP7_75t_L g753 ( .A(n_621), .Y(n_753) );
O2A1O1Ixp33_ASAP7_75t_L g754 ( .A1(n_639), .A2(n_18), .B(n_21), .C(n_22), .Y(n_754) );
BUFx6f_ASAP7_75t_L g755 ( .A(n_727), .Y(n_755) );
INVx4_ASAP7_75t_SL g756 ( .A(n_621), .Y(n_756) );
OAI21xp5_ASAP7_75t_L g757 ( .A1(n_644), .A2(n_472), .B(n_86), .Y(n_757) );
OAI21x1_ASAP7_75t_L g758 ( .A1(n_697), .A2(n_521), .B(n_493), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_702), .A2(n_521), .B1(n_495), .B2(n_493), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_625), .Y(n_760) );
BUFx8_ASAP7_75t_L g761 ( .A(n_635), .Y(n_761) );
OR2x6_ASAP7_75t_L g762 ( .A(n_679), .B(n_21), .Y(n_762) );
BUFx8_ASAP7_75t_L g763 ( .A(n_674), .Y(n_763) );
INVx2_ASAP7_75t_L g764 ( .A(n_624), .Y(n_764) );
INVx3_ASAP7_75t_L g765 ( .A(n_676), .Y(n_765) );
OAI21x1_ASAP7_75t_L g766 ( .A1(n_633), .A2(n_493), .B(n_484), .Y(n_766) );
OA21x2_ASAP7_75t_L g767 ( .A1(n_633), .A2(n_493), .B(n_484), .Y(n_767) );
INVx2_ASAP7_75t_L g768 ( .A(n_725), .Y(n_768) );
HB1xp67_ASAP7_75t_L g769 ( .A(n_621), .Y(n_769) );
O2A1O1Ixp33_ASAP7_75t_SL g770 ( .A1(n_719), .A2(n_139), .B(n_291), .C(n_290), .Y(n_770) );
AND2x2_ASAP7_75t_L g771 ( .A(n_653), .B(n_23), .Y(n_771) );
NAND3xp33_ASAP7_75t_L g772 ( .A(n_673), .B(n_493), .C(n_484), .Y(n_772) );
OAI21xp5_ASAP7_75t_L g773 ( .A1(n_644), .A2(n_90), .B(n_84), .Y(n_773) );
HB1xp67_ASAP7_75t_L g774 ( .A(n_640), .Y(n_774) );
OAI21x1_ASAP7_75t_L g775 ( .A1(n_694), .A2(n_521), .B(n_493), .Y(n_775) );
O2A1O1Ixp33_ASAP7_75t_L g776 ( .A1(n_648), .A2(n_23), .B(n_24), .C(n_25), .Y(n_776) );
OAI22x1_ASAP7_75t_L g777 ( .A1(n_637), .A2(n_24), .B1(n_25), .B2(n_26), .Y(n_777) );
OAI21x1_ASAP7_75t_L g778 ( .A1(n_694), .A2(n_495), .B(n_484), .Y(n_778) );
AOI22xp5_ASAP7_75t_L g779 ( .A1(n_698), .A2(n_521), .B1(n_495), .B2(n_484), .Y(n_779) );
CKINVDCx5p33_ASAP7_75t_R g780 ( .A(n_704), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_657), .Y(n_781) );
BUFx2_ASAP7_75t_L g782 ( .A(n_704), .Y(n_782) );
OR2x6_ASAP7_75t_L g783 ( .A(n_679), .B(n_27), .Y(n_783) );
INVx4_ASAP7_75t_L g784 ( .A(n_640), .Y(n_784) );
A2O1A1Ixp33_ASAP7_75t_L g785 ( .A1(n_710), .A2(n_521), .B(n_495), .C(n_31), .Y(n_785) );
NAND2x1p5_ASAP7_75t_L g786 ( .A(n_676), .B(n_29), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_740), .Y(n_787) );
OAI21x1_ASAP7_75t_SL g788 ( .A1(n_687), .A2(n_30), .B(n_31), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_740), .Y(n_789) );
AND2x2_ASAP7_75t_L g790 ( .A(n_617), .B(n_32), .Y(n_790) );
NAND2x1p5_ASAP7_75t_L g791 ( .A(n_640), .B(n_32), .Y(n_791) );
AND2x4_ASAP7_75t_L g792 ( .A(n_669), .B(n_33), .Y(n_792) );
AO21x2_ASAP7_75t_L g793 ( .A1(n_655), .A2(n_711), .B(n_656), .Y(n_793) );
AO31x2_ASAP7_75t_L g794 ( .A1(n_655), .A2(n_33), .A3(n_34), .B(n_35), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_629), .Y(n_795) );
BUFx3_ASAP7_75t_L g796 ( .A(n_666), .Y(n_796) );
AND2x4_ASAP7_75t_L g797 ( .A(n_620), .B(n_35), .Y(n_797) );
OAI21x1_ASAP7_75t_L g798 ( .A1(n_731), .A2(n_732), .B(n_667), .Y(n_798) );
OAI21x1_ASAP7_75t_L g799 ( .A1(n_731), .A2(n_92), .B(n_91), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_683), .B(n_36), .Y(n_800) );
OAI21x1_ASAP7_75t_L g801 ( .A1(n_734), .A2(n_100), .B(n_95), .Y(n_801) );
INVx2_ASAP7_75t_L g802 ( .A(n_665), .Y(n_802) );
INVx2_ASAP7_75t_L g803 ( .A(n_671), .Y(n_803) );
INVx4_ASAP7_75t_L g804 ( .A(n_666), .Y(n_804) );
OA21x2_ASAP7_75t_L g805 ( .A1(n_741), .A2(n_104), .B(n_101), .Y(n_805) );
OA21x2_ASAP7_75t_L g806 ( .A1(n_741), .A2(n_106), .B(n_105), .Y(n_806) );
OAI221xp5_ASAP7_75t_L g807 ( .A1(n_630), .A2(n_38), .B1(n_39), .B2(n_40), .C(n_41), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_703), .A2(n_38), .B1(n_39), .B2(n_41), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_705), .A2(n_42), .B1(n_43), .B2(n_45), .Y(n_809) );
OAI21x1_ASAP7_75t_L g810 ( .A1(n_706), .A2(n_109), .B(n_107), .Y(n_810) );
INVxp67_ASAP7_75t_SL g811 ( .A(n_664), .Y(n_811) );
OAI21x1_ASAP7_75t_L g812 ( .A1(n_706), .A2(n_112), .B(n_110), .Y(n_812) );
OAI22xp5_ASAP7_75t_L g813 ( .A1(n_743), .A2(n_43), .B1(n_45), .B2(n_46), .Y(n_813) );
CKINVDCx11_ASAP7_75t_R g814 ( .A(n_748), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_646), .A2(n_47), .B1(n_48), .B2(n_49), .Y(n_815) );
INVx2_ASAP7_75t_L g816 ( .A(n_675), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_678), .Y(n_817) );
AND2x4_ASAP7_75t_L g818 ( .A(n_622), .B(n_50), .Y(n_818) );
INVx2_ASAP7_75t_L g819 ( .A(n_680), .Y(n_819) );
INVxp33_ASAP7_75t_L g820 ( .A(n_632), .Y(n_820) );
OAI22x1_ASAP7_75t_L g821 ( .A1(n_685), .A2(n_51), .B1(n_52), .B2(n_53), .Y(n_821) );
NOR2xp33_ASAP7_75t_L g822 ( .A(n_638), .B(n_51), .Y(n_822) );
OAI22xp5_ASAP7_75t_L g823 ( .A1(n_743), .A2(n_53), .B1(n_54), .B2(n_55), .Y(n_823) );
OA21x2_ASAP7_75t_L g824 ( .A1(n_729), .A2(n_184), .B(n_285), .Y(n_824) );
AND2x2_ASAP7_75t_L g825 ( .A(n_673), .B(n_56), .Y(n_825) );
INVx6_ASAP7_75t_L g826 ( .A(n_666), .Y(n_826) );
OAI21x1_ASAP7_75t_SL g827 ( .A1(n_744), .A2(n_57), .B(n_58), .Y(n_827) );
INVx2_ASAP7_75t_SL g828 ( .A(n_628), .Y(n_828) );
NOR2xp33_ASAP7_75t_L g829 ( .A(n_638), .B(n_57), .Y(n_829) );
OAI21x1_ASAP7_75t_L g830 ( .A1(n_658), .A2(n_187), .B(n_284), .Y(n_830) );
OA21x2_ASAP7_75t_L g831 ( .A1(n_658), .A2(n_182), .B(n_283), .Y(n_831) );
OAI21xp5_ASAP7_75t_L g832 ( .A1(n_721), .A2(n_181), .B(n_282), .Y(n_832) );
OAI21x1_ASAP7_75t_L g833 ( .A1(n_645), .A2(n_180), .B(n_280), .Y(n_833) );
OAI21x1_ASAP7_75t_L g834 ( .A1(n_645), .A2(n_179), .B(n_277), .Y(n_834) );
HB1xp67_ASAP7_75t_L g835 ( .A(n_650), .Y(n_835) );
CKINVDCx5p33_ASAP7_75t_R g836 ( .A(n_692), .Y(n_836) );
OR2x6_ASAP7_75t_L g837 ( .A(n_724), .B(n_59), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_744), .Y(n_838) );
INVx2_ASAP7_75t_L g839 ( .A(n_727), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_646), .A2(n_60), .B1(n_61), .B2(n_62), .Y(n_840) );
HB1xp67_ASAP7_75t_L g841 ( .A(n_650), .Y(n_841) );
NOR2xp33_ASAP7_75t_L g842 ( .A(n_677), .B(n_62), .Y(n_842) );
OAI21x1_ASAP7_75t_L g843 ( .A1(n_647), .A2(n_190), .B(n_273), .Y(n_843) );
AND2x4_ASAP7_75t_L g844 ( .A(n_746), .B(n_63), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_659), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_681), .Y(n_846) );
INVx6_ASAP7_75t_L g847 ( .A(n_715), .Y(n_847) );
AND2x2_ASAP7_75t_L g848 ( .A(n_619), .B(n_63), .Y(n_848) );
OAI21x1_ASAP7_75t_L g849 ( .A1(n_647), .A2(n_192), .B(n_272), .Y(n_849) );
CKINVDCx20_ASAP7_75t_R g850 ( .A(n_699), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_686), .Y(n_851) );
OAI21xp5_ASAP7_75t_L g852 ( .A1(n_722), .A2(n_188), .B(n_271), .Y(n_852) );
OAI21x1_ASAP7_75t_L g853 ( .A1(n_718), .A2(n_174), .B(n_270), .Y(n_853) );
AO31x2_ASAP7_75t_L g854 ( .A1(n_713), .A2(n_64), .A3(n_65), .B(n_66), .Y(n_854) );
AND2x2_ASAP7_75t_L g855 ( .A(n_745), .B(n_64), .Y(n_855) );
BUFx3_ASAP7_75t_L g856 ( .A(n_700), .Y(n_856) );
CKINVDCx11_ASAP7_75t_R g857 ( .A(n_700), .Y(n_857) );
AOI22xp33_ASAP7_75t_SL g858 ( .A1(n_632), .A2(n_65), .B1(n_67), .B2(n_68), .Y(n_858) );
OAI21x1_ASAP7_75t_L g859 ( .A1(n_663), .A2(n_196), .B(n_269), .Y(n_859) );
INVx2_ASAP7_75t_L g860 ( .A(n_727), .Y(n_860) );
OAI21x1_ASAP7_75t_L g861 ( .A1(n_682), .A2(n_172), .B(n_267), .Y(n_861) );
OAI22xp33_ASAP7_75t_L g862 ( .A1(n_649), .A2(n_67), .B1(n_69), .B2(n_71), .Y(n_862) );
AOI22xp5_ASAP7_75t_L g863 ( .A1(n_616), .A2(n_69), .B1(n_72), .B2(n_73), .Y(n_863) );
OAI21xp5_ASAP7_75t_L g864 ( .A1(n_643), .A2(n_200), .B(n_266), .Y(n_864) );
OR2x6_ASAP7_75t_L g865 ( .A(n_634), .B(n_73), .Y(n_865) );
OAI21x1_ASAP7_75t_L g866 ( .A1(n_736), .A2(n_199), .B(n_265), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_649), .A2(n_74), .B1(n_75), .B2(n_76), .Y(n_867) );
BUFx3_ASAP7_75t_L g868 ( .A(n_700), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_668), .B(n_74), .Y(n_869) );
OAI21x1_ASAP7_75t_L g870 ( .A1(n_693), .A2(n_203), .B(n_113), .Y(n_870) );
OAI21x1_ASAP7_75t_L g871 ( .A1(n_696), .A2(n_205), .B(n_117), .Y(n_871) );
BUFx2_ASAP7_75t_L g872 ( .A(n_723), .Y(n_872) );
OAI21x1_ASAP7_75t_L g873 ( .A1(n_689), .A2(n_206), .B(n_118), .Y(n_873) );
OAI21x1_ASAP7_75t_L g874 ( .A1(n_690), .A2(n_207), .B(n_119), .Y(n_874) );
BUFx2_ASAP7_75t_L g875 ( .A(n_723), .Y(n_875) );
AND2x4_ASAP7_75t_L g876 ( .A(n_709), .B(n_120), .Y(n_876) );
AOI221xp5_ASAP7_75t_L g877 ( .A1(n_654), .A2(n_289), .B1(n_124), .B2(n_125), .C(n_126), .Y(n_877) );
INVx2_ASAP7_75t_L g878 ( .A(n_738), .Y(n_878) );
INVx2_ASAP7_75t_L g879 ( .A(n_747), .Y(n_879) );
OAI21x1_ASAP7_75t_L g880 ( .A1(n_739), .A2(n_121), .B(n_127), .Y(n_880) );
NAND2xp33_ASAP7_75t_R g881 ( .A(n_723), .B(n_129), .Y(n_881) );
OAI21x1_ASAP7_75t_SL g882 ( .A1(n_636), .A2(n_135), .B(n_136), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_643), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_662), .A2(n_137), .B1(n_141), .B2(n_143), .Y(n_884) );
OAI21x1_ASAP7_75t_L g885 ( .A1(n_712), .A2(n_144), .B(n_145), .Y(n_885) );
BUFx3_ASAP7_75t_L g886 ( .A(n_726), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g887 ( .A(n_636), .B(n_147), .Y(n_887) );
AO21x2_ASAP7_75t_L g888 ( .A1(n_716), .A2(n_148), .B(n_158), .Y(n_888) );
OAI21x1_ASAP7_75t_L g889 ( .A1(n_712), .A2(n_159), .B(n_160), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_662), .B(n_162), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_660), .Y(n_891) );
AOI21xp5_ASAP7_75t_L g892 ( .A1(n_717), .A2(n_165), .B(n_166), .Y(n_892) );
HB1xp67_ASAP7_75t_L g893 ( .A(n_714), .Y(n_893) );
INVx2_ASAP7_75t_L g894 ( .A(n_749), .Y(n_894) );
AOI22x1_ASAP7_75t_L g895 ( .A1(n_733), .A2(n_168), .B1(n_171), .B2(n_208), .Y(n_895) );
AOI22xp5_ASAP7_75t_L g896 ( .A1(n_825), .A2(n_684), .B1(n_701), .B2(n_631), .Y(n_896) );
OAI221xp5_ASAP7_75t_L g897 ( .A1(n_845), .A2(n_651), .B1(n_670), .B2(n_626), .C(n_691), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_772), .A2(n_631), .B1(n_684), .B2(n_623), .Y(n_898) );
AOI21xp33_ASAP7_75t_SL g899 ( .A1(n_780), .A2(n_661), .B(n_660), .Y(n_899) );
OAI221xp5_ASAP7_75t_L g900 ( .A1(n_842), .A2(n_672), .B1(n_720), .B2(n_627), .C(n_618), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_842), .A2(n_730), .B1(n_652), .B2(n_641), .Y(n_901) );
OR2x2_ASAP7_75t_L g902 ( .A(n_782), .B(n_728), .Y(n_902) );
INVx3_ASAP7_75t_L g903 ( .A(n_784), .Y(n_903) );
INVx2_ASAP7_75t_L g904 ( .A(n_781), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_750), .A2(n_695), .B1(n_707), .B2(n_688), .Y(n_905) );
CKINVDCx5p33_ASAP7_75t_R g906 ( .A(n_763), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_750), .A2(n_715), .B1(n_726), .B2(n_737), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_751), .B(n_733), .Y(n_908) );
AOI21x1_ASAP7_75t_L g909 ( .A1(n_766), .A2(n_735), .B(n_212), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_795), .B(n_735), .Y(n_910) );
A2O1A1Ixp33_ASAP7_75t_L g911 ( .A1(n_822), .A2(n_210), .B(n_213), .C(n_218), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_817), .Y(n_912) );
OAI221xp5_ASAP7_75t_SL g913 ( .A1(n_863), .A2(n_220), .B1(n_221), .B2(n_223), .C(n_225), .Y(n_913) );
OAI21x1_ASAP7_75t_L g914 ( .A1(n_758), .A2(n_227), .B(n_231), .Y(n_914) );
INVx1_ASAP7_75t_L g915 ( .A(n_851), .Y(n_915) );
BUFx6f_ASAP7_75t_L g916 ( .A(n_857), .Y(n_916) );
OAI211xp5_ASAP7_75t_L g917 ( .A1(n_809), .A2(n_232), .B(n_235), .C(n_236), .Y(n_917) );
INVx2_ASAP7_75t_L g918 ( .A(n_781), .Y(n_918) );
AO31x2_ASAP7_75t_L g919 ( .A1(n_785), .A2(n_240), .A3(n_243), .B(n_245), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_829), .A2(n_246), .B1(n_248), .B2(n_249), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_829), .A2(n_251), .B1(n_254), .B2(n_257), .Y(n_921) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_838), .A2(n_258), .B1(n_260), .B2(n_261), .Y(n_922) );
OAI22xp5_ASAP7_75t_L g923 ( .A1(n_837), .A2(n_787), .B1(n_789), .B2(n_792), .Y(n_923) );
AOI221xp5_ASAP7_75t_L g924 ( .A1(n_862), .A2(n_752), .B1(n_807), .B2(n_771), .C(n_800), .Y(n_924) );
OAI211xp5_ASAP7_75t_L g925 ( .A1(n_808), .A2(n_858), .B(n_840), .C(n_867), .Y(n_925) );
AOI21xp5_ASAP7_75t_L g926 ( .A1(n_811), .A2(n_887), .B(n_778), .Y(n_926) );
AOI21xp5_ASAP7_75t_L g927 ( .A1(n_811), .A2(n_775), .B(n_890), .Y(n_927) );
AOI221xp5_ASAP7_75t_L g928 ( .A1(n_862), .A2(n_752), .B1(n_807), .B2(n_754), .C(n_776), .Y(n_928) );
INVx2_ASAP7_75t_L g929 ( .A(n_768), .Y(n_929) );
AOI21xp5_ASAP7_75t_L g930 ( .A1(n_757), .A2(n_770), .B(n_767), .Y(n_930) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_802), .B(n_803), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_816), .Y(n_932) );
AO31x2_ASAP7_75t_L g933 ( .A1(n_785), .A2(n_892), .A3(n_891), .B(n_883), .Y(n_933) );
AOI222xp33_ASAP7_75t_L g934 ( .A1(n_814), .A2(n_821), .B1(n_777), .B2(n_840), .C1(n_867), .C2(n_815), .Y(n_934) );
AND2x2_ASAP7_75t_L g935 ( .A(n_893), .B(n_762), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_819), .B(n_848), .Y(n_936) );
INVx2_ASAP7_75t_L g937 ( .A(n_768), .Y(n_937) );
BUFx2_ASAP7_75t_L g938 ( .A(n_837), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_846), .Y(n_939) );
AOI22xp33_ASAP7_75t_SL g940 ( .A1(n_837), .A2(n_783), .B1(n_762), .B2(n_844), .Y(n_940) );
OR2x2_ASAP7_75t_L g941 ( .A(n_836), .B(n_828), .Y(n_941) );
OAI22xp5_ASAP7_75t_L g942 ( .A1(n_872), .A2(n_875), .B1(n_820), .B2(n_783), .Y(n_942) );
INVx2_ASAP7_75t_L g943 ( .A(n_764), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_865), .A2(n_869), .B1(n_790), .B2(n_818), .Y(n_944) );
OR2x6_ASAP7_75t_L g945 ( .A(n_783), .B(n_786), .Y(n_945) );
AOI222xp33_ASAP7_75t_L g946 ( .A1(n_814), .A2(n_844), .B1(n_818), .B2(n_797), .C1(n_815), .C2(n_763), .Y(n_946) );
OAI22xp5_ASAP7_75t_L g947 ( .A1(n_820), .A2(n_786), .B1(n_797), .B2(n_808), .Y(n_947) );
AOI22xp5_ASAP7_75t_L g948 ( .A1(n_881), .A2(n_865), .B1(n_813), .B2(n_823), .Y(n_948) );
INVx3_ASAP7_75t_L g949 ( .A(n_784), .Y(n_949) );
OR2x2_ASAP7_75t_L g950 ( .A(n_835), .B(n_841), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_764), .Y(n_951) );
OAI211xp5_ASAP7_75t_SL g952 ( .A1(n_776), .A2(n_857), .B(n_877), .C(n_892), .Y(n_952) );
OA21x2_ASAP7_75t_L g953 ( .A1(n_885), .A2(n_889), .B(n_773), .Y(n_953) );
AND2x4_ASAP7_75t_L g954 ( .A(n_756), .B(n_804), .Y(n_954) );
INVx2_ASAP7_75t_L g955 ( .A(n_760), .Y(n_955) );
OAI22xp5_ASAP7_75t_L g956 ( .A1(n_835), .A2(n_841), .B1(n_791), .B2(n_855), .Y(n_956) );
AND2x4_ASAP7_75t_L g957 ( .A(n_756), .B(n_804), .Y(n_957) );
OAI22xp33_ASAP7_75t_SL g958 ( .A1(n_791), .A2(n_847), .B1(n_864), .B2(n_895), .Y(n_958) );
OAI21xp33_ASAP7_75t_L g959 ( .A1(n_877), .A2(n_759), .B(n_884), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_876), .A2(n_793), .B1(n_827), .B2(n_765), .Y(n_960) );
AOI21xp5_ASAP7_75t_L g961 ( .A1(n_770), .A2(n_767), .B(n_759), .Y(n_961) );
INVx1_ASAP7_75t_L g962 ( .A(n_794), .Y(n_962) );
INVx2_ASAP7_75t_L g963 ( .A(n_878), .Y(n_963) );
INVx1_ASAP7_75t_L g964 ( .A(n_794), .Y(n_964) );
OAI21xp5_ASAP7_75t_L g965 ( .A1(n_779), .A2(n_798), .B(n_801), .Y(n_965) );
OAI21xp5_ASAP7_75t_L g966 ( .A1(n_879), .A2(n_894), .B(n_830), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_876), .A2(n_793), .B1(n_765), .B2(n_847), .Y(n_967) );
AND2x2_ASAP7_75t_L g968 ( .A(n_753), .B(n_769), .Y(n_968) );
OR2x2_ASAP7_75t_L g969 ( .A(n_753), .B(n_769), .Y(n_969) );
AOI22xp5_ASAP7_75t_L g970 ( .A1(n_847), .A2(n_806), .B1(n_805), .B2(n_826), .Y(n_970) );
NAND2xp5_ASAP7_75t_SL g971 ( .A(n_756), .B(n_796), .Y(n_971) );
AOI21xp5_ASAP7_75t_R g972 ( .A1(n_761), .A2(n_850), .B(n_854), .Y(n_972) );
O2A1O1Ixp33_ASAP7_75t_L g973 ( .A1(n_788), .A2(n_882), .B(n_852), .C(n_832), .Y(n_973) );
AND2x4_ASAP7_75t_L g974 ( .A(n_856), .B(n_868), .Y(n_974) );
AOI221xp5_ASAP7_75t_L g975 ( .A1(n_774), .A2(n_886), .B1(n_856), .B2(n_868), .C(n_888), .Y(n_975) );
OR2x6_ASAP7_75t_L g976 ( .A(n_826), .B(n_886), .Y(n_976) );
AND2x2_ASAP7_75t_L g977 ( .A(n_854), .B(n_794), .Y(n_977) );
OAI21xp5_ASAP7_75t_L g978 ( .A1(n_880), .A2(n_853), .B(n_866), .Y(n_978) );
NAND2xp5_ASAP7_75t_L g979 ( .A(n_794), .B(n_854), .Y(n_979) );
INVx8_ASAP7_75t_L g980 ( .A(n_755), .Y(n_980) );
AOI21xp5_ASAP7_75t_L g981 ( .A1(n_755), .A2(n_839), .B(n_860), .Y(n_981) );
OAI221xp5_ASAP7_75t_L g982 ( .A1(n_805), .A2(n_806), .B1(n_831), .B2(n_860), .C(n_839), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_761), .A2(n_805), .B1(n_806), .B2(n_831), .Y(n_983) );
BUFx6f_ASAP7_75t_L g984 ( .A(n_755), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_831), .A2(n_755), .B1(n_810), .B2(n_812), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g986 ( .A1(n_824), .A2(n_833), .B1(n_834), .B2(n_843), .Y(n_986) );
AND2x4_ASAP7_75t_L g987 ( .A(n_849), .B(n_799), .Y(n_987) );
NAND2xp5_ASAP7_75t_L g988 ( .A(n_874), .B(n_873), .Y(n_988) );
AOI221xp5_ASAP7_75t_L g989 ( .A1(n_859), .A2(n_861), .B1(n_870), .B2(n_871), .C(n_824), .Y(n_989) );
HB1xp67_ASAP7_75t_L g990 ( .A(n_824), .Y(n_990) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_825), .A2(n_561), .B1(n_616), .B2(n_703), .Y(n_991) );
AND2x2_ASAP7_75t_L g992 ( .A(n_825), .B(n_531), .Y(n_992) );
NAND3xp33_ASAP7_75t_L g993 ( .A(n_785), .B(n_772), .C(n_877), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_751), .Y(n_994) );
BUFx2_ASAP7_75t_L g995 ( .A(n_837), .Y(n_995) );
AOI222xp33_ASAP7_75t_L g996 ( .A1(n_825), .A2(n_561), .B1(n_464), .B2(n_548), .C1(n_544), .C2(n_530), .Y(n_996) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_751), .B(n_544), .Y(n_997) );
OAI21x1_ASAP7_75t_L g998 ( .A1(n_758), .A2(n_766), .B(n_775), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_825), .A2(n_561), .B1(n_616), .B2(n_703), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g1000 ( .A(n_751), .B(n_544), .Y(n_1000) );
AOI222xp33_ASAP7_75t_L g1001 ( .A1(n_825), .A2(n_561), .B1(n_464), .B2(n_454), .C1(n_408), .C2(n_548), .Y(n_1001) );
OAI221xp5_ASAP7_75t_SL g1002 ( .A1(n_750), .A2(n_530), .B1(n_536), .B2(n_544), .C(n_673), .Y(n_1002) );
AOI21xp5_ASAP7_75t_L g1003 ( .A1(n_811), .A2(n_644), .B(n_633), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_825), .B(n_531), .Y(n_1004) );
AND2x4_ASAP7_75t_L g1005 ( .A(n_756), .B(n_669), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_825), .A2(n_561), .B1(n_616), .B2(n_703), .Y(n_1006) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_825), .A2(n_561), .B1(n_616), .B2(n_703), .Y(n_1007) );
INVx1_ASAP7_75t_L g1008 ( .A(n_751), .Y(n_1008) );
HB1xp67_ASAP7_75t_L g1009 ( .A(n_837), .Y(n_1009) );
OAI22x1_ASAP7_75t_L g1010 ( .A1(n_782), .A2(n_470), .B1(n_536), .B2(n_575), .Y(n_1010) );
INVx2_ASAP7_75t_SL g1011 ( .A(n_782), .Y(n_1011) );
INVx2_ASAP7_75t_L g1012 ( .A(n_781), .Y(n_1012) );
NAND2xp5_ASAP7_75t_L g1013 ( .A(n_751), .B(n_544), .Y(n_1013) );
AO31x2_ASAP7_75t_L g1014 ( .A1(n_785), .A2(n_644), .A3(n_633), .B(n_694), .Y(n_1014) );
OR2x2_ASAP7_75t_L g1015 ( .A(n_782), .B(n_531), .Y(n_1015) );
INVx4_ASAP7_75t_L g1016 ( .A(n_857), .Y(n_1016) );
BUFx6f_ASAP7_75t_L g1017 ( .A(n_857), .Y(n_1017) );
INVx1_ASAP7_75t_L g1018 ( .A(n_951), .Y(n_1018) );
INVx1_ASAP7_75t_L g1019 ( .A(n_904), .Y(n_1019) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_918), .B(n_1012), .Y(n_1020) );
OA21x2_ASAP7_75t_L g1021 ( .A1(n_930), .A2(n_961), .B(n_998), .Y(n_1021) );
BUFx3_ASAP7_75t_L g1022 ( .A(n_1005), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_929), .Y(n_1023) );
NAND2xp5_ASAP7_75t_L g1024 ( .A(n_996), .B(n_992), .Y(n_1024) );
AND2x4_ASAP7_75t_L g1025 ( .A(n_945), .B(n_1005), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_937), .Y(n_1026) );
HB1xp67_ASAP7_75t_L g1027 ( .A(n_950), .Y(n_1027) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_943), .B(n_932), .Y(n_1028) );
NOR2xp33_ASAP7_75t_L g1029 ( .A(n_1002), .B(n_1015), .Y(n_1029) );
AND2x4_ASAP7_75t_L g1030 ( .A(n_945), .B(n_954), .Y(n_1030) );
BUFx2_ASAP7_75t_L g1031 ( .A(n_945), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_955), .B(n_912), .Y(n_1032) );
INVx2_ASAP7_75t_SL g1033 ( .A(n_980), .Y(n_1033) );
AND2x4_ASAP7_75t_L g1034 ( .A(n_954), .B(n_957), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_994), .B(n_1008), .Y(n_1035) );
AND2x4_ASAP7_75t_L g1036 ( .A(n_957), .B(n_974), .Y(n_1036) );
AND2x4_ASAP7_75t_L g1037 ( .A(n_974), .B(n_968), .Y(n_1037) );
INVx1_ASAP7_75t_L g1038 ( .A(n_962), .Y(n_1038) );
INVx2_ASAP7_75t_L g1039 ( .A(n_909), .Y(n_1039) );
INVx2_ASAP7_75t_L g1040 ( .A(n_914), .Y(n_1040) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_939), .B(n_977), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g1042 ( .A(n_1004), .B(n_1001), .Y(n_1042) );
NAND2xp5_ASAP7_75t_L g1043 ( .A(n_1001), .B(n_991), .Y(n_1043) );
OR2x2_ASAP7_75t_SL g1044 ( .A(n_1009), .B(n_916), .Y(n_1044) );
BUFx3_ASAP7_75t_L g1045 ( .A(n_980), .Y(n_1045) );
AND2x2_ASAP7_75t_L g1046 ( .A(n_963), .B(n_915), .Y(n_1046) );
INVx1_ASAP7_75t_L g1047 ( .A(n_964), .Y(n_1047) );
NAND2xp5_ASAP7_75t_L g1048 ( .A(n_999), .B(n_1006), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_979), .Y(n_1049) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_931), .B(n_940), .Y(n_1050) );
INVx2_ASAP7_75t_L g1051 ( .A(n_984), .Y(n_1051) );
OAI21x1_ASAP7_75t_L g1052 ( .A1(n_965), .A2(n_988), .B(n_978), .Y(n_1052) );
HB1xp67_ASAP7_75t_L g1053 ( .A(n_902), .Y(n_1053) );
OAI321xp33_ASAP7_75t_L g1054 ( .A1(n_952), .A2(n_947), .A3(n_948), .B1(n_913), .B2(n_923), .C(n_983), .Y(n_1054) );
INVx2_ASAP7_75t_L g1055 ( .A(n_984), .Y(n_1055) );
INVxp67_ASAP7_75t_SL g1056 ( .A(n_956), .Y(n_1056) );
AND2x2_ASAP7_75t_L g1057 ( .A(n_934), .B(n_936), .Y(n_1057) );
OAI221xp5_ASAP7_75t_L g1058 ( .A1(n_1007), .A2(n_896), .B1(n_944), .B2(n_948), .C(n_946), .Y(n_1058) );
INVx1_ASAP7_75t_L g1059 ( .A(n_933), .Y(n_1059) );
NOR2xp33_ASAP7_75t_L g1060 ( .A(n_938), .B(n_995), .Y(n_1060) );
OR2x2_ASAP7_75t_L g1061 ( .A(n_969), .B(n_997), .Y(n_1061) );
OR2x2_ASAP7_75t_L g1062 ( .A(n_1000), .B(n_1013), .Y(n_1062) );
NOR2xp67_ASAP7_75t_L g1063 ( .A(n_1016), .B(n_906), .Y(n_1063) );
INVx3_ASAP7_75t_L g1064 ( .A(n_980), .Y(n_1064) );
BUFx3_ASAP7_75t_L g1065 ( .A(n_916), .Y(n_1065) );
AND2x4_ASAP7_75t_L g1066 ( .A(n_903), .B(n_949), .Y(n_1066) );
OR2x2_ASAP7_75t_L g1067 ( .A(n_942), .B(n_896), .Y(n_1067) );
BUFx2_ASAP7_75t_L g1068 ( .A(n_970), .Y(n_1068) );
HB1xp67_ASAP7_75t_L g1069 ( .A(n_935), .Y(n_1069) );
NAND2xp5_ASAP7_75t_L g1070 ( .A(n_934), .B(n_1010), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_903), .B(n_949), .Y(n_1071) );
INVx1_ASAP7_75t_L g1072 ( .A(n_908), .Y(n_1072) );
AOI22xp33_ASAP7_75t_L g1073 ( .A1(n_928), .A2(n_924), .B1(n_897), .B2(n_959), .Y(n_1073) );
NAND2xp5_ASAP7_75t_L g1074 ( .A(n_899), .B(n_905), .Y(n_1074) );
INVx2_ASAP7_75t_L g1075 ( .A(n_1014), .Y(n_1075) );
NAND2xp5_ASAP7_75t_L g1076 ( .A(n_1011), .B(n_925), .Y(n_1076) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_898), .B(n_901), .Y(n_1077) );
INVx2_ASAP7_75t_L g1078 ( .A(n_1014), .Y(n_1078) );
OAI211xp5_ASAP7_75t_L g1079 ( .A1(n_907), .A2(n_960), .B(n_972), .C(n_967), .Y(n_1079) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_976), .B(n_910), .Y(n_1080) );
INVx2_ASAP7_75t_L g1081 ( .A(n_1014), .Y(n_1081) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_976), .B(n_919), .Y(n_1082) );
INVx2_ASAP7_75t_L g1083 ( .A(n_987), .Y(n_1083) );
AND2x4_ASAP7_75t_L g1084 ( .A(n_976), .B(n_971), .Y(n_1084) );
INVx8_ASAP7_75t_L g1085 ( .A(n_1017), .Y(n_1085) );
AND2x2_ASAP7_75t_L g1086 ( .A(n_919), .B(n_966), .Y(n_1086) );
INVx2_ASAP7_75t_L g1087 ( .A(n_987), .Y(n_1087) );
INVxp67_ASAP7_75t_L g1088 ( .A(n_941), .Y(n_1088) );
AND2x2_ASAP7_75t_L g1089 ( .A(n_919), .B(n_970), .Y(n_1089) );
NAND2xp5_ASAP7_75t_L g1090 ( .A(n_993), .B(n_900), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_993), .B(n_1003), .Y(n_1091) );
INVx1_ASAP7_75t_L g1092 ( .A(n_982), .Y(n_1092) );
INVx1_ASAP7_75t_L g1093 ( .A(n_990), .Y(n_1093) );
HB1xp67_ASAP7_75t_L g1094 ( .A(n_981), .Y(n_1094) );
NAND3xp33_ASAP7_75t_L g1095 ( .A(n_975), .B(n_911), .C(n_973), .Y(n_1095) );
NOR2xp33_ASAP7_75t_L g1096 ( .A(n_917), .B(n_958), .Y(n_1096) );
NAND2xp5_ASAP7_75t_L g1097 ( .A(n_920), .B(n_921), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1098 ( .A(n_922), .B(n_953), .Y(n_1098) );
AND2x4_ASAP7_75t_L g1099 ( .A(n_985), .B(n_926), .Y(n_1099) );
BUFx3_ASAP7_75t_L g1100 ( .A(n_958), .Y(n_1100) );
INVx1_ASAP7_75t_L g1101 ( .A(n_986), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_927), .B(n_989), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_1041), .B(n_1091), .Y(n_1103) );
BUFx3_ASAP7_75t_L g1104 ( .A(n_1045), .Y(n_1104) );
INVxp67_ASAP7_75t_L g1105 ( .A(n_1053), .Y(n_1105) );
AOI221xp5_ASAP7_75t_L g1106 ( .A1(n_1058), .A2(n_1043), .B1(n_1024), .B2(n_1048), .C(n_1042), .Y(n_1106) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_1057), .A2(n_1067), .B1(n_1070), .B2(n_1029), .Y(n_1107) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1038), .Y(n_1108) );
OR2x2_ASAP7_75t_L g1109 ( .A(n_1067), .B(n_1027), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1035), .Y(n_1110) );
OR2x2_ASAP7_75t_L g1111 ( .A(n_1049), .B(n_1038), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_1020), .B(n_1049), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_1020), .B(n_1047), .Y(n_1113) );
AOI22xp5_ASAP7_75t_L g1114 ( .A1(n_1050), .A2(n_1073), .B1(n_1074), .B2(n_1076), .Y(n_1114) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_1028), .B(n_1032), .Y(n_1115) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_1028), .B(n_1032), .Y(n_1116) );
NOR2xp33_ASAP7_75t_R g1117 ( .A(n_1022), .B(n_1064), .Y(n_1117) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1093), .Y(n_1118) );
HB1xp67_ASAP7_75t_L g1119 ( .A(n_1046), .Y(n_1119) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_1046), .B(n_1019), .Y(n_1120) );
AND2x2_ASAP7_75t_L g1121 ( .A(n_1019), .B(n_1101), .Y(n_1121) );
OAI31xp33_ASAP7_75t_L g1122 ( .A1(n_1079), .A2(n_1031), .A3(n_1077), .B(n_1090), .Y(n_1122) );
AND2x2_ASAP7_75t_L g1123 ( .A(n_1101), .B(n_1023), .Y(n_1123) );
AND2x2_ASAP7_75t_L g1124 ( .A(n_1023), .B(n_1026), .Y(n_1124) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1018), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_1026), .B(n_1092), .Y(n_1126) );
AOI221xp5_ASAP7_75t_L g1127 ( .A1(n_1072), .A2(n_1054), .B1(n_1088), .B2(n_1060), .C(n_1056), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1128 ( .A(n_1061), .B(n_1062), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1129 ( .A(n_1092), .B(n_1078), .Y(n_1129) );
HB1xp67_ASAP7_75t_L g1130 ( .A(n_1071), .Y(n_1130) );
NAND3xp33_ASAP7_75t_SL g1131 ( .A(n_1071), .B(n_1096), .C(n_1095), .Y(n_1131) );
NAND2xp5_ASAP7_75t_L g1132 ( .A(n_1037), .B(n_1069), .Y(n_1132) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_1075), .B(n_1078), .Y(n_1133) );
OAI22xp33_ASAP7_75t_SL g1134 ( .A1(n_1025), .A2(n_1030), .B1(n_1022), .B2(n_1066), .Y(n_1134) );
AND2x4_ASAP7_75t_L g1135 ( .A(n_1083), .B(n_1087), .Y(n_1135) );
INVx2_ASAP7_75t_SL g1136 ( .A(n_1025), .Y(n_1136) );
INVx5_ASAP7_75t_SL g1137 ( .A(n_1025), .Y(n_1137) );
OR2x6_ASAP7_75t_L g1138 ( .A(n_1068), .B(n_1030), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1081), .B(n_1089), .Y(n_1139) );
AOI22xp5_ASAP7_75t_L g1140 ( .A1(n_1097), .A2(n_1030), .B1(n_1080), .B2(n_1063), .Y(n_1140) );
INVx5_ASAP7_75t_SL g1141 ( .A(n_1034), .Y(n_1141) );
HB1xp67_ASAP7_75t_L g1142 ( .A(n_1066), .Y(n_1142) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1059), .Y(n_1143) );
NAND3xp33_ASAP7_75t_L g1144 ( .A(n_1094), .B(n_1102), .C(n_1082), .Y(n_1144) );
BUFx2_ASAP7_75t_L g1145 ( .A(n_1044), .Y(n_1145) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1044), .Y(n_1146) );
INVx1_ASAP7_75t_SL g1147 ( .A(n_1045), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_1037), .B(n_1086), .Y(n_1148) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1108), .Y(n_1149) );
OAI211xp5_ASAP7_75t_L g1150 ( .A1(n_1122), .A2(n_1085), .B(n_1100), .C(n_1065), .Y(n_1150) );
INVx1_ASAP7_75t_SL g1151 ( .A(n_1117), .Y(n_1151) );
NAND2x1p5_ASAP7_75t_L g1152 ( .A(n_1104), .B(n_1034), .Y(n_1152) );
NAND2xp5_ASAP7_75t_L g1153 ( .A(n_1115), .B(n_1080), .Y(n_1153) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_1103), .B(n_1100), .Y(n_1154) );
NAND3xp33_ASAP7_75t_L g1155 ( .A(n_1127), .B(n_1106), .C(n_1114), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1156 ( .A(n_1139), .B(n_1099), .Y(n_1156) );
HB1xp67_ASAP7_75t_L g1157 ( .A(n_1119), .Y(n_1157) );
AND2x2_ASAP7_75t_L g1158 ( .A(n_1139), .B(n_1099), .Y(n_1158) );
AND2x4_ASAP7_75t_L g1159 ( .A(n_1135), .B(n_1099), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_1148), .B(n_1052), .Y(n_1160) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_1148), .B(n_1052), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_1129), .B(n_1098), .Y(n_1162) );
HB1xp67_ASAP7_75t_L g1163 ( .A(n_1130), .Y(n_1163) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1129), .B(n_1098), .Y(n_1164) );
INVx1_ASAP7_75t_SL g1165 ( .A(n_1147), .Y(n_1165) );
INVx1_ASAP7_75t_SL g1166 ( .A(n_1104), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_1113), .B(n_1021), .Y(n_1167) );
AND2x2_ASAP7_75t_L g1168 ( .A(n_1113), .B(n_1051), .Y(n_1168) );
AOI211xp5_ASAP7_75t_L g1169 ( .A1(n_1134), .A2(n_1036), .B(n_1084), .C(n_1033), .Y(n_1169) );
OAI21xp5_ASAP7_75t_L g1170 ( .A1(n_1131), .A2(n_1084), .B(n_1033), .Y(n_1170) );
O2A1O1Ixp33_ASAP7_75t_L g1171 ( .A1(n_1105), .A2(n_1064), .B(n_1039), .C(n_1051), .Y(n_1171) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1143), .Y(n_1172) );
OR2x2_ASAP7_75t_L g1173 ( .A(n_1109), .B(n_1036), .Y(n_1173) );
OR2x2_ASAP7_75t_L g1174 ( .A(n_1109), .B(n_1036), .Y(n_1174) );
BUFx2_ASAP7_75t_L g1175 ( .A(n_1138), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1116), .B(n_1055), .Y(n_1176) );
OR2x2_ASAP7_75t_L g1177 ( .A(n_1111), .B(n_1085), .Y(n_1177) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1111), .Y(n_1178) );
INVx4_ASAP7_75t_L g1179 ( .A(n_1138), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1112), .B(n_1123), .Y(n_1180) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1125), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1112), .B(n_1040), .Y(n_1182) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_1157), .B(n_1110), .Y(n_1183) );
NAND2xp5_ASAP7_75t_L g1184 ( .A(n_1180), .B(n_1120), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1160), .B(n_1161), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1160), .B(n_1138), .Y(n_1186) );
INVx1_ASAP7_75t_SL g1187 ( .A(n_1165), .Y(n_1187) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1149), .Y(n_1188) );
AND2x2_ASAP7_75t_L g1189 ( .A(n_1161), .B(n_1138), .Y(n_1189) );
INVxp67_ASAP7_75t_L g1190 ( .A(n_1165), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1156), .B(n_1133), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1158), .B(n_1135), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1162), .B(n_1123), .Y(n_1193) );
NAND2xp5_ASAP7_75t_L g1194 ( .A(n_1178), .B(n_1107), .Y(n_1194) );
INVx1_ASAP7_75t_SL g1195 ( .A(n_1166), .Y(n_1195) );
NOR2xp67_ASAP7_75t_L g1196 ( .A(n_1179), .B(n_1146), .Y(n_1196) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1172), .Y(n_1197) );
NAND2xp5_ASAP7_75t_L g1198 ( .A(n_1163), .B(n_1126), .Y(n_1198) );
NAND2xp5_ASAP7_75t_SL g1199 ( .A(n_1151), .B(n_1145), .Y(n_1199) );
OR2x2_ASAP7_75t_L g1200 ( .A(n_1162), .B(n_1118), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1164), .B(n_1121), .Y(n_1201) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1172), .Y(n_1202) );
AND2x2_ASAP7_75t_SL g1203 ( .A(n_1179), .B(n_1142), .Y(n_1203) );
AND2x2_ASAP7_75t_L g1204 ( .A(n_1164), .B(n_1121), .Y(n_1204) );
INVxp67_ASAP7_75t_SL g1205 ( .A(n_1171), .Y(n_1205) );
AOI22xp5_ASAP7_75t_L g1206 ( .A1(n_1155), .A2(n_1128), .B1(n_1140), .B2(n_1132), .Y(n_1206) );
NAND2xp5_ASAP7_75t_L g1207 ( .A(n_1176), .B(n_1153), .Y(n_1207) );
NAND2xp5_ASAP7_75t_L g1208 ( .A(n_1176), .B(n_1124), .Y(n_1208) );
INVx4_ASAP7_75t_L g1209 ( .A(n_1152), .Y(n_1209) );
OAI22xp5_ASAP7_75t_L g1210 ( .A1(n_1206), .A2(n_1151), .B1(n_1169), .B2(n_1155), .Y(n_1210) );
HB1xp67_ASAP7_75t_L g1211 ( .A(n_1195), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g1212 ( .A(n_1193), .B(n_1167), .Y(n_1212) );
INVx3_ASAP7_75t_L g1213 ( .A(n_1209), .Y(n_1213) );
AOI21xp5_ASAP7_75t_L g1214 ( .A1(n_1203), .A2(n_1169), .B(n_1170), .Y(n_1214) );
AND2x4_ASAP7_75t_L g1215 ( .A(n_1196), .B(n_1179), .Y(n_1215) );
OAI21xp5_ASAP7_75t_L g1216 ( .A1(n_1205), .A2(n_1166), .B(n_1150), .Y(n_1216) );
AND2x2_ASAP7_75t_L g1217 ( .A(n_1185), .B(n_1154), .Y(n_1217) );
OAI32xp33_ASAP7_75t_L g1218 ( .A1(n_1187), .A2(n_1152), .A3(n_1179), .B1(n_1177), .B2(n_1174), .Y(n_1218) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1200), .Y(n_1219) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1200), .Y(n_1220) );
INVxp33_ASAP7_75t_L g1221 ( .A(n_1196), .Y(n_1221) );
OAI22xp33_ASAP7_75t_L g1222 ( .A1(n_1209), .A2(n_1177), .B1(n_1175), .B2(n_1173), .Y(n_1222) );
AOI222xp33_ASAP7_75t_L g1223 ( .A1(n_1194), .A2(n_1167), .B1(n_1175), .B2(n_1144), .C1(n_1182), .C2(n_1181), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1183), .Y(n_1224) );
NAND2xp5_ASAP7_75t_L g1225 ( .A(n_1193), .B(n_1168), .Y(n_1225) );
NOR2xp33_ASAP7_75t_L g1226 ( .A(n_1190), .B(n_1173), .Y(n_1226) );
NAND2xp5_ASAP7_75t_L g1227 ( .A(n_1201), .B(n_1168), .Y(n_1227) );
NAND2xp5_ASAP7_75t_L g1228 ( .A(n_1201), .B(n_1182), .Y(n_1228) );
AND2x2_ASAP7_75t_L g1229 ( .A(n_1185), .B(n_1159), .Y(n_1229) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1188), .Y(n_1230) );
OAI22xp5_ASAP7_75t_L g1231 ( .A1(n_1209), .A2(n_1152), .B1(n_1141), .B2(n_1137), .Y(n_1231) );
NOR2xp33_ASAP7_75t_L g1232 ( .A(n_1224), .B(n_1184), .Y(n_1232) );
O2A1O1Ixp5_ASAP7_75t_L g1233 ( .A1(n_1210), .A2(n_1199), .B(n_1209), .C(n_1198), .Y(n_1233) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1230), .Y(n_1234) );
NAND2xp5_ASAP7_75t_L g1235 ( .A(n_1223), .B(n_1204), .Y(n_1235) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1219), .Y(n_1236) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1220), .Y(n_1237) );
OR2x2_ASAP7_75t_L g1238 ( .A(n_1212), .B(n_1207), .Y(n_1238) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1225), .Y(n_1239) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1227), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1228), .Y(n_1241) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1211), .Y(n_1242) );
XNOR2xp5_ASAP7_75t_L g1243 ( .A(n_1214), .B(n_1208), .Y(n_1243) );
NAND2xp5_ASAP7_75t_L g1244 ( .A(n_1217), .B(n_1204), .Y(n_1244) );
OAI31xp33_ASAP7_75t_L g1245 ( .A1(n_1235), .A2(n_1222), .A3(n_1213), .B(n_1221), .Y(n_1245) );
INVxp67_ASAP7_75t_SL g1246 ( .A(n_1242), .Y(n_1246) );
O2A1O1Ixp33_ASAP7_75t_L g1247 ( .A1(n_1233), .A2(n_1216), .B(n_1218), .C(n_1213), .Y(n_1247) );
A2O1A1Ixp33_ASAP7_75t_L g1248 ( .A1(n_1235), .A2(n_1215), .B(n_1226), .C(n_1231), .Y(n_1248) );
AND2x2_ASAP7_75t_L g1249 ( .A(n_1239), .B(n_1229), .Y(n_1249) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1234), .Y(n_1250) );
NOR2x1_ASAP7_75t_L g1251 ( .A(n_1243), .B(n_1215), .Y(n_1251) );
AOI22xp33_ASAP7_75t_L g1252 ( .A1(n_1251), .A2(n_1232), .B1(n_1241), .B2(n_1240), .Y(n_1252) );
OAI21xp5_ASAP7_75t_L g1253 ( .A1(n_1247), .A2(n_1236), .B(n_1237), .Y(n_1253) );
O2A1O1Ixp33_ASAP7_75t_L g1254 ( .A1(n_1248), .A2(n_1244), .B(n_1238), .C(n_1136), .Y(n_1254) );
AOI211xp5_ASAP7_75t_L g1255 ( .A1(n_1245), .A2(n_1215), .B(n_1186), .C(n_1189), .Y(n_1255) );
AOI211xp5_ASAP7_75t_L g1256 ( .A1(n_1254), .A2(n_1246), .B(n_1250), .C(n_1249), .Y(n_1256) );
OAI22xp5_ASAP7_75t_L g1257 ( .A1(n_1252), .A2(n_1203), .B1(n_1137), .B2(n_1141), .Y(n_1257) );
OR2x2_ASAP7_75t_L g1258 ( .A(n_1253), .B(n_1191), .Y(n_1258) );
NOR3xp33_ASAP7_75t_SL g1259 ( .A(n_1257), .B(n_1255), .C(n_1252), .Y(n_1259) );
OAI22xp5_ASAP7_75t_L g1260 ( .A1(n_1259), .A2(n_1256), .B1(n_1258), .B2(n_1203), .Y(n_1260) );
INVx2_ASAP7_75t_L g1261 ( .A(n_1260), .Y(n_1261) );
XNOR2xp5_ASAP7_75t_L g1262 ( .A(n_1261), .B(n_1192), .Y(n_1262) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1262), .Y(n_1263) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1263), .Y(n_1264) );
AOI21xp5_ASAP7_75t_L g1265 ( .A1(n_1264), .A2(n_1202), .B(n_1197), .Y(n_1265) );
endmodule