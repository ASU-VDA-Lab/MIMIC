module fake_jpeg_9728_n_204 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_204);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_14;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_31),
.B(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_0),
.Y(n_33)
);

AND2x2_ASAP7_75t_SL g44 ( 
.A(n_33),
.B(n_25),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_21),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_35),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_44),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_27),
.A2(n_30),
.B1(n_29),
.B2(n_25),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_30),
.B1(n_27),
.B2(n_20),
.Y(n_55)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_53),
.Y(n_67)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_55),
.A2(n_56),
.B1(n_42),
.B2(n_22),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_36),
.A2(n_22),
.B1(n_23),
.B2(n_26),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_33),
.B(n_31),
.C(n_17),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_57),
.B(n_43),
.Y(n_74)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_59),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_44),
.B(n_33),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_28),
.Y(n_81)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_52),
.A2(n_40),
.B1(n_36),
.B2(n_26),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_68),
.A2(n_50),
.B1(n_23),
.B2(n_64),
.Y(n_97)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_71),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_61),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_73),
.A2(n_72),
.B1(n_70),
.B2(n_76),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_76),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_60),
.B(n_32),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_77),
.Y(n_87)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_60),
.B(n_16),
.Y(n_77)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_63),
.B(n_23),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_54),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_83),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_46),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_84),
.A2(n_97),
.B1(n_99),
.B2(n_28),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_83),
.A2(n_15),
.B1(n_21),
.B2(n_65),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_75),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_91),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_77),
.Y(n_105)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_67),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_92),
.B(n_93),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_66),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_95),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_66),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_98),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_68),
.A2(n_50),
.B1(n_28),
.B2(n_58),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_58),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_100),
.Y(n_115)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_74),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_102),
.B(n_106),
.Y(n_125)
);

AND2x6_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_81),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_103),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_105),
.A2(n_111),
.B(n_88),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_38),
.C(n_46),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_84),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_110),
.A2(n_111),
.B1(n_107),
.B2(n_108),
.Y(n_134)
);

NAND2x1p5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_38),
.Y(n_111)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_82),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_114),
.B(n_117),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_85),
.Y(n_116)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_0),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_106),
.B(n_117),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_112),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_126),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_104),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_90),
.Y(n_127)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_109),
.Y(n_135)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_130),
.Y(n_142)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_103),
.A2(n_87),
.B1(n_91),
.B2(n_49),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_131),
.A2(n_134),
.B1(n_110),
.B2(n_101),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_111),
.A2(n_87),
.B(n_2),
.C(n_3),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_102),
.Y(n_136)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_133),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_79),
.C(n_28),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_143),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_107),
.Y(n_140)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_141),
.Y(n_159)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_144),
.B(n_147),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_119),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_146),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_124),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_121),
.A2(n_113),
.B(n_2),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_149),
.Y(n_154)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_138),
.A2(n_125),
.B1(n_128),
.B2(n_118),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_150),
.A2(n_157),
.B1(n_1),
.B2(n_4),
.Y(n_168)
);

AO22x2_ASAP7_75t_L g151 ( 
.A1(n_146),
.A2(n_123),
.B1(n_132),
.B2(n_82),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_142),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_162),
.Y(n_163)
);

A2O1A1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_136),
.A2(n_123),
.B(n_3),
.C(n_4),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_160),
.C(n_144),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_79),
.C(n_18),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_11),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_140),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_164),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_167),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_161),
.A2(n_147),
.B1(n_139),
.B2(n_141),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_168),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_150),
.B(n_18),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_9),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_1),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_18),
.C(n_14),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_171),
.C(n_155),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_14),
.C(n_13),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_157),
.B(n_1),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_151),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_174),
.B(n_175),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_163),
.B(n_159),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_178),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_173),
.B(n_151),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_173),
.Y(n_180)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_180),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_4),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_177),
.Y(n_185)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_185),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_180),
.A2(n_154),
.B(n_178),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_188),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_151),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_189),
.B(n_5),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_6),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_187),
.A2(n_167),
.B(n_13),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_191),
.B(n_194),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_183),
.A2(n_13),
.B(n_14),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_195),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_184),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_196),
.A2(n_197),
.B(n_6),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_184),
.Y(n_197)
);

O2A1O1Ixp33_ASAP7_75t_SL g201 ( 
.A1(n_199),
.A2(n_7),
.B(n_8),
.C(n_198),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_201),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_202),
.A2(n_200),
.B(n_7),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_7),
.Y(n_204)
);


endmodule