module real_jpeg_9030_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_265, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_265;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_249;
wire n_78;
wire n_215;
wire n_176;
wire n_221;
wire n_166;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_1),
.A2(n_40),
.B1(n_42),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_1),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_1),
.A2(n_54),
.B1(n_55),
.B2(n_62),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_62),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_2),
.Y(n_26)
);

AOI21xp33_ASAP7_75t_L g205 ( 
.A1(n_2),
.A2(n_9),
.B(n_25),
.Y(n_205)
);

BUFx10_ASAP7_75t_L g82 ( 
.A(n_3),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_5),
.A2(n_54),
.B1(n_55),
.B2(n_58),
.Y(n_53)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_5),
.A2(n_40),
.B(n_53),
.C(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_5),
.B(n_40),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_5),
.A2(n_9),
.B(n_55),
.Y(n_147)
);

BUFx6f_ASAP7_75t_SL g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_8),
.A2(n_11),
.B1(n_20),
.B2(n_21),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_8),
.A2(n_20),
.B1(n_24),
.B2(n_25),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_8),
.A2(n_20),
.B1(n_40),
.B2(n_42),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_8),
.A2(n_20),
.B1(n_54),
.B2(n_55),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_9),
.A2(n_11),
.B1(n_21),
.B2(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_29),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_9),
.A2(n_29),
.B1(n_40),
.B2(n_42),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_9),
.A2(n_29),
.B1(n_54),
.B2(n_55),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_9),
.B(n_73),
.Y(n_165)
);

O2A1O1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_9),
.A2(n_24),
.B(n_39),
.C(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_9),
.B(n_22),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_37),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_10),
.A2(n_37),
.B1(n_40),
.B2(n_42),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_10),
.A2(n_37),
.B1(n_54),
.B2(n_55),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_11),
.Y(n_21)
);

A2O1A1Ixp33_ASAP7_75t_L g30 ( 
.A1(n_11),
.A2(n_23),
.B(n_26),
.C(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_11),
.B(n_26),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_11),
.A2(n_26),
.B(n_29),
.C(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_105),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_104),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_91),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_16),
.B(n_91),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_65),
.C(n_74),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_17),
.B(n_65),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_32),
.B1(n_33),
.B2(n_64),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_18),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_18),
.A2(n_64),
.B1(n_93),
.B2(n_102),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_18),
.A2(n_64),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_18),
.B(n_118),
.C(n_198),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_18),
.A2(n_64),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_18),
.B(n_229),
.C(n_231),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_22),
.B(n_27),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_19),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_23),
.B(n_30),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_23),
.A2(n_28),
.B1(n_30),
.B2(n_95),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_24),
.A2(n_38),
.B(n_39),
.C(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_24),
.B(n_39),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_28),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_29),
.A2(n_42),
.B(n_58),
.C(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_29),
.B(n_81),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_29),
.B(n_53),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_SL g176 ( 
.A1(n_29),
.A2(n_40),
.B(n_43),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_49),
.B1(n_50),
.B2(n_63),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_34),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_38),
.B(n_44),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_36),
.A2(n_71),
.B1(n_73),
.B2(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_39),
.Y(n_43)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_45),
.A2(n_70),
.B(n_73),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_46),
.B(n_233),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_47),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_49),
.A2(n_50),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_49),
.B(n_63),
.C(n_64),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_61),
.Y(n_50)
);

INVxp33_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_52),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_59),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_53),
.A2(n_59),
.B1(n_61),
.B2(n_67),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_53),
.A2(n_67),
.B(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_53),
.A2(n_59),
.B1(n_87),
.B2(n_117),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_53),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_54),
.B(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_81),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx24_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_65),
.A2(n_66),
.B(n_68),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_68),
.A2(n_69),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_68),
.A2(n_69),
.B1(n_94),
.B2(n_101),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_69),
.B(n_136),
.C(n_187),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_69),
.B(n_101),
.C(n_221),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_71),
.B(n_73),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_74),
.A2(n_75),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_83),
.B(n_88),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_76),
.A2(n_88),
.B1(n_123),
.B2(n_124),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_76),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_76),
.A2(n_84),
.B1(n_123),
.B2(n_249),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_78),
.B(n_140),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_79),
.A2(n_82),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_80),
.B(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_80),
.A2(n_81),
.B1(n_138),
.B2(n_140),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_81),
.A2(n_216),
.B(n_217),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_82),
.A2(n_137),
.B(n_139),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_83),
.B(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_84),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_86),
.A2(n_143),
.B(n_144),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_87),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_88),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_103),
.Y(n_91)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_96),
.B1(n_97),
.B2(n_101),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_94),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_94),
.A2(n_101),
.B1(n_118),
.B2(n_173),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_110),
.C(n_118),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_128),
.B(n_263),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_125),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_107),
.B(n_125),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_119),
.C(n_120),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_108),
.A2(n_109),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_110),
.A2(n_111),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_115),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_112),
.A2(n_115),
.B1(n_116),
.B2(n_227),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_112),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_113),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_115),
.A2(n_116),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_115),
.A2(n_116),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_116),
.B(n_156),
.C(n_164),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_116),
.B(n_183),
.C(n_190),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_118),
.A2(n_142),
.B1(n_148),
.B2(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_118),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_118),
.B(n_142),
.C(n_178),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_118),
.A2(n_173),
.B1(n_198),
.B2(n_200),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_119),
.A2(n_120),
.B1(n_121),
.B2(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_119),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_126),
.Y(n_127)
);

AOI321xp33_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_238),
.A3(n_251),
.B1(n_257),
.B2(n_262),
.C(n_265),
.Y(n_128)
);

NOR3xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_210),
.C(n_235),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_192),
.B(n_209),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_180),
.B(n_191),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_168),
.B(n_179),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_159),
.B(n_167),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_149),
.B(n_158),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_141),
.Y(n_135)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_136),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_136),
.B(n_141),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_136),
.A2(n_151),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_139),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_145),
.B1(n_146),
.B2(n_148),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_142),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_142),
.B(n_146),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_142),
.A2(n_148),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_148),
.B(n_215),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_154),
.B(n_157),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_155),
.B(n_156),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_156),
.A2(n_162),
.B1(n_163),
.B2(n_166),
.Y(n_161)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_156),
.A2(n_166),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_156),
.B(n_203),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_160),
.B(n_161),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_169),
.B(n_170),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_174),
.B2(n_178),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_174),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_177),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_181),
.B(n_182),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_188),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_189),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_193),
.B(n_194),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_201),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_195),
.B(n_202),
.C(n_208),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_198),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_202),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_206),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

AOI21xp33_ASAP7_75t_L g258 ( 
.A1(n_211),
.A2(n_259),
.B(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_222),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_212),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_212),
.B(n_222),
.Y(n_260)
);

FAx1_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_218),
.CI(n_219),
.CON(n_212),
.SN(n_212)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_225),
.B2(n_234),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_223),
.Y(n_234)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_228),
.C(n_234),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_237),
.Y(n_259)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_239),
.A2(n_258),
.B(n_261),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_240),
.B(n_241),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_250),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_247),
.B2(n_248),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_248),
.C(n_250),
.Y(n_252)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_253),
.Y(n_262)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);


endmodule