module fake_jpeg_31382_n_156 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_156);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_156;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_16),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_20),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_31),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx16f_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_1),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_71),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

CKINVDCx6p67_ASAP7_75t_R g72 ( 
.A(n_66),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_64),
.A2(n_60),
.B1(n_44),
.B2(n_58),
.Y(n_76)
);

AND2x4_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_45),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_42),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_83),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_82),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_71),
.B(n_57),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_58),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_84),
.A2(n_75),
.B1(n_81),
.B2(n_77),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_85),
.A2(n_86),
.B1(n_0),
.B2(n_1),
.Y(n_116)
);

AO22x2_ASAP7_75t_L g86 ( 
.A1(n_72),
.A2(n_62),
.B1(n_55),
.B2(n_58),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_78),
.B(n_43),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_52),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_72),
.A2(n_81),
.B1(n_77),
.B2(n_78),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_62),
.B1(n_55),
.B2(n_53),
.Y(n_105)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_90),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_56),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_48),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_82),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_94),
.B(n_95),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_82),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_98),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_3),
.Y(n_118)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_50),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_104),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_100),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_103),
.B(n_109),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_51),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_54),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_110),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_118),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_85),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_47),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_114),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_86),
.A2(n_49),
.B1(n_42),
.B2(n_2),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_113),
.A2(n_116),
.B1(n_4),
.B2(n_7),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_86),
.B(n_0),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_3),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_117),
.B(n_11),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_120),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_116),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_124),
.Y(n_140)
);

NOR4xp25_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_25),
.C(n_39),
.D(n_35),
.Y(n_126)
);

NAND3xp33_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_128),
.C(n_134),
.Y(n_139)
);

AO22x1_ASAP7_75t_L g128 ( 
.A1(n_113),
.A2(n_23),
.B1(n_32),
.B2(n_27),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_130),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_22),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_119),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_120),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_135)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_135),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_15),
.Y(n_136)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_132),
.Y(n_142)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_142),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_L g144 ( 
.A1(n_140),
.A2(n_128),
.B1(n_133),
.B2(n_121),
.Y(n_144)
);

OAI21x1_ASAP7_75t_L g149 ( 
.A1(n_144),
.A2(n_138),
.B(n_139),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_143),
.B(n_130),
.C(n_127),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_146),
.B(n_147),
.C(n_122),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_137),
.A2(n_129),
.B1(n_118),
.B2(n_111),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_148),
.A2(n_149),
.B(n_145),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_139),
.C(n_141),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_123),
.C(n_125),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_152),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);

BUFx24_ASAP7_75t_SL g155 ( 
.A(n_154),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_144),
.Y(n_156)
);


endmodule