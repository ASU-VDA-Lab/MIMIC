module fake_jpeg_14307_n_429 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_429);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_429;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_47),
.B(n_48),
.Y(n_94)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_23),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_50),
.B(n_56),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_22),
.B(n_32),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_53),
.B(n_66),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_22),
.B(n_18),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_54),
.B(n_60),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g57 ( 
.A(n_23),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_57),
.B(n_71),
.Y(n_132)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_18),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_61),
.B(n_75),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_40),
.B(n_18),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

INVx2_ASAP7_75t_R g71 ( 
.A(n_26),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_26),
.B(n_15),
.Y(n_75)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_42),
.B(n_0),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_84),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_40),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_80),
.B(n_81),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_41),
.B(n_16),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_41),
.B(n_16),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_86),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_49),
.A2(n_31),
.B1(n_29),
.B2(n_37),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_90),
.A2(n_92),
.B1(n_98),
.B2(n_130),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_29),
.B1(n_31),
.B2(n_37),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_52),
.A2(n_36),
.B1(n_37),
.B2(n_35),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_75),
.A2(n_36),
.B1(n_25),
.B2(n_44),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_104),
.A2(n_108),
.B1(n_112),
.B2(n_121),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_76),
.A2(n_25),
.B1(n_44),
.B2(n_20),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_73),
.A2(n_64),
.B1(n_59),
.B2(n_45),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_76),
.A2(n_25),
.B1(n_43),
.B2(n_33),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_119),
.B(n_1),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_73),
.A2(n_43),
.B1(n_27),
.B2(n_24),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_55),
.A2(n_28),
.B1(n_20),
.B2(n_27),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_125),
.A2(n_126),
.B1(n_129),
.B2(n_58),
.Y(n_163)
);

OA22x2_ASAP7_75t_L g126 ( 
.A1(n_71),
.A2(n_28),
.B1(n_27),
.B2(n_24),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_68),
.A2(n_24),
.B1(n_19),
.B2(n_33),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_62),
.A2(n_19),
.B1(n_14),
.B2(n_13),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_85),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_135),
.B(n_138),
.Y(n_176)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_136),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_98),
.A2(n_79),
.B1(n_82),
.B2(n_51),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_127),
.A2(n_19),
.B(n_57),
.C(n_14),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_139),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_87),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_140),
.B(n_141),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_77),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_0),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_142),
.B(n_149),
.Y(n_200)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_143),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_69),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_144),
.Y(n_194)
);

INVx11_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_145),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_94),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_146),
.B(n_151),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_106),
.Y(n_147)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_159),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_113),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_104),
.B(n_63),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_83),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_158),
.Y(n_187)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_105),
.Y(n_155)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_132),
.A2(n_126),
.B1(n_67),
.B2(n_70),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_156),
.A2(n_122),
.B1(n_107),
.B2(n_133),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_89),
.B(n_0),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_99),
.B(n_74),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_134),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_160),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_99),
.B(n_72),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_106),
.Y(n_162)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_163),
.A2(n_171),
.B1(n_172),
.B2(n_95),
.Y(n_188)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_88),
.Y(n_164)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_164),
.Y(n_201)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_88),
.Y(n_165)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_165),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_122),
.B(n_100),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_170),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_103),
.B(n_114),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_168),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_119),
.B(n_1),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_169),
.Y(n_199)
);

INVx4_ASAP7_75t_SL g170 ( 
.A(n_120),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_129),
.A2(n_65),
.B1(n_10),
.B2(n_9),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_166),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_L g225 ( 
.A1(n_183),
.A2(n_146),
.B(n_167),
.Y(n_225)
);

OAI22x1_ASAP7_75t_L g185 ( 
.A1(n_152),
.A2(n_121),
.B1(n_112),
.B2(n_133),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_185),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_188),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_195),
.A2(n_154),
.B1(n_155),
.B2(n_144),
.Y(n_215)
);

AOI32xp33_ASAP7_75t_L g196 ( 
.A1(n_149),
.A2(n_91),
.A3(n_107),
.B1(n_102),
.B2(n_111),
.Y(n_196)
);

A2O1A1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_196),
.A2(n_168),
.B(n_144),
.C(n_154),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_163),
.A2(n_131),
.B1(n_115),
.B2(n_97),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_198),
.A2(n_152),
.B1(n_137),
.B2(n_151),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_197),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_204),
.B(n_205),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_197),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_202),
.Y(n_206)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_206),
.Y(n_231)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_202),
.Y(n_207)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_207),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_135),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_227),
.C(n_187),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_197),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_209),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_140),
.Y(n_211)
);

XNOR2x1_ASAP7_75t_L g248 ( 
.A(n_211),
.B(n_145),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_213),
.A2(n_194),
.B1(n_196),
.B2(n_185),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_158),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_216),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_215),
.A2(n_159),
.B1(n_161),
.B2(n_155),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_180),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_179),
.B(n_142),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_222),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_191),
.B(n_141),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_218),
.B(n_176),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_186),
.Y(n_219)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_219),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_186),
.Y(n_220)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_177),
.Y(n_221)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_221),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_138),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_174),
.A2(n_172),
.B(n_160),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_223),
.A2(n_191),
.B(n_194),
.Y(n_237)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_177),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_224),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_201),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_226),
.A2(n_183),
.B1(n_181),
.B2(n_200),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_153),
.Y(n_227)
);

INVxp33_ASAP7_75t_L g228 ( 
.A(n_193),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_228),
.Y(n_239)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_192),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_229),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_230),
.A2(n_235),
.B1(n_242),
.B2(n_246),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_234),
.B(n_252),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_203),
.A2(n_176),
.B1(n_185),
.B2(n_188),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_237),
.A2(n_222),
.B(n_223),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_240),
.B(n_243),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_241),
.A2(n_220),
.B(n_209),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_203),
.A2(n_198),
.B1(n_195),
.B2(n_184),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_212),
.A2(n_184),
.B1(n_173),
.B2(n_189),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_250),
.C(n_208),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_211),
.B(n_227),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_216),
.B(n_201),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_212),
.A2(n_173),
.B1(n_192),
.B2(n_175),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_254),
.A2(n_199),
.B1(n_210),
.B2(n_175),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_217),
.Y(n_268)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_256),
.Y(n_257)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_257),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_258),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_235),
.A2(n_230),
.B1(n_241),
.B2(n_247),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_259),
.B(n_266),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_219),
.Y(n_260)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_260),
.Y(n_289)
);

NAND2x1p5_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_264),
.Y(n_292)
);

INVxp33_ASAP7_75t_L g263 ( 
.A(n_249),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_263),
.A2(n_279),
.B1(n_238),
.B2(n_233),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_237),
.A2(n_213),
.B(n_204),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_264),
.A2(n_271),
.B(n_277),
.Y(n_310)
);

NAND4xp25_ASAP7_75t_SL g265 ( 
.A(n_253),
.B(n_170),
.C(n_95),
.D(n_147),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_265),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_247),
.A2(n_215),
.B1(n_214),
.B2(n_213),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_256),
.Y(n_267)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_267),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_268),
.A2(n_286),
.B1(n_236),
.B2(n_178),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_227),
.Y(n_269)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_269),
.Y(n_293)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_231),
.Y(n_270)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_270),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_244),
.A2(n_218),
.B(n_224),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_232),
.Y(n_299)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_231),
.Y(n_273)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_273),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_207),
.Y(n_274)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_274),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_251),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_275),
.B(n_278),
.Y(n_297)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_233),
.Y(n_276)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_276),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_245),
.A2(n_229),
.B(n_206),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_242),
.A2(n_226),
.B1(n_221),
.B2(n_208),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_239),
.B(n_210),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_280),
.B(n_282),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_243),
.A2(n_190),
.B(n_164),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_281),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_236),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_251),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_283),
.B(n_285),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_238),
.A2(n_165),
.B(n_190),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_254),
.A2(n_157),
.B1(n_150),
.B2(n_139),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_274),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_288),
.B(n_292),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_250),
.C(n_240),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_295),
.B(n_305),
.C(n_309),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_248),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_298),
.B(n_299),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_303),
.A2(n_307),
.B1(n_285),
.B2(n_282),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_232),
.C(n_246),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_269),
.B(n_143),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_266),
.B(n_199),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_312),
.C(n_281),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_278),
.B(n_178),
.C(n_169),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_289),
.B(n_284),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_315),
.B(n_318),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_262),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_316),
.B(n_321),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_293),
.B(n_284),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_304),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_319),
.B(n_327),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_295),
.B(n_259),
.C(n_258),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_322),
.B(n_329),
.C(n_331),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_297),
.B(n_280),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_323),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_291),
.A2(n_275),
.B1(n_283),
.B2(n_268),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_324),
.Y(n_351)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_313),
.Y(n_325)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_325),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_300),
.A2(n_260),
.B(n_271),
.Y(n_326)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_326),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_308),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_300),
.A2(n_261),
.B1(n_279),
.B2(n_286),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_328),
.A2(n_296),
.B1(n_308),
.B2(n_310),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_305),
.B(n_298),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_293),
.B(n_261),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_330),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_302),
.B(n_309),
.C(n_292),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_292),
.B(n_277),
.C(n_267),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_333),
.B(n_337),
.C(n_338),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_291),
.A2(n_276),
.B1(n_273),
.B2(n_270),
.Y(n_334)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_334),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_297),
.B(n_257),
.Y(n_335)
);

INVx13_ASAP7_75t_L g340 ( 
.A(n_335),
.Y(n_340)
);

XNOR2x1_ASAP7_75t_L g339 ( 
.A(n_336),
.B(n_307),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_312),
.B(n_265),
.C(n_139),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_311),
.B(n_150),
.C(n_157),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_339),
.B(n_170),
.Y(n_368)
);

BUFx12f_ASAP7_75t_SL g341 ( 
.A(n_322),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g374 ( 
.A(n_341),
.B(n_162),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_352),
.A2(n_353),
.B1(n_334),
.B2(n_333),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_328),
.A2(n_296),
.B1(n_310),
.B2(n_313),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_317),
.B(n_314),
.C(n_306),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_354),
.B(n_357),
.Y(n_367)
);

BUFx12_ASAP7_75t_L g355 ( 
.A(n_332),
.Y(n_355)
);

CKINVDCx14_ASAP7_75t_R g376 ( 
.A(n_355),
.Y(n_376)
);

XNOR2x1_ASAP7_75t_L g356 ( 
.A(n_316),
.B(n_331),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g373 ( 
.A(n_356),
.B(n_347),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_317),
.B(n_320),
.C(n_329),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_320),
.B(n_294),
.C(n_290),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_359),
.B(n_321),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_360),
.B(n_362),
.Y(n_386)
);

AO21x1_ASAP7_75t_L g379 ( 
.A1(n_361),
.A2(n_344),
.B(n_352),
.Y(n_379)
);

BUFx24_ASAP7_75t_SL g362 ( 
.A(n_342),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_346),
.Y(n_363)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_363),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_354),
.B(n_301),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_364),
.B(n_365),
.Y(n_388)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_345),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_350),
.A2(n_338),
.B1(n_337),
.B2(n_323),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_366),
.A2(n_369),
.B1(n_370),
.B2(n_368),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_368),
.B(n_373),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_349),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_351),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_357),
.B(n_97),
.C(n_131),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_371),
.B(n_372),
.C(n_375),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_359),
.B(n_96),
.C(n_115),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_374),
.A2(n_358),
.B(n_353),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_343),
.B(n_348),
.C(n_347),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_377),
.A2(n_371),
.B(n_105),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_379),
.B(n_91),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_376),
.A2(n_351),
.B1(n_344),
.B2(n_348),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_380),
.A2(n_101),
.B1(n_111),
.B2(n_102),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_361),
.A2(n_340),
.B1(n_339),
.B2(n_355),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_382),
.B(n_383),
.Y(n_399)
);

OAI321xp33_ASAP7_75t_L g385 ( 
.A1(n_374),
.A2(n_340),
.A3(n_355),
.B1(n_341),
.B2(n_356),
.C(n_343),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_385),
.B(n_389),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_375),
.B(n_367),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_387),
.B(n_390),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_373),
.B(n_109),
.C(n_136),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_372),
.A2(n_136),
.B1(n_147),
.B2(n_109),
.Y(n_390)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_391),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_392),
.B(n_393),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_387),
.B(n_10),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_386),
.A2(n_91),
.B(n_101),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_394),
.A2(n_398),
.B(n_377),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_381),
.B(n_10),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_395),
.B(n_396),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_378),
.B(n_1),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_397),
.B(n_400),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_380),
.A2(n_2),
.B(n_3),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_388),
.B(n_8),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_401),
.B(n_381),
.Y(n_403)
);

OR2x2_ASAP7_75t_L g415 ( 
.A(n_403),
.B(n_407),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_404),
.B(n_2),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_402),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_399),
.B(n_395),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_409),
.B(n_405),
.Y(n_417)
);

A2O1A1Ixp33_ASAP7_75t_L g410 ( 
.A1(n_396),
.A2(n_379),
.B(n_389),
.C(n_384),
.Y(n_410)
);

AO221x1_ASAP7_75t_L g419 ( 
.A1(n_410),
.A2(n_411),
.B1(n_412),
.B2(n_4),
.C(n_5),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_391),
.B(n_384),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_408),
.A2(n_8),
.B(n_3),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_413),
.A2(n_416),
.B(n_418),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_406),
.B(n_8),
.C(n_3),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_414),
.B(n_417),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_411),
.A2(n_7),
.B(n_4),
.Y(n_416)
);

AO21x1_ASAP7_75t_L g423 ( 
.A1(n_419),
.A2(n_7),
.B(n_5),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_415),
.A2(n_2),
.B(n_4),
.Y(n_421)
);

AOI21x1_ASAP7_75t_L g426 ( 
.A1(n_421),
.A2(n_6),
.B(n_420),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_419),
.B(n_2),
.C(n_5),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_422),
.B(n_423),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_426),
.B(n_6),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_427),
.A2(n_425),
.B(n_424),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_428),
.B(n_6),
.Y(n_429)
);


endmodule