module real_aes_10314_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_92;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_658;
wire n_676;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_456;
wire n_156;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_646;
wire n_650;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
NAND2xp5_ASAP7_75t_L g122 ( .A(n_0), .B(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g560 ( .A(n_1), .Y(n_560) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_1), .Y(n_574) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_2), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_3), .B(n_120), .Y(n_119) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_3), .Y(n_667) );
INVx2_ASAP7_75t_L g476 ( .A(n_4), .Y(n_476) );
BUFx2_ASAP7_75t_L g462 ( .A(n_5), .Y(n_462) );
INVx1_ASAP7_75t_L g556 ( .A(n_5), .Y(n_556) );
BUFx2_ASAP7_75t_L g585 ( .A(n_5), .Y(n_585) );
INVx1_ASAP7_75t_L g505 ( .A(n_6), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_6), .A2(n_57), .B1(n_531), .B2(n_539), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_7), .B(n_151), .Y(n_188) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_8), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g117 ( .A(n_9), .B(n_118), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_10), .B(n_112), .Y(n_183) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_11), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_12), .A2(n_65), .B1(n_513), .B2(n_515), .Y(n_512) );
AOI22xp33_ASAP7_75t_SL g568 ( .A1(n_12), .A2(n_65), .B1(n_546), .B2(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_13), .B(n_118), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_14), .A2(n_454), .B1(n_455), .B2(n_456), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_14), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_15), .B(n_169), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_16), .A2(n_66), .B1(n_478), .B2(n_486), .Y(n_477) );
OAI22xp33_ASAP7_75t_L g596 ( .A1(n_16), .A2(n_66), .B1(n_597), .B2(n_601), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_17), .B(n_118), .Y(n_202) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_18), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_19), .B(n_151), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_20), .B(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_21), .B(n_169), .Y(n_238) );
BUFx6f_ASAP7_75t_L g90 ( .A(n_22), .Y(n_90) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_23), .B(n_112), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_24), .B(n_185), .Y(n_233) );
INVx1_ASAP7_75t_L g460 ( .A(n_25), .Y(n_460) );
INVx1_ASAP7_75t_L g665 ( .A(n_25), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_26), .A2(n_46), .B1(n_515), .B2(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g618 ( .A(n_26), .Y(n_618) );
NAND2xp33_ASAP7_75t_SL g218 ( .A(n_27), .B(n_89), .Y(n_218) );
AOI22xp33_ASAP7_75t_SL g517 ( .A1(n_28), .A2(n_42), .B1(n_518), .B2(n_520), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_28), .A2(n_42), .B1(n_563), .B2(n_564), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_29), .B(n_172), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_30), .B(n_114), .Y(n_187) );
OAI21x1_ASAP7_75t_L g106 ( .A1(n_31), .A2(n_52), .B(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_32), .B(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g465 ( .A(n_33), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_33), .A2(n_55), .B1(n_546), .B2(n_550), .Y(n_545) );
AND2x6_ASAP7_75t_L g83 ( .A(n_34), .B(n_84), .Y(n_83) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_34), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_34), .B(n_625), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_35), .B(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_36), .B(n_143), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_37), .B(n_133), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_38), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_39), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_40), .Y(n_113) );
INVx1_ASAP7_75t_L g84 ( .A(n_41), .Y(n_84) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_41), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_43), .B(n_138), .Y(n_137) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_43), .Y(n_633) );
NAND2xp33_ASAP7_75t_L g216 ( .A(n_44), .B(n_89), .Y(n_216) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_45), .A2(n_68), .B1(n_581), .B2(n_583), .Y(n_580) );
INVx1_ASAP7_75t_L g608 ( .A(n_45), .Y(n_608) );
INVx1_ASAP7_75t_L g590 ( .A(n_46), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_47), .B(n_169), .Y(n_168) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_48), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_49), .B(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_50), .B(n_139), .Y(n_152) );
INVx2_ASAP7_75t_L g538 ( .A(n_51), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_53), .B(n_112), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_54), .B(n_133), .Y(n_165) );
INVx1_ASAP7_75t_L g491 ( .A(n_55), .Y(n_491) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_56), .Y(n_643) );
INVx1_ASAP7_75t_L g501 ( .A(n_57), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_58), .B(n_172), .Y(n_190) );
BUFx10_ASAP7_75t_L g659 ( .A(n_59), .Y(n_659) );
INVx2_ASAP7_75t_L g559 ( .A(n_60), .Y(n_559) );
INVx1_ASAP7_75t_L g575 ( .A(n_60), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g134 ( .A(n_61), .B(n_112), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_62), .B(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_63), .B(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_64), .B(n_118), .Y(n_164) );
INVx2_ASAP7_75t_L g107 ( .A(n_67), .Y(n_107) );
INVx1_ASAP7_75t_L g612 ( .A(n_68), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_69), .B(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_70), .B(n_185), .Y(n_184) );
CKINVDCx5p33_ASAP7_75t_R g635 ( .A(n_71), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_72), .B(n_151), .Y(n_157) );
INVx2_ASAP7_75t_L g535 ( .A(n_73), .Y(n_535) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_74), .Y(n_200) );
BUFx3_ASAP7_75t_L g470 ( .A(n_75), .Y(n_470) );
INVx1_ASAP7_75t_L g509 ( .A(n_75), .Y(n_509) );
BUFx3_ASAP7_75t_L g471 ( .A(n_76), .Y(n_471) );
INVx1_ASAP7_75t_L g504 ( .A(n_76), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_94), .B(n_452), .Y(n_77) );
BUFx3_ASAP7_75t_L g78 ( .A(n_79), .Y(n_78) );
AND2x2_ASAP7_75t_L g79 ( .A(n_80), .B(n_85), .Y(n_79) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
INVx2_ASAP7_75t_SL g141 ( .A(n_82), .Y(n_141) );
INVx8_ASAP7_75t_L g189 ( .A(n_82), .Y(n_189) );
INVx8_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
A2O1A1Ixp33_ASAP7_75t_L g108 ( .A1(n_83), .A2(n_109), .B(n_111), .C(n_116), .Y(n_108) );
OAI21x1_ASAP7_75t_SL g148 ( .A1(n_83), .A2(n_149), .B(n_154), .Y(n_148) );
OAI21x1_ASAP7_75t_L g162 ( .A1(n_83), .A2(n_163), .B(n_166), .Y(n_162) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_86), .Y(n_85) );
AO21x1_ASAP7_75t_L g676 ( .A1(n_86), .A2(n_677), .B(n_678), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g86 ( .A(n_87), .B(n_91), .Y(n_86) );
HB1xp67_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx2_ASAP7_75t_L g156 ( .A(n_89), .Y(n_156) );
BUFx6f_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
BUFx6f_ASAP7_75t_L g112 ( .A(n_90), .Y(n_112) );
INVx2_ASAP7_75t_L g114 ( .A(n_90), .Y(n_114) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_90), .Y(n_118) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_90), .Y(n_121) );
INVx1_ASAP7_75t_L g140 ( .A(n_90), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_92), .Y(n_91) );
AOI21xp5_ASAP7_75t_L g116 ( .A1(n_92), .A2(n_117), .B(n_119), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_92), .A2(n_155), .B(n_157), .Y(n_154) );
BUFx12f_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx5_ASAP7_75t_L g110 ( .A(n_93), .Y(n_110) );
INVx5_ASAP7_75t_L g153 ( .A(n_93), .Y(n_153) );
BUFx3_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
BUFx2_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
NAND3x2_ASAP7_75t_L g96 ( .A(n_97), .B(n_327), .C(n_406), .Y(n_96) );
AND2x2_ASAP7_75t_L g97 ( .A(n_98), .B(n_280), .Y(n_97) );
AOI211xp5_ASAP7_75t_SL g98 ( .A1(n_99), .A2(n_174), .B(n_221), .C(n_271), .Y(n_98) );
AND2x2_ASAP7_75t_L g99 ( .A(n_100), .B(n_125), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_101), .B(n_248), .Y(n_381) );
AND2x2_ASAP7_75t_L g412 ( .A(n_101), .B(n_145), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_101), .B(n_301), .Y(n_415) );
INVx4_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
NAND2x1_ASAP7_75t_L g247 ( .A(n_102), .B(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g299 ( .A(n_102), .B(n_260), .Y(n_299) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x2_ASAP7_75t_L g224 ( .A(n_103), .B(n_147), .Y(n_224) );
INVx3_ASAP7_75t_L g259 ( .A(n_103), .Y(n_259) );
AND2x2_ASAP7_75t_L g279 ( .A(n_103), .B(n_127), .Y(n_279) );
OA21x2_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_108), .B(n_122), .Y(n_103) );
OAI21x1_ASAP7_75t_L g180 ( .A1(n_104), .A2(n_181), .B(n_190), .Y(n_180) );
OAI21x1_ASAP7_75t_L g193 ( .A1(n_104), .A2(n_194), .B(n_203), .Y(n_193) );
OAI21x1_ASAP7_75t_L g230 ( .A1(n_104), .A2(n_231), .B(n_239), .Y(n_230) );
BUFx5_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g144 ( .A(n_105), .Y(n_144) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_105), .Y(n_240) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g124 ( .A(n_106), .Y(n_124) );
AOI21x1_ASAP7_75t_L g135 ( .A1(n_109), .A2(n_136), .B(n_137), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_109), .A2(n_218), .B(n_219), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_109), .A2(n_236), .B(n_238), .Y(n_235) );
INVx2_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g131 ( .A1(n_110), .A2(n_132), .B(n_134), .Y(n_131) );
INVx2_ASAP7_75t_SL g170 ( .A(n_110), .Y(n_170) );
O2A1O1Ixp33_ASAP7_75t_L g213 ( .A1(n_110), .A2(n_214), .B(n_215), .C(n_216), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_110), .A2(n_233), .B(n_234), .Y(n_232) );
OAI22xp33_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_113), .B1(n_114), .B2(n_115), .Y(n_111) );
INVx1_ASAP7_75t_L g215 ( .A(n_114), .Y(n_215) );
INVx2_ASAP7_75t_L g237 ( .A(n_114), .Y(n_237) );
INVx5_ASAP7_75t_L g133 ( .A(n_118), .Y(n_133) );
INVx1_ASAP7_75t_L g201 ( .A(n_120), .Y(n_201) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g169 ( .A(n_121), .Y(n_169) );
INVx2_ASAP7_75t_L g185 ( .A(n_121), .Y(n_185) );
INVx2_ASAP7_75t_L g197 ( .A(n_121), .Y(n_197) );
BUFx4f_ASAP7_75t_L g129 ( .A(n_123), .Y(n_129) );
OAI21x1_ASAP7_75t_L g147 ( .A1(n_123), .A2(n_148), .B(n_158), .Y(n_147) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g173 ( .A(n_124), .Y(n_173) );
INVx2_ASAP7_75t_L g390 ( .A(n_125), .Y(n_390) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_145), .Y(n_125) );
AND2x2_ASAP7_75t_L g223 ( .A(n_126), .B(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g315 ( .A(n_126), .Y(n_315) );
AND2x2_ASAP7_75t_L g411 ( .A(n_126), .B(n_412), .Y(n_411) );
INVx2_ASAP7_75t_SL g126 ( .A(n_127), .Y(n_126) );
AND2x4_ASAP7_75t_L g248 ( .A(n_127), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g258 ( .A(n_127), .B(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVxp67_ASAP7_75t_R g309 ( .A(n_128), .Y(n_309) );
OAI21x1_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_130), .B(n_142), .Y(n_128) );
OAI21xp5_ASAP7_75t_L g293 ( .A1(n_129), .A2(n_130), .B(n_142), .Y(n_293) );
OAI21x1_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_135), .B(n_141), .Y(n_130) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g151 ( .A(n_140), .Y(n_151) );
OAI21xp5_ASAP7_75t_L g194 ( .A1(n_141), .A2(n_195), .B(n_199), .Y(n_194) );
OAI21x1_ASAP7_75t_L g212 ( .A1(n_141), .A2(n_213), .B(n_217), .Y(n_212) );
OAI21x1_ASAP7_75t_L g161 ( .A1(n_143), .A2(n_162), .B(n_171), .Y(n_161) );
OAI21x1_ASAP7_75t_L g211 ( .A1(n_143), .A2(n_212), .B(n_220), .Y(n_211) );
INVx2_ASAP7_75t_SL g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g159 ( .A(n_144), .Y(n_159) );
AND2x2_ASAP7_75t_L g308 ( .A(n_145), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_160), .Y(n_145) );
INVx2_ASAP7_75t_SL g261 ( .A(n_146), .Y(n_261) );
INVx1_ASAP7_75t_L g267 ( .A(n_146), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_146), .B(n_259), .Y(n_288) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_146), .Y(n_320) );
INVx1_ASAP7_75t_L g366 ( .A(n_146), .Y(n_366) );
AND2x2_ASAP7_75t_L g387 ( .A(n_146), .B(n_340), .Y(n_387) );
INVxp67_ASAP7_75t_SL g402 ( .A(n_146), .Y(n_402) );
INVx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
O2A1O1Ixp33_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_151), .B(n_152), .C(n_153), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_153), .A2(n_164), .B(n_165), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_153), .A2(n_187), .B(n_188), .Y(n_186) );
O2A1O1Ixp5_ASAP7_75t_L g199 ( .A1(n_153), .A2(n_200), .B(n_201), .C(n_202), .Y(n_199) );
INVx1_ASAP7_75t_L g249 ( .A(n_160), .Y(n_249) );
AND2x2_ASAP7_75t_L g260 ( .A(n_160), .B(n_261), .Y(n_260) );
NOR2xp67_ASAP7_75t_L g266 ( .A(n_160), .B(n_267), .Y(n_266) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_160), .Y(n_278) );
AND2x2_ASAP7_75t_L g333 ( .A(n_160), .B(n_293), .Y(n_333) );
INVx1_ASAP7_75t_L g341 ( .A(n_160), .Y(n_341) );
INVx1_ASAP7_75t_L g403 ( .A(n_160), .Y(n_403) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_L g301 ( .A(n_161), .B(n_293), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_168), .B(n_170), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_170), .A2(n_183), .B(n_184), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_170), .A2(n_196), .B(n_198), .Y(n_195) );
INVx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_175), .B(n_204), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_176), .B(n_253), .Y(n_417) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g389 ( .A(n_177), .Y(n_389) );
OR2x2_ASAP7_75t_L g428 ( .A(n_177), .B(n_376), .Y(n_428) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AND2x2_ASAP7_75t_L g283 ( .A(n_178), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g360 ( .A(n_178), .B(n_312), .Y(n_360) );
AND2x2_ASAP7_75t_L g178 ( .A(n_179), .B(n_191), .Y(n_178) );
INVx2_ASAP7_75t_L g246 ( .A(n_179), .Y(n_246) );
AND2x2_ASAP7_75t_L g252 ( .A(n_179), .B(n_192), .Y(n_252) );
INVx1_ASAP7_75t_L g264 ( .A(n_179), .Y(n_264) );
INVx1_ASAP7_75t_L g375 ( .A(n_179), .Y(n_375) );
INVx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
OAI21x1_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_186), .B(n_189), .Y(n_181) );
OAI21x1_ASAP7_75t_L g231 ( .A1(n_189), .A2(n_232), .B(n_235), .Y(n_231) );
INVx1_ASAP7_75t_L g205 ( .A(n_191), .Y(n_205) );
AND2x2_ASAP7_75t_L g269 ( .A(n_191), .B(n_264), .Y(n_269) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_191), .Y(n_353) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx1_ASAP7_75t_L g326 ( .A(n_192), .Y(n_326) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g241 ( .A(n_193), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
AND2x2_ASAP7_75t_L g430 ( .A(n_206), .B(n_362), .Y(n_430) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx1_ASAP7_75t_L g274 ( .A(n_208), .Y(n_274) );
INVx1_ASAP7_75t_L g284 ( .A(n_208), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_208), .B(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g270 ( .A(n_209), .B(n_229), .Y(n_270) );
AND2x2_ASAP7_75t_L g410 ( .A(n_209), .B(n_245), .Y(n_410) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g244 ( .A(n_210), .Y(n_244) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_210), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_210), .B(n_229), .Y(n_348) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g322 ( .A(n_211), .B(n_246), .Y(n_322) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_211), .Y(n_422) );
OAI221xp5_ASAP7_75t_SL g221 ( .A1(n_222), .A2(n_225), .B1(n_247), .B2(n_250), .C(n_256), .Y(n_221) );
OAI32xp33_ASAP7_75t_L g424 ( .A1(n_222), .A2(n_322), .A3(n_425), .B1(n_427), .B2(n_428), .Y(n_424) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g358 ( .A(n_224), .B(n_333), .Y(n_358) );
AND2x2_ASAP7_75t_L g362 ( .A(n_224), .B(n_254), .Y(n_362) );
INVx1_ASAP7_75t_L g449 ( .A(n_224), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_226), .B(n_242), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_226), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g427 ( .A(n_226), .Y(n_427) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
OR2x2_ASAP7_75t_L g330 ( .A(n_227), .B(n_296), .Y(n_330) );
NAND2x1p5_ASAP7_75t_L g227 ( .A(n_228), .B(n_241), .Y(n_227) );
BUFx2_ASAP7_75t_L g262 ( .A(n_228), .Y(n_262) );
INVx2_ASAP7_75t_L g305 ( .A(n_228), .Y(n_305) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g255 ( .A(n_230), .Y(n_255) );
INVx2_ASAP7_75t_L g371 ( .A(n_241), .Y(n_371) );
INVx1_ASAP7_75t_L g302 ( .A(n_242), .Y(n_302) );
AOI322xp5_ASAP7_75t_L g343 ( .A1(n_242), .A2(n_344), .A3(n_346), .B1(n_347), .B2(n_349), .C1(n_350), .C2(n_351), .Y(n_343) );
AND2x4_ASAP7_75t_SL g439 ( .A(n_242), .B(n_376), .Y(n_439) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
OR2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
INVx1_ASAP7_75t_L g296 ( .A(n_244), .Y(n_296) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g426 ( .A(n_248), .Y(n_426) );
OAI221xp5_ASAP7_75t_L g306 ( .A1(n_250), .A2(n_307), .B1(n_310), .B2(n_313), .C(n_316), .Y(n_306) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
AND2x2_ASAP7_75t_L g273 ( .A(n_252), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g342 ( .A(n_252), .B(n_296), .Y(n_342) );
INVx1_ASAP7_75t_L g445 ( .A(n_252), .Y(n_445) );
INVx1_ASAP7_75t_L g282 ( .A(n_253), .Y(n_282) );
AND2x2_ASAP7_75t_L g380 ( .A(n_253), .B(n_269), .Y(n_380) );
BUFx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_254), .B(n_326), .Y(n_345) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
BUFx3_ASAP7_75t_L g324 ( .A(n_255), .Y(n_324) );
AOI32xp33_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_262), .A3(n_263), .B1(n_265), .B2(n_268), .Y(n_256) );
INVx1_ASAP7_75t_L g378 ( .A(n_257), .Y(n_378) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_260), .Y(n_257) );
AND2x4_ASAP7_75t_L g265 ( .A(n_258), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g404 ( .A(n_258), .Y(n_404) );
AND2x2_ASAP7_75t_L g335 ( .A(n_259), .B(n_261), .Y(n_335) );
INVx1_ASAP7_75t_L g340 ( .A(n_259), .Y(n_340) );
AND2x2_ASAP7_75t_L g451 ( .A(n_260), .B(n_279), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_262), .A2(n_272), .B(n_275), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_262), .B(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_263), .B(n_305), .Y(n_304) );
NAND2x1_ASAP7_75t_L g405 ( .A(n_263), .B(n_323), .Y(n_405) );
BUFx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g361 ( .A1(n_265), .A2(n_289), .B(n_362), .Y(n_361) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_267), .Y(n_276) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVx1_ASAP7_75t_L g297 ( .A(n_269), .Y(n_297) );
AND2x2_ASAP7_75t_L g311 ( .A(n_269), .B(n_312), .Y(n_311) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_269), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_269), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND3xp33_ASAP7_75t_SL g367 ( .A(n_275), .B(n_368), .C(n_372), .Y(n_367) );
INVx2_ASAP7_75t_L g392 ( .A(n_275), .Y(n_392) );
OR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
OR2x2_ASAP7_75t_L g425 ( .A(n_276), .B(n_426), .Y(n_425) );
BUFx3_ASAP7_75t_L g303 ( .A(n_277), .Y(n_303) );
NAND2x1_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
AOI311xp33_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_285), .A3(n_289), .B(n_294), .C(n_306), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
BUFx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_287), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g314 ( .A(n_287), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_288), .B(n_315), .Y(n_349) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g399 ( .A(n_291), .B(n_387), .Y(n_399) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g365 ( .A(n_292), .B(n_366), .Y(n_365) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_292), .Y(n_448) );
BUFx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OAI222xp33_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_298), .B1(n_300), .B2(n_302), .C1(n_303), .C2(n_304), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
OR2x2_ASAP7_75t_L g356 ( .A(n_296), .B(n_345), .Y(n_356) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_301), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g350 ( .A(n_301), .B(n_320), .Y(n_350) );
AND2x2_ASAP7_75t_L g386 ( .A(n_301), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g396 ( .A(n_301), .B(n_335), .Y(n_396) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OAI21xp5_ASAP7_75t_L g316 ( .A1(n_308), .A2(n_317), .B(n_321), .Y(n_316) );
AND2x2_ASAP7_75t_L g337 ( .A(n_309), .B(n_335), .Y(n_337) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVxp67_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_322), .B(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g436 ( .A(n_322), .B(n_437), .Y(n_436) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_322), .Y(n_450) );
INVxp67_ASAP7_75t_SL g384 ( .A(n_323), .Y(n_384) );
AND2x4_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx3_ASAP7_75t_L g376 ( .A(n_324), .Y(n_376) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_324), .Y(n_437) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND3x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_363), .C(n_391), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_329), .B(n_355), .Y(n_328) );
OAI211xp5_ASAP7_75t_SL g329 ( .A1(n_330), .A2(n_331), .B(n_336), .C(n_343), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_331), .B(n_447), .Y(n_446) );
OR2x6_ASAP7_75t_L g331 ( .A(n_332), .B(n_334), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g346 ( .A(n_334), .Y(n_346) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OAI21xp33_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_338), .B(n_342), .Y(n_336) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g364 ( .A(n_339), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_341), .Y(n_433) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_347), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVxp67_ASAP7_75t_L g354 ( .A(n_348), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_350), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_354), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_357), .B1(n_359), .B2(n_361), .Y(n_355) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AOI211xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_367), .B(n_377), .C(n_382), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_368), .A2(n_378), .B1(n_379), .B2(n_381), .Y(n_377) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_376), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OR2x2_ASAP7_75t_L g421 ( .A(n_375), .B(n_422), .Y(n_421) );
INVx2_ASAP7_75t_SL g395 ( .A(n_376), .Y(n_395) );
NOR2x1_ASAP7_75t_L g444 ( .A(n_376), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OAI22xp33_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_385), .B1(n_388), .B2(n_390), .Y(n_382) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_393), .B1(n_394), .B2(n_396), .C(n_397), .Y(n_391) );
AOI21xp33_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_400), .B(n_405), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
OR2x6_ASAP7_75t_L g400 ( .A(n_401), .B(n_404), .Y(n_400) );
INVxp67_ASAP7_75t_SL g423 ( .A(n_401), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
AND4x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_413), .C(n_429), .D(n_441), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_408), .B(n_411), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g440 ( .A(n_412), .Y(n_440) );
AOI221xp5_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_416), .B1(n_418), .B2(n_423), .C(n_424), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVxp67_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AOI21xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_431), .B(n_434), .Y(n_429) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AOI21xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_438), .B(n_440), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_446), .B1(n_450), .B2(n_451), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OR2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
OAI221xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_455), .B1(n_623), .B2(n_628), .C(n_670), .Y(n_452) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_455), .A2(n_667), .B1(n_671), .B2(n_675), .Y(n_670) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AO211x2_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_463), .B(n_510), .C(n_588), .Y(n_457) );
AND2x4_ASAP7_75t_L g458 ( .A(n_459), .B(n_461), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g528 ( .A(n_460), .B(n_476), .Y(n_528) );
AND2x4_ASAP7_75t_L g586 ( .A(n_460), .B(n_587), .Y(n_586) );
BUFx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g526 ( .A(n_462), .Y(n_526) );
NAND3xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_490), .C(n_500), .Y(n_463) );
AOI211xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_466), .B(n_472), .C(n_477), .Y(n_464) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND2x4_ASAP7_75t_L g472 ( .A(n_468), .B(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g516 ( .A(n_468), .Y(n_516) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
INVx2_ASAP7_75t_L g489 ( .A(n_470), .Y(n_489) );
AND2x4_ASAP7_75t_L g503 ( .A(n_470), .B(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g485 ( .A(n_471), .Y(n_485) );
AND2x4_ASAP7_75t_L g508 ( .A(n_471), .B(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x6_ASAP7_75t_L g502 ( .A(n_474), .B(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x6_ASAP7_75t_L g487 ( .A(n_475), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_476), .Y(n_481) );
INVx1_ASAP7_75t_L g494 ( .A(n_476), .Y(n_494) );
INVx2_ASAP7_75t_L g587 ( .A(n_476), .Y(n_587) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x4_ASAP7_75t_L g479 ( .A(n_480), .B(n_482), .Y(n_479) );
AND2x4_ASAP7_75t_L g499 ( .A(n_480), .B(n_497), .Y(n_499) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g657 ( .A(n_484), .Y(n_657) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x4_ASAP7_75t_L g497 ( .A(n_485), .B(n_489), .Y(n_497) );
INVx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_492), .B1(n_498), .B2(n_499), .Y(n_490) );
AND2x4_ASAP7_75t_L g492 ( .A(n_493), .B(n_495), .Y(n_492) );
AND2x6_ASAP7_75t_L g506 ( .A(n_493), .B(n_507), .Y(n_506) );
INVx1_ASAP7_75t_SL g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx2_ASAP7_75t_L g514 ( .A(n_496), .Y(n_514) );
BUFx6f_ASAP7_75t_L g579 ( .A(n_496), .Y(n_579) );
INVx6_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AOI22xp33_ASAP7_75t_SL g613 ( .A1(n_498), .A2(n_614), .B1(n_618), .B2(n_619), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_502), .B1(n_505), .B2(n_506), .Y(n_500) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_503), .Y(n_519) );
INVx2_ASAP7_75t_SL g582 ( .A(n_503), .Y(n_582) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g523 ( .A(n_508), .Y(n_523) );
NAND4xp25_ASAP7_75t_L g510 ( .A(n_511), .B(n_529), .C(n_561), .D(n_576), .Y(n_510) );
NAND3xp33_ASAP7_75t_L g511 ( .A(n_512), .B(n_517), .C(n_524), .Y(n_511) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx3_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx4f_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g583 ( .A(n_521), .Y(n_583) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
AND2x4_ASAP7_75t_L g571 ( .A(n_526), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_SL g653 ( .A(n_528), .Y(n_653) );
NAND3xp33_ASAP7_75t_L g529 ( .A(n_530), .B(n_545), .C(n_553), .Y(n_529) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
BUFx2_ASAP7_75t_L g563 ( .A(n_533), .Y(n_563) );
AND2x4_ASAP7_75t_L g605 ( .A(n_533), .B(n_606), .Y(n_605) );
AND2x4_ASAP7_75t_L g533 ( .A(n_534), .B(n_536), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AND2x4_ASAP7_75t_L g543 ( .A(n_535), .B(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g549 ( .A(n_535), .B(n_538), .Y(n_549) );
INVx1_ASAP7_75t_L g552 ( .A(n_535), .Y(n_552) );
INVx1_ASAP7_75t_L g603 ( .A(n_535), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_535), .B(n_538), .Y(n_617) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g544 ( .A(n_538), .Y(n_544) );
INVx1_ASAP7_75t_L g600 ( .A(n_538), .Y(n_600) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx3_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx3_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g567 ( .A(n_543), .Y(n_567) );
INVx1_ASAP7_75t_L g611 ( .A(n_543), .Y(n_611) );
AND2x4_ASAP7_75t_L g551 ( .A(n_544), .B(n_552), .Y(n_551) );
BUFx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
INVx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx2_ASAP7_75t_SL g592 ( .A(n_550), .Y(n_592) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_551), .Y(n_570) );
AND2x4_ASAP7_75t_L g593 ( .A(n_551), .B(n_594), .Y(n_593) );
INVx5_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
OR2x6_ASAP7_75t_L g554 ( .A(n_555), .B(n_557), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2x1p5_ASAP7_75t_L g557 ( .A(n_558), .B(n_560), .Y(n_557) );
INVx1_ASAP7_75t_L g595 ( .A(n_558), .Y(n_595) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g607 ( .A(n_559), .Y(n_607) );
NAND3xp33_ASAP7_75t_L g561 ( .A(n_562), .B(n_568), .C(n_571), .Y(n_561) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_573), .Y(n_622) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx2_ASAP7_75t_SL g599 ( .A(n_575), .Y(n_599) );
OR2x2_ASAP7_75t_L g601 ( .A(n_575), .B(n_602), .Y(n_601) );
NAND3xp33_ASAP7_75t_L g576 ( .A(n_577), .B(n_580), .C(n_584), .Y(n_576) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x4_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
OR2x6_ASAP7_75t_L g621 ( .A(n_585), .B(n_622), .Y(n_621) );
AND2x4_ASAP7_75t_L g663 ( .A(n_587), .B(n_664), .Y(n_663) );
AOI31xp33_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_604), .A3(n_613), .B(n_621), .Y(n_588) );
AOI211xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B(n_593), .C(n_596), .Y(n_589) );
INVx2_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x4_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
OR2x6_ASAP7_75t_L g615 ( .A(n_599), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AOI22xp33_ASAP7_75t_SL g604 ( .A1(n_605), .A2(n_608), .B1(n_609), .B2(n_612), .Y(n_604) );
AND2x4_ASAP7_75t_L g609 ( .A(n_606), .B(n_610), .Y(n_609) );
OR2x6_ASAP7_75t_L g620 ( .A(n_606), .B(n_616), .Y(n_620) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx8_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
BUFx6f_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx5_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
BUFx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_625), .B(n_627), .Y(n_649) );
INVx1_ASAP7_75t_SL g677 ( .A(n_625), .Y(n_677) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_645), .B1(n_667), .B2(n_668), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_629), .A2(n_667), .B1(n_672), .B2(n_673), .Y(n_671) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_631), .B1(n_636), .B2(n_637), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_633), .B1(n_634), .B2(n_635), .Y(n_631) );
CKINVDCx5p33_ASAP7_75t_R g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_639), .B1(n_640), .B2(n_644), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g644 ( .A(n_640), .Y(n_644) );
XNOR2xp5_ASAP7_75t_SL g640 ( .A(n_641), .B(n_642), .Y(n_640) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx8_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx8_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
CKINVDCx20_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
BUFx6f_ASAP7_75t_L g672 ( .A(n_648), .Y(n_672) );
OR2x6_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
OR2x4_ASAP7_75t_L g669 ( .A(n_649), .B(n_651), .Y(n_669) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AOI31xp33_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_654), .A3(n_658), .B(n_660), .Y(n_651) );
BUFx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVxp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g666 ( .A(n_657), .Y(n_666) );
INVx6_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVxp67_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
INVx2_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
AND2x4_ASAP7_75t_L g662 ( .A(n_663), .B(n_666), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx8_ASAP7_75t_L g674 ( .A(n_669), .Y(n_674) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
BUFx2_ASAP7_75t_SL g675 ( .A(n_676), .Y(n_675) );
endmodule