module fake_jpeg_30329_n_105 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_105);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_105;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_10),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_22),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_24),
.A2(n_28),
.B1(n_5),
.B2(n_7),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_20),
.B(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_16),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_1),
.C(n_3),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_32),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_20),
.A2(n_22),
.B1(n_15),
.B2(n_16),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_1),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_31),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_9),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_37),
.Y(n_43)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

AOI21xp33_ASAP7_75t_SL g36 ( 
.A1(n_23),
.A2(n_5),
.B(n_6),
.Y(n_36)
);

AOI21xp33_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_13),
.B(n_6),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_46),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_36),
.A2(n_21),
.B1(n_12),
.B2(n_18),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_14),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_56),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_30),
.A2(n_21),
.B1(n_12),
.B2(n_18),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_SL g62 ( 
.A(n_48),
.B(n_49),
.C(n_54),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_30),
.A2(n_21),
.B1(n_14),
.B2(n_13),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_52),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_26),
.B(n_27),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_32),
.B1(n_39),
.B2(n_56),
.Y(n_70)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_59),
.B(n_61),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_24),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_SL g63 ( 
.A(n_44),
.B(n_25),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_63),
.B(n_64),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_32),
.C(n_8),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_7),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_69),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_8),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_67),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_9),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_53),
.B1(n_41),
.B2(n_56),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_32),
.Y(n_71)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_68),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_77),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_78),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_71),
.B1(n_62),
.B2(n_61),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_80),
.Y(n_85)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_60),
.C(n_63),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_74),
.C(n_79),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_77),
.A2(n_58),
.B(n_67),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_85),
.Y(n_96)
);

OAI22x1_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_64),
.B1(n_57),
.B2(n_41),
.Y(n_88)
);

AOI21xp33_ASAP7_75t_L g92 ( 
.A1(n_88),
.A2(n_74),
.B(n_78),
.Y(n_92)
);

AO21x1_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_38),
.B(n_51),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_75),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_91),
.B(n_92),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_86),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_93),
.B(n_94),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_73),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_95),
.A2(n_96),
.B1(n_88),
.B2(n_90),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_98),
.A2(n_99),
.B1(n_95),
.B2(n_50),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_94),
.A2(n_90),
.B1(n_89),
.B2(n_72),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_100),
.A2(n_98),
.B(n_97),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_101),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_99),
.Y(n_104)
);

AOI322xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_38),
.A3(n_40),
.B1(n_53),
.B2(n_102),
.C1(n_101),
.C2(n_100),
.Y(n_105)
);


endmodule