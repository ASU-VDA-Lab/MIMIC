module fake_jpeg_11731_n_38 (n_3, n_2, n_1, n_0, n_4, n_5, n_38);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_38;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NAND2xp5_ASAP7_75t_L g6 ( 
.A(n_2),
.B(n_5),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_0),
.Y(n_7)
);

BUFx2_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g13 ( 
.A(n_8),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_17),
.Y(n_18)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_15),
.B(n_1),
.Y(n_22)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_6),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_6),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_7),
.Y(n_26)
);

NAND3xp33_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_1),
.C(n_3),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_17),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_11),
.B(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_11),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_24),
.A2(n_25),
.B(n_26),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_25),
.A2(n_15),
.B(n_20),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_29),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_16),
.B1(n_14),
.B2(n_20),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_30),
.A2(n_13),
.B(n_19),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_13),
.B(n_31),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_7),
.Y(n_33)
);

AOI31xp67_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_10),
.A3(n_8),
.B(n_9),
.Y(n_35)
);

AOI31xp67_ASAP7_75t_SL g36 ( 
.A1(n_34),
.A2(n_35),
.A3(n_14),
.B(n_16),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_10),
.B(n_4),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_4),
.Y(n_38)
);


endmodule