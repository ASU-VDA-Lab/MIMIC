module fake_jpeg_23440_n_136 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_136);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx2_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_10),
.B(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_25),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_30),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_27),
.B(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_18),
.B(n_2),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_13),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_35),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_12),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_36),
.B(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_20),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_24),
.B1(n_23),
.B2(n_26),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_54),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_50),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_24),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_51),
.B(n_31),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_19),
.Y(n_52)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_33),
.A2(n_23),
.B(n_11),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_53),
.A2(n_38),
.B(n_14),
.Y(n_63)
);

OA21x2_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_24),
.B(n_29),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_56),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_67),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_41),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_66),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_49),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_43),
.B(n_37),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_43),
.B1(n_48),
.B2(n_46),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_51),
.B(n_34),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_71),
.B(n_75),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_78),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_54),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_58),
.A2(n_54),
.B1(n_49),
.B2(n_11),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_34),
.B1(n_38),
.B2(n_60),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_49),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_79),
.A2(n_21),
.B(n_14),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_56),
.Y(n_81)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_78),
.A2(n_67),
.B1(n_34),
.B2(n_66),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_83),
.A2(n_59),
.B1(n_38),
.B2(n_76),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_66),
.C(n_65),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_85),
.C(n_79),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_57),
.C(n_63),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_88),
.B1(n_75),
.B2(n_71),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_77),
.A2(n_60),
.B1(n_48),
.B2(n_62),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_91),
.Y(n_96)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_89),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_94),
.Y(n_109)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_36),
.C(n_13),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_29),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_87),
.A2(n_62),
.B1(n_18),
.B2(n_19),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_100),
.A2(n_101),
.B1(n_16),
.B2(n_21),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_83),
.B1(n_84),
.B2(n_90),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_37),
.Y(n_102)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_106),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_99),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_21),
.C(n_50),
.Y(n_115)
);

AOI321xp33_ASAP7_75t_L g108 ( 
.A1(n_97),
.A2(n_16),
.A3(n_21),
.B1(n_9),
.B2(n_10),
.C(n_8),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_111),
.Y(n_113)
);

AOI322xp5_ASAP7_75t_L g112 ( 
.A1(n_104),
.A2(n_96),
.A3(n_101),
.B1(n_98),
.B2(n_93),
.C1(n_100),
.C2(n_92),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_115),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_68),
.B1(n_50),
.B2(n_5),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_111),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_3),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_117),
.B(n_103),
.Y(n_121)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_118),
.B(n_21),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_121),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_107),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_122),
.A2(n_114),
.B(n_115),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_108),
.Y(n_123)
);

NOR2xp67_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_4),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_6),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_128),
.C(n_129),
.Y(n_131)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_126),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_120),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_119),
.C(n_5),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_132),
.B(n_4),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_134),
.Y(n_135)
);

INVxp33_ASAP7_75t_SL g134 ( 
.A(n_131),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_130),
.Y(n_136)
);


endmodule