module fake_jpeg_3510_n_147 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_147);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_147;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

CKINVDCx9p33_ASAP7_75t_R g54 ( 
.A(n_44),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_54),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_56),
.B(n_57),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_47),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_60),
.B(n_43),
.Y(n_79)
);

NOR2x1_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_49),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_56),
.A2(n_50),
.B1(n_45),
.B2(n_41),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_63),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_57),
.A2(n_41),
.B1(n_50),
.B2(n_42),
.Y(n_63)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_60),
.B(n_49),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_69),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_48),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_61),
.B(n_40),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_78),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_77),
.Y(n_88)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

OAI32xp33_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_37),
.A3(n_38),
.B1(n_18),
.B2(n_36),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_66),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_81),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_38),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_62),
.B(n_1),
.C(n_2),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_69),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_82),
.B(n_70),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_72),
.A2(n_64),
.B1(n_67),
.B2(n_59),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_94),
.Y(n_103)
);

AOI32xp33_ASAP7_75t_L g89 ( 
.A1(n_68),
.A2(n_67),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_73),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_72),
.A2(n_37),
.B1(n_3),
.B2(n_4),
.Y(n_90)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_72),
.A2(n_0),
.B1(n_4),
.B2(n_6),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_86),
.B(n_68),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_97),
.B(n_100),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_99),
.Y(n_114)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_87),
.B(n_80),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_87),
.B(n_8),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_102),
.Y(n_116)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_105),
.Y(n_117)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_95),
.A2(n_81),
.B(n_77),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_106),
.A2(n_88),
.B(n_9),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_75),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_108),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_85),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_76),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_21),
.C(n_34),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_110),
.B(n_10),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_108),
.A2(n_88),
.B(n_20),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_121),
.B(n_11),
.Y(n_131)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_119),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_8),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_120),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_10),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_107),
.C(n_22),
.Y(n_126)
);

INVxp33_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_123),
.A2(n_111),
.B1(n_117),
.B2(n_119),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_124),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_131),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_129),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_19),
.C(n_33),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_122),
.C(n_114),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_135),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_125),
.A2(n_111),
.B1(n_115),
.B2(n_116),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_134),
.A2(n_136),
.B1(n_130),
.B2(n_126),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_132),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_135)
);

OA21x2_ASAP7_75t_SL g138 ( 
.A1(n_136),
.A2(n_127),
.B(n_137),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_138),
.B(n_140),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_26),
.C(n_16),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_141),
.A2(n_32),
.B(n_17),
.C(n_25),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_143),
.B(n_28),
.Y(n_144)
);

OAI21x1_ASAP7_75t_SL g145 ( 
.A1(n_144),
.A2(n_35),
.B(n_142),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_14),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_139),
.Y(n_147)
);


endmodule