module fake_jpeg_7506_n_83 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_83);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_83;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_48;
wire n_46;
wire n_62;
wire n_43;
wire n_82;

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

CKINVDCx12_ASAP7_75t_R g47 ( 
.A(n_20),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_30),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_53),
.B(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_0),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_56),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_1),
.B(n_2),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_59),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_52),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_1),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_61),
.Y(n_67)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_3),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_42),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_54),
.A2(n_45),
.B1(n_51),
.B2(n_44),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_63),
.A2(n_69),
.B1(n_46),
.B2(n_39),
.Y(n_71)
);

OA21x2_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_11),
.B(n_14),
.Y(n_72)
);

AO22x1_ASAP7_75t_SL g69 ( 
.A1(n_53),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_15),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_67),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_75),
.B(n_66),
.Y(n_76)
);

A2O1A1O1Ixp25_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_69),
.B(n_65),
.C(n_73),
.D(n_68),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_77),
.B(n_72),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_78),
.A2(n_64),
.B1(n_18),
.B2(n_22),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_17),
.B(n_23),
.Y(n_80)
);

BUFx24_ASAP7_75t_SL g81 ( 
.A(n_80),
.Y(n_81)
);

MAJx2_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_24),
.C(n_25),
.Y(n_82)
);

AOI322xp5_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_26),
.A3(n_28),
.B1(n_31),
.B2(n_32),
.C1(n_33),
.C2(n_34),
.Y(n_83)
);


endmodule