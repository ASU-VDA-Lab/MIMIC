module real_jpeg_25716_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_1),
.A2(n_48),
.B1(n_56),
.B2(n_144),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_1),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_1),
.A2(n_51),
.B1(n_54),
.B2(n_144),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_144),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_1),
.A2(n_25),
.B1(n_28),
.B2(n_144),
.Y(n_272)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_3),
.A2(n_51),
.B1(n_54),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_3),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_72),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_3),
.A2(n_25),
.B1(n_28),
.B2(n_72),
.Y(n_132)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_5),
.A2(n_48),
.B1(n_56),
.B2(n_160),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_5),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_5),
.A2(n_51),
.B1(n_54),
.B2(n_160),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_160),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_5),
.A2(n_25),
.B1(n_28),
.B2(n_160),
.Y(n_285)
);

INVx8_ASAP7_75t_SL g47 ( 
.A(n_6),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_7),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_7),
.A2(n_41),
.B1(n_51),
.B2(n_54),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_41),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_7),
.A2(n_25),
.B1(n_28),
.B2(n_41),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_8),
.A2(n_35),
.B1(n_51),
.B2(n_54),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_8),
.A2(n_25),
.B1(n_28),
.B2(n_35),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_9),
.Y(n_66)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_11),
.A2(n_51),
.B1(n_54),
.B2(n_62),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_11),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_11),
.A2(n_39),
.B1(n_62),
.B2(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_62),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_11),
.A2(n_25),
.B1(n_28),
.B2(n_62),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_12),
.B(n_56),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_12),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_12),
.B(n_50),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_12),
.B(n_32),
.C(n_66),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_12),
.A2(n_51),
.B1(n_54),
.B2(n_211),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_12),
.B(n_69),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_211),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_12),
.B(n_25),
.C(n_27),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_12),
.A2(n_101),
.B(n_273),
.Y(n_298)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_14),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_14),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_14),
.A2(n_51),
.B1(n_54),
.B2(n_58),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_58),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_14),
.A2(n_25),
.B1(n_28),
.B2(n_58),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_15),
.A2(n_48),
.B1(n_56),
.B2(n_116),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_15),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_15),
.A2(n_51),
.B1(n_54),
.B2(n_116),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_116),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_15),
.A2(n_25),
.B1(n_28),
.B2(n_116),
.Y(n_243)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_16),
.Y(n_102)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_16),
.Y(n_105)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_16),
.Y(n_221)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_16),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_119),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_117),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_86),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_20),
.B(n_86),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_73),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_36),
.C(n_59),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_22),
.A2(n_81),
.B1(n_82),
.B2(n_84),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_22),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_22),
.A2(n_59),
.B1(n_84),
.B2(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_29),
.B(n_33),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_23),
.A2(n_29),
.B1(n_98),
.B2(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_23),
.A2(n_29),
.B1(n_110),
.B2(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_23),
.A2(n_29),
.B1(n_245),
.B2(n_247),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_23),
.B(n_207),
.Y(n_261)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_24),
.A2(n_34),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_24),
.A2(n_96),
.B1(n_138),
.B2(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_24),
.A2(n_170),
.B(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_24),
.A2(n_206),
.B(n_246),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_24),
.B(n_211),
.Y(n_292)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_24)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_25),
.B(n_102),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_28),
.B(n_297),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_29),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_29),
.B(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_31),
.A2(n_32),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_32),
.B(n_280),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_36),
.A2(n_74),
.B1(n_75),
.B2(n_85),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_36),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_36),
.A2(n_85),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_42),
.B1(n_49),
.B2(n_55),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_37),
.A2(n_49),
.B(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_44)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_42),
.A2(n_49),
.B1(n_55),
.B2(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_42),
.A2(n_142),
.B(n_145),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_43),
.B(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_43),
.A2(n_50),
.B1(n_143),
.B2(n_159),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_43),
.A2(n_146),
.B(n_209),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_49),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_46),
.B1(n_51),
.B2(n_54),
.Y(n_50)
);

NAND2xp33_ASAP7_75t_SL g187 ( 
.A(n_45),
.B(n_51),
.Y(n_187)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI32xp33_ASAP7_75t_L g185 ( 
.A1(n_46),
.A2(n_48),
.A3(n_54),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_49),
.B(n_115),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_49),
.A2(n_113),
.B(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_54),
.B1(n_66),
.B2(n_67),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_51),
.B(n_236),
.Y(n_235)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_63),
.B1(n_69),
.B2(n_70),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_61),
.A2(n_64),
.B1(n_65),
.B2(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_63),
.B(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_63),
.A2(n_69),
.B1(n_178),
.B2(n_203),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_64),
.A2(n_65),
.B1(n_71),
.B2(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_64),
.A2(n_65),
.B1(n_94),
.B2(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_64),
.A2(n_177),
.B(n_179),
.Y(n_176)
);

OAI21xp33_ASAP7_75t_L g249 ( 
.A1(n_64),
.A2(n_179),
.B(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_68),
.Y(n_64)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_65),
.A2(n_140),
.B(n_163),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_65),
.A2(n_163),
.B(n_216),
.Y(n_215)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_69),
.B(n_164),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_80),
.Y(n_75)
);

INVx8_ASAP7_75t_L g210 ( 
.A(n_78),
.Y(n_210)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_91),
.C(n_99),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_87),
.A2(n_91),
.B1(n_92),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_87),
.Y(n_149)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_92),
.A2(n_93),
.B(n_95),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_96),
.A2(n_260),
.B(n_261),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_96),
.A2(n_261),
.B(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_99),
.B(n_148),
.Y(n_147)
);

AOI21xp33_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_107),
.B(n_111),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_111),
.B1(n_112),
.B2(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_100),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_100),
.A2(n_108),
.B1(n_109),
.B2(n_124),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_103),
.B(n_106),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_101),
.A2(n_106),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_101),
.A2(n_103),
.B1(n_132),
.B2(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_101),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_101),
.A2(n_184),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_101),
.B(n_243),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_101),
.A2(n_272),
.B(n_273),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_103),
.B(n_211),
.Y(n_297)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_150),
.B(n_329),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_147),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_121),
.B(n_147),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_125),
.C(n_127),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_122),
.A2(n_125),
.B1(n_126),
.B2(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_122),
.Y(n_325)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_127),
.A2(n_128),
.B1(n_324),
.B2(n_326),
.Y(n_323)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_139),
.C(n_141),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_129),
.A2(n_130),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_131),
.A2(n_135),
.B1(n_136),
.B2(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_131),
.Y(n_172)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_134),
.A2(n_168),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_134),
.B(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_139),
.B(n_141),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_322),
.B(n_328),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_195),
.B(n_321),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_188),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_153),
.B(n_188),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_171),
.C(n_173),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_154),
.A2(n_155),
.B1(n_171),
.B2(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_165),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_161),
.B2(n_162),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_158),
.B(n_161),
.C(n_165),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_159),
.Y(n_175)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_166),
.B(n_169),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_171),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_173),
.B(n_318),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.C(n_180),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_174),
.B(n_176),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_180),
.B(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_185),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_185),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_182),
.A2(n_284),
.B1(n_286),
.B2(n_287),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVxp33_ASAP7_75t_L g212 ( 
.A(n_186),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_194),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_190),
.B(n_191),
.C(n_194),
.Y(n_327)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

O2A1O1Ixp33_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_228),
.B(n_315),
.C(n_320),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_222),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_222),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_213),
.C(n_214),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_198),
.A2(n_199),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_208),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_204),
.B2(n_205),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_204),
.C(n_208),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_203),
.Y(n_216)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI21xp33_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B(n_212),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_213),
.B(n_214),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_217),
.C(n_219),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_215),
.B(n_254),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_217),
.A2(n_218),
.B1(n_219),
.B2(n_255),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_219),
.Y(n_255)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_221),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_223),
.B(n_226),
.C(n_227),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_309),
.B(n_314),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_262),
.B(n_308),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_251),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_233),
.B(n_251),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_244),
.C(n_248),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_234),
.B(n_304),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_237),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B(n_242),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_241),
.A2(n_285),
.B(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_242),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_243),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_244),
.A2(n_248),
.B1(n_249),
.B2(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_244),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_247),
.Y(n_260)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_256),
.B2(n_257),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_252),
.B(n_258),
.C(n_259),
.Y(n_313)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_302),
.B(n_307),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_281),
.B(n_301),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_275),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_265),
.B(n_275),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_271),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_267),
.B(n_270),
.C(n_271),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_272),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_279),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_276),
.A2(n_277),
.B1(n_279),
.B2(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_279),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_290),
.B(n_300),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_288),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_288),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_291),
.A2(n_295),
.B(n_299),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_293),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_298),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_306),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_303),
.B(n_306),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_313),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_313),
.Y(n_314)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_317),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_327),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_327),
.Y(n_328)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_324),
.Y(n_326)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);


endmodule