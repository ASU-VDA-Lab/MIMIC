module fake_jpeg_29129_n_178 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_178);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx12_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_9),
.Y(n_62)
);

INVx8_ASAP7_75t_SL g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_44),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_17),
.B(n_6),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_1),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_76),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_22),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_62),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_52),
.B(n_54),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_80),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

BUFx4f_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_89),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_77),
.A2(n_56),
.B1(n_69),
.B2(n_59),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_88),
.B1(n_57),
.B2(n_76),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_72),
.A2(n_56),
.B1(n_59),
.B2(n_60),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_85),
.A2(n_87),
.B1(n_65),
.B2(n_50),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_79),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_67),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_58),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_94),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_74),
.B(n_70),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_93),
.B(n_96),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_66),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_66),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_55),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_99),
.B(n_106),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_111),
.B1(n_114),
.B2(n_48),
.Y(n_123)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_87),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_102),
.B(n_2),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_87),
.A2(n_80),
.B1(n_75),
.B2(n_55),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_103),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_126)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_51),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g107 ( 
.A(n_91),
.B(n_26),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_5),
.C(n_7),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_68),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_109),
.B(n_115),
.Y(n_129)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

INVxp67_ASAP7_75t_SL g121 ( 
.A(n_112),
.Y(n_121)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_113),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_86),
.A2(n_48),
.B1(n_3),
.B2(n_4),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_48),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_2),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_119),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_3),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_124),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_123),
.A2(n_126),
.B1(n_136),
.B2(n_43),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_4),
.Y(n_124)
);

BUFx24_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_125),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_25),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_128),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_9),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_132),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_10),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_126),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_103),
.A2(n_113),
.B(n_108),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_135),
.A2(n_137),
.B(n_15),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_100),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_109),
.A2(n_12),
.B(n_13),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_146),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_131),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_142),
.B(n_144),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_120),
.B(n_14),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_154),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_16),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_128),
.B(n_19),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_148),
.B(n_155),
.Y(n_164)
);

A2O1A1Ixp33_ASAP7_75t_SL g149 ( 
.A1(n_133),
.A2(n_47),
.B(n_23),
.C(n_27),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_149),
.A2(n_151),
.B(n_152),
.Y(n_160)
);

A2O1A1O1Ixp25_ASAP7_75t_L g151 ( 
.A1(n_127),
.A2(n_20),
.B(n_30),
.C(n_32),
.D(n_33),
.Y(n_151)
);

AOI32xp33_ASAP7_75t_L g152 ( 
.A1(n_118),
.A2(n_34),
.A3(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_153),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_138),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_46),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_125),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_125),
.C(n_121),
.Y(n_157)
);

FAx1_ASAP7_75t_SL g168 ( 
.A(n_157),
.B(n_163),
.CI(n_150),
.CON(n_168),
.SN(n_168)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_121),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_165),
.B(n_141),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_166),
.B(n_167),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_159),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_168),
.A2(n_169),
.B(n_160),
.Y(n_171)
);

A2O1A1O1Ixp25_ASAP7_75t_L g169 ( 
.A1(n_158),
.A2(n_140),
.B(n_139),
.C(n_143),
.D(n_151),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_171),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_166),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_170),
.C(n_161),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_164),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_162),
.C(n_157),
.Y(n_176)
);

OAI21x1_ASAP7_75t_L g177 ( 
.A1(n_176),
.A2(n_162),
.B(n_149),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_149),
.Y(n_178)
);


endmodule