module fake_jpeg_8449_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx8_ASAP7_75t_SL g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

BUFx2_ASAP7_75t_SL g64 ( 
.A(n_36),
.Y(n_64)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_0),
.Y(n_63)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_17),
.B(n_14),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_39),
.B(n_47),
.Y(n_50)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_46),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_21),
.Y(n_47)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_59),
.Y(n_71)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_16),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_58),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_32),
.B1(n_30),
.B2(n_29),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_57),
.A2(n_32),
.B1(n_29),
.B2(n_30),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_16),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_23),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_40),
.A2(n_18),
.B1(n_27),
.B2(n_24),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_68),
.B1(n_17),
.B2(n_25),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_16),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_63),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_40),
.A2(n_30),
.B1(n_29),
.B2(n_25),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVxp67_ASAP7_75t_SL g118 ( 
.A(n_69),
.Y(n_118)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_72),
.Y(n_100)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_73),
.A2(n_35),
.B1(n_27),
.B2(n_54),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_58),
.B(n_41),
.Y(n_74)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_42),
.B(n_17),
.C(n_25),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_79),
.Y(n_111)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_80),
.A2(n_22),
.B(n_66),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_51),
.A2(n_42),
.B1(n_32),
.B2(n_47),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_81),
.A2(n_99),
.B1(n_49),
.B2(n_55),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_19),
.Y(n_84)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_87),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_19),
.Y(n_86)
);

OAI32xp33_ASAP7_75t_L g125 ( 
.A1(n_86),
.A2(n_94),
.A3(n_98),
.B1(n_44),
.B2(n_46),
.Y(n_125)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_50),
.B(n_46),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_88),
.A2(n_22),
.B(n_44),
.Y(n_127)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_91),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_18),
.B1(n_20),
.B2(n_24),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_92),
.A2(n_93),
.B1(n_35),
.B2(n_20),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_67),
.A2(n_18),
.B1(n_20),
.B2(n_24),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_33),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_95),
.Y(n_103)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_96),
.Y(n_112)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_26),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_48),
.Y(n_99)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_87),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_79),
.A2(n_54),
.B1(n_66),
.B2(n_48),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_104),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_105),
.A2(n_114),
.B(n_127),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_106),
.B(n_107),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_95),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_95),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_108),
.B(n_109),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_94),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_123),
.B1(n_70),
.B2(n_74),
.Y(n_131)
);

AND2x4_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_46),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_117),
.A2(n_125),
.B1(n_69),
.B2(n_77),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_85),
.A2(n_54),
.B1(n_53),
.B2(n_65),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_119),
.A2(n_91),
.B1(n_98),
.B2(n_72),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_75),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_121),
.B(n_112),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_78),
.A2(n_53),
.B1(n_65),
.B2(n_35),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_86),
.A2(n_53),
.B1(n_27),
.B2(n_33),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_126),
.A2(n_82),
.B1(n_33),
.B2(n_19),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_83),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_136),
.C(n_142),
.Y(n_160)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_137),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_131),
.A2(n_132),
.B1(n_110),
.B2(n_121),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_111),
.A2(n_83),
.B1(n_77),
.B2(n_89),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_133),
.A2(n_135),
.B1(n_146),
.B2(n_154),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_101),
.C(n_114),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_105),
.A2(n_88),
.B1(n_97),
.B2(n_71),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_139),
.A2(n_14),
.B1(n_12),
.B2(n_11),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_71),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_140),
.B(n_147),
.Y(n_171)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_141),
.A2(n_158),
.B1(n_128),
.B2(n_102),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_73),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_115),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_143),
.A2(n_34),
.B(n_1),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_101),
.B(n_99),
.C(n_90),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_113),
.C(n_100),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_111),
.A2(n_96),
.B1(n_82),
.B2(n_28),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_145),
.A2(n_107),
.B1(n_108),
.B2(n_103),
.Y(n_175)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_150),
.Y(n_180)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_116),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_153),
.Y(n_190)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_100),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_114),
.A2(n_43),
.B1(n_45),
.B2(n_33),
.Y(n_154)
);

AOI32xp33_ASAP7_75t_L g155 ( 
.A1(n_125),
.A2(n_45),
.A3(n_43),
.B1(n_76),
.B2(n_28),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_155),
.A2(n_104),
.B(n_117),
.Y(n_174)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_118),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_109),
.A2(n_26),
.B1(n_19),
.B2(n_45),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_159),
.A2(n_34),
.B1(n_1),
.B2(n_2),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_152),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_161),
.B(n_162),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_159),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_166),
.C(n_167),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_113),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_127),
.C(n_119),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_156),
.A2(n_120),
.B(n_126),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_168),
.A2(n_3),
.B(n_4),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_123),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_177),
.C(n_185),
.Y(n_204)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_141),
.Y(n_170)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_170),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_132),
.Y(n_172)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_106),
.Y(n_173)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_173),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_174),
.A2(n_178),
.B(n_181),
.Y(n_210)
);

OAI21xp33_ASAP7_75t_SL g217 ( 
.A1(n_175),
.A2(n_186),
.B(n_189),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_182),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_43),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_148),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_156),
.A2(n_103),
.B(n_22),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_112),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_112),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_183),
.B(n_188),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_134),
.B(n_116),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_155),
.A2(n_128),
.B1(n_26),
.B2(n_22),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_187),
.A2(n_130),
.B1(n_150),
.B2(n_151),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_26),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_137),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_191),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_149),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_154),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_139),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_205),
.C(n_207),
.Y(n_233)
);

AND2x6_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_160),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_199),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_200),
.B(n_209),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_188),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_202),
.B(n_206),
.Y(n_244)
);

NAND2x1_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_147),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_203),
.A2(n_221),
.B(n_3),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_166),
.B(n_144),
.C(n_131),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_146),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_169),
.B(n_158),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_187),
.C(n_194),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_191),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_211),
.A2(n_193),
.B1(n_192),
.B2(n_179),
.Y(n_231)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_165),
.Y(n_212)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_212),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_184),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_213),
.A2(n_173),
.B1(n_179),
.B2(n_183),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_174),
.A2(n_14),
.B1(n_12),
.B2(n_11),
.Y(n_214)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_214),
.Y(n_227)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_180),
.Y(n_215)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_215),
.Y(n_229)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_171),
.Y(n_220)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_220),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_167),
.B(n_2),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_178),
.B(n_3),
.Y(n_223)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_224),
.A2(n_189),
.B(n_181),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_228),
.A2(n_222),
.B1(n_202),
.B2(n_196),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_230),
.B(n_237),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_231),
.A2(n_234),
.B1(n_238),
.B2(n_240),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_164),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_235),
.C(n_239),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_201),
.A2(n_184),
.B1(n_163),
.B2(n_168),
.Y(n_234)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_203),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_217),
.A2(n_163),
.B1(n_170),
.B2(n_175),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_191),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_222),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_241),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_247),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_218),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_243),
.B(n_197),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_198),
.B(n_11),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_248),
.C(n_195),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_208),
.B(n_4),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_195),
.B(n_205),
.C(n_199),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_211),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_196),
.Y(n_267)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_251),
.Y(n_278)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_244),
.Y(n_255)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_255),
.Y(n_288)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_246),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_257),
.Y(n_277)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_269),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_250),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_262),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_207),
.C(n_219),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_245),
.C(n_247),
.Y(n_281)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_228),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_263),
.A2(n_264),
.B1(n_271),
.B2(n_235),
.Y(n_275)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_234),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_266),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_267),
.A2(n_219),
.B(n_223),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_225),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_268),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_210),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_233),
.B(n_210),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_232),
.Y(n_279)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_231),
.Y(n_271)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_273),
.Y(n_294)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_275),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_248),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_276),
.A2(n_5),
.B(n_6),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_283),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_262),
.A2(n_226),
.B1(n_227),
.B2(n_200),
.Y(n_280)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_280),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_286),
.C(n_6),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_258),
.A2(n_249),
.B(n_229),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_282),
.A2(n_221),
.B(n_6),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_230),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_252),
.B(n_224),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_251),
.A2(n_257),
.B1(n_236),
.B2(n_213),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_287),
.A2(n_221),
.B1(n_252),
.B2(n_7),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_284),
.B(n_265),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_298),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_278),
.A2(n_260),
.B1(n_265),
.B2(n_259),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_291),
.A2(n_302),
.B1(n_283),
.B2(n_282),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_272),
.B(n_261),
.Y(n_292)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_292),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_288),
.A2(n_270),
.B1(n_254),
.B2(n_253),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_293),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_253),
.Y(n_295)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_295),
.Y(n_307)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_296),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_276),
.Y(n_300)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_300),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_301),
.A2(n_273),
.B(n_277),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_285),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_281),
.C(n_288),
.Y(n_304)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_304),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_279),
.C(n_274),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_290),
.C(n_303),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_277),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_295),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_311),
.A2(n_298),
.B(n_299),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_294),
.A2(n_276),
.B(n_280),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_314),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_294),
.Y(n_316)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_316),
.Y(n_325)
);

INVx11_ASAP7_75t_L g317 ( 
.A(n_312),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_319),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_318),
.A2(n_323),
.B(n_324),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_322),
.A2(n_301),
.B1(n_310),
.B2(n_293),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_297),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_306),
.B(n_313),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_326),
.A2(n_329),
.B(n_320),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_317),
.A2(n_304),
.B1(n_310),
.B2(n_307),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_327),
.Y(n_332)
);

A2O1A1Ixp33_ASAP7_75t_L g329 ( 
.A1(n_322),
.A2(n_291),
.B(n_286),
.C(n_274),
.Y(n_329)
);

MAJx2_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_333),
.C(n_321),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_330),
.A2(n_321),
.B(n_318),
.Y(n_333)
);

O2A1O1Ixp33_ASAP7_75t_SL g335 ( 
.A1(n_334),
.A2(n_332),
.B(n_328),
.C(n_325),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_305),
.C(n_329),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_336),
.B(n_9),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_10),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_10),
.B(n_337),
.Y(n_339)
);


endmodule