module fake_jpeg_1382_n_67 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_67);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_67;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;
wire n_66;

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_10),
.B(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_19),
.B(n_22),
.Y(n_25)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_1),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_23),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_16),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_21),
.A2(n_17),
.B(n_13),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_27),
.A2(n_20),
.B1(n_11),
.B2(n_9),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_12),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_35),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_29),
.A2(n_18),
.B1(n_14),
.B2(n_3),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_26),
.Y(n_38)
);

NAND3xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_25),
.C(n_7),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_25),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_27),
.C(n_26),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_46),
.C(n_40),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_31),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_50),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_49),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_33),
.B1(n_32),
.B2(n_18),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_54),
.C(n_53),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_28),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_42),
.Y(n_55)
);

NAND3xp33_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_56),
.C(n_14),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_39),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_58),
.Y(n_63)
);

AOI221xp5_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_60),
.C(n_2),
.Y(n_61)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_28),
.C(n_3),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

A2O1A1O1Ixp25_ASAP7_75t_L g66 ( 
.A1(n_64),
.A2(n_63),
.B(n_5),
.C(n_6),
.D(n_2),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_65),
.Y(n_67)
);


endmodule