module fake_jpeg_12344_n_530 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_530);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_530;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx6_ASAP7_75t_SL g19 ( 
.A(n_17),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_10),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_7),
.B(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_56),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_58),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_59),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_30),
.Y(n_60)
);

INVx5_ASAP7_75t_SL g127 ( 
.A(n_60),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_61),
.Y(n_142)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_62),
.Y(n_137)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_64),
.Y(n_150)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_67),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_19),
.B(n_0),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_69),
.B(n_92),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_35),
.B(n_0),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_102),
.Y(n_108)
);

INVx6_ASAP7_75t_SL g71 ( 
.A(n_30),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_71),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_72),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_73),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_74),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_30),
.Y(n_79)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_83),
.Y(n_140)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_86),
.Y(n_138)
);

INVx4_ASAP7_75t_SL g87 ( 
.A(n_30),
.Y(n_87)
);

INVx5_ASAP7_75t_SL g156 ( 
.A(n_87),
.Y(n_156)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_88),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_89),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_91),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_35),
.B(n_1),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_95),
.Y(n_121)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

BUFx12_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_47),
.B(n_20),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_99),
.Y(n_131)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_21),
.Y(n_98)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_98),
.Y(n_158)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_100),
.B(n_101),
.Y(n_148)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_21),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_34),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_76),
.A2(n_34),
.B1(n_46),
.B2(n_47),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_105),
.A2(n_132),
.B1(n_161),
.B2(n_58),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_79),
.A2(n_34),
.B1(n_46),
.B2(n_44),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_107),
.A2(n_118),
.B(n_120),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_115),
.B(n_87),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_82),
.A2(n_44),
.B1(n_46),
.B2(n_48),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_80),
.A2(n_34),
.B1(n_44),
.B2(n_39),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_23),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_130),
.B(n_144),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_L g132 ( 
.A1(n_83),
.A2(n_39),
.B1(n_31),
.B2(n_29),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_89),
.A2(n_39),
.B1(n_21),
.B2(n_52),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_143),
.A2(n_21),
.B1(n_73),
.B2(n_72),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_69),
.B(n_23),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_60),
.B(n_52),
.C(n_27),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_149),
.A2(n_32),
.B(n_22),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_92),
.B(n_48),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_153),
.B(n_159),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_63),
.B(n_43),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_85),
.A2(n_103),
.B1(n_102),
.B2(n_75),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_162),
.B(n_164),
.Y(n_220)
);

O2A1O1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_127),
.A2(n_33),
.B(n_31),
.C(n_29),
.Y(n_163)
);

A2O1A1Ixp33_ASAP7_75t_L g251 ( 
.A1(n_163),
.A2(n_185),
.B(n_22),
.C(n_116),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_156),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_108),
.B(n_33),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_165),
.B(n_174),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_156),
.Y(n_166)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_166),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_127),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_168),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_148),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_169),
.B(n_173),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_126),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_170),
.Y(n_232)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_171),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_147),
.Y(n_172)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_172),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_121),
.B(n_24),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_131),
.B(n_24),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_176),
.Y(n_230)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_177),
.Y(n_248)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_122),
.Y(n_178)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_178),
.Y(n_218)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_179),
.Y(n_223)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_138),
.Y(n_180)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_180),
.Y(n_245)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_123),
.Y(n_181)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_131),
.B(n_21),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_182),
.B(n_154),
.C(n_141),
.Y(n_224)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_113),
.Y(n_183)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_183),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_148),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_184),
.B(n_192),
.Y(n_225)
);

A2O1A1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_106),
.A2(n_95),
.B(n_43),
.C(n_36),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_25),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_186),
.B(n_191),
.Y(n_239)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_152),
.Y(n_187)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_187),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_145),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_188),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_109),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_189),
.Y(n_250)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_128),
.Y(n_190)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_190),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_110),
.B(n_25),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_111),
.B(n_36),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_193),
.Y(n_256)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_124),
.Y(n_194)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_194),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_111),
.B(n_32),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_195),
.B(n_199),
.Y(n_244)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_134),
.Y(n_196)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_196),
.Y(n_260)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_158),
.Y(n_197)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_197),
.Y(n_243)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_104),
.Y(n_198)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_198),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_123),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_200),
.B(n_161),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_146),
.Y(n_201)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_201),
.Y(n_249)
);

BUFx4f_ASAP7_75t_L g202 ( 
.A(n_160),
.Y(n_202)
);

INVx11_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_126),
.Y(n_203)
);

NAND2xp33_ASAP7_75t_SL g258 ( 
.A(n_203),
.B(n_211),
.Y(n_258)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_112),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_205),
.B(n_212),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_125),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_206),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_207),
.A2(n_55),
.B1(n_74),
.B2(n_66),
.Y(n_247)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_104),
.Y(n_208)
);

INVx11_ASAP7_75t_L g259 ( 
.A(n_208),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_105),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_209),
.B(n_150),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_114),
.Y(n_210)
);

BUFx12f_ASAP7_75t_L g233 ( 
.A(n_210),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_155),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_132),
.B(n_1),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_117),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_213),
.Y(n_227)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_140),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_214),
.Y(n_231)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_160),
.Y(n_215)
);

NAND2xp33_ASAP7_75t_SL g261 ( 
.A(n_215),
.B(n_133),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_185),
.A2(n_143),
.B1(n_120),
.B2(n_107),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_217),
.A2(n_253),
.B1(n_256),
.B2(n_182),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_224),
.B(n_166),
.C(n_182),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_234),
.B(n_163),
.Y(n_274)
);

AOI32xp33_ASAP7_75t_L g238 ( 
.A1(n_165),
.A2(n_111),
.A3(n_116),
.B1(n_112),
.B2(n_135),
.Y(n_238)
);

A2O1A1Ixp33_ASAP7_75t_L g277 ( 
.A1(n_238),
.A2(n_255),
.B(n_205),
.C(n_198),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_247),
.A2(n_136),
.B1(n_117),
.B2(n_119),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_200),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_167),
.A2(n_54),
.B1(n_57),
.B2(n_59),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_212),
.A2(n_157),
.B1(n_129),
.B2(n_135),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_254),
.A2(n_168),
.B1(n_167),
.B2(n_191),
.Y(n_266)
);

FAx1_ASAP7_75t_SL g255 ( 
.A(n_174),
.B(n_1),
.CI(n_2),
.CON(n_255),
.SN(n_255)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_186),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_175),
.Y(n_281)
);

NAND2xp33_ASAP7_75t_SL g273 ( 
.A(n_261),
.B(n_203),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_263),
.Y(n_290)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_226),
.Y(n_264)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_264),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_265),
.B(n_270),
.C(n_286),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_266),
.A2(n_283),
.B1(n_298),
.B2(n_228),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_267),
.A2(n_273),
.B(n_274),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_268),
.A2(n_292),
.B1(n_297),
.B2(n_301),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_256),
.A2(n_162),
.B(n_170),
.Y(n_269)
);

A2O1A1Ixp33_ASAP7_75t_SL g328 ( 
.A1(n_269),
.A2(n_275),
.B(n_304),
.C(n_216),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_224),
.B(n_162),
.C(n_194),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_226),
.Y(n_271)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_271),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_239),
.B(n_204),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_272),
.B(n_277),
.Y(n_318)
);

OA21x2_ASAP7_75t_L g275 ( 
.A1(n_253),
.A2(n_172),
.B(n_206),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_259),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_276),
.B(n_281),
.Y(n_317)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_236),
.Y(n_278)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_278),
.Y(n_322)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_236),
.Y(n_279)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_279),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_234),
.B(n_220),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_280),
.Y(n_319)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_249),
.Y(n_282)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_282),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_240),
.A2(n_129),
.B1(n_157),
.B2(n_150),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_249),
.Y(n_284)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_284),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_240),
.B(n_183),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_285),
.B(n_289),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_237),
.B(n_180),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_258),
.A2(n_208),
.B(n_181),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_287),
.A2(n_291),
.B(n_232),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_239),
.B(n_196),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_288),
.B(n_295),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_254),
.B(n_214),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_258),
.B(n_231),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_237),
.A2(n_177),
.B1(n_142),
.B2(n_136),
.Y(n_292)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_293),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_229),
.B(n_178),
.C(n_213),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_294),
.B(n_300),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_244),
.B(n_215),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_218),
.Y(n_296)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_296),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_251),
.A2(n_142),
.B1(n_119),
.B2(n_133),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_222),
.A2(n_64),
.B1(n_61),
.B2(n_210),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_255),
.B(n_179),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_299),
.B(n_245),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_225),
.B(n_190),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_255),
.A2(n_202),
.B1(n_4),
.B2(n_5),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_259),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_302),
.B(n_305),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_261),
.A2(n_202),
.B(n_6),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_303),
.A2(n_273),
.B(n_269),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_242),
.A2(n_16),
.B(n_6),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_228),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_241),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_306),
.A2(n_260),
.B1(n_246),
.B2(n_221),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_308),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_295),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_309),
.B(n_310),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_288),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_312),
.B(n_338),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_266),
.A2(n_227),
.B1(n_248),
.B2(n_230),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_313),
.A2(n_315),
.B1(n_324),
.B2(n_332),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_314),
.A2(n_328),
.B(n_334),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_275),
.A2(n_274),
.B1(n_267),
.B2(n_280),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_299),
.A2(n_250),
.B(n_216),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_320),
.A2(n_329),
.B(n_333),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_291),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_321),
.B(n_337),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_275),
.A2(n_248),
.B1(n_243),
.B2(n_219),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_287),
.A2(n_219),
.B(n_235),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_331),
.A2(n_289),
.B1(n_283),
.B2(n_271),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_275),
.A2(n_242),
.B1(n_245),
.B2(n_260),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_291),
.A2(n_223),
.B(n_252),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_280),
.A2(n_223),
.B(n_252),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_276),
.Y(n_337)
);

OAI32xp33_ASAP7_75t_L g338 ( 
.A1(n_277),
.A2(n_272),
.A3(n_274),
.B1(n_268),
.B2(n_285),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_341),
.B(n_290),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_303),
.A2(n_262),
.B(n_246),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_342),
.Y(n_352)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_264),
.Y(n_343)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_343),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_345),
.B(n_270),
.C(n_265),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_347),
.B(n_358),
.C(n_373),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_336),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_348),
.B(n_351),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_335),
.A2(n_302),
.B1(n_305),
.B2(n_278),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_349),
.A2(n_329),
.B(n_308),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_350),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_336),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_345),
.B(n_318),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_354),
.B(n_330),
.Y(n_400)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_317),
.Y(n_355)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_355),
.Y(n_390)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_307),
.Y(n_356)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_356),
.Y(n_397)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_307),
.Y(n_357)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_357),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_319),
.B(n_286),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_316),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_359),
.B(n_360),
.Y(n_387)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_316),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_311),
.A2(n_290),
.B1(n_285),
.B2(n_289),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_362),
.A2(n_368),
.B1(n_323),
.B2(n_322),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_310),
.B(n_279),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_363),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_365),
.B(n_375),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_311),
.A2(n_298),
.B1(n_297),
.B2(n_284),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_327),
.B(n_282),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_369),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_317),
.B(n_294),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_372),
.B(n_376),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_319),
.B(n_296),
.C(n_292),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_319),
.B(n_301),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_374),
.B(n_380),
.C(n_328),
.Y(n_395)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_322),
.Y(n_375)
);

OAI32xp33_ASAP7_75t_L g376 ( 
.A1(n_341),
.A2(n_218),
.A3(n_221),
.B1(n_304),
.B2(n_306),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_327),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_377),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_337),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_378),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_330),
.B(n_235),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_379),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_344),
.B(n_262),
.C(n_233),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_381),
.A2(n_383),
.B(n_394),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_367),
.A2(n_314),
.B(n_344),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_362),
.A2(n_315),
.B1(n_312),
.B2(n_313),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_385),
.A2(n_388),
.B1(n_392),
.B2(n_396),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_364),
.A2(n_324),
.B1(n_332),
.B2(n_321),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_377),
.A2(n_309),
.B1(n_318),
.B2(n_328),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_367),
.A2(n_333),
.B(n_320),
.Y(n_394)
);

XNOR2x1_ASAP7_75t_L g415 ( 
.A(n_395),
.B(n_380),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_363),
.A2(n_328),
.B1(n_342),
.B2(n_338),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_370),
.A2(n_328),
.B1(n_335),
.B2(n_334),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_399),
.A2(n_405),
.B1(n_407),
.B2(n_350),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g439 ( 
.A(n_400),
.B(n_353),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_354),
.B(n_340),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_401),
.B(n_409),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_361),
.A2(n_340),
.B(n_343),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_402),
.B(n_371),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_404),
.B(n_410),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_368),
.A2(n_346),
.B1(n_352),
.B2(n_369),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_346),
.A2(n_323),
.B1(n_326),
.B2(n_325),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_347),
.B(n_326),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_361),
.A2(n_325),
.B(n_339),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_358),
.B(n_339),
.C(n_331),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_412),
.B(n_348),
.C(n_351),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_413),
.B(n_427),
.C(n_429),
.Y(n_452)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_406),
.Y(n_414)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_414),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_415),
.B(n_430),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_403),
.B(n_378),
.Y(n_416)
);

NAND3xp33_ASAP7_75t_L g441 ( 
.A(n_416),
.B(n_422),
.C(n_428),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_406),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_417),
.B(n_419),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_409),
.B(n_389),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_418),
.B(n_426),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_387),
.Y(n_419)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_387),
.Y(n_421)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_421),
.Y(n_440)
);

NOR3xp33_ASAP7_75t_SL g422 ( 
.A(n_390),
.B(n_353),
.C(n_375),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_424),
.A2(n_383),
.B(n_394),
.Y(n_457)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_393),
.Y(n_425)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_425),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_389),
.B(n_374),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_400),
.B(n_366),
.C(n_373),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_403),
.B(n_359),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_401),
.B(n_412),
.C(n_395),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_398),
.B(n_366),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_402),
.B(n_392),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_431),
.B(n_439),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_410),
.B(n_352),
.C(n_370),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_432),
.B(n_435),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_408),
.B(n_360),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_434),
.B(n_411),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_408),
.B(n_357),
.C(n_356),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_436),
.A2(n_385),
.B1(n_405),
.B2(n_404),
.Y(n_443)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_393),
.Y(n_438)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_438),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_422),
.B(n_391),
.Y(n_442)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_442),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_443),
.A2(n_446),
.B1(n_448),
.B2(n_459),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_437),
.A2(n_382),
.B1(n_399),
.B2(n_391),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_445),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_420),
.A2(n_396),
.B1(n_407),
.B2(n_382),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_420),
.A2(n_388),
.B1(n_384),
.B2(n_386),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_437),
.A2(n_386),
.B1(n_384),
.B2(n_390),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_449),
.B(n_450),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_435),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_457),
.B(n_427),
.C(n_413),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_432),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_459),
.B(n_429),
.Y(n_466)
);

CKINVDCx16_ASAP7_75t_R g477 ( 
.A(n_460),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_420),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_461),
.B(n_411),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_452),
.B(n_418),
.C(n_426),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_462),
.B(n_467),
.Y(n_491)
);

XNOR2x1_ASAP7_75t_L g463 ( 
.A(n_447),
.B(n_415),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_SL g492 ( 
.A(n_463),
.B(n_466),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_464),
.B(n_468),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_452),
.B(n_423),
.C(n_431),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_444),
.B(n_423),
.C(n_439),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_469),
.A2(n_445),
.B1(n_456),
.B2(n_440),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_444),
.B(n_433),
.C(n_430),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_470),
.B(n_472),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_447),
.B(n_433),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_471),
.B(n_474),
.C(n_476),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_451),
.B(n_381),
.C(n_397),
.Y(n_472)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_473),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_457),
.B(n_376),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_455),
.B(n_397),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_477),
.B(n_454),
.Y(n_480)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_480),
.Y(n_497)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_481),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_475),
.B(n_441),
.Y(n_482)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_482),
.Y(n_505)
);

NOR2xp67_ASAP7_75t_L g484 ( 
.A(n_466),
.B(n_458),
.Y(n_484)
);

OAI21x1_ASAP7_75t_SL g495 ( 
.A1(n_484),
.A2(n_474),
.B(n_471),
.Y(n_495)
);

FAx1_ASAP7_75t_SL g485 ( 
.A(n_470),
.B(n_442),
.CI(n_448),
.CON(n_485),
.SN(n_485)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_485),
.B(n_486),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_465),
.B(n_458),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_462),
.B(n_453),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_487),
.A2(n_10),
.B(n_11),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_467),
.B(n_455),
.C(n_443),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_488),
.B(n_494),
.C(n_463),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_478),
.A2(n_440),
.B1(n_453),
.B2(n_446),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_490),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_476),
.B(n_233),
.C(n_7),
.Y(n_494)
);

NAND2xp33_ASAP7_75t_SL g513 ( 
.A(n_495),
.B(n_492),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_488),
.B(n_468),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_496),
.B(n_499),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_491),
.B(n_233),
.C(n_8),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_500),
.B(n_501),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_493),
.B(n_3),
.C(n_8),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_479),
.A2(n_3),
.B1(n_8),
.B2(n_10),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_503),
.B(n_504),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_483),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_506),
.B(n_11),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_497),
.B(n_485),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_508),
.B(n_511),
.Y(n_517)
);

AOI31xp67_ASAP7_75t_SL g509 ( 
.A1(n_505),
.A2(n_485),
.A3(n_490),
.B(n_481),
.Y(n_509)
);

AOI21x1_ASAP7_75t_L g521 ( 
.A1(n_509),
.A2(n_513),
.B(n_499),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_507),
.A2(n_489),
.B1(n_479),
.B2(n_494),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_514),
.B(n_501),
.Y(n_518)
);

AOI21xp33_ASAP7_75t_L g516 ( 
.A1(n_507),
.A2(n_492),
.B(n_14),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_516),
.A2(n_502),
.B(n_500),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_518),
.B(n_519),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_515),
.B(n_498),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_520),
.B(n_521),
.C(n_496),
.Y(n_524)
);

AO21x1_ASAP7_75t_L g522 ( 
.A1(n_517),
.A2(n_515),
.B(n_512),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_522),
.A2(n_524),
.B(n_13),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_523),
.B(n_510),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_525),
.A2(n_526),
.B1(n_13),
.B2(n_14),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_527),
.A2(n_13),
.B(n_15),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_528),
.A2(n_15),
.B(n_403),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_529),
.Y(n_530)
);


endmodule