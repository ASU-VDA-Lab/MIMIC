module fake_jpeg_4291_n_279 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx4f_ASAP7_75t_SL g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_19),
.B(n_14),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_36),
.Y(n_43)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_27),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_14),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_39),
.B(n_29),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_23),
.B1(n_29),
.B2(n_18),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_48),
.A2(n_23),
.B1(n_31),
.B2(n_20),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_22),
.B1(n_25),
.B2(n_15),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_26),
.B(n_16),
.C(n_38),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_18),
.B1(n_20),
.B2(n_15),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_50),
.A2(n_61),
.B1(n_64),
.B2(n_26),
.Y(n_73)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_53),
.B(n_59),
.Y(n_84)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_35),
.A2(n_25),
.B1(n_22),
.B2(n_31),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_42),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_31),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_63),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_15),
.B1(n_30),
.B2(n_22),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_66),
.A2(n_72),
.B1(n_78),
.B2(n_57),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_20),
.Y(n_70)
);

FAx1_ASAP7_75t_SL g103 ( 
.A(n_70),
.B(n_26),
.CI(n_16),
.CON(n_103),
.SN(n_103)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_71),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_52),
.A2(n_30),
.B1(n_12),
.B2(n_13),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_73),
.A2(n_79),
.B1(n_82),
.B2(n_26),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_54),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_81),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_86),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_46),
.A2(n_10),
.B1(n_8),
.B2(n_11),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_55),
.A2(n_24),
.B1(n_17),
.B2(n_38),
.Y(n_82)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_43),
.B(n_42),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_43),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_46),
.B1(n_58),
.B2(n_49),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_88),
.A2(n_93),
.B1(n_70),
.B2(n_82),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_107),
.Y(n_118)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_96),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_46),
.B1(n_62),
.B2(n_51),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_53),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_94),
.Y(n_112)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_99),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_51),
.C(n_63),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_98),
.A2(n_105),
.B(n_69),
.Y(n_116)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_100),
.A2(n_108),
.B1(n_75),
.B2(n_76),
.Y(n_114)
);

BUFx24_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_101),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_40),
.B1(n_54),
.B2(n_57),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_85),
.B1(n_95),
.B2(n_75),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_103),
.A2(n_47),
.B(n_16),
.Y(n_128)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_104),
.B(n_106),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_40),
.C(n_42),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_47),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_56),
.Y(n_109)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_109),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_67),
.B(n_80),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_110),
.B(n_13),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_107),
.A2(n_67),
.B1(n_74),
.B2(n_70),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_113),
.A2(n_120),
.B1(n_121),
.B2(n_125),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_114),
.A2(n_123),
.B1(n_124),
.B2(n_132),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_116),
.A2(n_133),
.B(n_100),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_90),
.A2(n_70),
.B1(n_85),
.B2(n_69),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_130),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_102),
.A2(n_56),
.B1(n_75),
.B2(n_86),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_102),
.A2(n_17),
.B1(n_24),
.B2(n_60),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_129),
.Y(n_136)
);

OAI32xp33_ASAP7_75t_L g127 ( 
.A1(n_102),
.A2(n_24),
.A3(n_17),
.B1(n_21),
.B2(n_65),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_128),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_104),
.B(n_0),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_88),
.A2(n_65),
.B1(n_60),
.B2(n_17),
.Y(n_132)
);

AOI32xp33_ASAP7_75t_L g133 ( 
.A1(n_103),
.A2(n_47),
.A3(n_44),
.B1(n_60),
.B2(n_65),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_98),
.C(n_91),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_144),
.C(n_148),
.Y(n_160)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_134),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_139),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_94),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_146),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_112),
.A2(n_95),
.B1(n_93),
.B2(n_103),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_126),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_105),
.C(n_109),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_97),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_99),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_158),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_96),
.C(n_92),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_68),
.Y(n_149)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_133),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_10),
.Y(n_178)
);

AO22x1_ASAP7_75t_L g151 ( 
.A1(n_127),
.A2(n_24),
.B1(n_44),
.B2(n_16),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_151),
.A2(n_152),
.B(n_125),
.Y(n_165)
);

NOR2x1_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_16),
.Y(n_153)
);

NAND3xp33_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_9),
.C(n_1),
.Y(n_182)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_119),
.Y(n_154)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_156),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_121),
.A2(n_68),
.B1(n_16),
.B2(n_101),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_157),
.A2(n_123),
.B1(n_132),
.B2(n_131),
.Y(n_162)
);

AND2x6_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_68),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_120),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_159),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_124),
.C(n_117),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_164),
.C(n_167),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_162),
.A2(n_180),
.B1(n_151),
.B2(n_135),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_172),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_112),
.C(n_115),
.Y(n_164)
);

NOR3xp33_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_182),
.C(n_153),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_115),
.C(n_129),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_169),
.Y(n_188)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_21),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_141),
.A2(n_101),
.B1(n_21),
.B2(n_2),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_173),
.A2(n_179),
.B1(n_9),
.B2(n_3),
.Y(n_202)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_177),
.B(n_136),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_145),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_158),
.A2(n_10),
.B1(n_9),
.B2(n_2),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_155),
.A2(n_101),
.B1(n_1),
.B2(n_2),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_176),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_184),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_168),
.B(n_135),
.Y(n_186)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_136),
.Y(n_189)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_189),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_152),
.C(n_155),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_198),
.C(n_200),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_192),
.A2(n_193),
.B1(n_201),
.B2(n_202),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_183),
.A2(n_151),
.B1(n_150),
.B2(n_145),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_203),
.Y(n_214)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_179),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_197),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_143),
.C(n_157),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_164),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_199),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_0),
.C(n_1),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_171),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_166),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_174),
.B(n_2),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_204),
.B(n_181),
.C(n_177),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_166),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_212),
.C(n_219),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_189),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_194),
.B(n_172),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_216),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_163),
.C(n_167),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_178),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_185),
.B(n_165),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_173),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_198),
.C(n_200),
.Y(n_226)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_227),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_209),
.Y(n_245)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_208),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_210),
.A2(n_188),
.B(n_193),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_228),
.A2(n_234),
.B(n_236),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_229),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_196),
.C(n_169),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_235),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_201),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_231),
.Y(n_238)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_222),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_233),
.Y(n_249)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_170),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_195),
.C(n_192),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_202),
.C(n_4),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_221),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_237),
.B(n_213),
.Y(n_240)
);

OAI21x1_ASAP7_75t_L g239 ( 
.A1(n_236),
.A2(n_210),
.B(n_216),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_219),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_240),
.Y(n_251)
);

NAND3xp33_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_218),
.C(n_217),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_241),
.A2(n_244),
.B(n_246),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_230),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_225),
.Y(n_256)
);

INVxp33_ASAP7_75t_L g246 ( 
.A(n_235),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_250),
.A2(n_3),
.B(n_4),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_214),
.Y(n_252)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_252),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_246),
.B(n_206),
.Y(n_253)
);

AOI221xp5_ASAP7_75t_L g262 ( 
.A1(n_253),
.A2(n_259),
.B1(n_248),
.B2(n_249),
.C(n_5),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_225),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_257),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_245),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_242),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_223),
.Y(n_258)
);

INVxp33_ASAP7_75t_L g266 ( 
.A(n_258),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_223),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_262),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_3),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_4),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_251),
.C(n_257),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_267),
.A2(n_268),
.B(n_269),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_255),
.C(n_250),
.Y(n_268)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_3),
.Y(n_269)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_270),
.Y(n_272)
);

O2A1O1Ixp33_ASAP7_75t_SL g273 ( 
.A1(n_270),
.A2(n_260),
.B(n_265),
.C(n_7),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_273),
.B(n_272),
.Y(n_275)
);

AOI322xp5_ASAP7_75t_L g277 ( 
.A1(n_275),
.A2(n_276),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_253),
.C2(n_272),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_271),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g278 ( 
.A(n_277),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_278),
.Y(n_279)
);


endmodule