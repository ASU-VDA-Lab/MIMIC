module fake_jpeg_5987_n_289 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_289);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_289;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

AOI21xp33_ASAP7_75t_L g30 ( 
.A1(n_14),
.A2(n_0),
.B(n_1),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_20),
.C(n_25),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_23),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_31),
.B(n_32),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_23),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_18),
.Y(n_35)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_30),
.B(n_27),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_48),
.Y(n_59)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_28),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_53),
.Y(n_80)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_55),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

NOR2x1_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_46),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_57),
.Y(n_83)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_31),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_61),
.B(n_65),
.Y(n_69)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_63),
.Y(n_76)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_31),
.Y(n_65)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_81),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_43),
.B1(n_48),
.B2(n_40),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_72),
.A2(n_29),
.B1(n_36),
.B2(n_33),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_43),
.Y(n_77)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_49),
.B1(n_16),
.B2(n_13),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_78),
.A2(n_79),
.B1(n_34),
.B2(n_19),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_49),
.B1(n_16),
.B2(n_32),
.Y(n_79)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_55),
.Y(n_106)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_75),
.A2(n_64),
.B1(n_44),
.B2(n_62),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_91),
.A2(n_93),
.B1(n_104),
.B2(n_70),
.Y(n_127)
);

AND2x6_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_37),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_96),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_75),
.A2(n_39),
.B1(n_51),
.B2(n_19),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_94),
.B(n_95),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_83),
.B(n_35),
.Y(n_95)
);

AND2x6_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_37),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_35),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_102),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_69),
.A2(n_37),
.B(n_33),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_99),
.C(n_105),
.Y(n_111)
);

AND2x6_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_39),
.Y(n_99)
);

NOR3xp33_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_32),
.C(n_34),
.Y(n_100)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

OA22x2_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_27),
.B1(n_16),
.B2(n_56),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_103),
.A2(n_105),
.B1(n_71),
.B2(n_42),
.Y(n_112)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_73),
.Y(n_120)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_109),
.B(n_110),
.Y(n_132)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_111),
.A2(n_116),
.B1(n_118),
.B2(n_127),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_113),
.Y(n_133)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_92),
.A2(n_13),
.B1(n_29),
.B2(n_87),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_119),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_96),
.A2(n_29),
.B1(n_42),
.B2(n_73),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_102),
.B(n_76),
.Y(n_119)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_126),
.Y(n_149)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_88),
.B(n_38),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_107),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_111),
.A2(n_110),
.B1(n_113),
.B2(n_115),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_129),
.A2(n_142),
.B1(n_18),
.B2(n_25),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_120),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_130),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_128),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_134),
.B(n_143),
.Y(n_158)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_118),
.A2(n_88),
.B1(n_97),
.B2(n_95),
.Y(n_138)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_141),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_98),
.Y(n_140)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_123),
.A2(n_97),
.B1(n_94),
.B2(n_86),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_108),
.B(n_114),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_144),
.B(n_151),
.Y(n_159)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_147),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_126),
.B1(n_125),
.B2(n_109),
.Y(n_146)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_150),
.Y(n_170)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_120),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_76),
.Y(n_152)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_152),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_27),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_156),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_27),
.Y(n_156)
);

AO22x1_ASAP7_75t_L g157 ( 
.A1(n_152),
.A2(n_24),
.B1(n_26),
.B2(n_14),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_157),
.A2(n_160),
.B(n_176),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_140),
.A2(n_101),
.B(n_67),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_147),
.B(n_85),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_148),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_151),
.Y(n_162)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_58),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_173),
.C(n_146),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_20),
.Y(n_166)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_168),
.A2(n_136),
.B1(n_15),
.B2(n_89),
.Y(n_191)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_132),
.B(n_58),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_130),
.B(n_14),
.Y(n_174)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_143),
.A2(n_15),
.B(n_14),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_175),
.A2(n_135),
.B(n_137),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_149),
.A2(n_52),
.B(n_28),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_169),
.A2(n_141),
.B1(n_134),
.B2(n_133),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_178),
.A2(n_181),
.B1(n_195),
.B2(n_175),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_168),
.A2(n_136),
.B1(n_138),
.B2(n_144),
.Y(n_179)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_179),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_177),
.A2(n_165),
.B1(n_172),
.B2(n_164),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_183),
.A2(n_188),
.B(n_193),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_170),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_194),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_196),
.C(n_198),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_150),
.Y(n_189)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_190),
.Y(n_207)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_71),
.Y(n_192)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_192),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_157),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_177),
.A2(n_155),
.B1(n_158),
.B2(n_153),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_162),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

INVxp67_ASAP7_75t_SL g200 ( 
.A(n_193),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_200),
.A2(n_213),
.B(n_58),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_156),
.C(n_163),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_218),
.C(n_197),
.Y(n_219)
);

AND2x2_ASAP7_75t_SL g202 ( 
.A(n_180),
.B(n_157),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_202),
.A2(n_217),
.B(n_26),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_154),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_209),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g205 ( 
.A(n_199),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_205),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_173),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_195),
.B(n_160),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_214),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_181),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_174),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_176),
.C(n_85),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_231),
.C(n_233),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_200),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_234),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_182),
.Y(n_223)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_204),
.A2(n_194),
.B1(n_191),
.B2(n_185),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_224),
.A2(n_227),
.B(n_229),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_183),
.C(n_188),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_228),
.C(n_203),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_213),
.A2(n_199),
.B(n_12),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_63),
.C(n_52),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_205),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_202),
.A2(n_0),
.B(n_1),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_202),
.A2(n_81),
.B(n_63),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_218),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_210),
.A2(n_0),
.B(n_1),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_206),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_211),
.A2(n_26),
.B1(n_24),
.B2(n_22),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_212),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_246),
.C(n_248),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_226),
.B(n_208),
.Y(n_237)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_237),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_243),
.Y(n_255)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_240),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_225),
.B(n_10),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_233),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_10),
.C(n_12),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_14),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_231),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_220),
.B(n_14),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_26),
.C(n_24),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_229),
.C(n_228),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_239),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_251),
.B(n_258),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_222),
.Y(n_252)
);

OAI211xp5_ASAP7_75t_L g265 ( 
.A1(n_252),
.A2(n_253),
.B(n_257),
.C(n_258),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_244),
.A2(n_242),
.B1(n_249),
.B2(n_235),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_254),
.A2(n_22),
.B1(n_3),
.B2(n_5),
.Y(n_269)
);

OAI21x1_ASAP7_75t_L g256 ( 
.A1(n_236),
.A2(n_225),
.B(n_232),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_256),
.A2(n_8),
.B(n_11),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_0),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_224),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_2),
.C(n_3),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_248),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_264),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_24),
.Y(n_264)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_265),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_2),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_268),
.C(n_271),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_250),
.A2(n_22),
.B(n_10),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_269),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_9),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_9),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_275),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_277),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_2),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_262),
.C(n_265),
.Y(n_280)
);

OAI21x1_ASAP7_75t_L g283 ( 
.A1(n_280),
.A2(n_282),
.B(n_5),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_278),
.B(n_272),
.C(n_275),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_283),
.A2(n_284),
.B(n_281),
.Y(n_285)
);

NAND2xp33_ASAP7_75t_L g284 ( 
.A(n_279),
.B(n_6),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_6),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_7),
.C(n_17),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_287),
.A2(n_7),
.B(n_17),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_7),
.Y(n_289)
);


endmodule