module fake_jpeg_226_n_132 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_132);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx3_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx6f_ASAP7_75t_SL g40 ( 
.A(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_27),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_60),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_49),
.B(n_44),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_54),
.A2(n_40),
.B1(n_35),
.B2(n_44),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_51),
.B1(n_53),
.B2(n_36),
.Y(n_73)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_67),
.Y(n_77)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_47),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_71),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_64),
.A2(n_52),
.B1(n_58),
.B2(n_63),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_69),
.A2(n_73),
.B1(n_61),
.B2(n_66),
.Y(n_81)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_70),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_42),
.Y(n_71)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_75),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_61),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_59),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_101)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_41),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_86),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_41),
.B(n_46),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_85),
.A2(n_88),
.B(n_0),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_38),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_45),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_87),
.B(n_8),
.Y(n_102)
);

OAI32xp33_ASAP7_75t_L g88 ( 
.A1(n_67),
.A2(n_59),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_85),
.A2(n_74),
.B1(n_72),
.B2(n_70),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_90),
.A2(n_101),
.B1(n_9),
.B2(n_10),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_17),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_100),
.Y(n_106)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_99),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_96),
.A2(n_97),
.B1(n_79),
.B2(n_88),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_89),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_97)
);

NOR2x1_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_5),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_102),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_6),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_20),
.C(n_33),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g104 ( 
.A(n_99),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_105),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_80),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_108),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_9),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_109),
.Y(n_117)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_112),
.C(n_114),
.Y(n_115)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_93),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_113),
.A2(n_14),
.B(n_15),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_13),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_116),
.A2(n_103),
.B(n_111),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_16),
.C(n_19),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_114),
.B(n_106),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_122),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_118),
.A2(n_104),
.B(n_22),
.Y(n_123)
);

OAI21xp33_ASAP7_75t_SL g125 ( 
.A1(n_123),
.A2(n_25),
.B(n_28),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_118),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_117),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_125),
.B(n_127),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_128),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_129),
.A2(n_126),
.B1(n_119),
.B2(n_115),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_29),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_31),
.C(n_34),
.Y(n_132)
);


endmodule