module real_jpeg_4513_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_188;
wire n_33;
wire n_65;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_262;
wire n_19;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_258;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g72 ( 
.A(n_0),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_1),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_19)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_1),
.A2(n_32),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_1),
.A2(n_91),
.B1(n_94),
.B2(n_95),
.Y(n_90)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_1),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_1),
.A2(n_94),
.B1(n_139),
.B2(n_142),
.Y(n_138)
);

O2A1O1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_1),
.A2(n_145),
.B(n_148),
.C(n_151),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_1),
.B(n_25),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_1),
.B(n_137),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_1),
.B(n_101),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_1),
.B(n_119),
.C(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_1),
.B(n_225),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_1),
.B(n_76),
.C(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_2),
.A2(n_174),
.B1(n_175),
.B2(n_177),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_2),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_3),
.Y(n_107)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_3),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_3),
.Y(n_136)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_5),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_5),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_5),
.Y(n_161)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_5),
.Y(n_179)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_6),
.Y(n_147)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_8),
.A2(n_20),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_8),
.A2(n_45),
.B1(n_81),
.B2(n_86),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_8),
.A2(n_45),
.B1(n_130),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_8),
.A2(n_45),
.B1(n_188),
.B2(n_191),
.Y(n_187)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_9),
.Y(n_153)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_10),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_10),
.Y(n_119)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_10),
.Y(n_121)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

OAI22xp5_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_196),
.B1(n_265),
.B2(n_266),
.Y(n_12)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_13),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_194),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_164),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_15),
.B(n_164),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_125),
.C(n_154),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_16),
.B(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_50),
.B2(n_51),
.Y(n_16)
);

INVx2_ASAP7_75t_SL g17 ( 
.A(n_18),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_18),
.B(n_53),
.C(n_89),
.Y(n_193)
);

OA22x2_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_24),
.B1(n_44),
.B2(n_49),
.Y(n_18)
);

OA22x2_ASAP7_75t_L g167 ( 
.A1(n_19),
.A2(n_24),
.B1(n_44),
.B2(n_49),
.Y(n_167)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_34),
.Y(n_24)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_32),
.Y(n_150)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_37),
.B1(n_40),
.B2(n_42),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_89),
.B2(n_124),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_52),
.A2(n_53),
.B1(n_183),
.B2(n_184),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_52),
.B(n_183),
.C(n_236),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_57),
.B1(n_68),
.B2(n_80),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g156 ( 
.A1(n_54),
.A2(n_57),
.B1(n_68),
.B2(n_80),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_L g148 ( 
.A1(n_55),
.A2(n_146),
.B(n_149),
.Y(n_148)
);

NAND2x1_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_68),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_63),
.B1(n_65),
.B2(n_67),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_64),
.Y(n_239)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_68),
.Y(n_225)
);

AOI22x1_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_73),
.B1(n_76),
.B2(n_78),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx8_ASAP7_75t_L g241 ( 
.A(n_74),
.Y(n_241)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_99),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_90),
.B(n_115),
.Y(n_185)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_90),
.Y(n_229)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_93),
.Y(n_190)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_93),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_93),
.Y(n_215)
);

INVx5_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_114),
.Y(n_99)
);

OA22x2_ASAP7_75t_L g227 ( 
.A1(n_100),
.A2(n_114),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_101),
.B(n_187),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NOR2x1_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_105),
.B1(n_108),
.B2(n_112),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

BUFx8_ASAP7_75t_L g176 ( 
.A(n_107),
.Y(n_176)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_120),
.B2(n_122),
.Y(n_116)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_125),
.A2(n_126),
.B1(n_154),
.B2(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_143),
.B2(n_144),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_144),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_127),
.A2(n_128),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_128),
.B(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_128),
.B(n_210),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_128),
.B(n_224),
.C(n_227),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_133),
.B1(n_137),
.B2(n_138),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_129),
.A2(n_133),
.B1(n_138),
.B2(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_129),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_130),
.Y(n_207)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_136),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_138),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_138),
.B(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_154),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.C(n_162),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_155),
.A2(n_156),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_155),
.A2(n_156),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_157),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_157),
.B(n_213),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_157),
.A2(n_158),
.B1(n_162),
.B2(n_163),
.Y(n_255)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_158),
.B(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_160),
.B(n_181),
.Y(n_243)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_170),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_167),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_193),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_183),
.B1(n_184),
.B2(n_192),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_178),
.B(n_180),
.Y(n_172)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_175),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_183),
.A2(n_184),
.B1(n_214),
.B2(n_218),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_183),
.B(n_218),
.Y(n_231)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

AND2x2_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_196),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_259),
.B(n_264),
.Y(n_197)
);

AOI21x1_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_247),
.B(n_258),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_233),
.B(n_246),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_220),
.B(n_232),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_212),
.B(n_219),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_209),
.B(n_211),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_207),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_214),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_231),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_231),
.Y(n_232)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_226),
.B1(n_227),
.B2(n_230),
.Y(n_223)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_224),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_226),
.A2(n_227),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_227),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_250),
.C(n_252),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_235),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_245),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_242),
.B2(n_244),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_244),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_242),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_257),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_257),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_252),
.B1(n_253),
.B2(n_256),
.Y(n_248)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_249),
.Y(n_256)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_250),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_261),
.Y(n_264)
);


endmodule