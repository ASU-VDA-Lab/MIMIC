module fake_jpeg_2433_n_465 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_465);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_465;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_46),
.B(n_61),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_19),
.B(n_16),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_47),
.B(n_55),
.Y(n_127)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_48),
.Y(n_128)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_20),
.B(n_0),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_28),
.B(n_0),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_56),
.B(n_73),
.Y(n_104)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_34),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_81),
.Y(n_93)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_63),
.Y(n_133)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

INVx2_ASAP7_75t_R g73 ( 
.A(n_37),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_76),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_35),
.B(n_16),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_77),
.B(n_78),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_38),
.B(n_16),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_38),
.B(n_0),
.Y(n_81)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_39),
.B(n_1),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_84),
.B(n_1),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_43),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_44),
.Y(n_100)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_21),
.C(n_43),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_92),
.B(n_66),
.C(n_76),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_46),
.A2(n_17),
.B1(n_21),
.B2(n_41),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_94),
.A2(n_119),
.B1(n_126),
.B2(n_145),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_100),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_45),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_106),
.B(n_108),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_51),
.B(n_45),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_58),
.B(n_33),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_115),
.B(n_118),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_61),
.A2(n_21),
.B1(n_41),
.B2(n_36),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_122),
.B1(n_73),
.B2(n_83),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_60),
.B(n_33),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_56),
.A2(n_17),
.B1(n_36),
.B2(n_41),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_56),
.A2(n_17),
.B1(n_32),
.B2(n_36),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_70),
.B(n_17),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_124),
.B(n_49),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_75),
.B(n_44),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_125),
.B(n_129),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_50),
.A2(n_42),
.B1(n_40),
.B2(n_27),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_50),
.A2(n_40),
.B1(n_27),
.B2(n_3),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_130),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_199)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_137),
.Y(n_190)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_48),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_138),
.B(n_140),
.Y(n_195)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_74),
.Y(n_139)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_79),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_72),
.Y(n_141)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_62),
.B(n_1),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_143),
.B(n_6),
.Y(n_201)
);

NAND3xp33_ASAP7_75t_L g180 ( 
.A(n_144),
.B(n_2),
.C(n_3),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_52),
.A2(n_27),
.B1(n_23),
.B2(n_4),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_92),
.B(n_85),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_148),
.B(n_161),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_126),
.A2(n_73),
.B1(n_83),
.B2(n_80),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_149),
.A2(n_150),
.B1(n_184),
.B2(n_199),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_117),
.A2(n_53),
.B1(n_80),
.B2(n_76),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_152),
.A2(n_135),
.B1(n_123),
.B2(n_101),
.Y(n_208)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_116),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_153),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_91),
.Y(n_154)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_154),
.Y(n_210)
);

A2O1A1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_127),
.A2(n_69),
.B(n_57),
.C(n_63),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g246 ( 
.A1(n_155),
.A2(n_156),
.B(n_180),
.Y(n_246)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_158),
.Y(n_245)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_159),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_104),
.B(n_52),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_160),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_90),
.B(n_71),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_116),
.Y(n_163)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_163),
.Y(n_215)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_107),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_164),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_146),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_165),
.B(n_169),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_104),
.B(n_71),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_166),
.B(n_191),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_96),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_167),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_146),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_171),
.B(n_192),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_93),
.A2(n_87),
.B1(n_82),
.B2(n_68),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_172),
.A2(n_194),
.B1(n_200),
.B2(n_7),
.Y(n_238)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_128),
.Y(n_173)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_173),
.Y(n_220)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_107),
.Y(n_174)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_174),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_88),
.B(n_57),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_175),
.B(n_176),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_95),
.B(n_57),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_134),
.Y(n_177)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_177),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_132),
.B(n_68),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_178),
.B(n_187),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_98),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_181),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_105),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_98),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_183),
.B(n_188),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_94),
.A2(n_67),
.B1(n_66),
.B2(n_54),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_105),
.B(n_111),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_185),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_97),
.Y(n_186)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_186),
.Y(n_227)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_122),
.A2(n_65),
.B(n_23),
.C(n_5),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_136),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_99),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_196),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_103),
.B(n_67),
.Y(n_191)
);

BUFx12f_ASAP7_75t_L g193 ( 
.A(n_111),
.Y(n_193)
);

INVx11_ASAP7_75t_L g214 ( 
.A(n_193),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_109),
.A2(n_112),
.B1(n_114),
.B2(n_141),
.Y(n_194)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_101),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_89),
.Y(n_197)
);

INVx11_ASAP7_75t_L g236 ( 
.A(n_197),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_130),
.A2(n_54),
.B(n_53),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_102),
.C(n_131),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_89),
.Y(n_200)
);

OAI211xp5_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_23),
.B(n_110),
.C(n_133),
.Y(n_222)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_137),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_120),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_148),
.A2(n_145),
.B1(n_135),
.B2(n_123),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_207),
.A2(n_216),
.B1(n_217),
.B2(n_233),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_208),
.A2(n_227),
.B1(n_245),
.B2(n_203),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_110),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_209),
.B(n_219),
.C(n_229),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_211),
.B(n_232),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_150),
.A2(n_97),
.B1(n_131),
.B2(n_102),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_166),
.B(n_133),
.C(n_113),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_222),
.B(n_163),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_195),
.Y(n_224)
);

OAI21xp33_ASAP7_75t_L g287 ( 
.A1(n_224),
.A2(n_239),
.B(n_244),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_162),
.B(n_113),
.C(n_142),
.Y(n_229)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_230),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_152),
.A2(n_142),
.B1(n_120),
.B2(n_23),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_231),
.A2(n_249),
.B1(n_175),
.B2(n_176),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_162),
.B(n_23),
.C(n_8),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_191),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_161),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_237),
.A2(n_173),
.B1(n_188),
.B2(n_177),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_238),
.A2(n_244),
.B1(n_215),
.B2(n_193),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_185),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_160),
.B(n_7),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_242),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_160),
.B(n_8),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_185),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_157),
.B(n_9),
.C(n_12),
.Y(n_248)
);

A2O1A1O1Ixp25_ASAP7_75t_L g271 ( 
.A1(n_248),
.A2(n_151),
.B(n_174),
.C(n_193),
.D(n_13),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_187),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_170),
.B(n_12),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_250),
.B(n_12),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_221),
.Y(n_252)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_252),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_253),
.A2(n_254),
.B1(n_259),
.B2(n_277),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_205),
.A2(n_198),
.B1(n_199),
.B2(n_196),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_226),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_256),
.B(n_269),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_205),
.B(n_182),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_257),
.B(n_268),
.Y(n_328)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_228),
.Y(n_258)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_258),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_213),
.A2(n_155),
.B1(n_189),
.B2(n_158),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_261),
.A2(n_263),
.B1(n_264),
.B2(n_283),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_235),
.A2(n_153),
.B(n_164),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_262),
.A2(n_223),
.B(n_215),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_239),
.A2(n_202),
.B1(n_147),
.B2(n_190),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_220),
.Y(n_265)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_265),
.Y(n_314)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_214),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_266),
.Y(n_317)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_227),
.Y(n_267)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_267),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_224),
.B(n_168),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_181),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_271),
.A2(n_276),
.B(n_236),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_204),
.Y(n_272)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_272),
.Y(n_324)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_220),
.Y(n_273)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_273),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_218),
.B(n_240),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_274),
.B(n_279),
.Y(n_315)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_225),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_275),
.B(n_278),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_246),
.A2(n_151),
.B(n_147),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_213),
.A2(n_167),
.B1(n_154),
.B2(n_186),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_225),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_218),
.A2(n_159),
.B1(n_190),
.B2(n_197),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_281),
.A2(n_286),
.B1(n_291),
.B2(n_293),
.Y(n_299)
);

BUFx8_ASAP7_75t_L g282 ( 
.A(n_214),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_282),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_211),
.A2(n_200),
.B1(n_13),
.B2(n_15),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_284),
.A2(n_234),
.B1(n_210),
.B2(n_248),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_212),
.B(n_219),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_285),
.B(n_290),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_212),
.A2(n_241),
.B1(n_231),
.B2(n_207),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_232),
.B(n_229),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_288),
.B(n_289),
.Y(n_319)
);

INVx13_ASAP7_75t_L g289 ( 
.A(n_243),
.Y(n_289)
);

A2O1A1Ixp33_ASAP7_75t_L g290 ( 
.A1(n_241),
.A2(n_242),
.B(n_217),
.C(n_209),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_243),
.A2(n_249),
.B1(n_216),
.B2(n_208),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_233),
.B(n_237),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_292),
.B(n_281),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_255),
.B(n_230),
.C(n_206),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_295),
.B(n_302),
.C(n_312),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_287),
.A2(n_206),
.B(n_223),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_296),
.B(n_297),
.Y(n_340)
);

AOI22x1_ASAP7_75t_L g300 ( 
.A1(n_259),
.A2(n_203),
.B1(n_234),
.B2(n_245),
.Y(n_300)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_300),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_255),
.B(n_247),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_304),
.B(n_305),
.Y(n_333)
);

OA22x2_ASAP7_75t_L g305 ( 
.A1(n_260),
.A2(n_210),
.B1(n_236),
.B2(n_251),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_306),
.B(n_282),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_290),
.A2(n_276),
.B(n_285),
.Y(n_307)
);

FAx1_ASAP7_75t_SL g336 ( 
.A(n_307),
.B(n_316),
.CI(n_313),
.CON(n_336),
.SN(n_336)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_262),
.A2(n_256),
.B(n_284),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_308),
.B(n_326),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_280),
.B(n_251),
.C(n_272),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_280),
.B(n_258),
.C(n_286),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_313),
.B(n_320),
.Y(n_347)
);

MAJx2_ASAP7_75t_L g316 ( 
.A(n_257),
.B(n_274),
.C(n_270),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_260),
.A2(n_292),
.B1(n_254),
.B2(n_291),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_318),
.B(n_322),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_270),
.B(n_279),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_277),
.A2(n_293),
.B1(n_264),
.B2(n_253),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_323),
.B(n_327),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_265),
.A2(n_275),
.B1(n_278),
.B2(n_273),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_325),
.A2(n_282),
.B1(n_299),
.B2(n_294),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_289),
.B(n_271),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_326),
.B(n_330),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_267),
.B(n_266),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_282),
.B(n_267),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_332),
.A2(n_346),
.B(n_296),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_334),
.A2(n_337),
.B1(n_341),
.B2(n_360),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_309),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_335),
.B(n_336),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_294),
.A2(n_299),
.B1(n_323),
.B2(n_310),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_309),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_338),
.B(n_345),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_301),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g367 ( 
.A(n_339),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_310),
.A2(n_318),
.B1(n_307),
.B2(n_305),
.Y(n_341)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_325),
.Y(n_344)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_344),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_327),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_311),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_348),
.B(n_352),
.Y(n_377)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_314),
.Y(n_350)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_350),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_317),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_324),
.B(n_331),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_353),
.B(n_354),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_315),
.B(n_331),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_320),
.B(n_312),
.Y(n_355)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_355),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_321),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_356),
.Y(n_371)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_329),
.Y(n_357)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_357),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_295),
.B(n_319),
.Y(n_358)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_358),
.Y(n_384)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_305),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_359),
.B(n_300),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_305),
.A2(n_322),
.B1(n_306),
.B2(n_297),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_316),
.B(n_308),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_361),
.A2(n_349),
.B1(n_348),
.B2(n_354),
.Y(n_373)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_363),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_337),
.A2(n_342),
.B1(n_334),
.B2(n_360),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_365),
.A2(n_369),
.B1(n_364),
.B2(n_385),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_366),
.B(n_373),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_342),
.A2(n_298),
.B1(n_302),
.B2(n_304),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_347),
.B(n_330),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_370),
.B(n_376),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_362),
.B(n_300),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_362),
.B(n_303),
.C(n_317),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_378),
.B(n_388),
.C(n_340),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_347),
.B(n_349),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_380),
.B(n_381),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_341),
.B(n_336),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_SL g383 ( 
.A(n_336),
.B(n_343),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_383),
.B(n_387),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_351),
.A2(n_359),
.B1(n_333),
.B2(n_340),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_385),
.A2(n_335),
.B(n_352),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_343),
.B(n_333),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_340),
.B(n_344),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_389),
.B(n_393),
.C(n_383),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_363),
.B(n_351),
.Y(n_390)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_390),
.Y(n_427)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_384),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_391),
.B(n_392),
.Y(n_425)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_377),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_378),
.B(n_380),
.C(n_376),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_395),
.A2(n_365),
.B1(n_369),
.B2(n_379),
.Y(n_416)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_375),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_396),
.B(n_397),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_375),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_388),
.A2(n_345),
.B(n_338),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_398),
.A2(n_403),
.B(n_394),
.Y(n_411)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_372),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_402),
.B(n_404),
.Y(n_421)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_382),
.Y(n_404)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_387),
.Y(n_406)
);

INVx13_ASAP7_75t_L g414 ( 
.A(n_406),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_368),
.B(n_356),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_407),
.A2(n_409),
.B1(n_398),
.B2(n_404),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_367),
.B(n_350),
.Y(n_408)
);

INVx13_ASAP7_75t_L g417 ( 
.A(n_408),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_371),
.Y(n_409)
);

INVx13_ASAP7_75t_L g419 ( 
.A(n_409),
.Y(n_419)
);

A2O1A1Ixp33_ASAP7_75t_L g410 ( 
.A1(n_396),
.A2(n_374),
.B(n_363),
.C(n_381),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_410),
.A2(n_411),
.B(n_412),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_403),
.A2(n_366),
.B(n_364),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g413 ( 
.A(n_401),
.B(n_370),
.Y(n_413)
);

XNOR2x1_ASAP7_75t_L g437 ( 
.A(n_413),
.B(n_424),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_415),
.B(n_401),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_416),
.A2(n_422),
.B1(n_400),
.B2(n_405),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_393),
.B(n_386),
.C(n_371),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_420),
.B(n_426),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_395),
.A2(n_357),
.B1(n_394),
.B2(n_390),
.Y(n_422)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_423),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_390),
.A2(n_399),
.B(n_389),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_406),
.A2(n_391),
.B1(n_407),
.B2(n_402),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_421),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_429),
.B(n_430),
.Y(n_447)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_431),
.Y(n_445)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_421),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_432),
.B(n_439),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_420),
.B(n_400),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_433),
.B(n_435),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_411),
.A2(n_412),
.B(n_418),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_416),
.A2(n_405),
.B1(n_422),
.B2(n_418),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_438),
.A2(n_427),
.B1(n_410),
.B2(n_419),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_425),
.B(n_426),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_433),
.B(n_425),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_442),
.B(n_443),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_436),
.B(n_424),
.C(n_415),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_444),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_430),
.B(n_427),
.C(n_423),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_446),
.B(n_434),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_435),
.B(n_410),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_448),
.B(n_434),
.C(n_438),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_449),
.A2(n_454),
.B(n_443),
.Y(n_457)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_440),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_451),
.A2(n_441),
.B1(n_445),
.B2(n_417),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_453),
.A2(n_441),
.B1(n_431),
.B2(n_446),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_447),
.B(n_428),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_455),
.B(n_456),
.C(n_457),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_450),
.A2(n_448),
.B(n_414),
.Y(n_458)
);

AO221x1_ASAP7_75t_L g460 ( 
.A1(n_458),
.A2(n_417),
.B1(n_419),
.B2(n_414),
.C(n_421),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_460),
.A2(n_452),
.B(n_437),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_461),
.A2(n_459),
.B(n_452),
.Y(n_462)
);

A2O1A1Ixp33_ASAP7_75t_L g463 ( 
.A1(n_462),
.A2(n_419),
.B(n_417),
.C(n_414),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_463),
.B(n_437),
.C(n_413),
.Y(n_464)
);

FAx1_ASAP7_75t_SL g465 ( 
.A(n_464),
.B(n_413),
.CI(n_459),
.CON(n_465),
.SN(n_465)
);


endmodule