module real_jpeg_23282_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_0),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_0),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_0),
.A2(n_22),
.B1(n_27),
.B2(n_82),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_0),
.A2(n_64),
.B1(n_66),
.B2(n_82),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_0),
.A2(n_52),
.B1(n_59),
.B2(n_82),
.Y(n_232)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_2),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_2),
.B(n_21),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_2),
.B(n_64),
.C(n_93),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_2),
.A2(n_22),
.B1(n_27),
.B2(n_194),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_2),
.B(n_135),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_2),
.A2(n_64),
.B1(n_66),
.B2(n_194),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_2),
.B(n_52),
.C(n_69),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_2),
.A2(n_51),
.B(n_281),
.Y(n_311)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_4),
.A2(n_30),
.B1(n_33),
.B2(n_170),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_4),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_4),
.A2(n_22),
.B1(n_27),
.B2(n_170),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_4),
.A2(n_64),
.B1(n_66),
.B2(n_170),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_4),
.A2(n_52),
.B1(n_59),
.B2(n_170),
.Y(n_294)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_7),
.A2(n_36),
.B1(n_52),
.B2(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_7),
.A2(n_36),
.B1(n_64),
.B2(n_66),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_7),
.A2(n_22),
.B1(n_27),
.B2(n_36),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_120),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_8),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_8),
.A2(n_22),
.B1(n_27),
.B2(n_120),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_8),
.A2(n_64),
.B1(n_66),
.B2(n_120),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_8),
.A2(n_52),
.B1(n_59),
.B2(n_120),
.Y(n_280)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_9),
.Y(n_93)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_11),
.A2(n_22),
.B1(n_27),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_11),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_11),
.A2(n_64),
.B1(n_66),
.B2(n_97),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_11),
.A2(n_32),
.B1(n_81),
.B2(n_97),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_11),
.A2(n_52),
.B1(n_59),
.B2(n_97),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_13),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_13),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_13),
.A2(n_22),
.B1(n_27),
.B2(n_63),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_13),
.A2(n_33),
.B1(n_63),
.B2(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_13),
.A2(n_52),
.B1(n_59),
.B2(n_63),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_14),
.A2(n_40),
.B1(n_64),
.B2(n_66),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_14),
.A2(n_40),
.B1(n_52),
.B2(n_59),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_14),
.A2(n_22),
.B1(n_27),
.B2(n_40),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_15),
.A2(n_81),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_15),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_15),
.A2(n_22),
.B1(n_27),
.B2(n_87),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_15),
.A2(n_64),
.B1(n_66),
.B2(n_87),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_15),
.A2(n_52),
.B1(n_59),
.B2(n_87),
.Y(n_251)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_16),
.Y(n_110)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_16),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_43),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_41),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_37),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_20),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_28),
.B(n_35),
.Y(n_20)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_21),
.A2(n_28),
.B1(n_35),
.B2(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_21),
.A2(n_28),
.B1(n_119),
.B2(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_21),
.A2(n_28),
.B1(n_39),
.B2(n_353),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_21)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_22),
.A2(n_27),
.B1(n_93),
.B2(n_94),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g192 ( 
.A1(n_22),
.A2(n_26),
.B(n_193),
.C(n_195),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_22),
.B(n_247),
.Y(n_246)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_26),
.B1(n_30),
.B2(n_33),
.Y(n_29)
);

NAND3xp33_ASAP7_75t_SL g195 ( 
.A(n_25),
.B(n_27),
.C(n_33),
.Y(n_195)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_28),
.B(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_28),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_28),
.A2(n_123),
.B(n_222),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_34),
.Y(n_28)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_33),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_34),
.A2(n_78),
.B(n_83),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_34),
.B(n_85),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_34),
.A2(n_78),
.B1(n_121),
.B2(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_34),
.A2(n_121),
.B1(n_143),
.B2(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_34),
.A2(n_83),
.B(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_38),
.B(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_38),
.B(n_359),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_358),
.B(n_360),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_346),
.B(n_357),
.Y(n_44)
);

OAI31xp33_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_145),
.A3(n_160),
.B(n_343),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_124),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_47),
.B(n_124),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_88),
.C(n_104),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_48),
.A2(n_88),
.B1(n_89),
.B2(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_48),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_74),
.Y(n_48)
);

AOI21xp33_ASAP7_75t_L g125 ( 
.A1(n_49),
.A2(n_50),
.B(n_76),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_60),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_50),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_50),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_50),
.A2(n_60),
.B1(n_61),
.B2(n_75),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_55),
.B(n_58),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_51),
.A2(n_58),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_51),
.A2(n_109),
.B1(n_110),
.B2(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_51),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_51),
.A2(n_110),
.B1(n_199),
.B2(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_51),
.B(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_51),
.A2(n_280),
.B(n_281),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_54),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_52),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_52),
.A2(n_59),
.B1(n_69),
.B2(n_70),
.Y(n_71)
);

BUFx4f_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_54),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g304 ( 
.A(n_54),
.Y(n_304)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_56),
.A2(n_249),
.B(n_250),
.Y(n_248)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_59),
.B(n_308),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_67),
.B1(n_72),
.B2(n_73),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_62),
.A2(n_67),
.B1(n_73),
.B2(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_64),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_64),
.A2(n_66),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_64),
.A2(n_66),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_64),
.B(n_289),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_67),
.A2(n_73),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_67),
.B(n_220),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_67),
.A2(n_73),
.B1(n_253),
.B2(n_255),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_71),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_71),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_71),
.A2(n_100),
.B1(n_114),
.B2(n_180),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_71),
.A2(n_180),
.B(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_71),
.A2(n_219),
.B(n_254),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_71),
.B(n_194),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_72),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_73),
.B(n_220),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g193 ( 
.A(n_80),
.B(n_194),
.Y(n_193)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_SL g222 ( 
.A1(n_81),
.A2(n_193),
.B(n_194),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_99),
.B(n_103),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_99),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_96),
.B2(n_98),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_91),
.A2(n_92),
.B1(n_96),
.B2(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_91),
.A2(n_92),
.B1(n_137),
.B2(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_91),
.A2(n_187),
.B(n_189),
.Y(n_186)
);

OAI21xp33_ASAP7_75t_L g257 ( 
.A1(n_91),
.A2(n_189),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_92),
.A2(n_116),
.B(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_92),
.A2(n_173),
.B(n_228),
.Y(n_227)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_98),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_100),
.A2(n_268),
.B(n_269),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_100),
.A2(n_269),
.B(n_287),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_102),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_104),
.A2(n_105),
.B1(n_338),
.B2(n_340),
.Y(n_337)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_115),
.C(n_117),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_106),
.A2(n_107),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_111),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_108),
.A2(n_111),
.B1(n_112),
.B2(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_108),
.Y(n_182)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_110),
.Y(n_200)
);

INVx5_ASAP7_75t_L g310 ( 
.A(n_110),
.Y(n_310)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_115),
.B(n_117),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_121),
.B(n_122),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_127),
.C(n_129),
.Y(n_159)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_142),
.B2(n_144),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_138),
.B1(n_139),
.B2(n_141),
.Y(n_131)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_132),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_139),
.C(n_142),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_134),
.A2(n_135),
.B1(n_188),
.B2(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_134),
.A2(n_135),
.B(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_135),
.B(n_174),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_138),
.A2(n_139),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_139),
.B(n_152),
.C(n_157),
.Y(n_356)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_142),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_142),
.A2(n_144),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_142),
.B(n_148),
.C(n_151),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_146),
.A2(n_344),
.B(n_345),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_159),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_147),
.B(n_159),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_153),
.Y(n_353)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_158),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_336),
.B(n_342),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_208),
.B(n_335),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_201),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_163),
.B(n_201),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_181),
.C(n_183),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_164),
.A2(n_165),
.B1(n_181),
.B2(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_175),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_171),
.B2(n_172),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_171),
.C(n_175),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_169),
.Y(n_185)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_179),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_176),
.B(n_179),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_178),
.A2(n_197),
.B1(n_198),
.B2(n_200),
.Y(n_196)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_181),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_183),
.B(n_332),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.C(n_190),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_184),
.B(n_186),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_190),
.B(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_196),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_191),
.A2(n_192),
.B1(n_196),
.B2(n_225),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_194),
.B(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_196),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_197),
.A2(n_293),
.B1(n_295),
.B2(n_297),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_207),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_203),
.B(n_204),
.C(n_207),
.Y(n_341)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

O2A1O1Ixp33_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_239),
.B(n_329),
.C(n_334),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_233),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_233),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_223),
.C(n_226),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_211),
.A2(n_212),
.B1(n_324),
.B2(n_325),
.Y(n_323)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_221),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_217),
.B2(n_218),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_217),
.C(n_221),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_216),
.Y(n_228)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_223),
.A2(n_224),
.B1(n_226),
.B2(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_226),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.C(n_231),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_227),
.B(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_229),
.A2(n_230),
.B1(n_231),
.B2(n_263),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_231),
.Y(n_263)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_234),
.B(n_237),
.C(n_238),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_322),
.B(n_328),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_270),
.B(n_321),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_259),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_244),
.B(n_259),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_252),
.C(n_256),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_245),
.B(n_317),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_248),
.Y(n_266)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_250),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_251),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_252),
.A2(n_256),
.B1(n_257),
.B2(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_252),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_255),
.Y(n_268)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_264),
.B2(n_265),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_260),
.B(n_266),
.C(n_267),
.Y(n_327)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_315),
.B(n_320),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_290),
.B(n_314),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_284),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_273),
.B(n_284),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_279),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_275),
.B(n_278),
.C(n_279),
.Y(n_319)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_288),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_285),
.A2(n_286),
.B1(n_288),
.B2(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_288),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_300),
.B(n_313),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_298),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_292),
.B(n_298),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_294),
.A2(n_304),
.B(n_305),
.Y(n_303)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_306),
.B(n_312),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_303),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_311),
.Y(n_306)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_319),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_319),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_327),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_327),
.Y(n_328)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_330),
.B(n_331),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_337),
.B(n_341),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_337),
.B(n_341),
.Y(n_342)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_338),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_347),
.B(n_348),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_356),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_350),
.A2(n_352),
.B1(n_354),
.B2(n_355),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_350),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_352),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_352),
.B(n_354),
.C(n_356),
.Y(n_359)
);


endmodule