module fake_jpeg_32112_n_38 (n_3, n_2, n_1, n_0, n_4, n_5, n_38);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_38;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_3),
.Y(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

BUFx5_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_6),
.B(n_0),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_19),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_15)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_15),
.A2(n_18),
.B(n_6),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_7),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_16),
.A2(n_15),
.B1(n_12),
.B2(n_10),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_4),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_12),
.C(n_10),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_8),
.A2(n_5),
.B(n_11),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_23),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_25),
.Y(n_26)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_29),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_24),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_32),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_20),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_27),
.B(n_26),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_26),
.B1(n_25),
.B2(n_17),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_35),
.A2(n_22),
.B(n_23),
.Y(n_36)
);

OAI32xp33_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_34),
.A3(n_30),
.B1(n_13),
.B2(n_16),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_12),
.B1(n_19),
.B2(n_5),
.Y(n_38)
);


endmodule