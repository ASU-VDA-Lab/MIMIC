module fake_aes_501_n_20 (n_1, n_2, n_0, n_20);
input n_1;
input n_2;
input n_0;
output n_20;
wire n_5;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_3;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_6;
wire n_4;
wire n_7;
INVx2_ASAP7_75t_L g3 ( .A(n_0), .Y(n_3) );
NAND2xp5_ASAP7_75t_SL g4 ( .A(n_2), .B(n_1), .Y(n_4) );
NAND2xp5_ASAP7_75t_SL g5 ( .A(n_0), .B(n_1), .Y(n_5) );
NOR2xp33_ASAP7_75t_L g6 ( .A(n_3), .B(n_0), .Y(n_6) );
INVxp67_ASAP7_75t_L g7 ( .A(n_4), .Y(n_7) );
AOI21xp5_ASAP7_75t_L g8 ( .A1(n_5), .A2(n_0), .B(n_1), .Y(n_8) );
OR2x2_ASAP7_75t_L g9 ( .A(n_7), .B(n_0), .Y(n_9) );
INVx2_ASAP7_75t_L g10 ( .A(n_6), .Y(n_10) );
BUFx6f_ASAP7_75t_L g11 ( .A(n_8), .Y(n_11) );
AND2x2_ASAP7_75t_L g12 ( .A(n_10), .B(n_8), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_11), .Y(n_13) );
OAI221xp5_ASAP7_75t_L g14 ( .A1(n_12), .A2(n_9), .B1(n_10), .B2(n_11), .C(n_2), .Y(n_14) );
OA211x2_ASAP7_75t_L g15 ( .A1(n_12), .A2(n_11), .B(n_1), .C(n_2), .Y(n_15) );
OAI22x1_ASAP7_75t_L g16 ( .A1(n_15), .A2(n_12), .B1(n_13), .B2(n_1), .Y(n_16) );
NOR5xp2_ASAP7_75t_SL g17 ( .A(n_15), .B(n_2), .C(n_11), .D(n_13), .E(n_14), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_16), .Y(n_18) );
AO22x2_ASAP7_75t_L g19 ( .A1(n_17), .A2(n_2), .B1(n_13), .B2(n_16), .Y(n_19) );
OAI21x1_ASAP7_75t_L g20 ( .A1(n_18), .A2(n_17), .B(n_19), .Y(n_20) );
endmodule