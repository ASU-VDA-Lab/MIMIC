module fake_jpeg_5907_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_59;
wire n_20;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_9),
.B(n_3),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_8),
.B(n_4),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

HAxp5_ASAP7_75t_SL g19 ( 
.A(n_2),
.B(n_1),
.CON(n_19),
.SN(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVxp33_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_23),
.B(n_25),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_19),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_24),
.A2(n_19),
.B1(n_14),
.B2(n_16),
.Y(n_30)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_12),
.B(n_3),
.Y(n_28)
);

BUFx24_ASAP7_75t_SL g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2x1_ASAP7_75t_R g48 ( 
.A(n_30),
.B(n_17),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_23),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_34),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_28),
.Y(n_35)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_16),
.B(n_11),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_42),
.C(n_45),
.Y(n_50)
);

BUFx24_ASAP7_75t_SL g42 ( 
.A(n_38),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_21),
.C(n_22),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_21),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_49),
.C(n_34),
.Y(n_52)
);

AO22x1_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_18),
.B1(n_10),
.B2(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_56),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_29),
.C(n_22),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_54),
.C(n_44),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_29),
.C(n_37),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_SL g59 ( 
.A(n_55),
.B(n_46),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_35),
.B1(n_25),
.B2(n_26),
.Y(n_56)
);

NAND3xp33_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_43),
.C(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_58),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_36),
.B1(n_25),
.B2(n_18),
.Y(n_64)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_60),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_SL g62 ( 
.A(n_51),
.B(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_4),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_65),
.A2(n_57),
.B(n_61),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_66),
.B(n_65),
.C(n_63),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_69),
.A2(n_70),
.B(n_5),
.Y(n_71)
);

OAI21x1_ASAP7_75t_SL g70 ( 
.A1(n_68),
.A2(n_20),
.B(n_5),
.Y(n_70)
);

AO21x1_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_7),
.B(n_20),
.Y(n_72)
);


endmodule