module fake_jpeg_24577_n_103 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_103);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_103;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx6_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_24),
.B(n_23),
.Y(n_33)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_28),
.Y(n_40)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_0),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_31),
.B(n_32),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_24),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_21),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_11),
.B1(n_18),
.B2(n_16),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_11),
.B1(n_14),
.B2(n_30),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_31),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_24),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_53),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_44),
.B(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_51),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_47),
.B(n_50),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_32),
.B1(n_26),
.B2(n_30),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_52),
.B(n_57),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_49),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_16),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_25),
.B1(n_27),
.B2(n_15),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_1),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_25),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_19),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_55),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_21),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_27),
.B1(n_23),
.B2(n_19),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_38),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_12),
.B1(n_17),
.B2(n_35),
.Y(n_57)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_60),
.Y(n_76)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

NOR3xp33_ASAP7_75t_SL g61 ( 
.A(n_57),
.B(n_17),
.C(n_12),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_67),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_56),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_38),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_67),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_72),
.B(n_68),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_64),
.A2(n_48),
.B(n_52),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_63),
.A2(n_58),
.B1(n_65),
.B2(n_60),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_69),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_74),
.B(n_75),
.Y(n_82)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_48),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_48),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_78),
.B(n_61),
.Y(n_80)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_80),
.Y(n_89)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_70),
.Y(n_84)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_85),
.A2(n_73),
.B1(n_78),
.B2(n_77),
.Y(n_88)
);

INVxp33_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_83),
.Y(n_94)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

OR2x2_ASAP7_75t_SL g92 ( 
.A(n_87),
.B(n_71),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_93),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_89),
.Y(n_93)
);

AOI322xp5_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_90),
.A3(n_86),
.B1(n_83),
.B2(n_81),
.C1(n_13),
.C2(n_20),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_97),
.Y(n_98)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g97 ( 
.A1(n_92),
.A2(n_44),
.B(n_2),
.C(n_1),
.D(n_8),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_91),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_99),
.A2(n_7),
.B(n_2),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_98),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_100)
);

NAND3xp33_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_101),
.C(n_2),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_99),
.Y(n_103)
);


endmodule