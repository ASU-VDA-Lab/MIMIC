module fake_jpeg_13863_n_29 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_29);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_29;

wire n_13;
wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_15;

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_7),
.B(n_9),
.Y(n_11)
);

INVx5_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx13_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

NAND2xp33_ASAP7_75t_SL g20 ( 
.A(n_15),
.B(n_17),
.Y(n_20)
);

OA22x2_ASAP7_75t_L g16 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_16),
.B(n_3),
.Y(n_18)
);

AO22x2_ASAP7_75t_SL g17 ( 
.A1(n_13),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_18),
.A2(n_19),
.B(n_12),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_15),
.B(n_12),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_21),
.A2(n_23),
.B(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_19),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_11),
.C(n_13),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_6),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_25),
.A2(n_13),
.B(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_27),
.C(n_10),
.Y(n_29)
);


endmodule