module fake_ariane_2878_n_2350 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2350);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2350;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_373;
wire n_2135;
wire n_2334;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_2207;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_2248;
wire n_813;
wire n_419;
wire n_1985;
wire n_2288;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_2322;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_1944;
wire n_331;
wire n_559;
wire n_2233;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_2332;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_249;
wire n_1108;
wire n_355;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_2185;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_967;
wire n_1083;
wire n_274;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_382;
wire n_489;
wire n_2294;
wire n_2274;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_307;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_2328;
wire n_347;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_479;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_299;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_2262;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_2168;
wire n_552;
wire n_348;
wire n_2312;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_502;
wire n_2194;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_2218;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_2184;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_321;
wire n_221;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_2300;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_2266;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2211;
wire n_2292;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_2306;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_2348;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2320;
wire n_979;
wire n_2329;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2314;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_2285;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_2173;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_330;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2331;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_601;
wire n_236;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2196;
wire n_1038;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_2303;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_223;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2270;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_2251;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2321;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_399;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_2212;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_2268;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2252;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2260;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_2206;
wire n_997;
wire n_635;
wire n_1902;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_2339;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_371;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_2209;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_2318;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_1010;
wire n_882;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_2336;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

BUFx8_ASAP7_75t_SL g219 ( 
.A(n_77),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_152),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_173),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_23),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_29),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_67),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_166),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_153),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_105),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_175),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_106),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_149),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_44),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_53),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_116),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_143),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_183),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_9),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_130),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_41),
.Y(n_238)
);

INVxp67_ASAP7_75t_SL g239 ( 
.A(n_38),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_161),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_19),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_214),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_108),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_97),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_205),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_186),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_93),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_177),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_140),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_78),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_36),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_216),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_90),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_92),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_194),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_204),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_4),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_42),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_0),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_197),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_75),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_32),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_39),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_90),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_120),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_85),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_1),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_200),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_127),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_3),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_193),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_14),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_168),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_151),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_179),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_78),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_124),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_70),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_134),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_154),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_190),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_70),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_6),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_86),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_189),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_158),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_82),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_29),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_31),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_65),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_79),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_23),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_12),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_2),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_136),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_89),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_18),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_69),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_34),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_69),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_30),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_180),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_169),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_165),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_76),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_163),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_104),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_67),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_103),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_16),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_82),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_199),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_88),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_44),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_156),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_133),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_203),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_8),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_159),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_9),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_75),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_46),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_7),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_97),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_63),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_181),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_12),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_36),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_174),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_195),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_217),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_182),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_210),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_207),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_31),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_110),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_60),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_15),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_46),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_94),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_113),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_45),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_32),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_66),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_147),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_184),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g347 ( 
.A(n_187),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_202),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_54),
.Y(n_349)
);

BUFx2_ASAP7_75t_SL g350 ( 
.A(n_191),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_80),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_122),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_96),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_57),
.Y(n_354)
);

BUFx10_ASAP7_75t_L g355 ( 
.A(n_155),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_43),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_94),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_83),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_66),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_20),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_54),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_176),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_93),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_138),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_92),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_85),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_129),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_59),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_119),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_86),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_208),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_22),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_81),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_212),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_34),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_3),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_213),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_74),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_20),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_22),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_142),
.Y(n_381)
);

INVxp33_ASAP7_75t_L g382 ( 
.A(n_101),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_59),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_27),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_28),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_11),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_131),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_51),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_24),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_218),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_209),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_198),
.Y(n_392)
);

BUFx10_ASAP7_75t_L g393 ( 
.A(n_7),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_49),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_135),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_5),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_58),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_172),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_72),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_2),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_79),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_80),
.Y(n_402)
);

INVx2_ASAP7_75t_SL g403 ( 
.A(n_71),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_0),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_39),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_112),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_89),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_43),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_50),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_13),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_77),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_115),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_45),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_61),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_13),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_88),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_87),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_6),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_96),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_4),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_100),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_81),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_60),
.Y(n_423)
);

BUFx10_ASAP7_75t_L g424 ( 
.A(n_15),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_201),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_157),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_25),
.Y(n_427)
);

BUFx10_ASAP7_75t_L g428 ( 
.A(n_42),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_19),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_188),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_196),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_237),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_273),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_351),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_351),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_219),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_230),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_248),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_279),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_306),
.Y(n_440)
);

INVxp67_ASAP7_75t_SL g441 ( 
.A(n_223),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_237),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_240),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_316),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_240),
.B(n_1),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_252),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g447 ( 
.A(n_276),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_331),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_252),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_222),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_260),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_260),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_268),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_352),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_268),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_381),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_303),
.B(n_5),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_430),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_277),
.B(n_8),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_232),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_241),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_301),
.Y(n_462)
);

INVxp67_ASAP7_75t_SL g463 ( 
.A(n_223),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_277),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_238),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_284),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_244),
.Y(n_467)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_301),
.B(n_10),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_247),
.Y(n_469)
);

NOR2xp67_ASAP7_75t_L g470 ( 
.A(n_403),
.B(n_10),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_250),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_315),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_315),
.B(n_11),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_319),
.B(n_14),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_261),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_251),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_253),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_319),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_324),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_325),
.Y(n_480)
);

NOR2xp67_ASAP7_75t_L g481 ( 
.A(n_403),
.B(n_16),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_357),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_257),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_329),
.B(n_17),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_329),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_259),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_333),
.Y(n_487)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_273),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_263),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_376),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_301),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_333),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_264),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_266),
.Y(n_494)
);

INVxp67_ASAP7_75t_SL g495 ( 
.A(n_224),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_341),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_341),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_267),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_270),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_345),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_345),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_346),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_278),
.Y(n_503)
);

INVx1_ASAP7_75t_SL g504 ( 
.A(n_276),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_346),
.B(n_17),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_362),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_379),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_261),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_362),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_282),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_377),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_377),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_406),
.Y(n_513)
);

INVxp33_ASAP7_75t_SL g514 ( 
.A(n_288),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_404),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_406),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_412),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_412),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_421),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_421),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_426),
.Y(n_521)
);

BUFx6f_ASAP7_75t_SL g522 ( 
.A(n_355),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_293),
.Y(n_523)
);

INVxp33_ASAP7_75t_SL g524 ( 
.A(n_297),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_305),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_426),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_409),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_382),
.B(n_18),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_R g529 ( 
.A(n_246),
.B(n_98),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_409),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_409),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_308),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_313),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_265),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_261),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_261),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_314),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_261),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_265),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_261),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_272),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_318),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_320),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_405),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_321),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_536),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_475),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_475),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_475),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_508),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_438),
.Y(n_551)
);

NAND2xp33_ASAP7_75t_L g552 ( 
.A(n_459),
.B(n_272),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_508),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_461),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_536),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_466),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_538),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_534),
.B(n_347),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_538),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_534),
.B(n_233),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_508),
.Y(n_561)
);

OA21x2_ASAP7_75t_L g562 ( 
.A1(n_540),
.A2(n_541),
.B(n_535),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_439),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_540),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_541),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_527),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_527),
.Y(n_567)
);

NAND2x1_ASAP7_75t_L g568 ( 
.A(n_432),
.B(n_225),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_447),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_530),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_530),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_479),
.Y(n_572)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_447),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_535),
.Y(n_574)
);

BUFx3_ASAP7_75t_L g575 ( 
.A(n_534),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_531),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_531),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_535),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_432),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_480),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_440),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_504),
.A2(n_435),
.B1(n_488),
.B2(n_433),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_442),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_504),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_442),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_443),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_443),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_482),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_435),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_444),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_446),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_448),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_446),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_456),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_458),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_539),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_449),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_437),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_449),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_451),
.Y(n_600)
);

INVxp67_ASAP7_75t_L g601 ( 
.A(n_450),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_451),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_454),
.Y(n_603)
);

INVxp67_ASAP7_75t_SL g604 ( 
.A(n_452),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_452),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_453),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_453),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_462),
.B(n_355),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_529),
.B(n_272),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_539),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_539),
.B(n_272),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_455),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_455),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_464),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_490),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_464),
.Y(n_616)
);

AND2x6_ASAP7_75t_L g617 ( 
.A(n_472),
.B(n_225),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_472),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_478),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_478),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_485),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_485),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_487),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_487),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_465),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_492),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_492),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_496),
.Y(n_628)
);

AND2x2_ASAP7_75t_SL g629 ( 
.A(n_468),
.B(n_225),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_462),
.B(n_355),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_491),
.B(n_355),
.Y(n_631)
);

NOR2xp67_ASAP7_75t_L g632 ( 
.A(n_496),
.B(n_317),
.Y(n_632)
);

AND2x6_ASAP7_75t_L g633 ( 
.A(n_497),
.B(n_226),
.Y(n_633)
);

OA21x2_ASAP7_75t_L g634 ( 
.A1(n_497),
.A2(n_256),
.B(n_226),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_500),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_562),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_625),
.B(n_433),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_626),
.Y(n_638)
);

AND2x4_ASAP7_75t_L g639 ( 
.A(n_604),
.B(n_441),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_604),
.B(n_488),
.Y(n_640)
);

INVx4_ASAP7_75t_L g641 ( 
.A(n_626),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_562),
.Y(n_642)
);

BUFx2_ASAP7_75t_L g643 ( 
.A(n_584),
.Y(n_643)
);

AND2x2_ASAP7_75t_SL g644 ( 
.A(n_629),
.B(n_468),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_562),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_626),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_629),
.B(n_500),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_575),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_608),
.B(n_441),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_562),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_626),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_629),
.B(n_501),
.Y(n_652)
);

AO22x2_ASAP7_75t_L g653 ( 
.A1(n_608),
.A2(n_630),
.B1(n_631),
.B2(n_568),
.Y(n_653)
);

AND3x4_ASAP7_75t_L g654 ( 
.A(n_632),
.B(n_481),
.C(n_470),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_626),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_575),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_551),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_626),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_626),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_563),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_626),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_629),
.B(n_467),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_562),
.Y(n_663)
);

INVx4_ASAP7_75t_L g664 ( 
.A(n_610),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_608),
.B(n_630),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_562),
.Y(n_666)
);

BUFx10_ASAP7_75t_L g667 ( 
.A(n_581),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_560),
.B(n_501),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_630),
.B(n_491),
.Y(n_669)
);

BUFx2_ASAP7_75t_L g670 ( 
.A(n_584),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_549),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_590),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_560),
.B(n_502),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_558),
.B(n_514),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_631),
.A2(n_457),
.B1(n_473),
.B2(n_445),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_549),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_596),
.B(n_558),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_579),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_579),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_596),
.B(n_502),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_579),
.Y(n_681)
);

HB1xp67_ASAP7_75t_L g682 ( 
.A(n_584),
.Y(n_682)
);

BUFx3_ASAP7_75t_L g683 ( 
.A(n_575),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_631),
.B(n_463),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_596),
.B(n_506),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_610),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_596),
.B(n_506),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_579),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_575),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_597),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_597),
.Y(n_691)
);

INVx4_ASAP7_75t_L g692 ( 
.A(n_610),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_597),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_549),
.Y(n_694)
);

OR2x2_ASAP7_75t_L g695 ( 
.A(n_569),
.B(n_434),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_597),
.Y(n_696)
);

INVx6_ASAP7_75t_L g697 ( 
.A(n_611),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_612),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_592),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_612),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_569),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_573),
.B(n_463),
.Y(n_702)
);

AND2x6_ASAP7_75t_L g703 ( 
.A(n_611),
.B(n_612),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_601),
.B(n_524),
.Y(n_704)
);

INVx4_ASAP7_75t_L g705 ( 
.A(n_610),
.Y(n_705)
);

INVxp67_ASAP7_75t_SL g706 ( 
.A(n_573),
.Y(n_706)
);

INVxp67_ASAP7_75t_SL g707 ( 
.A(n_596),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_612),
.Y(n_708)
);

INVx5_ASAP7_75t_L g709 ( 
.A(n_617),
.Y(n_709)
);

INVx1_ASAP7_75t_SL g710 ( 
.A(n_554),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_550),
.Y(n_711)
);

AND2x2_ASAP7_75t_SL g712 ( 
.A(n_552),
.B(n_226),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_583),
.B(n_495),
.Y(n_713)
);

BUFx2_ASAP7_75t_L g714 ( 
.A(n_594),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_601),
.B(n_469),
.Y(n_715)
);

NOR3xp33_ASAP7_75t_L g716 ( 
.A(n_589),
.B(n_457),
.C(n_528),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_583),
.B(n_471),
.Y(n_717)
);

INVx4_ASAP7_75t_L g718 ( 
.A(n_610),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_619),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_595),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_610),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_585),
.B(n_476),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_632),
.B(n_495),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_585),
.B(n_477),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_610),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_619),
.Y(n_726)
);

AND2x4_ASAP7_75t_L g727 ( 
.A(n_586),
.B(n_470),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_586),
.B(n_509),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_619),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_587),
.B(n_509),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_587),
.B(n_511),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_619),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_610),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_621),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_582),
.B(n_483),
.Y(n_735)
);

INVx8_ASAP7_75t_L g736 ( 
.A(n_611),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_554),
.Y(n_737)
);

BUFx3_ASAP7_75t_L g738 ( 
.A(n_611),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_591),
.B(n_511),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_591),
.B(n_486),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_611),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_550),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_593),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_578),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_634),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_568),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_621),
.Y(n_747)
);

HB1xp67_ASAP7_75t_L g748 ( 
.A(n_589),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_621),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_593),
.B(n_481),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_621),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_550),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_623),
.Y(n_753)
);

INVx3_ASAP7_75t_L g754 ( 
.A(n_634),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_623),
.Y(n_755)
);

BUFx4f_ASAP7_75t_L g756 ( 
.A(n_617),
.Y(n_756)
);

OAI22xp5_ASAP7_75t_L g757 ( 
.A1(n_582),
.A2(n_505),
.B1(n_459),
.B2(n_337),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_623),
.Y(n_758)
);

OAI22xp5_ASAP7_75t_L g759 ( 
.A1(n_599),
.A2(n_505),
.B1(n_337),
.B2(n_484),
.Y(n_759)
);

INVx4_ASAP7_75t_L g760 ( 
.A(n_634),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_599),
.B(n_600),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_600),
.B(n_512),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_598),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_623),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_602),
.B(n_512),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_602),
.B(n_513),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_578),
.Y(n_767)
);

INVx1_ASAP7_75t_SL g768 ( 
.A(n_556),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_553),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_605),
.B(n_513),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_624),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_634),
.Y(n_772)
);

AND2x4_ASAP7_75t_L g773 ( 
.A(n_605),
.B(n_516),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_553),
.Y(n_774)
);

INVx5_ASAP7_75t_L g775 ( 
.A(n_617),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_607),
.B(n_516),
.Y(n_776)
);

BUFx6f_ASAP7_75t_SL g777 ( 
.A(n_617),
.Y(n_777)
);

INVx1_ASAP7_75t_SL g778 ( 
.A(n_556),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_634),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_607),
.B(n_517),
.Y(n_780)
);

NAND3x1_ASAP7_75t_L g781 ( 
.A(n_613),
.B(n_474),
.C(n_231),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_553),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_624),
.Y(n_783)
);

OR2x6_ASAP7_75t_L g784 ( 
.A(n_568),
.B(n_606),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_578),
.Y(n_785)
);

INVx3_ASAP7_75t_L g786 ( 
.A(n_634),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_613),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_614),
.Y(n_788)
);

INVx1_ASAP7_75t_SL g789 ( 
.A(n_572),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_574),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_644),
.B(n_723),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_644),
.B(n_614),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_671),
.Y(n_793)
);

NAND2xp33_ASAP7_75t_L g794 ( 
.A(n_642),
.B(n_616),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_657),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_671),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_644),
.B(n_616),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_647),
.B(n_620),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_652),
.B(n_620),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_736),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_723),
.B(n_622),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_736),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_743),
.Y(n_803)
);

OAI21xp5_ASAP7_75t_L g804 ( 
.A1(n_745),
.A2(n_552),
.B(n_622),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_736),
.Y(n_805)
);

OR2x2_ASAP7_75t_L g806 ( 
.A(n_643),
.B(n_603),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_743),
.Y(n_807)
);

OR2x2_ASAP7_75t_L g808 ( 
.A(n_643),
.B(n_460),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_723),
.B(n_627),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_677),
.A2(n_707),
.B(n_685),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_723),
.B(n_627),
.Y(n_811)
);

OR2x2_ASAP7_75t_L g812 ( 
.A(n_670),
.B(n_489),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_639),
.B(n_628),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_649),
.B(n_628),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_639),
.B(n_635),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_757),
.A2(n_609),
.B1(n_522),
.B2(n_420),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_639),
.B(n_649),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_743),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_639),
.B(n_635),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_649),
.B(n_665),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_649),
.B(n_606),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_668),
.B(n_606),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_676),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_673),
.B(n_665),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_746),
.B(n_624),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_660),
.Y(n_826)
);

NAND2xp33_ASAP7_75t_L g827 ( 
.A(n_642),
.B(n_624),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_684),
.B(n_618),
.Y(n_828)
);

NOR2xp67_ASAP7_75t_L g829 ( 
.A(n_672),
.B(n_436),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_684),
.B(n_618),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_746),
.B(n_642),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_787),
.Y(n_832)
);

AND2x6_ASAP7_75t_SL g833 ( 
.A(n_704),
.B(n_224),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_R g834 ( 
.A(n_699),
.B(n_572),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_701),
.B(n_493),
.Y(n_835)
);

AND2x6_ASAP7_75t_SL g836 ( 
.A(n_715),
.B(n_231),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_717),
.B(n_618),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_676),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_712),
.A2(n_609),
.B1(n_522),
.B2(n_410),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_712),
.A2(n_522),
.B1(n_517),
.B2(n_519),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_722),
.B(n_494),
.Y(n_841)
);

OAI221xp5_ASAP7_75t_L g842 ( 
.A1(n_675),
.A2(n_239),
.B1(n_375),
.B2(n_365),
.C(n_363),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_787),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_SL g844 ( 
.A1(n_710),
.A2(n_515),
.B1(n_544),
.B2(n_507),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_701),
.B(n_498),
.Y(n_845)
);

OR2x6_ASAP7_75t_L g846 ( 
.A(n_736),
.B(n_566),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_642),
.B(n_499),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_680),
.A2(n_567),
.B(n_566),
.Y(n_848)
);

OAI22xp5_ASAP7_75t_L g849 ( 
.A1(n_662),
.A2(n_328),
.B1(n_335),
.B2(n_327),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_640),
.B(n_503),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_724),
.B(n_510),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_740),
.B(n_525),
.Y(n_852)
);

O2A1O1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_759),
.A2(n_570),
.B(n_571),
.C(n_567),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_712),
.A2(n_522),
.B1(n_519),
.B2(n_520),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_670),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_674),
.B(n_532),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_642),
.B(n_533),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_787),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_788),
.Y(n_859)
);

A2O1A1Ixp33_ASAP7_75t_SL g860 ( 
.A1(n_716),
.A2(n_571),
.B(n_576),
.C(n_570),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_706),
.B(n_537),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_762),
.B(n_542),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_762),
.B(n_543),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_735),
.B(n_545),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_653),
.A2(n_304),
.B1(n_617),
.B2(n_633),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_788),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_788),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_682),
.B(n_523),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_762),
.B(n_576),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_654),
.A2(n_520),
.B1(n_521),
.B2(n_518),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_694),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_738),
.B(n_518),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_694),
.Y(n_873)
);

INVx8_ASAP7_75t_L g874 ( 
.A(n_736),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_654),
.A2(n_526),
.B1(n_521),
.B2(n_617),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_653),
.A2(n_304),
.B1(n_633),
.B2(n_617),
.Y(n_876)
);

AOI22xp5_ASAP7_75t_L g877 ( 
.A1(n_653),
.A2(n_617),
.B1(n_633),
.B2(n_526),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_762),
.B(n_577),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_761),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_738),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_748),
.B(n_580),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_770),
.B(n_577),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_642),
.B(n_256),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_770),
.B(n_617),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_650),
.B(n_256),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_687),
.A2(n_555),
.B(n_546),
.Y(n_886)
);

INVx1_ASAP7_75t_SL g887 ( 
.A(n_737),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_770),
.B(n_617),
.Y(n_888)
);

AOI221xp5_ASAP7_75t_L g889 ( 
.A1(n_702),
.A2(n_669),
.B1(n_653),
.B2(n_258),
.C(n_262),
.Y(n_889)
);

NAND2xp33_ASAP7_75t_L g890 ( 
.A(n_650),
.B(n_663),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_770),
.B(n_633),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_650),
.B(n_309),
.Y(n_892)
);

BUFx2_ASAP7_75t_L g893 ( 
.A(n_763),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_773),
.B(n_633),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_773),
.B(n_633),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_637),
.B(n_580),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_713),
.A2(n_340),
.B1(n_343),
.B2(n_338),
.Y(n_897)
);

AND2x6_ASAP7_75t_SL g898 ( 
.A(n_720),
.B(n_236),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_702),
.B(n_588),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_695),
.B(n_588),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_761),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_711),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_738),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_711),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_650),
.B(n_309),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_695),
.B(n_669),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_742),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_773),
.B(n_713),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_697),
.B(n_615),
.Y(n_909)
);

INVx5_ASAP7_75t_L g910 ( 
.A(n_650),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_742),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_650),
.B(n_663),
.Y(n_912)
);

OR2x6_ASAP7_75t_L g913 ( 
.A(n_784),
.B(n_350),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_768),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_654),
.A2(n_727),
.B1(n_750),
.B2(n_703),
.Y(n_915)
);

NOR3xp33_ASAP7_75t_L g916 ( 
.A(n_714),
.B(n_254),
.C(n_236),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_741),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_663),
.B(n_309),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_773),
.B(n_633),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_727),
.A2(n_633),
.B1(n_350),
.B2(n_221),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_727),
.B(n_633),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_727),
.A2(n_633),
.B1(n_227),
.B2(n_228),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_741),
.Y(n_923)
);

AND2x6_ASAP7_75t_SL g924 ( 
.A(n_714),
.B(n_254),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_741),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_663),
.B(n_326),
.Y(n_926)
);

OR2x6_ASAP7_75t_L g927 ( 
.A(n_784),
.B(n_258),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_663),
.B(n_326),
.Y(n_928)
);

AOI22xp33_ASAP7_75t_L g929 ( 
.A1(n_750),
.A2(n_393),
.B1(n_428),
.B2(n_424),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_750),
.B(n_262),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_752),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_697),
.B(n_615),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_SL g933 ( 
.A(n_667),
.B(n_393),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_663),
.B(n_326),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_752),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_750),
.B(n_546),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_728),
.B(n_555),
.Y(n_937)
);

NOR2x2_ASAP7_75t_L g938 ( 
.A(n_784),
.B(n_393),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_697),
.B(n_349),
.Y(n_939)
);

INVx2_ASAP7_75t_SL g940 ( 
.A(n_697),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_728),
.B(n_557),
.Y(n_941)
);

BUFx3_ASAP7_75t_L g942 ( 
.A(n_703),
.Y(n_942)
);

AOI22xp33_ASAP7_75t_L g943 ( 
.A1(n_636),
.A2(n_428),
.B1(n_424),
.B2(n_393),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_667),
.B(n_354),
.Y(n_944)
);

AOI22xp33_ASAP7_75t_L g945 ( 
.A1(n_636),
.A2(n_428),
.B1(n_424),
.B2(n_565),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_739),
.B(n_557),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_739),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_730),
.B(n_559),
.Y(n_948)
);

NAND2x1p5_ASAP7_75t_L g949 ( 
.A(n_756),
.B(n_547),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_667),
.B(n_356),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_667),
.B(n_358),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_778),
.B(n_359),
.Y(n_952)
);

AOI22xp33_ASAP7_75t_L g953 ( 
.A1(n_645),
.A2(n_428),
.B1(n_424),
.B2(n_565),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_760),
.B(n_398),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_789),
.B(n_361),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_760),
.B(n_366),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_769),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_678),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_731),
.B(n_559),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_760),
.B(n_398),
.Y(n_960)
);

O2A1O1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_765),
.A2(n_416),
.B(n_298),
.C(n_296),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_769),
.Y(n_962)
);

NAND2xp33_ASAP7_75t_SL g963 ( 
.A(n_805),
.B(n_800),
.Y(n_963)
);

AND2x6_ASAP7_75t_SL g964 ( 
.A(n_881),
.B(n_283),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_855),
.Y(n_965)
);

BUFx4_ASAP7_75t_SL g966 ( 
.A(n_795),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_793),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_846),
.B(n_703),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_793),
.Y(n_969)
);

OR2x4_ASAP7_75t_L g970 ( 
.A(n_856),
.B(n_766),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_850),
.B(n_776),
.Y(n_971)
);

INVx2_ASAP7_75t_SL g972 ( 
.A(n_874),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_872),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_914),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_872),
.Y(n_975)
);

HB1xp67_ASAP7_75t_L g976 ( 
.A(n_887),
.Y(n_976)
);

BUFx3_ASAP7_75t_L g977 ( 
.A(n_795),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_846),
.B(n_703),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_800),
.Y(n_979)
);

AOI22xp5_ASAP7_75t_L g980 ( 
.A1(n_791),
.A2(n_703),
.B1(n_781),
.B2(n_784),
.Y(n_980)
);

BUFx2_ASAP7_75t_L g981 ( 
.A(n_834),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_841),
.B(n_760),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_846),
.B(n_703),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_826),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_872),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_817),
.B(n_780),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_879),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_796),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_800),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_796),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_901),
.Y(n_991)
);

AND2x6_ASAP7_75t_L g992 ( 
.A(n_942),
.B(n_645),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_823),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_846),
.B(n_703),
.Y(n_994)
);

BUFx4f_ASAP7_75t_L g995 ( 
.A(n_874),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_L g996 ( 
.A1(n_861),
.A2(n_781),
.B1(n_784),
.B2(n_754),
.Y(n_996)
);

INVx6_ASAP7_75t_L g997 ( 
.A(n_800),
.Y(n_997)
);

INVxp67_ASAP7_75t_L g998 ( 
.A(n_806),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_823),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_958),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_851),
.B(n_678),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_838),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_852),
.B(n_824),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_802),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_927),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_947),
.Y(n_1006)
);

INVx1_ASAP7_75t_SL g1007 ( 
.A(n_808),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_942),
.B(n_648),
.Y(n_1008)
);

AOI211xp5_ASAP7_75t_L g1009 ( 
.A1(n_845),
.A2(n_287),
.B(n_289),
.C(n_283),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_900),
.B(n_648),
.Y(n_1010)
);

INVx1_ASAP7_75t_SL g1011 ( 
.A(n_812),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_903),
.Y(n_1012)
);

BUFx8_ASAP7_75t_L g1013 ( 
.A(n_893),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_908),
.B(n_820),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_917),
.Y(n_1015)
);

AOI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_889),
.A2(n_666),
.B1(n_754),
.B2(n_745),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_820),
.B(n_679),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_910),
.B(n_641),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_870),
.A2(n_875),
.B1(n_792),
.B2(n_797),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_906),
.B(n_679),
.Y(n_1020)
);

INVx3_ASAP7_75t_L g1021 ( 
.A(n_802),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_802),
.B(n_648),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_835),
.B(n_656),
.Y(n_1023)
);

BUFx2_ASAP7_75t_L g1024 ( 
.A(n_927),
.Y(n_1024)
);

INVx5_ASAP7_75t_L g1025 ( 
.A(n_874),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_814),
.B(n_681),
.Y(n_1026)
);

INVxp67_ASAP7_75t_SL g1027 ( 
.A(n_890),
.Y(n_1027)
);

BUFx6f_ASAP7_75t_L g1028 ( 
.A(n_802),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_923),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_838),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_910),
.B(n_641),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_927),
.B(n_681),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_954),
.A2(n_754),
.B(n_745),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_925),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_821),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_937),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_941),
.Y(n_1037)
);

NAND2xp33_ASAP7_75t_SL g1038 ( 
.A(n_805),
.B(n_688),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_871),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_909),
.B(n_656),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_927),
.B(n_656),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_899),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_910),
.B(n_641),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_946),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_814),
.B(n_688),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_828),
.B(n_690),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_R g1047 ( 
.A(n_826),
.B(n_777),
.Y(n_1047)
);

OAI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_954),
.A2(n_754),
.B(n_745),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_813),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_815),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_874),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_819),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_871),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_830),
.Y(n_1054)
);

AND2x4_ASAP7_75t_L g1055 ( 
.A(n_915),
.B(n_683),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_801),
.Y(n_1056)
);

AOI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_862),
.A2(n_863),
.B1(n_864),
.B2(n_913),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_837),
.B(n_690),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_880),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_930),
.B(n_691),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_R g1061 ( 
.A(n_933),
.B(n_777),
.Y(n_1061)
);

BUFx12f_ASAP7_75t_L g1062 ( 
.A(n_898),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_R g1063 ( 
.A(n_932),
.B(n_777),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_873),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_880),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_809),
.B(n_691),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_880),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_811),
.B(n_693),
.Y(n_1068)
);

O2A1O1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_860),
.A2(n_696),
.B(n_698),
.C(n_693),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_873),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_913),
.B(n_683),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_869),
.Y(n_1072)
);

NOR3xp33_ASAP7_75t_SL g1073 ( 
.A(n_944),
.B(n_370),
.C(n_368),
.Y(n_1073)
);

BUFx2_ASAP7_75t_L g1074 ( 
.A(n_913),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_878),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_882),
.Y(n_1076)
);

INVx2_ASAP7_75t_SL g1077 ( 
.A(n_913),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_R g1078 ( 
.A(n_950),
.B(n_777),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_902),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_880),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_902),
.Y(n_1081)
);

BUFx4f_ASAP7_75t_L g1082 ( 
.A(n_940),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_930),
.B(n_696),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_930),
.B(n_698),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_L g1085 ( 
.A1(n_842),
.A2(n_666),
.B1(n_779),
.B2(n_772),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_951),
.B(n_700),
.Y(n_1086)
);

AND2x4_ASAP7_75t_L g1087 ( 
.A(n_940),
.B(n_683),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_904),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_R g1089 ( 
.A(n_896),
.B(n_772),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_949),
.Y(n_1090)
);

AOI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_939),
.A2(n_890),
.B1(n_956),
.B2(n_839),
.Y(n_1091)
);

INVx2_ASAP7_75t_SL g1092 ( 
.A(n_910),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_910),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_844),
.Y(n_1094)
);

INVx1_ASAP7_75t_SL g1095 ( 
.A(n_938),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_822),
.B(n_700),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_884),
.B(n_689),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_816),
.B(n_708),
.Y(n_1098)
);

NOR3xp33_ASAP7_75t_SL g1099 ( 
.A(n_868),
.B(n_373),
.C(n_372),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_877),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_949),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_904),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_907),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_R g1104 ( 
.A(n_794),
.B(n_772),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_803),
.Y(n_1105)
);

INVx3_ASAP7_75t_L g1106 ( 
.A(n_807),
.Y(n_1106)
);

BUFx2_ASAP7_75t_L g1107 ( 
.A(n_888),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_798),
.B(n_708),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_912),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_952),
.B(n_689),
.Y(n_1110)
);

INVx3_ASAP7_75t_L g1111 ( 
.A(n_818),
.Y(n_1111)
);

BUFx3_ASAP7_75t_L g1112 ( 
.A(n_832),
.Y(n_1112)
);

NOR3xp33_ASAP7_75t_SL g1113 ( 
.A(n_849),
.B(n_380),
.C(n_378),
.Y(n_1113)
);

HB1xp67_ASAP7_75t_L g1114 ( 
.A(n_829),
.Y(n_1114)
);

BUFx2_ASAP7_75t_L g1115 ( 
.A(n_891),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_R g1116 ( 
.A(n_794),
.B(n_924),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_798),
.B(n_719),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_907),
.Y(n_1118)
);

BUFx8_ASAP7_75t_L g1119 ( 
.A(n_843),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_912),
.Y(n_1120)
);

O2A1O1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_860),
.A2(n_726),
.B(n_729),
.C(n_719),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_911),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_911),
.Y(n_1123)
);

INVx5_ASAP7_75t_L g1124 ( 
.A(n_931),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_931),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_916),
.B(n_865),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_876),
.B(n_726),
.Y(n_1127)
);

AND2x6_ASAP7_75t_SL g1128 ( 
.A(n_955),
.B(n_287),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_799),
.B(n_729),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_831),
.B(n_689),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_R g1131 ( 
.A(n_827),
.B(n_772),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_858),
.Y(n_1132)
);

INVx3_ASAP7_75t_L g1133 ( 
.A(n_859),
.Y(n_1133)
);

OAI221xp5_ASAP7_75t_L g1134 ( 
.A1(n_929),
.A2(n_418),
.B1(n_383),
.B2(n_384),
.C(n_385),
.Y(n_1134)
);

BUFx2_ASAP7_75t_L g1135 ( 
.A(n_894),
.Y(n_1135)
);

INVx5_ASAP7_75t_L g1136 ( 
.A(n_935),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_935),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_957),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_957),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_962),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_R g1141 ( 
.A(n_827),
.B(n_779),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_799),
.B(n_732),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_962),
.Y(n_1143)
);

AOI21xp33_ASAP7_75t_L g1144 ( 
.A1(n_921),
.A2(n_734),
.B(n_732),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_936),
.Y(n_1145)
);

INVx3_ASAP7_75t_L g1146 ( 
.A(n_866),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_867),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_948),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_959),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_895),
.B(n_779),
.Y(n_1150)
);

NOR3xp33_ASAP7_75t_SL g1151 ( 
.A(n_897),
.B(n_397),
.C(n_388),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_825),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_919),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_833),
.Y(n_1154)
);

INVx3_ASAP7_75t_L g1155 ( 
.A(n_836),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_840),
.B(n_734),
.Y(n_1156)
);

OA21x2_ASAP7_75t_L g1157 ( 
.A1(n_1091),
.A2(n_857),
.B(n_847),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1033),
.A2(n_1048),
.B(n_1069),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1006),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_974),
.Y(n_1160)
);

AO31x2_ASAP7_75t_L g1161 ( 
.A1(n_982),
.A2(n_848),
.A3(n_810),
.B(n_886),
.Y(n_1161)
);

AOI211x1_ASAP7_75t_L g1162 ( 
.A1(n_1003),
.A2(n_804),
.B(n_825),
.C(n_290),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_987),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1042),
.B(n_943),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_967),
.Y(n_1165)
);

OAI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_971),
.A2(n_854),
.B1(n_920),
.B2(n_922),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_991),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1014),
.A2(n_1148),
.B1(n_1149),
.B2(n_996),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_1121),
.A2(n_885),
.B(n_883),
.Y(n_1169)
);

OR2x6_ASAP7_75t_L g1170 ( 
.A(n_968),
.B(n_831),
.Y(n_1170)
);

O2A1O1Ixp5_ASAP7_75t_L g1171 ( 
.A1(n_1086),
.A2(n_857),
.B(n_847),
.C(n_960),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1000),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_1057),
.B(n_960),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1020),
.B(n_945),
.Y(n_1174)
);

OR2x2_ASAP7_75t_L g1175 ( 
.A(n_1007),
.B(n_747),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1027),
.A2(n_885),
.B(n_883),
.Y(n_1176)
);

AO31x2_ASAP7_75t_L g1177 ( 
.A1(n_1130),
.A2(n_749),
.A3(n_751),
.B(n_747),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1096),
.A2(n_905),
.B(n_892),
.Y(n_1178)
);

O2A1O1Ixp5_ASAP7_75t_L g1179 ( 
.A1(n_1038),
.A2(n_905),
.B(n_918),
.C(n_892),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1012),
.Y(n_1180)
);

OAI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1144),
.A2(n_926),
.B(n_918),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1058),
.A2(n_928),
.B(n_926),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1015),
.Y(n_1183)
);

NAND2x1p5_ASAP7_75t_L g1184 ( 
.A(n_968),
.B(n_756),
.Y(n_1184)
);

INVx2_ASAP7_75t_SL g1185 ( 
.A(n_1013),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1020),
.B(n_953),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1109),
.B(n_744),
.Y(n_1187)
);

O2A1O1Ixp5_ASAP7_75t_L g1188 ( 
.A1(n_1038),
.A2(n_934),
.B(n_928),
.C(n_751),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_1093),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_1109),
.B(n_744),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1156),
.A2(n_934),
.B(n_1108),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1017),
.A2(n_786),
.B(n_779),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1001),
.A2(n_786),
.B(n_692),
.Y(n_1193)
);

OR2x2_ASAP7_75t_L g1194 ( 
.A(n_1011),
.B(n_749),
.Y(n_1194)
);

BUFx3_ASAP7_75t_L g1195 ( 
.A(n_1013),
.Y(n_1195)
);

AO21x1_ASAP7_75t_L g1196 ( 
.A1(n_1009),
.A2(n_853),
.B(n_755),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_998),
.B(n_641),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1046),
.A2(n_786),
.B(n_692),
.Y(n_1198)
);

NAND2x1p5_ASAP7_75t_L g1199 ( 
.A(n_968),
.B(n_756),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_1013),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1110),
.A2(n_1068),
.B(n_1066),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1029),
.Y(n_1202)
);

NAND3xp33_ASAP7_75t_SL g1203 ( 
.A(n_1010),
.B(n_961),
.C(n_400),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1036),
.B(n_753),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_995),
.Y(n_1205)
);

A2O1A1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1126),
.A2(n_755),
.B(n_758),
.C(n_753),
.Y(n_1206)
);

NAND3x1_ASAP7_75t_L g1207 ( 
.A(n_1126),
.B(n_938),
.C(n_290),
.Y(n_1207)
);

AOI21xp33_ASAP7_75t_L g1208 ( 
.A1(n_1083),
.A2(n_764),
.B(n_758),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1018),
.A2(n_786),
.B(n_725),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_986),
.A2(n_646),
.B(n_638),
.Y(n_1210)
);

A2O1A1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1037),
.A2(n_764),
.B(n_783),
.C(n_771),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1018),
.A2(n_725),
.B(n_721),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1044),
.B(n_771),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_995),
.A2(n_692),
.B(n_664),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1049),
.B(n_783),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1050),
.B(n_774),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1052),
.B(n_774),
.Y(n_1217)
);

AOI21xp33_ASAP7_75t_L g1218 ( 
.A1(n_1084),
.A2(n_790),
.B(n_782),
.Y(n_1218)
);

OR2x2_ASAP7_75t_L g1219 ( 
.A(n_1042),
.B(n_790),
.Y(n_1219)
);

AO21x1_ASAP7_75t_L g1220 ( 
.A1(n_1040),
.A2(n_1098),
.B(n_1055),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1031),
.A2(n_725),
.B(n_721),
.Y(n_1221)
);

BUFx5_ASAP7_75t_L g1222 ( 
.A(n_992),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1031),
.A2(n_725),
.B(n_721),
.Y(n_1223)
);

AO21x2_ASAP7_75t_L g1224 ( 
.A1(n_1131),
.A2(n_646),
.B(n_638),
.Y(n_1224)
);

O2A1O1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1023),
.A2(n_298),
.B(n_296),
.C(n_299),
.Y(n_1225)
);

NAND3xp33_ASAP7_75t_SL g1226 ( 
.A(n_1113),
.B(n_402),
.C(n_399),
.Y(n_1226)
);

INVx1_ASAP7_75t_SL g1227 ( 
.A(n_976),
.Y(n_1227)
);

NAND2xp33_ASAP7_75t_L g1228 ( 
.A(n_1025),
.B(n_651),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1043),
.A2(n_721),
.B(n_655),
.Y(n_1229)
);

AO31x2_ASAP7_75t_L g1230 ( 
.A1(n_1100),
.A2(n_969),
.A3(n_988),
.B(n_967),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_970),
.B(n_651),
.Y(n_1231)
);

OAI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1150),
.A2(n_658),
.B(n_655),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1043),
.A2(n_659),
.B(n_658),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1117),
.A2(n_1142),
.B(n_1129),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_995),
.A2(n_692),
.B(n_664),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1072),
.B(n_782),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_969),
.A2(n_661),
.B(n_659),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1075),
.B(n_661),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_963),
.A2(n_705),
.B(n_664),
.Y(n_1239)
);

OR2x2_ASAP7_75t_L g1240 ( 
.A(n_965),
.B(n_289),
.Y(n_1240)
);

BUFx2_ASAP7_75t_L g1241 ( 
.A(n_977),
.Y(n_1241)
);

OAI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1150),
.A2(n_705),
.B(n_664),
.Y(n_1242)
);

OR2x2_ASAP7_75t_L g1243 ( 
.A(n_1094),
.B(n_291),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1034),
.Y(n_1244)
);

INVx3_ASAP7_75t_SL g1245 ( 
.A(n_984),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_SL g1246 ( 
.A(n_984),
.B(n_709),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1155),
.B(n_408),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1076),
.B(n_411),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1019),
.A2(n_396),
.B1(n_322),
.B2(n_291),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1056),
.B(n_413),
.Y(n_1250)
);

HB1xp67_ASAP7_75t_L g1251 ( 
.A(n_973),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_988),
.A2(n_564),
.B(n_548),
.Y(n_1252)
);

INVx4_ASAP7_75t_L g1253 ( 
.A(n_1025),
.Y(n_1253)
);

AO31x2_ASAP7_75t_L g1254 ( 
.A1(n_1100),
.A2(n_705),
.A3(n_718),
.B(n_564),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1054),
.B(n_1035),
.Y(n_1255)
);

OAI22x1_ASAP7_75t_L g1256 ( 
.A1(n_1094),
.A2(n_292),
.B1(n_294),
.B2(n_299),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_990),
.A2(n_548),
.B(n_574),
.Y(n_1257)
);

AOI211x1_ASAP7_75t_L g1258 ( 
.A1(n_1060),
.A2(n_292),
.B(n_294),
.C(n_300),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_990),
.A2(n_548),
.B(n_574),
.Y(n_1259)
);

AO32x2_ASAP7_75t_L g1260 ( 
.A1(n_1077),
.A2(n_705),
.A3(n_718),
.B1(n_310),
.B2(n_396),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1147),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1150),
.A2(n_718),
.B(n_733),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_993),
.A2(n_548),
.B(n_547),
.Y(n_1263)
);

NAND3xp33_ASAP7_75t_L g1264 ( 
.A(n_1151),
.B(n_415),
.C(n_414),
.Y(n_1264)
);

OA21x2_ASAP7_75t_L g1265 ( 
.A1(n_993),
.A2(n_398),
.B(n_310),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1145),
.B(n_417),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_999),
.A2(n_561),
.B(n_547),
.Y(n_1267)
);

O2A1O1Ixp5_ASAP7_75t_L g1268 ( 
.A1(n_1105),
.A2(n_718),
.B(n_300),
.C(n_311),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_999),
.A2(n_561),
.B(n_547),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_975),
.B(n_419),
.Y(n_1270)
);

BUFx2_ASAP7_75t_L g1271 ( 
.A(n_977),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1147),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1002),
.Y(n_1273)
);

CKINVDCx20_ASAP7_75t_R g1274 ( 
.A(n_981),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1002),
.A2(n_1039),
.B(n_1030),
.Y(n_1275)
);

AO21x1_ASAP7_75t_L g1276 ( 
.A1(n_1055),
.A2(n_322),
.B(n_311),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_985),
.B(n_1060),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_963),
.A2(n_733),
.B(n_686),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1030),
.A2(n_561),
.B(n_547),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1127),
.B(n_1089),
.Y(n_1280)
);

AO22x2_ASAP7_75t_L g1281 ( 
.A1(n_1077),
.A2(n_407),
.B1(n_323),
.B2(n_342),
.Y(n_1281)
);

OAI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1026),
.A2(n_733),
.B(n_709),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1082),
.A2(n_686),
.B(n_744),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1127),
.B(n_423),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1082),
.A2(n_686),
.B(n_744),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_966),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1079),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1082),
.A2(n_686),
.B(n_744),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1103),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1123),
.Y(n_1290)
);

NAND2x1_ASAP7_75t_L g1291 ( 
.A(n_1051),
.B(n_744),
.Y(n_1291)
);

INVx3_ASAP7_75t_L g1292 ( 
.A(n_1025),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1089),
.B(n_429),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_970),
.B(n_323),
.Y(n_1294)
);

NOR2xp67_ASAP7_75t_L g1295 ( 
.A(n_1114),
.B(n_561),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1039),
.A2(n_561),
.B(n_342),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1005),
.B(n_339),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_SL g1298 ( 
.A(n_1109),
.B(n_767),
.Y(n_1298)
);

INVx2_ASAP7_75t_SL g1299 ( 
.A(n_981),
.Y(n_1299)
);

INVxp67_ASAP7_75t_L g1300 ( 
.A(n_1032),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1005),
.B(n_339),
.Y(n_1301)
);

HB1xp67_ASAP7_75t_L g1302 ( 
.A(n_1032),
.Y(n_1302)
);

O2A1O1Ixp5_ASAP7_75t_L g1303 ( 
.A1(n_1105),
.A2(n_389),
.B(n_344),
.C(n_363),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_SL g1304 ( 
.A1(n_1092),
.A2(n_353),
.B(n_344),
.Y(n_1304)
);

AOI21x1_ASAP7_75t_SL g1305 ( 
.A1(n_1045),
.A2(n_686),
.B(n_767),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1095),
.B(n_1024),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1053),
.A2(n_360),
.B(n_353),
.Y(n_1307)
);

AND2x4_ASAP7_75t_L g1308 ( 
.A(n_978),
.B(n_709),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_SL g1309 ( 
.A1(n_1092),
.A2(n_365),
.B(n_360),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_980),
.A2(n_375),
.B1(n_394),
.B2(n_386),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_978),
.A2(n_427),
.B1(n_389),
.B2(n_401),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1155),
.B(n_386),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1024),
.B(n_1107),
.Y(n_1313)
);

A2O1A1Ixp33_ASAP7_75t_SL g1314 ( 
.A1(n_1105),
.A2(n_422),
.B(n_401),
.C(n_407),
.Y(n_1314)
);

OA21x2_ASAP7_75t_L g1315 ( 
.A1(n_1053),
.A2(n_394),
.B(n_416),
.Y(n_1315)
);

OAI21xp33_ASAP7_75t_L g1316 ( 
.A1(n_1099),
.A2(n_422),
.B(n_427),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1025),
.A2(n_686),
.B(n_767),
.Y(n_1317)
);

INVx3_ASAP7_75t_L g1318 ( 
.A(n_1025),
.Y(n_1318)
);

O2A1O1Ixp33_ASAP7_75t_SL g1319 ( 
.A1(n_1152),
.A2(n_21),
.B(n_24),
.C(n_25),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1107),
.B(n_785),
.Y(n_1320)
);

AOI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1055),
.A2(n_785),
.B1(n_767),
.B2(n_312),
.Y(n_1321)
);

AO31x2_ASAP7_75t_L g1322 ( 
.A1(n_1064),
.A2(n_578),
.A3(n_785),
.B(n_767),
.Y(n_1322)
);

OAI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1085),
.A2(n_709),
.B(n_775),
.Y(n_1323)
);

NAND2xp33_ASAP7_75t_L g1324 ( 
.A(n_1222),
.B(n_1078),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1165),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_SL g1326 ( 
.A(n_1280),
.B(n_1041),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1230),
.Y(n_1327)
);

CKINVDCx14_ASAP7_75t_R g1328 ( 
.A(n_1286),
.Y(n_1328)
);

CKINVDCx16_ASAP7_75t_R g1329 ( 
.A(n_1274),
.Y(n_1329)
);

BUFx8_ASAP7_75t_L g1330 ( 
.A(n_1200),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_1286),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1305),
.A2(n_1070),
.B(n_1064),
.Y(n_1332)
);

AO21x2_ASAP7_75t_L g1333 ( 
.A1(n_1173),
.A2(n_1141),
.B(n_1131),
.Y(n_1333)
);

OAI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1243),
.A2(n_1155),
.B1(n_1154),
.B2(n_1134),
.Y(n_1334)
);

OAI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1284),
.A2(n_1154),
.B1(n_1074),
.B2(n_1128),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1305),
.A2(n_1081),
.B(n_1070),
.Y(n_1336)
);

OA21x2_ASAP7_75t_L g1337 ( 
.A1(n_1171),
.A2(n_1138),
.B(n_1125),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1209),
.A2(n_1088),
.B(n_1081),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1201),
.A2(n_978),
.B1(n_983),
.B2(n_994),
.Y(n_1339)
);

AO32x2_ASAP7_75t_L g1340 ( 
.A1(n_1168),
.A2(n_1074),
.A3(n_1073),
.B1(n_1116),
.B2(n_972),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1165),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1268),
.A2(n_1087),
.B(n_1097),
.Y(n_1342)
);

INVx3_ASAP7_75t_SL g1343 ( 
.A(n_1245),
.Y(n_1343)
);

OAI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1268),
.A2(n_1087),
.B(n_1097),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_1245),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1228),
.A2(n_1093),
.B(n_994),
.Y(n_1346)
);

O2A1O1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1203),
.A2(n_1146),
.B(n_1111),
.C(n_1106),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1169),
.A2(n_1102),
.B(n_1088),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1179),
.A2(n_1087),
.B(n_1097),
.Y(n_1349)
);

NAND2x1p5_ASAP7_75t_L g1350 ( 
.A(n_1189),
.B(n_1093),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1158),
.A2(n_1178),
.B(n_1191),
.Y(n_1351)
);

OAI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1197),
.A2(n_983),
.B1(n_994),
.B2(n_1041),
.Y(n_1352)
);

BUFx2_ASAP7_75t_SL g1353 ( 
.A(n_1274),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1273),
.Y(n_1354)
);

OA21x2_ASAP7_75t_L g1355 ( 
.A1(n_1171),
.A2(n_1140),
.B(n_1139),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1255),
.B(n_1116),
.Y(n_1356)
);

O2A1O1Ixp33_ASAP7_75t_SL g1357 ( 
.A1(n_1206),
.A2(n_972),
.B(n_1051),
.C(n_1021),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1230),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1249),
.A2(n_1153),
.B1(n_1132),
.B2(n_1112),
.Y(n_1359)
);

OR2x6_ASAP7_75t_L g1360 ( 
.A(n_1170),
.B(n_1071),
.Y(n_1360)
);

A2O1A1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1225),
.A2(n_1112),
.B(n_1132),
.C(n_1115),
.Y(n_1361)
);

OA21x2_ASAP7_75t_L g1362 ( 
.A1(n_1191),
.A2(n_1143),
.B(n_1118),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1178),
.A2(n_1118),
.B(n_1102),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1269),
.A2(n_1137),
.B(n_1122),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1269),
.A2(n_1137),
.B(n_1122),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_L g1366 ( 
.A(n_1160),
.B(n_964),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1300),
.B(n_1062),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1230),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1273),
.Y(n_1369)
);

INVx6_ASAP7_75t_L g1370 ( 
.A(n_1308),
.Y(n_1370)
);

AO21x1_ASAP7_75t_L g1371 ( 
.A1(n_1173),
.A2(n_1166),
.B(n_1210),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1227),
.B(n_1119),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1275),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1279),
.A2(n_1111),
.B(n_1106),
.Y(n_1374)
);

NAND2x1p5_ASAP7_75t_L g1375 ( 
.A(n_1189),
.B(n_1093),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1279),
.A2(n_1111),
.B(n_1106),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1230),
.Y(n_1377)
);

INVx8_ASAP7_75t_L g1378 ( 
.A(n_1170),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1261),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1175),
.B(n_1119),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1307),
.A2(n_1146),
.B(n_1133),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1194),
.B(n_1119),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1272),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_SL g1384 ( 
.A1(n_1196),
.A2(n_1016),
.B(n_1104),
.Y(n_1384)
);

INVxp67_ASAP7_75t_L g1385 ( 
.A(n_1241),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1287),
.Y(n_1386)
);

NAND2x1p5_ASAP7_75t_L g1387 ( 
.A(n_1189),
.B(n_1109),
.Y(n_1387)
);

OAI211xp5_ASAP7_75t_L g1388 ( 
.A1(n_1316),
.A2(n_1047),
.B(n_272),
.C(n_1146),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1302),
.Y(n_1389)
);

BUFx12f_ASAP7_75t_L g1390 ( 
.A(n_1185),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1197),
.A2(n_983),
.B1(n_1041),
.B2(n_1133),
.Y(n_1391)
);

AO21x2_ASAP7_75t_L g1392 ( 
.A1(n_1220),
.A2(n_1141),
.B(n_1104),
.Y(n_1392)
);

AO31x2_ASAP7_75t_L g1393 ( 
.A1(n_1206),
.A2(n_1182),
.A3(n_1276),
.B(n_1176),
.Y(n_1393)
);

AO21x2_ASAP7_75t_L g1394 ( 
.A1(n_1181),
.A2(n_1078),
.B(n_1063),
.Y(n_1394)
);

AOI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1157),
.A2(n_1071),
.B(n_1115),
.Y(n_1395)
);

OA21x2_ASAP7_75t_L g1396 ( 
.A1(n_1179),
.A2(n_1135),
.B(n_1071),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1289),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_SL g1398 ( 
.A(n_1195),
.B(n_1062),
.Y(n_1398)
);

OAI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1188),
.A2(n_1133),
.B(n_1135),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1307),
.A2(n_1101),
.B(n_1021),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1302),
.B(n_1047),
.Y(n_1401)
);

AOI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1228),
.A2(n_1120),
.B(n_1124),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1300),
.B(n_1008),
.Y(n_1403)
);

INVx3_ASAP7_75t_L g1404 ( 
.A(n_1253),
.Y(n_1404)
);

OAI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1188),
.A2(n_1303),
.B(n_1293),
.Y(n_1405)
);

OAI221xp5_ASAP7_75t_L g1406 ( 
.A1(n_1294),
.A2(n_1101),
.B1(n_1153),
.B2(n_1090),
.C(n_1021),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1277),
.B(n_1008),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1170),
.B(n_1153),
.Y(n_1408)
);

INVxp67_ASAP7_75t_L g1409 ( 
.A(n_1271),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1290),
.Y(n_1410)
);

CKINVDCx20_ASAP7_75t_R g1411 ( 
.A(n_1195),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1164),
.B(n_1153),
.Y(n_1412)
);

AND2x4_ASAP7_75t_L g1413 ( 
.A(n_1308),
.B(n_1008),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1251),
.B(n_1059),
.Y(n_1414)
);

NAND3xp33_ASAP7_75t_SL g1415 ( 
.A(n_1247),
.B(n_1061),
.C(n_229),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1315),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1315),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1281),
.A2(n_992),
.B1(n_1063),
.B2(n_1061),
.Y(n_1418)
);

BUFx3_ASAP7_75t_L g1419 ( 
.A(n_1299),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1308),
.B(n_1090),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_SL g1421 ( 
.A1(n_1232),
.A2(n_1120),
.B(n_992),
.Y(n_1421)
);

INVx1_ASAP7_75t_SL g1422 ( 
.A(n_1306),
.Y(n_1422)
);

AOI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1207),
.A2(n_992),
.B1(n_1022),
.B2(n_1101),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1315),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_1256),
.Y(n_1425)
);

CKINVDCx6p67_ASAP7_75t_R g1426 ( 
.A(n_1312),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1237),
.A2(n_1051),
.B(n_1120),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1322),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1313),
.B(n_1059),
.Y(n_1429)
);

CKINVDCx11_ASAP7_75t_R g1430 ( 
.A(n_1189),
.Y(n_1430)
);

INVx3_ASAP7_75t_L g1431 ( 
.A(n_1253),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1212),
.A2(n_1120),
.B(n_992),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1177),
.Y(n_1433)
);

OA21x2_ASAP7_75t_L g1434 ( 
.A1(n_1296),
.A2(n_1234),
.B(n_1263),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1221),
.A2(n_992),
.B(n_1124),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1322),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1251),
.B(n_1059),
.Y(n_1437)
);

OAI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1303),
.A2(n_1022),
.B(n_1124),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1223),
.A2(n_1124),
.B(n_1136),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1322),
.Y(n_1440)
);

BUFx2_ASAP7_75t_L g1441 ( 
.A(n_1224),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1219),
.Y(n_1442)
);

INVx2_ASAP7_75t_SL g1443 ( 
.A(n_1205),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1172),
.B(n_1059),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1322),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1252),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1267),
.A2(n_1136),
.B(n_1124),
.Y(n_1447)
);

CKINVDCx20_ASAP7_75t_R g1448 ( 
.A(n_1240),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1233),
.A2(n_1136),
.B(n_1080),
.Y(n_1449)
);

AOI221xp5_ASAP7_75t_L g1450 ( 
.A1(n_1310),
.A2(n_272),
.B1(n_1022),
.B2(n_265),
.C(n_1065),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1177),
.Y(n_1451)
);

OA21x2_ASAP7_75t_L g1452 ( 
.A1(n_1211),
.A2(n_364),
.B(n_234),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1177),
.B(n_1065),
.Y(n_1453)
);

NAND2x1p5_ASAP7_75t_L g1454 ( 
.A(n_1187),
.B(n_1136),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1226),
.B(n_1065),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1159),
.B(n_1065),
.Y(n_1456)
);

INVx4_ASAP7_75t_L g1457 ( 
.A(n_1205),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1163),
.B(n_1067),
.Y(n_1458)
);

BUFx3_ASAP7_75t_L g1459 ( 
.A(n_1184),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1281),
.A2(n_1136),
.B1(n_1080),
.B2(n_1067),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1281),
.A2(n_1080),
.B1(n_1067),
.B2(n_997),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1257),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1259),
.Y(n_1463)
);

AND2x4_ASAP7_75t_L g1464 ( 
.A(n_1292),
.B(n_1067),
.Y(n_1464)
);

AO21x2_ASAP7_75t_L g1465 ( 
.A1(n_1224),
.A2(n_1080),
.B(n_785),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_1184),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1177),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1229),
.A2(n_1193),
.B(n_1198),
.Y(n_1468)
);

AND2x4_ASAP7_75t_L g1469 ( 
.A(n_1292),
.B(n_979),
.Y(n_1469)
);

CKINVDCx6p67_ASAP7_75t_R g1470 ( 
.A(n_1297),
.Y(n_1470)
);

OA21x2_ASAP7_75t_L g1471 ( 
.A1(n_1211),
.A2(n_220),
.B(n_235),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1167),
.B(n_979),
.Y(n_1472)
);

AOI21x1_ASAP7_75t_L g1473 ( 
.A1(n_1157),
.A2(n_785),
.B(n_767),
.Y(n_1473)
);

NAND3xp33_ASAP7_75t_L g1474 ( 
.A(n_1162),
.B(n_1028),
.C(n_1004),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1180),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1278),
.A2(n_785),
.B(n_997),
.Y(n_1476)
);

INVx2_ASAP7_75t_SL g1477 ( 
.A(n_1318),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1203),
.A2(n_997),
.B1(n_1004),
.B2(n_1028),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1183),
.Y(n_1479)
);

OAI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1248),
.A2(n_997),
.B1(n_1004),
.B2(n_1028),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1202),
.Y(n_1481)
);

INVx4_ASAP7_75t_L g1482 ( 
.A(n_1199),
.Y(n_1482)
);

OA21x2_ASAP7_75t_L g1483 ( 
.A1(n_1218),
.A2(n_242),
.B(n_243),
.Y(n_1483)
);

AOI221xp5_ASAP7_75t_L g1484 ( 
.A1(n_1311),
.A2(n_348),
.B1(n_249),
.B2(n_255),
.C(n_269),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1226),
.B(n_979),
.Y(n_1485)
);

AOI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1207),
.A2(n_1004),
.B1(n_989),
.B2(n_979),
.Y(n_1486)
);

AND2x4_ASAP7_75t_L g1487 ( 
.A(n_1318),
.B(n_989),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1244),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1265),
.Y(n_1489)
);

AND2x4_ASAP7_75t_L g1490 ( 
.A(n_1295),
.B(n_989),
.Y(n_1490)
);

OAI21x1_ASAP7_75t_L g1491 ( 
.A1(n_1187),
.A2(n_1028),
.B(n_989),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1265),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1301),
.B(n_578),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1265),
.Y(n_1494)
);

BUFx6f_ASAP7_75t_L g1495 ( 
.A(n_1199),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1320),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1216),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1254),
.Y(n_1498)
);

NAND2x1p5_ASAP7_75t_L g1499 ( 
.A(n_1190),
.B(n_709),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1217),
.Y(n_1500)
);

OA21x2_ASAP7_75t_L g1501 ( 
.A1(n_1282),
.A2(n_245),
.B(n_271),
.Y(n_1501)
);

INVx4_ASAP7_75t_L g1502 ( 
.A(n_1222),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_L g1503 ( 
.A1(n_1448),
.A2(n_1186),
.B1(n_1174),
.B2(n_1231),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1426),
.B(n_1412),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1442),
.B(n_1254),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1448),
.A2(n_1231),
.B1(n_1157),
.B2(n_1266),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1408),
.B(n_1190),
.Y(n_1507)
);

OAI211xp5_ASAP7_75t_L g1508 ( 
.A1(n_1356),
.A2(n_1319),
.B(n_1264),
.C(n_1250),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1470),
.A2(n_1321),
.B1(n_1204),
.B2(n_1213),
.Y(n_1509)
);

INVx4_ASAP7_75t_L g1510 ( 
.A(n_1430),
.Y(n_1510)
);

AOI221xp5_ASAP7_75t_L g1511 ( 
.A1(n_1334),
.A2(n_1319),
.B1(n_1258),
.B2(n_1270),
.C(n_1314),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_1331),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1389),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1470),
.B(n_1215),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1385),
.A2(n_1238),
.B1(n_1298),
.B2(n_1192),
.Y(n_1515)
);

OR2x6_ASAP7_75t_L g1516 ( 
.A(n_1378),
.B(n_1298),
.Y(n_1516)
);

AND2x4_ASAP7_75t_L g1517 ( 
.A(n_1408),
.B(n_1254),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1425),
.A2(n_1208),
.B1(n_1236),
.B2(n_1309),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1425),
.A2(n_1335),
.B1(n_1426),
.B2(n_1371),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1412),
.B(n_21),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1325),
.Y(n_1521)
);

OAI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1409),
.A2(n_1242),
.B1(n_1235),
.B2(n_1214),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1422),
.B(n_1475),
.Y(n_1523)
);

INVxp67_ASAP7_75t_L g1524 ( 
.A(n_1353),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1419),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1475),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1479),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_1331),
.Y(n_1528)
);

OAI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1391),
.A2(n_1352),
.B1(n_1361),
.B2(n_1418),
.Y(n_1529)
);

OAI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1366),
.A2(n_1246),
.B1(n_1262),
.B2(n_1323),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_SL g1531 ( 
.A1(n_1384),
.A2(n_1222),
.B1(n_1304),
.B2(n_1260),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1341),
.Y(n_1532)
);

OAI221xp5_ASAP7_75t_L g1533 ( 
.A1(n_1405),
.A2(n_1314),
.B1(n_1288),
.B2(n_1285),
.C(n_1283),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1479),
.B(n_1254),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_SL g1535 ( 
.A1(n_1384),
.A2(n_1222),
.B1(n_1260),
.B2(n_336),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_SL g1536 ( 
.A1(n_1333),
.A2(n_1222),
.B1(n_1260),
.B2(n_336),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1481),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1371),
.A2(n_1222),
.B1(n_578),
.B2(n_336),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1341),
.Y(n_1539)
);

INVx2_ASAP7_75t_SL g1540 ( 
.A(n_1330),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1354),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1481),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1353),
.B(n_26),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1326),
.A2(n_578),
.B1(n_336),
.B2(n_1260),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1360),
.B(n_1291),
.Y(n_1545)
);

AOI221xp5_ASAP7_75t_L g1546 ( 
.A1(n_1484),
.A2(n_369),
.B1(n_275),
.B2(n_280),
.C(n_281),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1339),
.A2(n_1239),
.B1(n_1317),
.B2(n_374),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1389),
.B(n_26),
.Y(n_1548)
);

O2A1O1Ixp33_ASAP7_75t_L g1549 ( 
.A1(n_1357),
.A2(n_1161),
.B(n_28),
.C(n_30),
.Y(n_1549)
);

BUFx6f_ASAP7_75t_L g1550 ( 
.A(n_1413),
.Y(n_1550)
);

BUFx3_ASAP7_75t_L g1551 ( 
.A(n_1419),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1354),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_1328),
.Y(n_1553)
);

AOI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1380),
.A2(n_371),
.B1(n_285),
.B2(n_286),
.Y(n_1554)
);

OAI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1359),
.A2(n_387),
.B1(n_295),
.B2(n_302),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1369),
.Y(n_1556)
);

AO21x2_ASAP7_75t_L g1557 ( 
.A1(n_1416),
.A2(n_1161),
.B(n_775),
.Y(n_1557)
);

INVx1_ASAP7_75t_SL g1558 ( 
.A(n_1329),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1488),
.Y(n_1559)
);

NOR3xp33_ASAP7_75t_SL g1560 ( 
.A(n_1345),
.B(n_274),
.C(n_307),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1360),
.B(n_1161),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1367),
.B(n_27),
.Y(n_1562)
);

INVx4_ASAP7_75t_L g1563 ( 
.A(n_1457),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_1345),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1456),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1456),
.Y(n_1566)
);

OAI21x1_ASAP7_75t_L g1567 ( 
.A1(n_1473),
.A2(n_1161),
.B(n_578),
.Y(n_1567)
);

OAI22xp33_ASAP7_75t_L g1568 ( 
.A1(n_1382),
.A2(n_391),
.B1(n_332),
.B2(n_431),
.Y(n_1568)
);

OAI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1398),
.A2(n_390),
.B1(n_334),
.B2(n_425),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1488),
.B(n_33),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1386),
.B(n_33),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_SL g1572 ( 
.A1(n_1333),
.A2(n_336),
.B1(n_395),
.B2(n_392),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1360),
.B(n_99),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_SL g1574 ( 
.A1(n_1333),
.A2(n_336),
.B1(n_367),
.B2(n_330),
.Y(n_1574)
);

NAND3xp33_ASAP7_75t_SL g1575 ( 
.A(n_1411),
.B(n_35),
.C(n_37),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1386),
.B(n_35),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1360),
.B(n_102),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1413),
.B(n_37),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_1390),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1414),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1397),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1407),
.B(n_38),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1413),
.B(n_1472),
.Y(n_1583)
);

BUFx4f_ASAP7_75t_SL g1584 ( 
.A(n_1411),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_SL g1585 ( 
.A1(n_1392),
.A2(n_775),
.B1(n_709),
.B2(n_47),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1397),
.Y(n_1586)
);

NAND3xp33_ASAP7_75t_SL g1587 ( 
.A(n_1372),
.B(n_1485),
.C(n_1455),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1472),
.B(n_1414),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1450),
.A2(n_775),
.B1(n_41),
.B2(n_47),
.Y(n_1589)
);

OAI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1423),
.A2(n_775),
.B1(n_48),
.B2(n_49),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1437),
.B(n_40),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1410),
.Y(n_1592)
);

BUFx3_ASAP7_75t_L g1593 ( 
.A(n_1330),
.Y(n_1593)
);

CKINVDCx6p67_ASAP7_75t_R g1594 ( 
.A(n_1343),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1437),
.B(n_40),
.Y(n_1595)
);

INVx4_ASAP7_75t_L g1596 ( 
.A(n_1457),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1343),
.B(n_48),
.Y(n_1597)
);

OAI21xp33_ASAP7_75t_L g1598 ( 
.A1(n_1478),
.A2(n_50),
.B(n_51),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1410),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1383),
.B(n_52),
.Y(n_1600)
);

O2A1O1Ixp33_ASAP7_75t_SL g1601 ( 
.A1(n_1347),
.A2(n_52),
.B(n_53),
.C(n_55),
.Y(n_1601)
);

O2A1O1Ixp33_ASAP7_75t_L g1602 ( 
.A1(n_1388),
.A2(n_55),
.B(n_56),
.C(n_57),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_L g1603 ( 
.A(n_1403),
.B(n_56),
.Y(n_1603)
);

A2O1A1Ixp33_ASAP7_75t_L g1604 ( 
.A1(n_1349),
.A2(n_775),
.B(n_61),
.C(n_62),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1392),
.A2(n_58),
.B1(n_62),
.B2(n_63),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1362),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1383),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1379),
.Y(n_1608)
);

CKINVDCx9p33_ASAP7_75t_R g1609 ( 
.A(n_1401),
.Y(n_1609)
);

OAI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1474),
.A2(n_64),
.B1(n_65),
.B2(n_68),
.Y(n_1610)
);

OAI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1486),
.A2(n_64),
.B1(n_68),
.B2(n_71),
.Y(n_1611)
);

O2A1O1Ixp33_ASAP7_75t_SL g1612 ( 
.A1(n_1399),
.A2(n_72),
.B(n_73),
.C(n_74),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1496),
.B(n_73),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1392),
.A2(n_1415),
.B1(n_1461),
.B2(n_1471),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_SL g1615 ( 
.A1(n_1501),
.A2(n_76),
.B1(n_83),
.B2(n_84),
.Y(n_1615)
);

OAI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1390),
.A2(n_84),
.B1(n_87),
.B2(n_91),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1362),
.Y(n_1617)
);

A2O1A1Ixp33_ASAP7_75t_L g1618 ( 
.A1(n_1342),
.A2(n_91),
.B(n_95),
.C(n_107),
.Y(n_1618)
);

OAI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1378),
.A2(n_95),
.B1(n_109),
.B2(n_111),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1452),
.A2(n_215),
.B1(n_117),
.B2(n_118),
.Y(n_1620)
);

AO31x2_ASAP7_75t_L g1621 ( 
.A1(n_1433),
.A2(n_114),
.A3(n_121),
.B(n_123),
.Y(n_1621)
);

OAI211xp5_ASAP7_75t_SL g1622 ( 
.A1(n_1443),
.A2(n_125),
.B(n_126),
.C(n_128),
.Y(n_1622)
);

OAI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1378),
.A2(n_132),
.B1(n_137),
.B2(n_139),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1370),
.B(n_1420),
.Y(n_1624)
);

A2O1A1Ixp33_ASAP7_75t_L g1625 ( 
.A1(n_1344),
.A2(n_141),
.B(n_144),
.C(n_145),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1420),
.B(n_146),
.Y(n_1626)
);

AND2x2_ASAP7_75t_SL g1627 ( 
.A(n_1324),
.B(n_148),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1452),
.A2(n_150),
.B1(n_160),
.B2(n_162),
.Y(n_1628)
);

OAI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1457),
.A2(n_164),
.B1(n_167),
.B2(n_170),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1370),
.B(n_171),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1379),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1429),
.B(n_211),
.Y(n_1632)
);

OAI21x1_ASAP7_75t_L g1633 ( 
.A1(n_1473),
.A2(n_178),
.B(n_185),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1370),
.B(n_192),
.Y(n_1634)
);

OR2x6_ASAP7_75t_L g1635 ( 
.A(n_1378),
.B(n_206),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1497),
.B(n_1500),
.Y(n_1636)
);

NAND2xp33_ASAP7_75t_SL g1637 ( 
.A(n_1443),
.B(n_1394),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1444),
.Y(n_1638)
);

BUFx10_ASAP7_75t_L g1639 ( 
.A(n_1469),
.Y(n_1639)
);

AOI21xp33_ASAP7_75t_L g1640 ( 
.A1(n_1452),
.A2(n_1471),
.B(n_1501),
.Y(n_1640)
);

OAI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1460),
.A2(n_1471),
.B1(n_1452),
.B2(n_1406),
.Y(n_1641)
);

BUFx2_ASAP7_75t_L g1642 ( 
.A(n_1330),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1370),
.B(n_1420),
.Y(n_1643)
);

OAI21x1_ASAP7_75t_L g1644 ( 
.A1(n_1468),
.A2(n_1351),
.B(n_1476),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1340),
.B(n_1458),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1340),
.B(n_1387),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1340),
.B(n_1387),
.Y(n_1647)
);

NAND3xp33_ASAP7_75t_L g1648 ( 
.A(n_1471),
.B(n_1501),
.C(n_1483),
.Y(n_1648)
);

HB1xp67_ASAP7_75t_L g1649 ( 
.A(n_1453),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1497),
.B(n_1500),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1501),
.A2(n_1433),
.B1(n_1451),
.B2(n_1467),
.Y(n_1651)
);

INVx3_ASAP7_75t_L g1652 ( 
.A(n_1350),
.Y(n_1652)
);

NOR2x1p5_ASAP7_75t_L g1653 ( 
.A(n_1459),
.B(n_1466),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_1459),
.Y(n_1654)
);

AOI21xp5_ASAP7_75t_L g1655 ( 
.A1(n_1324),
.A2(n_1346),
.B(n_1402),
.Y(n_1655)
);

OAI22xp5_ASAP7_75t_L g1656 ( 
.A1(n_1438),
.A2(n_1480),
.B1(n_1453),
.B2(n_1482),
.Y(n_1656)
);

NAND2x1_ASAP7_75t_L g1657 ( 
.A(n_1404),
.B(n_1431),
.Y(n_1657)
);

OAI221xp5_ASAP7_75t_SL g1658 ( 
.A1(n_1340),
.A2(n_1467),
.B1(n_1451),
.B2(n_1498),
.C(n_1493),
.Y(n_1658)
);

INVx6_ASAP7_75t_L g1659 ( 
.A(n_1495),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1387),
.Y(n_1660)
);

OAI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1482),
.A2(n_1431),
.B1(n_1404),
.B2(n_1477),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1441),
.B(n_1498),
.Y(n_1662)
);

AND2x4_ASAP7_75t_L g1663 ( 
.A(n_1466),
.B(n_1464),
.Y(n_1663)
);

CKINVDCx9p33_ASAP7_75t_R g1664 ( 
.A(n_1441),
.Y(n_1664)
);

INVx3_ASAP7_75t_L g1665 ( 
.A(n_1350),
.Y(n_1665)
);

AND2x4_ASAP7_75t_L g1666 ( 
.A(n_1464),
.B(n_1469),
.Y(n_1666)
);

BUFx12f_ASAP7_75t_L g1667 ( 
.A(n_1350),
.Y(n_1667)
);

INVx4_ASAP7_75t_L g1668 ( 
.A(n_1464),
.Y(n_1668)
);

AOI22xp33_ASAP7_75t_L g1669 ( 
.A1(n_1483),
.A2(n_1327),
.B1(n_1377),
.B2(n_1368),
.Y(n_1669)
);

INVx8_ASAP7_75t_L g1670 ( 
.A(n_1469),
.Y(n_1670)
);

INVx4_ASAP7_75t_SL g1671 ( 
.A(n_1495),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1327),
.Y(n_1672)
);

INVx8_ASAP7_75t_L g1673 ( 
.A(n_1487),
.Y(n_1673)
);

INVx3_ASAP7_75t_L g1674 ( 
.A(n_1375),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1477),
.B(n_1417),
.Y(n_1675)
);

INVxp67_ASAP7_75t_SL g1676 ( 
.A(n_1428),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1340),
.B(n_1487),
.Y(n_1677)
);

OAI221xp5_ASAP7_75t_L g1678 ( 
.A1(n_1483),
.A2(n_1454),
.B1(n_1499),
.B2(n_1396),
.C(n_1482),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1362),
.Y(n_1679)
);

BUFx2_ASAP7_75t_L g1680 ( 
.A(n_1375),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1358),
.Y(n_1681)
);

INVx4_ASAP7_75t_L g1682 ( 
.A(n_1487),
.Y(n_1682)
);

HB1xp67_ASAP7_75t_L g1683 ( 
.A(n_1396),
.Y(n_1683)
);

INVx6_ASAP7_75t_L g1684 ( 
.A(n_1495),
.Y(n_1684)
);

BUFx2_ASAP7_75t_SL g1685 ( 
.A(n_1490),
.Y(n_1685)
);

HB1xp67_ASAP7_75t_L g1686 ( 
.A(n_1396),
.Y(n_1686)
);

OAI22x1_ASAP7_75t_L g1687 ( 
.A1(n_1483),
.A2(n_1396),
.B1(n_1395),
.B2(n_1454),
.Y(n_1687)
);

OAI221xp5_ASAP7_75t_L g1688 ( 
.A1(n_1519),
.A2(n_1605),
.B1(n_1618),
.B2(n_1615),
.C(n_1604),
.Y(n_1688)
);

AOI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1519),
.A2(n_1495),
.B1(n_1394),
.B2(n_1490),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1581),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1588),
.B(n_1445),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1513),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1503),
.A2(n_1377),
.B1(n_1368),
.B2(n_1394),
.Y(n_1693)
);

AND2x4_ASAP7_75t_L g1694 ( 
.A(n_1561),
.B(n_1465),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1586),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1503),
.A2(n_1421),
.B1(n_1495),
.B2(n_1416),
.Y(n_1696)
);

AOI22xp33_ASAP7_75t_SL g1697 ( 
.A1(n_1627),
.A2(n_1421),
.B1(n_1465),
.B2(n_1417),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1592),
.Y(n_1698)
);

AOI222xp33_ASAP7_75t_L g1699 ( 
.A1(n_1575),
.A2(n_1424),
.B1(n_1489),
.B2(n_1494),
.C1(n_1492),
.C2(n_1490),
.Y(n_1699)
);

BUFx2_ASAP7_75t_L g1700 ( 
.A(n_1664),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1599),
.Y(n_1701)
);

AO21x2_ASAP7_75t_L g1702 ( 
.A1(n_1640),
.A2(n_1494),
.B(n_1489),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1517),
.A2(n_1506),
.B1(n_1598),
.B2(n_1605),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1517),
.A2(n_1424),
.B1(n_1465),
.B2(n_1436),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1580),
.B(n_1428),
.Y(n_1705)
);

AOI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1529),
.A2(n_1454),
.B1(n_1445),
.B2(n_1440),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1517),
.A2(n_1506),
.B1(n_1509),
.B2(n_1561),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1607),
.Y(n_1708)
);

BUFx2_ASAP7_75t_L g1709 ( 
.A(n_1664),
.Y(n_1709)
);

OAI221xp5_ASAP7_75t_SL g1710 ( 
.A1(n_1618),
.A2(n_1436),
.B1(n_1440),
.B2(n_1492),
.C(n_1446),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1561),
.A2(n_1337),
.B1(n_1355),
.B2(n_1373),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_L g1712 ( 
.A1(n_1511),
.A2(n_1337),
.B1(n_1355),
.B2(n_1373),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1548),
.B(n_1355),
.Y(n_1713)
);

OA21x2_ASAP7_75t_L g1714 ( 
.A1(n_1644),
.A2(n_1351),
.B(n_1468),
.Y(n_1714)
);

AOI222xp33_ASAP7_75t_L g1715 ( 
.A1(n_1616),
.A2(n_1363),
.B1(n_1364),
.B2(n_1365),
.C1(n_1348),
.C2(n_1332),
.Y(n_1715)
);

OAI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1604),
.A2(n_1491),
.B(n_1381),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1526),
.Y(n_1717)
);

AOI221xp5_ASAP7_75t_L g1718 ( 
.A1(n_1612),
.A2(n_1446),
.B1(n_1463),
.B2(n_1462),
.C(n_1393),
.Y(n_1718)
);

NOR2xp33_ASAP7_75t_L g1719 ( 
.A(n_1584),
.B(n_1404),
.Y(n_1719)
);

NAND2x1_ASAP7_75t_L g1720 ( 
.A(n_1563),
.B(n_1431),
.Y(n_1720)
);

AOI221xp5_ASAP7_75t_L g1721 ( 
.A1(n_1612),
.A2(n_1462),
.B1(n_1463),
.B2(n_1393),
.C(n_1502),
.Y(n_1721)
);

OAI221xp5_ASAP7_75t_L g1722 ( 
.A1(n_1508),
.A2(n_1337),
.B1(n_1355),
.B2(n_1499),
.C(n_1375),
.Y(n_1722)
);

AND2x4_ASAP7_75t_L g1723 ( 
.A(n_1507),
.B(n_1395),
.Y(n_1723)
);

INVx3_ASAP7_75t_L g1724 ( 
.A(n_1563),
.Y(n_1724)
);

OAI211xp5_ASAP7_75t_L g1725 ( 
.A1(n_1603),
.A2(n_1601),
.B(n_1549),
.C(n_1514),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1591),
.B(n_1337),
.Y(n_1726)
);

AOI221xp5_ASAP7_75t_L g1727 ( 
.A1(n_1601),
.A2(n_1603),
.B1(n_1611),
.B2(n_1658),
.C(n_1610),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1595),
.B(n_1393),
.Y(n_1728)
);

AOI22xp33_ASAP7_75t_L g1729 ( 
.A1(n_1587),
.A2(n_1363),
.B1(n_1400),
.B2(n_1348),
.Y(n_1729)
);

OAI211xp5_ASAP7_75t_L g1730 ( 
.A1(n_1554),
.A2(n_1491),
.B(n_1381),
.C(n_1434),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1649),
.B(n_1393),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1648),
.A2(n_1400),
.B1(n_1502),
.B2(n_1364),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1672),
.Y(n_1733)
);

AOI221xp5_ASAP7_75t_L g1734 ( 
.A1(n_1641),
.A2(n_1393),
.B1(n_1502),
.B2(n_1499),
.C(n_1332),
.Y(n_1734)
);

OAI221xp5_ASAP7_75t_L g1735 ( 
.A1(n_1620),
.A2(n_1434),
.B1(n_1336),
.B2(n_1432),
.C(n_1427),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1527),
.Y(n_1736)
);

OAI211xp5_ASAP7_75t_L g1737 ( 
.A1(n_1620),
.A2(n_1434),
.B(n_1427),
.C(n_1336),
.Y(n_1737)
);

AOI22xp33_ASAP7_75t_L g1738 ( 
.A1(n_1677),
.A2(n_1365),
.B1(n_1338),
.B2(n_1434),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1505),
.B(n_1374),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1537),
.Y(n_1740)
);

OAI211xp5_ASAP7_75t_L g1741 ( 
.A1(n_1628),
.A2(n_1374),
.B(n_1376),
.C(n_1476),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_SL g1742 ( 
.A1(n_1627),
.A2(n_1432),
.B1(n_1435),
.B2(n_1449),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1542),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1559),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1507),
.A2(n_1338),
.B1(n_1376),
.B2(n_1435),
.Y(n_1745)
);

OAI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1589),
.A2(n_1449),
.B1(n_1439),
.B2(n_1447),
.Y(n_1746)
);

BUFx2_ASAP7_75t_L g1747 ( 
.A(n_1646),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1507),
.A2(n_1439),
.B1(n_1447),
.B2(n_1530),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1565),
.B(n_1566),
.Y(n_1749)
);

NAND3xp33_ASAP7_75t_L g1750 ( 
.A(n_1628),
.B(n_1582),
.C(n_1613),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1645),
.B(n_1647),
.Y(n_1751)
);

AOI22xp33_ASAP7_75t_L g1752 ( 
.A1(n_1518),
.A2(n_1535),
.B1(n_1589),
.B2(n_1536),
.Y(n_1752)
);

OAI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1625),
.A2(n_1538),
.B1(n_1518),
.B2(n_1590),
.Y(n_1753)
);

AOI221xp5_ASAP7_75t_L g1754 ( 
.A1(n_1568),
.A2(n_1569),
.B1(n_1600),
.B2(n_1602),
.C(n_1619),
.Y(n_1754)
);

AO31x2_ASAP7_75t_L g1755 ( 
.A1(n_1687),
.A2(n_1617),
.A3(n_1606),
.B(n_1679),
.Y(n_1755)
);

AOI22xp33_ASAP7_75t_L g1756 ( 
.A1(n_1650),
.A2(n_1520),
.B1(n_1614),
.B2(n_1636),
.Y(n_1756)
);

AOI22xp33_ASAP7_75t_L g1757 ( 
.A1(n_1614),
.A2(n_1538),
.B1(n_1635),
.B2(n_1631),
.Y(n_1757)
);

AOI22xp33_ASAP7_75t_L g1758 ( 
.A1(n_1635),
.A2(n_1608),
.B1(n_1504),
.B2(n_1523),
.Y(n_1758)
);

AOI221xp5_ASAP7_75t_L g1759 ( 
.A1(n_1571),
.A2(n_1515),
.B1(n_1546),
.B2(n_1555),
.C(n_1562),
.Y(n_1759)
);

AOI22xp33_ASAP7_75t_L g1760 ( 
.A1(n_1635),
.A2(n_1577),
.B1(n_1573),
.B2(n_1544),
.Y(n_1760)
);

NOR2x1_ASAP7_75t_SL g1761 ( 
.A(n_1516),
.B(n_1667),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1681),
.Y(n_1762)
);

AOI21xp5_ASAP7_75t_L g1763 ( 
.A1(n_1655),
.A2(n_1625),
.B(n_1522),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1584),
.B(n_1512),
.Y(n_1764)
);

OAI21x1_ASAP7_75t_L g1765 ( 
.A1(n_1644),
.A2(n_1567),
.B(n_1633),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1675),
.Y(n_1766)
);

AOI22xp33_ASAP7_75t_L g1767 ( 
.A1(n_1573),
.A2(n_1577),
.B1(n_1544),
.B2(n_1585),
.Y(n_1767)
);

AOI22xp33_ASAP7_75t_L g1768 ( 
.A1(n_1573),
.A2(n_1577),
.B1(n_1638),
.B2(n_1653),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1534),
.Y(n_1769)
);

INVx3_ASAP7_75t_L g1770 ( 
.A(n_1563),
.Y(n_1770)
);

AOI21xp5_ASAP7_75t_SL g1771 ( 
.A1(n_1626),
.A2(n_1547),
.B(n_1545),
.Y(n_1771)
);

OAI221xp5_ASAP7_75t_L g1772 ( 
.A1(n_1572),
.A2(n_1574),
.B1(n_1560),
.B2(n_1531),
.C(n_1570),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1583),
.B(n_1525),
.Y(n_1773)
);

AOI22xp33_ASAP7_75t_L g1774 ( 
.A1(n_1663),
.A2(n_1626),
.B1(n_1662),
.B2(n_1637),
.Y(n_1774)
);

OAI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1524),
.A2(n_1558),
.B1(n_1551),
.B2(n_1525),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1521),
.Y(n_1776)
);

AO221x2_ASAP7_75t_L g1777 ( 
.A1(n_1656),
.A2(n_1623),
.B1(n_1629),
.B2(n_1609),
.C(n_1661),
.Y(n_1777)
);

OAI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1551),
.A2(n_1510),
.B1(n_1564),
.B2(n_1579),
.Y(n_1778)
);

AOI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1663),
.A2(n_1626),
.B1(n_1637),
.B2(n_1539),
.Y(n_1779)
);

HB1xp67_ASAP7_75t_L g1780 ( 
.A(n_1660),
.Y(n_1780)
);

AOI22xp33_ASAP7_75t_L g1781 ( 
.A1(n_1663),
.A2(n_1541),
.B1(n_1552),
.B2(n_1539),
.Y(n_1781)
);

AOI22xp33_ASAP7_75t_SL g1782 ( 
.A1(n_1543),
.A2(n_1576),
.B1(n_1678),
.B2(n_1685),
.Y(n_1782)
);

AND2x4_ASAP7_75t_L g1783 ( 
.A(n_1666),
.B(n_1671),
.Y(n_1783)
);

AOI22xp33_ASAP7_75t_L g1784 ( 
.A1(n_1532),
.A2(n_1541),
.B1(n_1552),
.B2(n_1556),
.Y(n_1784)
);

CKINVDCx20_ASAP7_75t_R g1785 ( 
.A(n_1553),
.Y(n_1785)
);

AOI22xp33_ASAP7_75t_SL g1786 ( 
.A1(n_1654),
.A2(n_1510),
.B1(n_1578),
.B2(n_1670),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1556),
.Y(n_1787)
);

INVx3_ASAP7_75t_L g1788 ( 
.A(n_1596),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1651),
.B(n_1606),
.Y(n_1789)
);

AOI22xp33_ASAP7_75t_L g1790 ( 
.A1(n_1651),
.A2(n_1669),
.B1(n_1622),
.B2(n_1659),
.Y(n_1790)
);

AOI21xp5_ASAP7_75t_L g1791 ( 
.A1(n_1533),
.A2(n_1657),
.B(n_1632),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1666),
.B(n_1686),
.Y(n_1792)
);

AOI22xp5_ASAP7_75t_L g1793 ( 
.A1(n_1654),
.A2(n_1516),
.B1(n_1666),
.B2(n_1545),
.Y(n_1793)
);

AOI222xp33_ASAP7_75t_L g1794 ( 
.A1(n_1597),
.A2(n_1510),
.B1(n_1669),
.B2(n_1593),
.C1(n_1642),
.C2(n_1643),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1512),
.B(n_1528),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1683),
.B(n_1668),
.Y(n_1796)
);

AOI21xp5_ASAP7_75t_L g1797 ( 
.A1(n_1516),
.A2(n_1596),
.B(n_1545),
.Y(n_1797)
);

OAI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1579),
.A2(n_1593),
.B1(n_1540),
.B2(n_1550),
.Y(n_1798)
);

OAI22xp33_ASAP7_75t_L g1799 ( 
.A1(n_1550),
.A2(n_1668),
.B1(n_1682),
.B2(n_1673),
.Y(n_1799)
);

OAI21xp33_ASAP7_75t_L g1800 ( 
.A1(n_1564),
.A2(n_1528),
.B(n_1553),
.Y(n_1800)
);

AOI211xp5_ASAP7_75t_L g1801 ( 
.A1(n_1630),
.A2(n_1634),
.B(n_1624),
.C(n_1609),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1668),
.B(n_1682),
.Y(n_1802)
);

AOI22xp33_ASAP7_75t_L g1803 ( 
.A1(n_1659),
.A2(n_1684),
.B1(n_1673),
.B2(n_1670),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1682),
.B(n_1557),
.Y(n_1804)
);

AOI22xp33_ASAP7_75t_SL g1805 ( 
.A1(n_1670),
.A2(n_1673),
.B1(n_1684),
.B2(n_1659),
.Y(n_1805)
);

AOI221xp5_ASAP7_75t_L g1806 ( 
.A1(n_1557),
.A2(n_1652),
.B1(n_1674),
.B2(n_1665),
.C(n_1676),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1567),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_1594),
.Y(n_1808)
);

OAI21xp5_ASAP7_75t_SL g1809 ( 
.A1(n_1550),
.A2(n_1680),
.B(n_1665),
.Y(n_1809)
);

AND2x4_ASAP7_75t_L g1810 ( 
.A(n_1671),
.B(n_1674),
.Y(n_1810)
);

OAI21xp5_ASAP7_75t_L g1811 ( 
.A1(n_1633),
.A2(n_1596),
.B(n_1652),
.Y(n_1811)
);

OAI22xp33_ASAP7_75t_L g1812 ( 
.A1(n_1550),
.A2(n_1667),
.B1(n_1684),
.B2(n_1621),
.Y(n_1812)
);

OAI21x1_ASAP7_75t_L g1813 ( 
.A1(n_1621),
.A2(n_1671),
.B(n_1639),
.Y(n_1813)
);

AOI22xp33_ASAP7_75t_L g1814 ( 
.A1(n_1639),
.A2(n_1094),
.B1(n_844),
.B2(n_1519),
.Y(n_1814)
);

AOI22xp33_ASAP7_75t_L g1815 ( 
.A1(n_1639),
.A2(n_1094),
.B1(n_844),
.B2(n_1519),
.Y(n_1815)
);

OAI22xp33_ASAP7_75t_L g1816 ( 
.A1(n_1621),
.A2(n_933),
.B1(n_1426),
.B2(n_1057),
.Y(n_1816)
);

O2A1O1Ixp33_ASAP7_75t_L g1817 ( 
.A1(n_1621),
.A2(n_856),
.B(n_841),
.C(n_852),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1588),
.B(n_1442),
.Y(n_1818)
);

AOI22xp33_ASAP7_75t_SL g1819 ( 
.A1(n_1627),
.A2(n_1094),
.B1(n_1281),
.B2(n_454),
.Y(n_1819)
);

AOI22xp33_ASAP7_75t_L g1820 ( 
.A1(n_1519),
.A2(n_1094),
.B1(n_844),
.B2(n_556),
.Y(n_1820)
);

AOI21xp5_ASAP7_75t_L g1821 ( 
.A1(n_1627),
.A2(n_1228),
.B(n_1201),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1581),
.Y(n_1822)
);

OAI211xp5_ASAP7_75t_L g1823 ( 
.A1(n_1519),
.A2(n_856),
.B(n_851),
.C(n_852),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1588),
.B(n_1442),
.Y(n_1824)
);

AOI22xp33_ASAP7_75t_SL g1825 ( 
.A1(n_1627),
.A2(n_1094),
.B1(n_1281),
.B2(n_454),
.Y(n_1825)
);

OAI22xp33_ASAP7_75t_L g1826 ( 
.A1(n_1529),
.A2(n_933),
.B1(n_1426),
.B2(n_1057),
.Y(n_1826)
);

AOI21xp33_ASAP7_75t_L g1827 ( 
.A1(n_1648),
.A2(n_1508),
.B(n_856),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_SL g1828 ( 
.A(n_1627),
.B(n_1519),
.Y(n_1828)
);

INVx5_ASAP7_75t_SL g1829 ( 
.A(n_1609),
.Y(n_1829)
);

AOI221xp5_ASAP7_75t_L g1830 ( 
.A1(n_1575),
.A2(n_856),
.B1(n_842),
.B2(n_1009),
.C(n_757),
.Y(n_1830)
);

OAI221xp5_ASAP7_75t_L g1831 ( 
.A1(n_1519),
.A2(n_856),
.B1(n_1009),
.B2(n_852),
.C(n_851),
.Y(n_1831)
);

AOI22xp33_ASAP7_75t_L g1832 ( 
.A1(n_1519),
.A2(n_1094),
.B1(n_844),
.B2(n_556),
.Y(n_1832)
);

OAI22xp5_ASAP7_75t_L g1833 ( 
.A1(n_1519),
.A2(n_856),
.B1(n_1618),
.B2(n_1207),
.Y(n_1833)
);

OR2x2_ASAP7_75t_L g1834 ( 
.A(n_1649),
.B(n_1505),
.Y(n_1834)
);

AOI21xp5_ASAP7_75t_SL g1835 ( 
.A1(n_1618),
.A2(n_1604),
.B(n_1625),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1519),
.A2(n_1094),
.B1(n_844),
.B2(n_556),
.Y(n_1836)
);

AOI21xp33_ASAP7_75t_SL g1837 ( 
.A1(n_1553),
.A2(n_826),
.B(n_795),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1588),
.B(n_1442),
.Y(n_1838)
);

AOI22xp33_ASAP7_75t_L g1839 ( 
.A1(n_1519),
.A2(n_1094),
.B1(n_844),
.B2(n_556),
.Y(n_1839)
);

BUFx2_ASAP7_75t_L g1840 ( 
.A(n_1513),
.Y(n_1840)
);

AOI222xp33_ASAP7_75t_L g1841 ( 
.A1(n_1519),
.A2(n_757),
.B1(n_1256),
.B2(n_1094),
.C1(n_1126),
.C2(n_1249),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1588),
.B(n_1580),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1588),
.B(n_1580),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1581),
.Y(n_1844)
);

AOI22xp33_ASAP7_75t_L g1845 ( 
.A1(n_1519),
.A2(n_1094),
.B1(n_844),
.B2(n_556),
.Y(n_1845)
);

AOI221xp5_ASAP7_75t_L g1846 ( 
.A1(n_1575),
.A2(n_856),
.B1(n_842),
.B2(n_1009),
.C(n_757),
.Y(n_1846)
);

OAI22xp33_ASAP7_75t_L g1847 ( 
.A1(n_1529),
.A2(n_933),
.B1(n_1426),
.B2(n_1057),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1733),
.Y(n_1848)
);

NAND2x1p5_ASAP7_75t_L g1849 ( 
.A(n_1813),
.B(n_1828),
.Y(n_1849)
);

HB1xp67_ASAP7_75t_L g1850 ( 
.A(n_1840),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1747),
.B(n_1751),
.Y(n_1851)
);

HB1xp67_ASAP7_75t_L g1852 ( 
.A(n_1840),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1733),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1762),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1751),
.B(n_1747),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1690),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1695),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1834),
.B(n_1728),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1792),
.B(n_1842),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1792),
.B(n_1842),
.Y(n_1860)
);

HB1xp67_ASAP7_75t_L g1861 ( 
.A(n_1692),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1698),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1701),
.Y(n_1863)
);

HB1xp67_ASAP7_75t_L g1864 ( 
.A(n_1749),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1708),
.Y(n_1865)
);

INVx2_ASAP7_75t_SL g1866 ( 
.A(n_1796),
.Y(n_1866)
);

INVx2_ASAP7_75t_SL g1867 ( 
.A(n_1796),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1822),
.Y(n_1868)
);

OAI33xp33_ASAP7_75t_L g1869 ( 
.A1(n_1833),
.A2(n_1753),
.A3(n_1847),
.B1(n_1826),
.B2(n_1816),
.B3(n_1750),
.Y(n_1869)
);

INVxp67_ASAP7_75t_L g1870 ( 
.A(n_1780),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1843),
.B(n_1691),
.Y(n_1871)
);

NOR2x1_ASAP7_75t_L g1872 ( 
.A(n_1771),
.B(n_1835),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1844),
.Y(n_1873)
);

OR2x2_ASAP7_75t_SL g1874 ( 
.A(n_1713),
.B(n_1726),
.Y(n_1874)
);

INVx3_ASAP7_75t_L g1875 ( 
.A(n_1714),
.Y(n_1875)
);

HB1xp67_ASAP7_75t_L g1876 ( 
.A(n_1749),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1843),
.B(n_1691),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1717),
.Y(n_1878)
);

BUFx2_ASAP7_75t_L g1879 ( 
.A(n_1700),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1834),
.B(n_1731),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1736),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1740),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1743),
.Y(n_1883)
);

INVx2_ASAP7_75t_SL g1884 ( 
.A(n_1723),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1769),
.B(n_1766),
.Y(n_1885)
);

HB1xp67_ASAP7_75t_L g1886 ( 
.A(n_1818),
.Y(n_1886)
);

HB1xp67_ASAP7_75t_L g1887 ( 
.A(n_1824),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1755),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1744),
.Y(n_1889)
);

HB1xp67_ASAP7_75t_L g1890 ( 
.A(n_1838),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1755),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1731),
.B(n_1739),
.Y(n_1892)
);

HB1xp67_ASAP7_75t_L g1893 ( 
.A(n_1755),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1755),
.Y(n_1894)
);

BUFx3_ASAP7_75t_L g1895 ( 
.A(n_1783),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1776),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1787),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1789),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1755),
.Y(n_1899)
);

OR2x2_ASAP7_75t_L g1900 ( 
.A(n_1739),
.B(n_1789),
.Y(n_1900)
);

AND2x4_ASAP7_75t_SL g1901 ( 
.A(n_1783),
.B(n_1723),
.Y(n_1901)
);

INVx4_ASAP7_75t_R g1902 ( 
.A(n_1829),
.Y(n_1902)
);

BUFx12f_ASAP7_75t_L g1903 ( 
.A(n_1808),
.Y(n_1903)
);

NAND2x1p5_ASAP7_75t_L g1904 ( 
.A(n_1813),
.B(n_1828),
.Y(n_1904)
);

INVxp67_ASAP7_75t_L g1905 ( 
.A(n_1723),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1705),
.B(n_1700),
.Y(n_1906)
);

AOI22xp33_ASAP7_75t_L g1907 ( 
.A1(n_1819),
.A2(n_1825),
.B1(n_1688),
.B2(n_1845),
.Y(n_1907)
);

BUFx6f_ASAP7_75t_L g1908 ( 
.A(n_1810),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1804),
.B(n_1705),
.Y(n_1909)
);

HB1xp67_ASAP7_75t_L g1910 ( 
.A(n_1773),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1694),
.B(n_1709),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1694),
.B(n_1709),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1763),
.B(n_1712),
.Y(n_1913)
);

INVxp67_ASAP7_75t_SL g1914 ( 
.A(n_1711),
.Y(n_1914)
);

INVxp67_ASAP7_75t_L g1915 ( 
.A(n_1722),
.Y(n_1915)
);

OAI22xp33_ASAP7_75t_L g1916 ( 
.A1(n_1831),
.A2(n_1772),
.B1(n_1727),
.B2(n_1759),
.Y(n_1916)
);

AND2x4_ASAP7_75t_L g1917 ( 
.A(n_1783),
.B(n_1810),
.Y(n_1917)
);

BUFx2_ASAP7_75t_L g1918 ( 
.A(n_1716),
.Y(n_1918)
);

OR2x2_ASAP7_75t_L g1919 ( 
.A(n_1707),
.B(n_1702),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1702),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1748),
.B(n_1699),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1702),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1738),
.B(n_1704),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1784),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1774),
.B(n_1829),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1745),
.B(n_1706),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1807),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1807),
.Y(n_1928)
);

OR2x2_ASAP7_75t_L g1929 ( 
.A(n_1829),
.B(n_1777),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1765),
.Y(n_1930)
);

NOR2x1_ASAP7_75t_L g1931 ( 
.A(n_1771),
.B(n_1835),
.Y(n_1931)
);

BUFx2_ASAP7_75t_L g1932 ( 
.A(n_1811),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1765),
.Y(n_1933)
);

INVxp33_ASAP7_75t_L g1934 ( 
.A(n_1764),
.Y(n_1934)
);

AOI22xp33_ASAP7_75t_SL g1935 ( 
.A1(n_1777),
.A2(n_1823),
.B1(n_1725),
.B2(n_1829),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1781),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1718),
.Y(n_1937)
);

AOI33xp33_ASAP7_75t_L g1938 ( 
.A1(n_1916),
.A2(n_1846),
.A3(n_1830),
.B1(n_1836),
.B2(n_1832),
.B3(n_1820),
.Y(n_1938)
);

INVxp67_ASAP7_75t_SL g1939 ( 
.A(n_1893),
.Y(n_1939)
);

INVxp67_ASAP7_75t_L g1940 ( 
.A(n_1861),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_SL g1941 ( 
.A(n_1872),
.B(n_1801),
.Y(n_1941)
);

CKINVDCx6p67_ASAP7_75t_R g1942 ( 
.A(n_1903),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1848),
.Y(n_1943)
);

AOI22xp33_ASAP7_75t_SL g1944 ( 
.A1(n_1921),
.A2(n_1777),
.B1(n_1761),
.B2(n_1814),
.Y(n_1944)
);

AOI22xp33_ASAP7_75t_L g1945 ( 
.A1(n_1907),
.A2(n_1841),
.B1(n_1815),
.B2(n_1703),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1888),
.Y(n_1946)
);

OAI31xp33_ASAP7_75t_L g1947 ( 
.A1(n_1921),
.A2(n_1839),
.A3(n_1827),
.B(n_1710),
.Y(n_1947)
);

INVx2_ASAP7_75t_SL g1948 ( 
.A(n_1850),
.Y(n_1948)
);

OR2x6_ASAP7_75t_L g1949 ( 
.A(n_1872),
.B(n_1797),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1848),
.Y(n_1950)
);

OR2x2_ASAP7_75t_L g1951 ( 
.A(n_1851),
.B(n_1775),
.Y(n_1951)
);

NAND4xp25_ASAP7_75t_L g1952 ( 
.A(n_1935),
.B(n_1719),
.C(n_1778),
.D(n_1754),
.Y(n_1952)
);

INVxp67_ASAP7_75t_L g1953 ( 
.A(n_1852),
.Y(n_1953)
);

AND2x2_ASAP7_75t_SL g1954 ( 
.A(n_1918),
.B(n_1760),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1855),
.B(n_1794),
.Y(n_1955)
);

OAI22xp5_ASAP7_75t_L g1956 ( 
.A1(n_1935),
.A2(n_1767),
.B1(n_1752),
.B2(n_1768),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1855),
.B(n_1795),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1871),
.B(n_1714),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1888),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1853),
.Y(n_1960)
);

AOI22xp33_ASAP7_75t_L g1961 ( 
.A1(n_1869),
.A2(n_1693),
.B1(n_1757),
.B2(n_1756),
.Y(n_1961)
);

OA21x2_ASAP7_75t_L g1962 ( 
.A1(n_1920),
.A2(n_1791),
.B(n_1806),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1888),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1853),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1854),
.Y(n_1965)
);

OAI221xp5_ASAP7_75t_SL g1966 ( 
.A1(n_1915),
.A2(n_1817),
.B1(n_1821),
.B2(n_1790),
.C(n_1782),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1891),
.Y(n_1967)
);

AND2x4_ASAP7_75t_L g1968 ( 
.A(n_1901),
.B(n_1793),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1886),
.B(n_1697),
.Y(n_1969)
);

AND2x4_ASAP7_75t_L g1970 ( 
.A(n_1901),
.B(n_1779),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1871),
.B(n_1714),
.Y(n_1971)
);

AOI221xp5_ASAP7_75t_L g1972 ( 
.A1(n_1915),
.A2(n_1812),
.B1(n_1758),
.B2(n_1798),
.C(n_1837),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1887),
.B(n_1802),
.Y(n_1973)
);

BUFx2_ASAP7_75t_L g1974 ( 
.A(n_1879),
.Y(n_1974)
);

OAI211xp5_ASAP7_75t_L g1975 ( 
.A1(n_1918),
.A2(n_1913),
.B(n_1931),
.C(n_1929),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1877),
.B(n_1786),
.Y(n_1976)
);

INVx1_ASAP7_75t_SL g1977 ( 
.A(n_1903),
.Y(n_1977)
);

NAND2xp33_ASAP7_75t_SL g1978 ( 
.A(n_1929),
.B(n_1785),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1854),
.Y(n_1979)
);

OAI33xp33_ASAP7_75t_L g1980 ( 
.A1(n_1937),
.A2(n_1800),
.A3(n_1799),
.B1(n_1808),
.B2(n_1746),
.B3(n_1785),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1890),
.B(n_1788),
.Y(n_1981)
);

AOI22xp33_ASAP7_75t_L g1982 ( 
.A1(n_1869),
.A2(n_1696),
.B1(n_1689),
.B2(n_1721),
.Y(n_1982)
);

OAI22xp5_ASAP7_75t_L g1983 ( 
.A1(n_1931),
.A2(n_1805),
.B1(n_1803),
.B2(n_1724),
.Y(n_1983)
);

OAI321xp33_ASAP7_75t_L g1984 ( 
.A1(n_1937),
.A2(n_1741),
.A3(n_1737),
.B1(n_1730),
.B2(n_1734),
.C(n_1735),
.Y(n_1984)
);

AOI22xp5_ASAP7_75t_L g1985 ( 
.A1(n_1926),
.A2(n_1923),
.B1(n_1914),
.B2(n_1913),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_R g1986 ( 
.A(n_1903),
.B(n_1788),
.Y(n_1986)
);

OA21x2_ASAP7_75t_L g1987 ( 
.A1(n_1920),
.A2(n_1809),
.B(n_1729),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1856),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1856),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1877),
.B(n_1788),
.Y(n_1990)
);

NAND4xp25_ASAP7_75t_L g1991 ( 
.A(n_1879),
.B(n_1870),
.C(n_1932),
.D(n_1875),
.Y(n_1991)
);

OAI221xp5_ASAP7_75t_L g1992 ( 
.A1(n_1914),
.A2(n_1742),
.B1(n_1732),
.B2(n_1715),
.C(n_1720),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1857),
.Y(n_1993)
);

AO21x2_ASAP7_75t_L g1994 ( 
.A1(n_1922),
.A2(n_1761),
.B(n_1810),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1857),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1862),
.Y(n_1996)
);

OAI22xp5_ASAP7_75t_L g1997 ( 
.A1(n_1851),
.A2(n_1724),
.B1(n_1770),
.B2(n_1720),
.Y(n_1997)
);

OAI211xp5_ASAP7_75t_L g1998 ( 
.A1(n_1932),
.A2(n_1724),
.B(n_1770),
.C(n_1870),
.Y(n_1998)
);

AOI211xp5_ASAP7_75t_L g1999 ( 
.A1(n_1919),
.A2(n_1770),
.B(n_1926),
.C(n_1923),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1862),
.Y(n_2000)
);

AND2x4_ASAP7_75t_L g2001 ( 
.A(n_1901),
.B(n_1895),
.Y(n_2001)
);

OAI221xp5_ASAP7_75t_L g2002 ( 
.A1(n_1849),
.A2(n_1904),
.B1(n_1919),
.B2(n_1893),
.C(n_1936),
.Y(n_2002)
);

OAI211xp5_ASAP7_75t_SL g2003 ( 
.A1(n_1875),
.A2(n_1905),
.B(n_1863),
.C(n_1873),
.Y(n_2003)
);

AOI22xp5_ASAP7_75t_L g2004 ( 
.A1(n_1936),
.A2(n_1925),
.B1(n_1849),
.B2(n_1904),
.Y(n_2004)
);

AOI21x1_ASAP7_75t_L g2005 ( 
.A1(n_1922),
.A2(n_1930),
.B(n_1933),
.Y(n_2005)
);

OR2x6_ASAP7_75t_L g2006 ( 
.A(n_1849),
.B(n_1904),
.Y(n_2006)
);

NAND3xp33_ASAP7_75t_L g2007 ( 
.A(n_1885),
.B(n_1905),
.C(n_1892),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1863),
.Y(n_2008)
);

AOI22xp33_ASAP7_75t_L g2009 ( 
.A1(n_1924),
.A2(n_1898),
.B1(n_1894),
.B2(n_1891),
.Y(n_2009)
);

AOI31xp67_ASAP7_75t_L g2010 ( 
.A1(n_1930),
.A2(n_1933),
.A3(n_1927),
.B(n_1928),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1859),
.B(n_1860),
.Y(n_2011)
);

CKINVDCx6p67_ASAP7_75t_R g2012 ( 
.A(n_1895),
.Y(n_2012)
);

OAI31xp33_ASAP7_75t_L g2013 ( 
.A1(n_1924),
.A2(n_1925),
.A3(n_1898),
.B(n_1885),
.Y(n_2013)
);

BUFx3_ASAP7_75t_L g2014 ( 
.A(n_1908),
.Y(n_2014)
);

AOI21xp33_ASAP7_75t_L g2015 ( 
.A1(n_1894),
.A2(n_1899),
.B(n_1878),
.Y(n_2015)
);

OAI221xp5_ASAP7_75t_L g2016 ( 
.A1(n_1900),
.A2(n_1881),
.B1(n_1878),
.B2(n_1882),
.C(n_1883),
.Y(n_2016)
);

AOI22xp33_ASAP7_75t_L g2017 ( 
.A1(n_1894),
.A2(n_1899),
.B1(n_1897),
.B2(n_1896),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1958),
.B(n_1859),
.Y(n_2018)
);

INVx1_ASAP7_75t_SL g2019 ( 
.A(n_1974),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1958),
.B(n_1900),
.Y(n_2020)
);

NOR2xp33_ASAP7_75t_L g2021 ( 
.A(n_1952),
.B(n_1934),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_2010),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1943),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1971),
.B(n_1860),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1950),
.Y(n_2025)
);

OR2x2_ASAP7_75t_L g2026 ( 
.A(n_1971),
.B(n_1874),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1960),
.Y(n_2027)
);

HB1xp67_ASAP7_75t_L g2028 ( 
.A(n_1953),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1964),
.Y(n_2029)
);

BUFx2_ASAP7_75t_L g2030 ( 
.A(n_2001),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_2005),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_2011),
.B(n_1884),
.Y(n_2032)
);

NOR3xp33_ASAP7_75t_L g2033 ( 
.A(n_1944),
.B(n_1875),
.C(n_1868),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1965),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1985),
.B(n_1858),
.Y(n_2035)
);

BUFx6f_ASAP7_75t_L g2036 ( 
.A(n_1962),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_2011),
.B(n_1884),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1979),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1988),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1989),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1946),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1993),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_1995),
.B(n_1858),
.Y(n_2043)
);

INVx1_ASAP7_75t_SL g2044 ( 
.A(n_1948),
.Y(n_2044)
);

OR2x2_ASAP7_75t_L g2045 ( 
.A(n_1991),
.B(n_1874),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1996),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_2000),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_1990),
.B(n_1884),
.Y(n_2048)
);

NAND2xp67_ASAP7_75t_L g2049 ( 
.A(n_1969),
.B(n_1899),
.Y(n_2049)
);

OR2x2_ASAP7_75t_L g2050 ( 
.A(n_2007),
.B(n_1880),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1959),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_2001),
.B(n_1866),
.Y(n_2052)
);

INVx3_ASAP7_75t_L g2053 ( 
.A(n_2001),
.Y(n_2053)
);

AOI22xp33_ASAP7_75t_L g2054 ( 
.A1(n_1945),
.A2(n_1889),
.B1(n_1882),
.B2(n_1881),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_1959),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1963),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_2008),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1963),
.Y(n_2058)
);

INVx1_ASAP7_75t_SL g2059 ( 
.A(n_1948),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1967),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1967),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_2013),
.B(n_1892),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_1955),
.B(n_1867),
.Y(n_2063)
);

AND2x4_ASAP7_75t_SL g2064 ( 
.A(n_1949),
.B(n_1917),
.Y(n_2064)
);

NAND2x1_ASAP7_75t_SL g2065 ( 
.A(n_2004),
.B(n_1917),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_2016),
.B(n_1880),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_1976),
.B(n_1867),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_2014),
.B(n_1867),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1939),
.B(n_1868),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2017),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_2014),
.B(n_1866),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_1940),
.B(n_1999),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_2012),
.B(n_1866),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_2012),
.B(n_1912),
.Y(n_2074)
);

OR2x2_ASAP7_75t_L g2075 ( 
.A(n_1973),
.B(n_1876),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1951),
.B(n_1912),
.Y(n_2076)
);

OR2x2_ASAP7_75t_L g2077 ( 
.A(n_1981),
.B(n_1864),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_2017),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1975),
.B(n_1873),
.Y(n_2079)
);

OR2x2_ASAP7_75t_L g2080 ( 
.A(n_1962),
.B(n_1906),
.Y(n_2080)
);

OAI22xp5_ASAP7_75t_L g2081 ( 
.A1(n_1945),
.A2(n_1906),
.B1(n_1910),
.B2(n_1895),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_1957),
.B(n_1911),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_2023),
.Y(n_2083)
);

OAI21xp33_ASAP7_75t_L g2084 ( 
.A1(n_2045),
.A2(n_2072),
.B(n_2033),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2023),
.Y(n_2085)
);

INVx1_ASAP7_75t_SL g2086 ( 
.A(n_2019),
.Y(n_2086)
);

OR2x2_ASAP7_75t_L g2087 ( 
.A(n_2050),
.B(n_1865),
.Y(n_2087)
);

OR2x2_ASAP7_75t_SL g2088 ( 
.A(n_2045),
.B(n_1962),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_2079),
.B(n_2028),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_2030),
.B(n_1911),
.Y(n_2090)
);

NAND3xp33_ASAP7_75t_L g2091 ( 
.A(n_2036),
.B(n_1947),
.C(n_1966),
.Y(n_2091)
);

OAI221xp5_ASAP7_75t_L g2092 ( 
.A1(n_2033),
.A2(n_2002),
.B1(n_1961),
.B2(n_1982),
.C(n_1956),
.Y(n_2092)
);

OR2x2_ASAP7_75t_L g2093 ( 
.A(n_2050),
.B(n_2066),
.Y(n_2093)
);

NOR2x1_ASAP7_75t_L g2094 ( 
.A(n_2045),
.B(n_1941),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_2031),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_2031),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2025),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_2031),
.Y(n_2098)
);

OAI31xp33_ASAP7_75t_L g2099 ( 
.A1(n_2070),
.A2(n_1941),
.A3(n_1992),
.B(n_1982),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_2030),
.B(n_1968),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2025),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_2030),
.B(n_1968),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_2079),
.B(n_1865),
.Y(n_2103)
);

AOI221xp5_ASAP7_75t_SL g2104 ( 
.A1(n_2072),
.A2(n_1972),
.B1(n_1977),
.B2(n_1997),
.C(n_1961),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_2028),
.B(n_1998),
.Y(n_2105)
);

NAND3xp33_ASAP7_75t_L g2106 ( 
.A(n_2036),
.B(n_2003),
.C(n_1987),
.Y(n_2106)
);

OR2x2_ASAP7_75t_L g2107 ( 
.A(n_2050),
.B(n_1889),
.Y(n_2107)
);

OAI322xp33_ASAP7_75t_L g2108 ( 
.A1(n_2080),
.A2(n_1954),
.A3(n_1883),
.B1(n_1980),
.B2(n_1983),
.C1(n_1984),
.C2(n_1938),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_2066),
.B(n_2075),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2027),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2027),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_2029),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_2053),
.B(n_1968),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2029),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2034),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_2053),
.B(n_1954),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_2075),
.B(n_1909),
.Y(n_2117)
);

AOI22xp5_ASAP7_75t_L g2118 ( 
.A1(n_2021),
.A2(n_1970),
.B1(n_1978),
.B2(n_2006),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_SL g2119 ( 
.A(n_2036),
.B(n_1978),
.Y(n_2119)
);

OR2x2_ASAP7_75t_L g2120 ( 
.A(n_2020),
.B(n_1987),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2034),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_2053),
.B(n_1970),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_2031),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_2036),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2038),
.Y(n_2125)
);

OR2x2_ASAP7_75t_L g2126 ( 
.A(n_2020),
.B(n_1987),
.Y(n_2126)
);

HB1xp67_ASAP7_75t_L g2127 ( 
.A(n_2069),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_2053),
.B(n_1970),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2053),
.B(n_1949),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_2075),
.B(n_1909),
.Y(n_2130)
);

OR2x2_ASAP7_75t_L g2131 ( 
.A(n_2026),
.B(n_1949),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2038),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_2062),
.B(n_1949),
.Y(n_2133)
);

NOR2xp33_ASAP7_75t_L g2134 ( 
.A(n_2021),
.B(n_1942),
.Y(n_2134)
);

NOR2xp33_ASAP7_75t_L g2135 ( 
.A(n_2019),
.B(n_1942),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_2100),
.B(n_2067),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2083),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2083),
.Y(n_2138)
);

NAND4xp25_ASAP7_75t_L g2139 ( 
.A(n_2091),
.B(n_1938),
.C(n_2022),
.D(n_2054),
.Y(n_2139)
);

INVxp67_ASAP7_75t_L g2140 ( 
.A(n_2094),
.Y(n_2140)
);

AND2x4_ASAP7_75t_L g2141 ( 
.A(n_2094),
.B(n_2064),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_2100),
.B(n_2067),
.Y(n_2142)
);

CKINVDCx5p33_ASAP7_75t_R g2143 ( 
.A(n_2134),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_2088),
.Y(n_2144)
);

INVxp67_ASAP7_75t_SL g2145 ( 
.A(n_2106),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_2104),
.B(n_2062),
.Y(n_2146)
);

AND2x4_ASAP7_75t_L g2147 ( 
.A(n_2102),
.B(n_2064),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2085),
.Y(n_2148)
);

OR2x2_ASAP7_75t_L g2149 ( 
.A(n_2109),
.B(n_2026),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_2103),
.B(n_2063),
.Y(n_2150)
);

OR2x2_ASAP7_75t_L g2151 ( 
.A(n_2087),
.B(n_2026),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_2102),
.B(n_2067),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_2099),
.B(n_2063),
.Y(n_2153)
);

NAND3xp33_ASAP7_75t_L g2154 ( 
.A(n_2084),
.B(n_2036),
.C(n_2022),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_2088),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_2124),
.Y(n_2156)
);

OR2x2_ASAP7_75t_L g2157 ( 
.A(n_2087),
.B(n_2080),
.Y(n_2157)
);

AOI22xp33_ASAP7_75t_L g2158 ( 
.A1(n_2092),
.A2(n_2070),
.B1(n_2078),
.B2(n_2036),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2085),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2097),
.Y(n_2160)
);

INVx3_ASAP7_75t_L g2161 ( 
.A(n_2124),
.Y(n_2161)
);

AOI22xp33_ASAP7_75t_L g2162 ( 
.A1(n_2108),
.A2(n_2078),
.B1(n_2036),
.B2(n_2054),
.Y(n_2162)
);

INVx3_ASAP7_75t_L g2163 ( 
.A(n_2122),
.Y(n_2163)
);

HB1xp67_ASAP7_75t_L g2164 ( 
.A(n_2127),
.Y(n_2164)
);

INVx3_ASAP7_75t_SL g2165 ( 
.A(n_2086),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_2089),
.B(n_2063),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_2133),
.B(n_2076),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2097),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2101),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2101),
.Y(n_2170)
);

NOR3xp33_ASAP7_75t_L g2171 ( 
.A(n_2105),
.B(n_2022),
.C(n_2081),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2110),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_2090),
.B(n_2018),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_2095),
.Y(n_2174)
);

NOR3xp33_ASAP7_75t_L g2175 ( 
.A(n_2095),
.B(n_2022),
.C(n_2081),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_2096),
.Y(n_2176)
);

NAND4xp25_ASAP7_75t_L g2177 ( 
.A(n_2135),
.B(n_2059),
.C(n_2044),
.D(n_2080),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_2093),
.B(n_2076),
.Y(n_2178)
);

BUFx2_ASAP7_75t_L g2179 ( 
.A(n_2110),
.Y(n_2179)
);

NAND2x1p5_ASAP7_75t_L g2180 ( 
.A(n_2119),
.B(n_2036),
.Y(n_2180)
);

AND2x2_ASAP7_75t_L g2181 ( 
.A(n_2090),
.B(n_2018),
.Y(n_2181)
);

INVx1_ASAP7_75t_SL g2182 ( 
.A(n_2116),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2111),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_2113),
.B(n_2018),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_2165),
.B(n_2129),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2179),
.Y(n_2186)
);

AOI211x1_ASAP7_75t_L g2187 ( 
.A1(n_2139),
.A2(n_2116),
.B(n_2128),
.C(n_2122),
.Y(n_2187)
);

OAI22xp5_ASAP7_75t_L g2188 ( 
.A1(n_2154),
.A2(n_2118),
.B1(n_2093),
.B2(n_2131),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_2146),
.B(n_2165),
.Y(n_2189)
);

NOR2xp33_ASAP7_75t_L g2190 ( 
.A(n_2165),
.B(n_2131),
.Y(n_2190)
);

AOI22xp5_ASAP7_75t_L g2191 ( 
.A1(n_2139),
.A2(n_2120),
.B1(n_2126),
.B2(n_2035),
.Y(n_2191)
);

CKINVDCx5p33_ASAP7_75t_R g2192 ( 
.A(n_2143),
.Y(n_2192)
);

AOI21xp5_ASAP7_75t_L g2193 ( 
.A1(n_2140),
.A2(n_2035),
.B(n_2126),
.Y(n_2193)
);

INVx1_ASAP7_75t_SL g2194 ( 
.A(n_2144),
.Y(n_2194)
);

INVx1_ASAP7_75t_SL g2195 ( 
.A(n_2144),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2179),
.Y(n_2196)
);

NAND3xp33_ASAP7_75t_SL g2197 ( 
.A(n_2171),
.B(n_2120),
.C(n_2129),
.Y(n_2197)
);

O2A1O1Ixp33_ASAP7_75t_L g2198 ( 
.A1(n_2144),
.A2(n_2096),
.B(n_2098),
.C(n_2123),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2137),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_2136),
.B(n_2113),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2137),
.Y(n_2201)
);

INVx1_ASAP7_75t_SL g2202 ( 
.A(n_2155),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_2163),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2138),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_2164),
.B(n_2107),
.Y(n_2205)
);

OR2x2_ASAP7_75t_L g2206 ( 
.A(n_2178),
.B(n_2107),
.Y(n_2206)
);

AND2x2_ASAP7_75t_L g2207 ( 
.A(n_2136),
.B(n_2128),
.Y(n_2207)
);

O2A1O1Ixp33_ASAP7_75t_SL g2208 ( 
.A1(n_2155),
.A2(n_2059),
.B(n_2044),
.C(n_2117),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2138),
.Y(n_2209)
);

AOI22xp5_ASAP7_75t_L g2210 ( 
.A1(n_2162),
.A2(n_2155),
.B1(n_2145),
.B2(n_2158),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_2142),
.B(n_2152),
.Y(n_2211)
);

AOI31xp33_ASAP7_75t_L g2212 ( 
.A1(n_2154),
.A2(n_2073),
.A3(n_2074),
.B(n_2076),
.Y(n_2212)
);

AOI22xp5_ASAP7_75t_L g2213 ( 
.A1(n_2175),
.A2(n_2006),
.B1(n_2123),
.B2(n_2098),
.Y(n_2213)
);

OAI21xp5_ASAP7_75t_L g2214 ( 
.A1(n_2177),
.A2(n_2065),
.B(n_2132),
.Y(n_2214)
);

OR2x2_ASAP7_75t_L g2215 ( 
.A(n_2149),
.B(n_2130),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2148),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2148),
.Y(n_2217)
);

OA22x2_ASAP7_75t_L g2218 ( 
.A1(n_2153),
.A2(n_2006),
.B1(n_2125),
.B2(n_2121),
.Y(n_2218)
);

NAND4xp25_ASAP7_75t_L g2219 ( 
.A(n_2177),
.B(n_2132),
.C(n_2125),
.D(n_2121),
.Y(n_2219)
);

AOI221xp5_ASAP7_75t_L g2220 ( 
.A1(n_2157),
.A2(n_2115),
.B1(n_2114),
.B2(n_2112),
.C(n_2111),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_2182),
.B(n_2112),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2159),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2159),
.Y(n_2223)
);

NAND3xp33_ASAP7_75t_L g2224 ( 
.A(n_2191),
.B(n_2141),
.C(n_2163),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2199),
.Y(n_2225)
);

AOI22xp5_ASAP7_75t_L g2226 ( 
.A1(n_2210),
.A2(n_2182),
.B1(n_2141),
.B2(n_2176),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_2187),
.B(n_2142),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_2185),
.B(n_2152),
.Y(n_2228)
);

AOI22xp5_ASAP7_75t_L g2229 ( 
.A1(n_2197),
.A2(n_2195),
.B1(n_2194),
.B2(n_2202),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2201),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2204),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2209),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_2203),
.Y(n_2233)
);

AOI22xp33_ASAP7_75t_L g2234 ( 
.A1(n_2189),
.A2(n_2176),
.B1(n_2174),
.B2(n_2141),
.Y(n_2234)
);

OAI22xp5_ASAP7_75t_L g2235 ( 
.A1(n_2212),
.A2(n_2141),
.B1(n_2147),
.B2(n_2180),
.Y(n_2235)
);

AOI22xp5_ASAP7_75t_L g2236 ( 
.A1(n_2218),
.A2(n_2190),
.B1(n_2188),
.B2(n_2219),
.Y(n_2236)
);

NAND3xp33_ASAP7_75t_L g2237 ( 
.A(n_2193),
.B(n_2163),
.C(n_2183),
.Y(n_2237)
);

XNOR2x2_ASAP7_75t_L g2238 ( 
.A(n_2190),
.B(n_2149),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_2186),
.B(n_2173),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_2196),
.B(n_2173),
.Y(n_2240)
);

A2O1A1Ixp33_ASAP7_75t_L g2241 ( 
.A1(n_2214),
.A2(n_2065),
.B(n_2157),
.C(n_2151),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2216),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2217),
.Y(n_2243)
);

OAI21xp5_ASAP7_75t_L g2244 ( 
.A1(n_2208),
.A2(n_2180),
.B(n_2163),
.Y(n_2244)
);

AOI21xp33_ASAP7_75t_L g2245 ( 
.A1(n_2218),
.A2(n_2176),
.B(n_2174),
.Y(n_2245)
);

AOI221xp5_ASAP7_75t_L g2246 ( 
.A1(n_2198),
.A2(n_2174),
.B1(n_2183),
.B2(n_2170),
.C(n_2160),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_2211),
.B(n_2181),
.Y(n_2247)
);

AOI221x1_ASAP7_75t_L g2248 ( 
.A1(n_2203),
.A2(n_2160),
.B1(n_2172),
.B2(n_2170),
.C(n_2169),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2222),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2223),
.Y(n_2250)
);

XNOR2xp5_ASAP7_75t_L g2251 ( 
.A(n_2192),
.B(n_2185),
.Y(n_2251)
);

OAI221xp5_ASAP7_75t_L g2252 ( 
.A1(n_2213),
.A2(n_2180),
.B1(n_2151),
.B2(n_2167),
.C(n_2166),
.Y(n_2252)
);

INVx4_ASAP7_75t_L g2253 ( 
.A(n_2233),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_2228),
.B(n_2211),
.Y(n_2254)
);

INVxp67_ASAP7_75t_L g2255 ( 
.A(n_2251),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_2247),
.B(n_2192),
.Y(n_2256)
);

AND2x2_ASAP7_75t_L g2257 ( 
.A(n_2234),
.B(n_2207),
.Y(n_2257)
);

INVx1_ASAP7_75t_SL g2258 ( 
.A(n_2238),
.Y(n_2258)
);

CKINVDCx5p33_ASAP7_75t_R g2259 ( 
.A(n_2238),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_2229),
.B(n_2207),
.Y(n_2260)
);

NOR2xp33_ASAP7_75t_L g2261 ( 
.A(n_2239),
.B(n_2215),
.Y(n_2261)
);

AND2x2_ASAP7_75t_L g2262 ( 
.A(n_2234),
.B(n_2200),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2248),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2225),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2240),
.B(n_2200),
.Y(n_2265)
);

OR2x2_ASAP7_75t_L g2266 ( 
.A(n_2227),
.B(n_2205),
.Y(n_2266)
);

INVx1_ASAP7_75t_SL g2267 ( 
.A(n_2226),
.Y(n_2267)
);

NOR3xp33_ASAP7_75t_L g2268 ( 
.A(n_2224),
.B(n_2208),
.C(n_2221),
.Y(n_2268)
);

NOR3xp33_ASAP7_75t_SL g2269 ( 
.A(n_2235),
.B(n_2220),
.C(n_2150),
.Y(n_2269)
);

AOI21xp5_ASAP7_75t_L g2270 ( 
.A1(n_2241),
.A2(n_2169),
.B(n_2168),
.Y(n_2270)
);

AOI21x1_ASAP7_75t_L g2271 ( 
.A1(n_2233),
.A2(n_2168),
.B(n_2172),
.Y(n_2271)
);

AND2x2_ASAP7_75t_L g2272 ( 
.A(n_2244),
.B(n_2147),
.Y(n_2272)
);

INVx1_ASAP7_75t_SL g2273 ( 
.A(n_2236),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_2230),
.B(n_2181),
.Y(n_2274)
);

AOI31xp33_ASAP7_75t_L g2275 ( 
.A1(n_2237),
.A2(n_2206),
.A3(n_2147),
.B(n_2184),
.Y(n_2275)
);

NAND3xp33_ASAP7_75t_L g2276 ( 
.A(n_2259),
.B(n_2246),
.C(n_2241),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_SL g2277 ( 
.A(n_2259),
.B(n_2147),
.Y(n_2277)
);

OR2x2_ASAP7_75t_L g2278 ( 
.A(n_2258),
.B(n_2231),
.Y(n_2278)
);

NOR4xp25_ASAP7_75t_L g2279 ( 
.A(n_2263),
.B(n_2242),
.C(n_2250),
.D(n_2249),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2253),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2253),
.Y(n_2281)
);

NAND4xp25_ASAP7_75t_SL g2282 ( 
.A(n_2268),
.B(n_2252),
.C(n_2243),
.D(n_2232),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2261),
.B(n_2184),
.Y(n_2283)
);

NOR2xp33_ASAP7_75t_L g2284 ( 
.A(n_2255),
.B(n_2114),
.Y(n_2284)
);

OAI21xp33_ASAP7_75t_SL g2285 ( 
.A1(n_2263),
.A2(n_2245),
.B(n_2161),
.Y(n_2285)
);

NOR2xp33_ASAP7_75t_L g2286 ( 
.A(n_2256),
.B(n_2161),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_2257),
.B(n_2262),
.Y(n_2287)
);

NAND5xp2_ASAP7_75t_L g2288 ( 
.A(n_2269),
.B(n_2073),
.C(n_2074),
.D(n_2052),
.E(n_2032),
.Y(n_2288)
);

NOR2x1p5_ASAP7_75t_L g2289 ( 
.A(n_2260),
.B(n_2161),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_L g2290 ( 
.A(n_2257),
.B(n_2115),
.Y(n_2290)
);

OAI221xp5_ASAP7_75t_L g2291 ( 
.A1(n_2276),
.A2(n_2273),
.B1(n_2267),
.B2(n_2270),
.C(n_2266),
.Y(n_2291)
);

NOR3xp33_ASAP7_75t_L g2292 ( 
.A(n_2285),
.B(n_2253),
.C(n_2262),
.Y(n_2292)
);

O2A1O1Ixp33_ASAP7_75t_SL g2293 ( 
.A1(n_2277),
.A2(n_2254),
.B(n_2265),
.C(n_2266),
.Y(n_2293)
);

AOI221xp5_ASAP7_75t_L g2294 ( 
.A1(n_2279),
.A2(n_2275),
.B1(n_2264),
.B2(n_2274),
.C(n_2272),
.Y(n_2294)
);

XNOR2x2_ASAP7_75t_SL g2295 ( 
.A(n_2278),
.B(n_2272),
.Y(n_2295)
);

AOI221xp5_ASAP7_75t_L g2296 ( 
.A1(n_2287),
.A2(n_2156),
.B1(n_2271),
.B2(n_2161),
.C(n_2069),
.Y(n_2296)
);

NOR2x1_ASAP7_75t_L g2297 ( 
.A(n_2280),
.B(n_2156),
.Y(n_2297)
);

OAI22xp33_ASAP7_75t_L g2298 ( 
.A1(n_2290),
.A2(n_2271),
.B1(n_2156),
.B2(n_2006),
.Y(n_2298)
);

AOI221x1_ASAP7_75t_L g2299 ( 
.A1(n_2281),
.A2(n_2039),
.B1(n_2057),
.B2(n_2047),
.C(n_2040),
.Y(n_2299)
);

AOI21xp5_ASAP7_75t_L g2300 ( 
.A1(n_2282),
.A2(n_2043),
.B(n_2064),
.Y(n_2300)
);

AOI21xp5_ASAP7_75t_L g2301 ( 
.A1(n_2288),
.A2(n_2043),
.B(n_2064),
.Y(n_2301)
);

AOI21xp5_ASAP7_75t_L g2302 ( 
.A1(n_2283),
.A2(n_2047),
.B(n_2039),
.Y(n_2302)
);

AOI211xp5_ASAP7_75t_L g2303 ( 
.A1(n_2284),
.A2(n_1986),
.B(n_2074),
.C(n_2073),
.Y(n_2303)
);

NAND4xp25_ASAP7_75t_SL g2304 ( 
.A(n_2289),
.B(n_2052),
.C(n_2032),
.D(n_2037),
.Y(n_2304)
);

INVx1_ASAP7_75t_SL g2305 ( 
.A(n_2286),
.Y(n_2305)
);

AOI222xp33_ASAP7_75t_L g2306 ( 
.A1(n_2286),
.A2(n_2009),
.B1(n_2055),
.B2(n_2058),
.C1(n_2056),
.C2(n_2041),
.Y(n_2306)
);

NOR2x1_ASAP7_75t_SL g2307 ( 
.A(n_2295),
.B(n_2082),
.Y(n_2307)
);

HB1xp67_ASAP7_75t_L g2308 ( 
.A(n_2305),
.Y(n_2308)
);

NAND3xp33_ASAP7_75t_L g2309 ( 
.A(n_2292),
.B(n_2057),
.C(n_2046),
.Y(n_2309)
);

INVx1_ASAP7_75t_SL g2310 ( 
.A(n_2297),
.Y(n_2310)
);

AOI21xp5_ASAP7_75t_L g2311 ( 
.A1(n_2293),
.A2(n_2291),
.B(n_2294),
.Y(n_2311)
);

XOR2xp5_ASAP7_75t_L g2312 ( 
.A(n_2300),
.B(n_1917),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_2299),
.Y(n_2313)
);

NOR2x1p5_ASAP7_75t_L g2314 ( 
.A(n_2304),
.B(n_2077),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2302),
.Y(n_2315)
);

AOI22xp5_ASAP7_75t_L g2316 ( 
.A1(n_2298),
.A2(n_2024),
.B1(n_1994),
.B2(n_2040),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2307),
.Y(n_2317)
);

NOR3xp33_ASAP7_75t_L g2318 ( 
.A(n_2308),
.B(n_2296),
.C(n_2301),
.Y(n_2318)
);

NAND4xp75_ASAP7_75t_L g2319 ( 
.A(n_2311),
.B(n_2315),
.C(n_2313),
.D(n_2316),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_2310),
.B(n_2303),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2309),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2309),
.Y(n_2322)
);

AND2x4_ASAP7_75t_L g2323 ( 
.A(n_2314),
.B(n_2082),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_2312),
.B(n_2306),
.Y(n_2324)
);

OR2x2_ASAP7_75t_L g2325 ( 
.A(n_2323),
.B(n_2317),
.Y(n_2325)
);

NOR2x1p5_ASAP7_75t_L g2326 ( 
.A(n_2319),
.B(n_2077),
.Y(n_2326)
);

AOI21xp5_ASAP7_75t_L g2327 ( 
.A1(n_2321),
.A2(n_2046),
.B(n_2042),
.Y(n_2327)
);

OAI22xp33_ASAP7_75t_L g2328 ( 
.A1(n_2322),
.A2(n_2077),
.B1(n_2042),
.B2(n_2055),
.Y(n_2328)
);

OAI22xp5_ASAP7_75t_L g2329 ( 
.A1(n_2320),
.A2(n_2024),
.B1(n_2032),
.B2(n_2037),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2323),
.B(n_2082),
.Y(n_2330)
);

AOI22xp5_ASAP7_75t_SL g2331 ( 
.A1(n_2324),
.A2(n_2024),
.B1(n_2037),
.B2(n_2052),
.Y(n_2331)
);

OAI222xp33_ASAP7_75t_L g2332 ( 
.A1(n_2318),
.A2(n_2009),
.B1(n_2049),
.B2(n_2068),
.C1(n_2071),
.C2(n_2061),
.Y(n_2332)
);

HB1xp67_ASAP7_75t_L g2333 ( 
.A(n_2326),
.Y(n_2333)
);

NOR3x2_ASAP7_75t_L g2334 ( 
.A(n_2325),
.B(n_1986),
.C(n_1902),
.Y(n_2334)
);

CKINVDCx5p33_ASAP7_75t_R g2335 ( 
.A(n_2331),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2330),
.Y(n_2336)
);

OR2x2_ASAP7_75t_L g2337 ( 
.A(n_2333),
.B(n_2329),
.Y(n_2337)
);

XNOR2xp5_ASAP7_75t_L g2338 ( 
.A(n_2335),
.B(n_2327),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_2338),
.B(n_2335),
.Y(n_2339)
);

AND2x4_ASAP7_75t_L g2340 ( 
.A(n_2337),
.B(n_2336),
.Y(n_2340)
);

INVxp67_ASAP7_75t_L g2341 ( 
.A(n_2340),
.Y(n_2341)
);

AOI22xp5_ASAP7_75t_L g2342 ( 
.A1(n_2339),
.A2(n_2328),
.B1(n_2334),
.B2(n_2332),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2340),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2343),
.Y(n_2344)
);

NAND3xp33_ASAP7_75t_L g2345 ( 
.A(n_2341),
.B(n_2041),
.C(n_2055),
.Y(n_2345)
);

AOI21xp5_ASAP7_75t_L g2346 ( 
.A1(n_2344),
.A2(n_2342),
.B(n_2048),
.Y(n_2346)
);

AOI22xp5_ASAP7_75t_L g2347 ( 
.A1(n_2345),
.A2(n_2071),
.B1(n_2068),
.B2(n_2048),
.Y(n_2347)
);

AOI22xp33_ASAP7_75t_SL g2348 ( 
.A1(n_2346),
.A2(n_1994),
.B1(n_2060),
.B2(n_2051),
.Y(n_2348)
);

AOI221xp5_ASAP7_75t_L g2349 ( 
.A1(n_2348),
.A2(n_2347),
.B1(n_1875),
.B2(n_2015),
.C(n_2068),
.Y(n_2349)
);

AOI211xp5_ASAP7_75t_L g2350 ( 
.A1(n_2349),
.A2(n_2071),
.B(n_1902),
.C(n_2048),
.Y(n_2350)
);


endmodule