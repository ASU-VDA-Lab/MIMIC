module fake_jpeg_28617_n_168 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_168);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_32),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_40),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_19),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_28),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_16),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_27),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_20),
.B(n_1),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_45),
.B(n_30),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_32),
.B1(n_28),
.B2(n_21),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_63),
.B(n_18),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_30),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_35),
.A2(n_36),
.B1(n_34),
.B2(n_33),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_55),
.A2(n_63),
.B1(n_58),
.B2(n_50),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_49),
.B1(n_41),
.B2(n_37),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_57),
.A2(n_43),
.B1(n_39),
.B2(n_22),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_35),
.A2(n_23),
.B1(n_22),
.B2(n_29),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_65),
.A2(n_39),
.B1(n_3),
.B2(n_4),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_70),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_68),
.B(n_15),
.Y(n_75)
);

OR2x2_ASAP7_75t_SL g70 ( 
.A(n_44),
.B(n_47),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_72),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_82),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_67),
.A2(n_38),
.B(n_43),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_74),
.A2(n_89),
.B(n_82),
.C(n_91),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_75),
.B(n_76),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_53),
.B(n_15),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_25),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_78),
.Y(n_93)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_92),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_57),
.A2(n_36),
.B1(n_47),
.B2(n_46),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_41),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_66),
.B(n_25),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_85),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_84),
.B(n_86),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_70),
.B(n_18),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_57),
.A2(n_46),
.B1(n_48),
.B2(n_43),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_69),
.B1(n_5),
.B2(n_51),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_39),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_55),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_2),
.C(n_4),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

OAI22x1_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_59),
.B1(n_92),
.B2(n_79),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_107),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_61),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_104),
.B(n_106),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_61),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_52),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_99),
.B(n_85),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_108),
.B(n_110),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_84),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_109),
.B(n_116),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_101),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_105),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_111),
.B(n_86),
.Y(n_124)
);

OA21x2_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_89),
.B(n_91),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_118),
.B(n_107),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_97),
.A2(n_87),
.B1(n_81),
.B2(n_89),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_97),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_74),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_103),
.A2(n_81),
.B(n_82),
.Y(n_118)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_105),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

AOI221xp5_ASAP7_75t_L g135 ( 
.A1(n_123),
.A2(n_125),
.B1(n_115),
.B2(n_113),
.C(n_117),
.Y(n_135)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_95),
.C(n_102),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_110),
.C(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_120),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_128),
.A2(n_115),
.B1(n_71),
.B2(n_72),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_112),
.B(n_94),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_118),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_137),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_135),
.A2(n_72),
.B1(n_79),
.B2(n_59),
.Y(n_148)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_131),
.A2(n_113),
.B1(n_108),
.B2(n_98),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_138),
.B(n_123),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_94),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_140),
.B(n_141),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_125),
.C(n_129),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_147),
.Y(n_153)
);

AOI211xp5_ASAP7_75t_SL g144 ( 
.A1(n_141),
.A2(n_131),
.B(n_122),
.C(n_83),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_144),
.Y(n_151)
);

AOI322xp5_ASAP7_75t_L g147 ( 
.A1(n_134),
.A2(n_62),
.A3(n_78),
.B1(n_7),
.B2(n_9),
.C1(n_11),
.C2(n_14),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_139),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_132),
.A2(n_62),
.B1(n_60),
.B2(n_11),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_149),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_132),
.C(n_133),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_145),
.C(n_148),
.Y(n_156)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_149),
.Y(n_154)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_154),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_155),
.A2(n_146),
.B1(n_142),
.B2(n_144),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_156),
.B(n_159),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_157),
.A2(n_151),
.B1(n_155),
.B2(n_153),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_6),
.Y(n_159)
);

NAND2xp33_ASAP7_75t_SL g160 ( 
.A(n_158),
.B(n_150),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_161),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_162),
.A2(n_6),
.B(n_12),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_13),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_161),
.C(n_163),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_5),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_5),
.Y(n_168)
);


endmodule