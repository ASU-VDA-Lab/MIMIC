module real_aes_1655_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_449;
wire n_417;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_456;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_L g329 ( .A(n_0), .B(n_239), .Y(n_329) );
AO22x2_ASAP7_75t_L g102 ( .A1(n_1), .A2(n_52), .B1(n_92), .B2(n_103), .Y(n_102) );
AOI22xp33_ASAP7_75t_R g80 ( .A1(n_2), .A2(n_81), .B1(n_177), .B2(n_178), .Y(n_80) );
INVx1_ASAP7_75t_L g177 ( .A(n_2), .Y(n_177) );
INVx1_ASAP7_75t_L g207 ( .A(n_3), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_4), .B(n_228), .Y(n_282) );
NAND2xp33_ASAP7_75t_SL g275 ( .A(n_5), .B(n_234), .Y(n_275) );
INVx1_ASAP7_75t_L g258 ( .A(n_6), .Y(n_258) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_7), .Y(n_159) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_8), .A2(n_22), .B1(n_92), .B2(n_100), .Y(n_99) );
AND2x2_ASAP7_75t_L g280 ( .A(n_9), .B(n_219), .Y(n_280) );
INVx2_ASAP7_75t_L g220 ( .A(n_10), .Y(n_220) );
INVx1_ASAP7_75t_L g104 ( .A(n_11), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_12), .Y(n_153) );
AOI221x1_ASAP7_75t_L g270 ( .A1(n_13), .A2(n_223), .B1(n_271), .B2(n_272), .C(n_274), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_14), .B(n_228), .Y(n_245) );
AOI221xp5_ASAP7_75t_SL g222 ( .A1(n_15), .A2(n_33), .B1(n_223), .B2(n_228), .C(n_235), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_16), .A2(n_223), .B(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_17), .B(n_239), .Y(n_285) );
AOI22xp5_ASAP7_75t_L g190 ( .A1(n_18), .A2(n_64), .B1(n_191), .B2(n_192), .Y(n_190) );
INVx1_ASAP7_75t_L g192 ( .A(n_18), .Y(n_192) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_19), .A2(n_81), .B1(n_178), .B2(n_538), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_19), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g120 ( .A1(n_20), .A2(n_62), .B1(n_121), .B2(n_125), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_21), .Y(n_170) );
OAI221xp5_ASAP7_75t_L g199 ( .A1(n_22), .A2(n_52), .B1(n_54), .B2(n_200), .C(n_202), .Y(n_199) );
OR2x2_ASAP7_75t_L g221 ( .A(n_23), .B(n_69), .Y(n_221) );
OA21x2_ASAP7_75t_L g251 ( .A1(n_23), .A2(n_69), .B(n_220), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_24), .B(n_237), .Y(n_249) );
INVxp67_ASAP7_75t_L g269 ( .A(n_25), .Y(n_269) );
CKINVDCx20_ASAP7_75t_R g141 ( .A(n_26), .Y(n_141) );
AND2x2_ASAP7_75t_L g318 ( .A(n_27), .B(n_218), .Y(n_318) );
INVx3_ASAP7_75t_L g92 ( .A(n_28), .Y(n_92) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_29), .A2(n_223), .B(n_328), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_29), .A2(n_81), .B1(n_178), .B2(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_29), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_30), .B(n_237), .Y(n_236) );
INVx1_ASAP7_75t_SL g93 ( .A(n_31), .Y(n_93) );
INVx1_ASAP7_75t_L g209 ( .A(n_32), .Y(n_209) );
AND2x2_ASAP7_75t_L g224 ( .A(n_32), .B(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g234 ( .A(n_32), .B(n_207), .Y(n_234) );
AOI22xp5_ASAP7_75t_L g302 ( .A1(n_34), .A2(n_60), .B1(n_223), .B2(n_264), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_35), .B(n_239), .Y(n_316) );
AO22x2_ASAP7_75t_L g95 ( .A1(n_36), .A2(n_54), .B1(n_92), .B2(n_96), .Y(n_95) );
AND2x2_ASAP7_75t_L g332 ( .A(n_37), .B(n_218), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_38), .B(n_218), .Y(n_241) );
INVx1_ASAP7_75t_L g227 ( .A(n_39), .Y(n_227) );
INVx1_ASAP7_75t_L g231 ( .A(n_39), .Y(n_231) );
INVx1_ASAP7_75t_L g94 ( .A(n_40), .Y(n_94) );
NAND2xp5_ASAP7_75t_SL g317 ( .A(n_41), .B(n_228), .Y(n_317) );
AND2x2_ASAP7_75t_L g296 ( .A(n_42), .B(n_218), .Y(n_296) );
CKINVDCx20_ASAP7_75t_R g148 ( .A(n_43), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_44), .B(n_237), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_45), .B(n_114), .Y(n_113) );
AND2x2_ASAP7_75t_SL g252 ( .A(n_46), .B(n_219), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_47), .B(n_239), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g313 ( .A1(n_48), .A2(n_223), .B(n_314), .Y(n_313) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_49), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_50), .B(n_237), .Y(n_286) );
AND2x2_ASAP7_75t_SL g303 ( .A(n_51), .B(n_250), .Y(n_303) );
INVxp33_ASAP7_75t_L g204 ( .A(n_52), .Y(n_204) );
INVx1_ASAP7_75t_L g225 ( .A(n_53), .Y(n_225) );
INVx1_ASAP7_75t_L g233 ( .A(n_53), .Y(n_233) );
INVxp67_ASAP7_75t_L g203 ( .A(n_54), .Y(n_203) );
AOI221xp5_ASAP7_75t_L g163 ( .A1(n_55), .A2(n_75), .B1(n_164), .B2(n_166), .C(n_169), .Y(n_163) );
INVx1_ASAP7_75t_L g183 ( .A(n_56), .Y(n_183) );
OAI22x1_ASAP7_75t_R g181 ( .A1(n_57), .A2(n_182), .B1(n_183), .B2(n_184), .Y(n_181) );
INVx1_ASAP7_75t_L g184 ( .A(n_57), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_58), .B(n_228), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g301 ( .A1(n_59), .A2(n_61), .B1(n_228), .B2(n_260), .Y(n_301) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_60), .A2(n_189), .B1(n_190), .B2(n_193), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_60), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g130 ( .A1(n_63), .A2(n_70), .B1(n_131), .B2(n_135), .Y(n_130) );
INVx1_ASAP7_75t_L g191 ( .A(n_64), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_65), .B(n_239), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_66), .B(n_239), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_67), .A2(n_223), .B(n_291), .Y(n_290) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_68), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_71), .B(n_237), .Y(n_292) );
INVxp67_ASAP7_75t_L g187 ( .A(n_72), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_73), .B(n_228), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_74), .B(n_237), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_76), .A2(n_223), .B(n_247), .Y(n_246) );
BUFx2_ASAP7_75t_SL g201 ( .A(n_77), .Y(n_201) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_196), .B1(n_210), .B2(n_525), .C(n_527), .Y(n_78) );
XOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_179), .Y(n_79) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
INVx2_ASAP7_75t_L g178 ( .A(n_82), .Y(n_178) );
AND3x2_ASAP7_75t_L g82 ( .A(n_83), .B(n_139), .C(n_163), .Y(n_82) );
NOR2xp33_ASAP7_75t_L g83 ( .A(n_84), .B(n_119), .Y(n_83) );
OAI221xp5_ASAP7_75t_L g84 ( .A1(n_85), .A2(n_104), .B1(n_105), .B2(n_112), .C(n_113), .Y(n_84) );
INVx1_ASAP7_75t_SL g85 ( .A(n_86), .Y(n_85) );
INVx4_ASAP7_75t_SL g86 ( .A(n_87), .Y(n_86) );
INVx6_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
AND2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_97), .Y(n_88) );
AND2x4_ASAP7_75t_L g127 ( .A(n_89), .B(n_128), .Y(n_127) );
AND2x4_ASAP7_75t_L g137 ( .A(n_89), .B(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g89 ( .A(n_90), .B(n_95), .Y(n_89) );
AND2x2_ASAP7_75t_L g110 ( .A(n_90), .B(n_111), .Y(n_110) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_90), .Y(n_118) );
INVx2_ASAP7_75t_L g134 ( .A(n_90), .Y(n_134) );
OAI22x1_ASAP7_75t_L g90 ( .A1(n_91), .A2(n_92), .B1(n_93), .B2(n_94), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx1_ASAP7_75t_L g96 ( .A(n_92), .Y(n_96) );
INVx2_ASAP7_75t_L g100 ( .A(n_92), .Y(n_100) );
INVx1_ASAP7_75t_L g103 ( .A(n_92), .Y(n_103) );
INVx2_ASAP7_75t_L g111 ( .A(n_95), .Y(n_111) );
AND2x2_ASAP7_75t_L g133 ( .A(n_95), .B(n_134), .Y(n_133) );
BUFx2_ASAP7_75t_L g151 ( .A(n_95), .Y(n_151) );
AND2x4_ASAP7_75t_L g157 ( .A(n_97), .B(n_158), .Y(n_157) );
AND2x2_ASAP7_75t_L g168 ( .A(n_97), .B(n_133), .Y(n_168) );
AND2x4_ASAP7_75t_L g172 ( .A(n_97), .B(n_110), .Y(n_172) );
AND2x4_ASAP7_75t_L g97 ( .A(n_98), .B(n_101), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
AND2x4_ASAP7_75t_L g109 ( .A(n_99), .B(n_101), .Y(n_109) );
AND2x2_ASAP7_75t_L g117 ( .A(n_99), .B(n_102), .Y(n_117) );
INVx1_ASAP7_75t_L g124 ( .A(n_99), .Y(n_124) );
INVxp67_ASAP7_75t_L g138 ( .A(n_101), .Y(n_138) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_L g123 ( .A(n_102), .B(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
BUFx6f_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
BUFx3_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
AND2x4_ASAP7_75t_L g132 ( .A(n_109), .B(n_133), .Y(n_132) );
AND2x4_ASAP7_75t_L g162 ( .A(n_109), .B(n_158), .Y(n_162) );
AND2x2_ASAP7_75t_L g122 ( .A(n_110), .B(n_123), .Y(n_122) );
AND2x4_ASAP7_75t_L g158 ( .A(n_111), .B(n_134), .Y(n_158) );
INVx3_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx3_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
AND2x4_ASAP7_75t_L g150 ( .A(n_117), .B(n_151), .Y(n_150) );
AND2x4_ASAP7_75t_L g165 ( .A(n_117), .B(n_158), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_130), .Y(n_119) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_L g147 ( .A(n_123), .B(n_133), .Y(n_147) );
AND2x4_ASAP7_75t_L g176 ( .A(n_123), .B(n_158), .Y(n_176) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_124), .Y(n_129) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx6_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g139 ( .A(n_140), .B(n_152), .Y(n_139) );
OAI22xp33_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_142), .B1(n_148), .B2(n_149), .Y(n_140) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx5_ASAP7_75t_SL g149 ( .A(n_150), .Y(n_149) );
OAI22xp33_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_154), .B1(n_159), .B2(n_160), .Y(n_152) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx4_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx8_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
BUFx2_ASAP7_75t_SL g164 ( .A(n_165), .Y(n_164) );
BUFx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
BUFx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
OAI22xp5_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B1(n_173), .B2(n_174), .Y(n_169) );
INVx6_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
HB1xp67_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx8_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B1(n_185), .B2(n_195), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g180 ( .A(n_181), .Y(n_180) );
INVx1_ASAP7_75t_SL g182 ( .A(n_183), .Y(n_182) );
CKINVDCx16_ASAP7_75t_R g195 ( .A(n_185), .Y(n_195) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B1(n_188), .B2(n_194), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_187), .B(n_259), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_188), .Y(n_194) );
INVx1_ASAP7_75t_L g193 ( .A(n_190), .Y(n_193) );
INVx1_ASAP7_75t_SL g196 ( .A(n_197), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g197 ( .A(n_198), .Y(n_197) );
AND3x1_ASAP7_75t_SL g198 ( .A(n_199), .B(n_205), .C(n_208), .Y(n_198) );
INVxp67_ASAP7_75t_L g535 ( .A(n_199), .Y(n_535) );
CKINVDCx8_ASAP7_75t_R g200 ( .A(n_201), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
CKINVDCx16_ASAP7_75t_R g533 ( .A(n_205), .Y(n_533) );
OAI21xp5_ASAP7_75t_L g543 ( .A1(n_205), .A2(n_544), .B(n_546), .Y(n_543) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g261 ( .A(n_206), .B(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_SL g541 ( .A(n_206), .B(n_208), .Y(n_541) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g226 ( .A(n_207), .B(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_208), .B(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NOR2x1p5_ASAP7_75t_L g265 ( .A(n_209), .B(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
OR2x6_ASAP7_75t_L g212 ( .A(n_213), .B(n_438), .Y(n_212) );
NAND3xp33_ASAP7_75t_SL g213 ( .A(n_214), .B(n_348), .C(n_388), .Y(n_213) );
O2A1O1Ixp33_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_253), .B(n_277), .C(n_304), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_215), .B(n_353), .Y(n_387) );
NOR2x1p5_ASAP7_75t_L g215 ( .A(n_216), .B(n_242), .Y(n_215) );
BUFx3_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g323 ( .A(n_217), .Y(n_323) );
INVx2_ASAP7_75t_L g339 ( .A(n_217), .Y(n_339) );
OR2x2_ASAP7_75t_L g351 ( .A(n_217), .B(n_243), .Y(n_351) );
AND2x2_ASAP7_75t_L g365 ( .A(n_217), .B(n_324), .Y(n_365) );
INVx1_ASAP7_75t_L g393 ( .A(n_217), .Y(n_393) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_217), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_217), .B(n_243), .Y(n_499) );
OA21x2_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_222), .B(n_241), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_218), .Y(n_295) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_SL g219 ( .A(n_220), .B(n_221), .Y(n_219) );
AND2x4_ASAP7_75t_L g259 ( .A(n_220), .B(n_221), .Y(n_259) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_223), .Y(n_526) );
AND2x6_ASAP7_75t_L g223 ( .A(n_224), .B(n_226), .Y(n_223) );
BUFx3_ASAP7_75t_L g263 ( .A(n_224), .Y(n_263) );
AND2x6_ASAP7_75t_L g239 ( .A(n_225), .B(n_230), .Y(n_239) );
INVx2_ASAP7_75t_L g267 ( .A(n_225), .Y(n_267) );
AND2x4_ASAP7_75t_L g264 ( .A(n_226), .B(n_265), .Y(n_264) );
AND2x4_ASAP7_75t_L g237 ( .A(n_227), .B(n_232), .Y(n_237) );
INVx2_ASAP7_75t_L g262 ( .A(n_227), .Y(n_262) );
AND2x4_ASAP7_75t_L g228 ( .A(n_229), .B(n_234), .Y(n_228) );
INVx1_ASAP7_75t_L g276 ( .A(n_229), .Y(n_276) );
AND2x4_ASAP7_75t_L g229 ( .A(n_230), .B(n_232), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx5_ASAP7_75t_L g240 ( .A(n_234), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_238), .B(n_240), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_240), .A2(n_248), .B(n_249), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_240), .A2(n_285), .B(n_286), .Y(n_284) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_240), .A2(n_292), .B(n_293), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_240), .A2(n_315), .B(n_316), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g328 ( .A1(n_240), .A2(n_329), .B(n_330), .Y(n_328) );
OR2x2_ASAP7_75t_L g320 ( .A(n_242), .B(n_321), .Y(n_320) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_242), .Y(n_455) );
AND2x2_ASAP7_75t_L g460 ( .A(n_242), .B(n_322), .Y(n_460) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x4_ASAP7_75t_L g253 ( .A(n_243), .B(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g319 ( .A(n_243), .B(n_255), .Y(n_319) );
OR2x2_ASAP7_75t_L g338 ( .A(n_243), .B(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g367 ( .A(n_243), .Y(n_367) );
AND2x4_ASAP7_75t_SL g406 ( .A(n_243), .B(n_255), .Y(n_406) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_243), .Y(n_410) );
OR2x2_ASAP7_75t_L g427 ( .A(n_243), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g437 ( .A(n_243), .B(n_344), .Y(n_437) );
INVx1_ASAP7_75t_L g466 ( .A(n_243), .Y(n_466) );
OR2x6_ASAP7_75t_L g243 ( .A(n_244), .B(n_252), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_246), .B(n_250), .Y(n_244) );
INVx2_ASAP7_75t_SL g299 ( .A(n_250), .Y(n_299) );
BUFx4f_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx3_ASAP7_75t_L g273 ( .A(n_251), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_253), .B(n_395), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_254), .B(n_324), .Y(n_341) );
AND2x2_ASAP7_75t_L g353 ( .A(n_254), .B(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g371 ( .A(n_254), .B(n_338), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_254), .B(n_392), .Y(n_391) );
INVx3_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x4_ASAP7_75t_L g344 ( .A(n_255), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g366 ( .A(n_255), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g401 ( .A(n_255), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_255), .B(n_324), .Y(n_425) );
AND2x4_ASAP7_75t_L g255 ( .A(n_256), .B(n_270), .Y(n_255) );
AOI22xp5_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_260), .B1(n_264), .B2(n_268), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_259), .B(n_269), .Y(n_268) );
NOR3xp33_ASAP7_75t_L g274 ( .A(n_259), .B(n_275), .C(n_276), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_259), .A2(n_282), .B(n_283), .Y(n_281) );
AND2x4_ASAP7_75t_L g260 ( .A(n_261), .B(n_263), .Y(n_260) );
INVx1_ASAP7_75t_L g546 ( .A(n_261), .Y(n_546) );
INVx1_ASAP7_75t_L g545 ( .A(n_263), .Y(n_545) );
INVx3_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx4_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AOI21x1_ASAP7_75t_L g325 ( .A1(n_273), .A2(n_326), .B(n_332), .Y(n_325) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_287), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_278), .B(n_357), .Y(n_356) );
AND2x4_ASAP7_75t_L g374 ( .A(n_278), .B(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_278), .B(n_288), .Y(n_379) );
NAND3xp33_ASAP7_75t_L g394 ( .A(n_278), .B(n_395), .C(n_396), .Y(n_394) );
AND2x2_ASAP7_75t_L g442 ( .A(n_278), .B(n_347), .Y(n_442) );
INVx5_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g309 ( .A(n_279), .B(n_310), .Y(n_309) );
AND2x4_ASAP7_75t_SL g346 ( .A(n_279), .B(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g362 ( .A(n_279), .Y(n_362) );
OR2x2_ASAP7_75t_L g385 ( .A(n_279), .B(n_375), .Y(n_385) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_279), .Y(n_402) );
AND2x2_ASAP7_75t_SL g420 ( .A(n_279), .B(n_308), .Y(n_420) );
AND2x4_ASAP7_75t_L g435 ( .A(n_279), .B(n_311), .Y(n_435) );
AND2x2_ASAP7_75t_L g449 ( .A(n_279), .B(n_288), .Y(n_449) );
OR2x2_ASAP7_75t_L g470 ( .A(n_279), .B(n_297), .Y(n_470) );
OR2x6_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
AND2x2_ASAP7_75t_L g524 ( .A(n_287), .B(n_402), .Y(n_524) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_297), .Y(n_287) );
AND2x4_ASAP7_75t_L g347 ( .A(n_288), .B(n_310), .Y(n_347) );
INVx2_ASAP7_75t_L g358 ( .A(n_288), .Y(n_358) );
AND2x2_ASAP7_75t_L g363 ( .A(n_288), .B(n_308), .Y(n_363) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_288), .Y(n_396) );
OR2x2_ASAP7_75t_L g419 ( .A(n_288), .B(n_311), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_288), .B(n_311), .Y(n_422) );
INVx1_ASAP7_75t_L g431 ( .A(n_288), .Y(n_431) );
AO21x2_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_295), .B(n_296), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_294), .Y(n_289) );
AO21x2_ASAP7_75t_L g311 ( .A1(n_295), .A2(n_312), .B(n_318), .Y(n_311) );
AO21x2_ASAP7_75t_L g375 ( .A1(n_295), .A2(n_312), .B(n_318), .Y(n_375) );
AND2x2_ASAP7_75t_L g334 ( .A(n_297), .B(n_311), .Y(n_334) );
BUFx2_ASAP7_75t_L g383 ( .A(n_297), .Y(n_383) );
AND2x2_ASAP7_75t_L g478 ( .A(n_297), .B(n_358), .Y(n_478) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_298), .Y(n_308) );
AOI21x1_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_300), .B(n_303), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
OAI221xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_319), .B1(n_320), .B2(n_333), .C(n_335), .Y(n_304) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
NOR2x1_ASAP7_75t_L g380 ( .A(n_307), .B(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_307), .B(n_374), .Y(n_414) );
OR2x2_ASAP7_75t_L g426 ( .A(n_307), .B(n_422), .Y(n_426) );
OR2x2_ASAP7_75t_L g429 ( .A(n_307), .B(n_430), .Y(n_429) );
OR2x2_ASAP7_75t_L g518 ( .A(n_307), .B(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x4_ASAP7_75t_L g357 ( .A(n_308), .B(n_358), .Y(n_357) );
OA33x2_ASAP7_75t_L g390 ( .A1(n_308), .A2(n_351), .A3(n_391), .B1(n_394), .B2(n_397), .B3(n_400), .Y(n_390) );
OR2x2_ASAP7_75t_L g421 ( .A(n_308), .B(n_422), .Y(n_421) );
OR2x2_ASAP7_75t_L g445 ( .A(n_308), .B(n_446), .Y(n_445) );
OR2x2_ASAP7_75t_L g453 ( .A(n_308), .B(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g473 ( .A(n_308), .B(n_347), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_308), .B(n_362), .Y(n_511) );
INVx2_ASAP7_75t_L g381 ( .A(n_309), .Y(n_381) );
AOI322xp5_ASAP7_75t_L g451 ( .A1(n_309), .A2(n_364), .A3(n_452), .B1(n_455), .B2(n_456), .C1(n_458), .C2(n_460), .Y(n_451) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_311), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_317), .Y(n_312) );
OR2x2_ASAP7_75t_L g433 ( .A(n_319), .B(n_412), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_319), .B(n_486), .Y(n_485) );
INVx1_ASAP7_75t_SL g506 ( .A(n_319), .Y(n_506) );
INVx1_ASAP7_75t_SL g372 ( .A(n_320), .Y(n_372) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g405 ( .A(n_322), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx2_ASAP7_75t_L g345 ( .A(n_324), .Y(n_345) );
INVx1_ASAP7_75t_L g354 ( .A(n_324), .Y(n_354) );
INVx1_ASAP7_75t_L g395 ( .A(n_324), .Y(n_395) );
OR2x2_ASAP7_75t_L g412 ( .A(n_324), .B(n_339), .Y(n_412) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_324), .Y(n_487) );
INVx3_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_331), .Y(n_326) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_SL g456 ( .A(n_334), .B(n_457), .Y(n_456) );
OAI21xp5_ASAP7_75t_SL g335 ( .A1(n_336), .A2(n_342), .B(n_346), .Y(n_335) );
A2O1A1Ixp33_ASAP7_75t_L g409 ( .A1(n_336), .A2(n_410), .B(n_411), .C(n_413), .Y(n_409) );
AND2x4_ASAP7_75t_L g336 ( .A(n_337), .B(n_340), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g474 ( .A(n_338), .B(n_475), .Y(n_474) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_339), .Y(n_343) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g498 ( .A(n_341), .B(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
AND2x2_ASAP7_75t_SL g467 ( .A(n_344), .B(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g475 ( .A(n_344), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_344), .B(n_466), .Y(n_483) );
INVx3_ASAP7_75t_SL g408 ( .A(n_347), .Y(n_408) );
AOI221xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_355), .B1(n_359), .B2(n_364), .C(n_368), .Y(n_348) );
INVx1_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_354), .Y(n_399) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_357), .A2(n_384), .B(n_456), .Y(n_462) );
AND2x2_ASAP7_75t_L g488 ( .A(n_357), .B(n_435), .Y(n_488) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_358), .Y(n_376) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_363), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_362), .B(n_478), .Y(n_477) );
OR2x2_ASAP7_75t_L g497 ( .A(n_362), .B(n_419), .Y(n_497) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
INVx2_ASAP7_75t_L g446 ( .A(n_365), .Y(n_446) );
OAI21xp33_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_373), .B(n_377), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_370), .B(n_372), .Y(n_369) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_376), .Y(n_373) );
INVx2_ASAP7_75t_L g519 ( .A(n_374), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_375), .B(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g448 ( .A(n_375), .B(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_376), .B(n_398), .Y(n_397) );
OAI31xp33_ASAP7_75t_SL g377 ( .A1(n_378), .A2(n_380), .A3(n_382), .B(n_386), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_381), .B(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
OR2x2_ASAP7_75t_L g459 ( .A(n_383), .B(n_385), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_383), .B(n_435), .Y(n_514) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NOR5xp2_ASAP7_75t_L g388 ( .A(n_389), .B(n_403), .C(n_415), .D(n_424), .E(n_432), .Y(n_388) );
INVxp67_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_393), .B(n_395), .Y(n_428) );
INVx1_ASAP7_75t_L g468 ( .A(n_393), .Y(n_468) );
INVxp67_ASAP7_75t_SL g505 ( .A(n_393), .Y(n_505) );
INVx1_ASAP7_75t_L g457 ( .A(n_396), .Y(n_457) );
INVxp67_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NAND2xp33_ASAP7_75t_SL g400 ( .A(n_401), .B(n_402), .Y(n_400) );
OAI321xp33_ASAP7_75t_L g440 ( .A1(n_401), .A2(n_441), .A3(n_443), .B1(n_447), .B2(n_450), .C(n_451), .Y(n_440) );
INVx1_ASAP7_75t_L g494 ( .A(n_402), .Y(n_494) );
OAI21xp33_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_407), .B(n_409), .Y(n_403) );
INVx1_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_405), .A2(n_478), .B1(n_485), .B2(n_488), .Y(n_484) );
AND2x2_ASAP7_75t_L g513 ( .A(n_406), .B(n_487), .Y(n_513) );
INVx1_ASAP7_75t_L g423 ( .A(n_411), .Y(n_423) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AOI21xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_421), .B(n_423), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_420), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_422), .A2(n_433), .B1(n_434), .B2(n_436), .Y(n_432) );
INVx1_ASAP7_75t_L g495 ( .A(n_422), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_426), .B1(n_427), .B2(n_429), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_431), .B(n_435), .Y(n_434) );
OAI221xp5_ASAP7_75t_L g509 ( .A1(n_433), .A2(n_510), .B1(n_512), .B2(n_514), .C(n_515), .Y(n_509) );
INVx1_ASAP7_75t_L g516 ( .A(n_433), .Y(n_516) );
OAI221xp5_ASAP7_75t_L g490 ( .A1(n_434), .A2(n_491), .B1(n_498), .B2(n_500), .C(n_501), .Y(n_490) );
OAI21xp5_ASAP7_75t_L g461 ( .A1(n_436), .A2(n_462), .B(n_463), .Y(n_461) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_439), .B(n_489), .Y(n_438) );
NOR3xp33_ASAP7_75t_L g439 ( .A(n_440), .B(n_461), .C(n_479), .Y(n_439) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_442), .Y(n_508) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx3_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g507 ( .A(n_450), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_452), .B(n_482), .Y(n_481) );
INVx1_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g500 ( .A(n_460), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_469), .B(n_471), .Y(n_463) );
INVxp67_ASAP7_75t_L g521 ( .A(n_464), .Y(n_521) );
AND2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_467), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_SL g476 ( .A(n_467), .Y(n_476) );
INVx1_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
OAI22xp33_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_474), .B1(n_476), .B2(n_477), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
OAI21xp33_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B(n_484), .Y(n_479) );
INVx1_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g522 ( .A(n_485), .Y(n_522) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NOR3xp33_ASAP7_75t_L g489 ( .A(n_490), .B(n_509), .C(n_520), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_492), .B(n_496), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_494), .B(n_495), .Y(n_493) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
OAI21xp5_ASAP7_75t_SL g501 ( .A1(n_502), .A2(n_507), .B(n_508), .Y(n_501) );
INVx1_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_506), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVxp67_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g515 ( .A1(n_513), .A2(n_516), .B(n_517), .Y(n_515) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AOI21xp33_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_522), .B(n_523), .Y(n_520) );
INVx1_ASAP7_75t_SL g523 ( .A(n_524), .Y(n_523) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OAI222xp33_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_529), .B1(n_530), .B2(n_536), .C1(n_539), .C2(n_542), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_531), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_532), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
CKINVDCx16_ASAP7_75t_R g536 ( .A(n_537), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_543), .Y(n_542) );
INVxp67_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
endmodule