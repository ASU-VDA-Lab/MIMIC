module real_aes_8361_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_502;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g245 ( .A1(n_0), .A2(n_246), .B(n_247), .C(n_251), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_1), .B(n_187), .Y(n_252) );
INVx1_ASAP7_75t_L g113 ( .A(n_2), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_3), .B(n_159), .Y(n_235) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_4), .A2(n_145), .B(n_150), .C(n_516), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_5), .A2(n_140), .B(n_554), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_6), .A2(n_140), .B(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_7), .B(n_187), .Y(n_560) );
AO21x2_ASAP7_75t_L g190 ( .A1(n_8), .A2(n_175), .B(n_191), .Y(n_190) );
AND2x6_ASAP7_75t_L g145 ( .A(n_9), .B(n_146), .Y(n_145) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_10), .A2(n_145), .B(n_150), .C(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g498 ( .A(n_11), .Y(n_498) );
INVx1_ASAP7_75t_L g110 ( .A(n_12), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_12), .B(n_41), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_13), .B(n_250), .Y(n_518) );
INVx1_ASAP7_75t_L g169 ( .A(n_14), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_15), .B(n_159), .Y(n_197) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_16), .A2(n_160), .B(n_506), .C(n_508), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_17), .B(n_187), .Y(n_509) );
AOI22xp5_ASAP7_75t_SL g473 ( .A1(n_18), .A2(n_467), .B1(n_474), .B2(n_755), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g126 ( .A1(n_19), .A2(n_47), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_19), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_19), .B(n_224), .Y(n_597) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_20), .A2(n_150), .B(n_201), .C(n_220), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_21), .A2(n_199), .B(n_249), .C(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_22), .B(n_250), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_23), .B(n_250), .Y(n_538) );
CKINVDCx16_ASAP7_75t_R g545 ( .A(n_24), .Y(n_545) );
INVx1_ASAP7_75t_L g537 ( .A(n_25), .Y(n_537) );
A2O1A1Ixp33_ASAP7_75t_L g193 ( .A1(n_26), .A2(n_150), .B(n_194), .C(n_201), .Y(n_193) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_27), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_28), .Y(n_514) );
INVx1_ASAP7_75t_L g594 ( .A(n_29), .Y(n_594) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_30), .A2(n_140), .B(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g143 ( .A(n_31), .Y(n_143) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_32), .A2(n_148), .B(n_163), .C(n_209), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_33), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_L g556 ( .A1(n_34), .A2(n_249), .B(n_557), .C(n_559), .Y(n_556) );
INVxp67_ASAP7_75t_L g595 ( .A(n_35), .Y(n_595) );
OAI22xp5_ASAP7_75t_SL g130 ( .A1(n_36), .A2(n_46), .B1(n_131), .B2(n_132), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_36), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_37), .B(n_196), .Y(n_195) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_38), .A2(n_150), .B(n_201), .C(n_536), .Y(n_535) );
CKINVDCx14_ASAP7_75t_R g555 ( .A(n_39), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g480 ( .A1(n_40), .A2(n_45), .B1(n_481), .B2(n_482), .Y(n_480) );
INVx1_ASAP7_75t_L g482 ( .A(n_40), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_41), .B(n_110), .Y(n_109) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_42), .A2(n_251), .B(n_496), .C(n_497), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_43), .B(n_218), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g265 ( .A(n_44), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_45), .Y(n_481) );
INVx1_ASAP7_75t_L g132 ( .A(n_46), .Y(n_132) );
INVx1_ASAP7_75t_L g128 ( .A(n_47), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_48), .B(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_49), .B(n_140), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_50), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g591 ( .A(n_51), .Y(n_591) );
A2O1A1Ixp33_ASAP7_75t_L g147 ( .A1(n_52), .A2(n_148), .B(n_153), .C(n_163), .Y(n_147) );
INVx1_ASAP7_75t_L g248 ( .A(n_53), .Y(n_248) );
INVx1_ASAP7_75t_L g154 ( .A(n_54), .Y(n_154) );
INVx1_ASAP7_75t_L g526 ( .A(n_55), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_56), .B(n_140), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_57), .Y(n_227) );
CKINVDCx14_ASAP7_75t_R g494 ( .A(n_58), .Y(n_494) );
INVx1_ASAP7_75t_L g146 ( .A(n_59), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_60), .B(n_140), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_61), .B(n_187), .Y(n_186) );
A2O1A1Ixp33_ASAP7_75t_L g180 ( .A1(n_62), .A2(n_181), .B(n_183), .C(n_185), .Y(n_180) );
INVx1_ASAP7_75t_L g168 ( .A(n_63), .Y(n_168) );
INVx1_ASAP7_75t_SL g558 ( .A(n_64), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_65), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_66), .B(n_159), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_67), .B(n_187), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_68), .B(n_160), .Y(n_262) );
INVx1_ASAP7_75t_L g548 ( .A(n_69), .Y(n_548) );
CKINVDCx16_ASAP7_75t_R g244 ( .A(n_70), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_71), .B(n_156), .Y(n_221) );
A2O1A1Ixp33_ASAP7_75t_L g232 ( .A1(n_72), .A2(n_150), .B(n_163), .C(n_233), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_73), .A2(n_105), .B1(n_118), .B2(n_760), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g179 ( .A(n_74), .Y(n_179) );
INVx1_ASAP7_75t_L g117 ( .A(n_75), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_76), .A2(n_140), .B(n_493), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_77), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_78), .A2(n_140), .B(n_503), .Y(n_502) );
OAI22xp5_ASAP7_75t_SL g475 ( .A1(n_79), .A2(n_476), .B1(n_477), .B2(n_483), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_79), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_80), .A2(n_218), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g504 ( .A(n_81), .Y(n_504) );
CKINVDCx16_ASAP7_75t_R g534 ( .A(n_82), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_83), .B(n_155), .Y(n_222) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_84), .A2(n_478), .B1(n_479), .B2(n_480), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_84), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_85), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_86), .A2(n_140), .B(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g507 ( .A(n_87), .Y(n_507) );
INVx2_ASAP7_75t_L g166 ( .A(n_88), .Y(n_166) );
INVx1_ASAP7_75t_L g517 ( .A(n_89), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_90), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_91), .B(n_250), .Y(n_263) );
INVx2_ASAP7_75t_L g114 ( .A(n_92), .Y(n_114) );
OR2x2_ASAP7_75t_L g466 ( .A(n_92), .B(n_467), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_L g546 ( .A1(n_93), .A2(n_150), .B(n_163), .C(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_94), .B(n_140), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_95), .B(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g210 ( .A(n_96), .Y(n_210) );
INVxp67_ASAP7_75t_L g184 ( .A(n_97), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_98), .B(n_175), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_99), .B(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g234 ( .A(n_100), .Y(n_234) );
INVx1_ASAP7_75t_L g258 ( .A(n_101), .Y(n_258) );
INVx2_ASAP7_75t_L g529 ( .A(n_102), .Y(n_529) );
AND2x2_ASAP7_75t_L g170 ( .A(n_103), .B(n_165), .Y(n_170) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g761 ( .A(n_106), .Y(n_761) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_111), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
CKINVDCx14_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
NAND3xp33_ASAP7_75t_SL g112 ( .A(n_113), .B(n_114), .C(n_115), .Y(n_112) );
AND2x2_ASAP7_75t_L g468 ( .A(n_113), .B(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g485 ( .A(n_114), .Y(n_485) );
INVx1_ASAP7_75t_L g754 ( .A(n_114), .Y(n_754) );
NOR2x2_ASAP7_75t_L g757 ( .A(n_114), .B(n_467), .Y(n_757) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
OA21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_124), .B(n_472), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
BUFx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_SL g759 ( .A(n_122), .Y(n_759) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI21xp5_ASAP7_75t_SL g124 ( .A1(n_125), .A2(n_463), .B(n_470), .Y(n_124) );
XNOR2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_129), .Y(n_125) );
XOR2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_133), .Y(n_129) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_133), .A2(n_485), .B1(n_486), .B2(n_753), .Y(n_484) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OR5x1_ASAP7_75t_L g134 ( .A(n_135), .B(n_336), .C(n_414), .D(n_438), .E(n_455), .Y(n_134) );
OAI211xp5_ASAP7_75t_SL g135 ( .A1(n_136), .A2(n_202), .B(n_253), .C(n_313), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_171), .Y(n_136) );
AND2x2_ASAP7_75t_L g267 ( .A(n_137), .B(n_173), .Y(n_267) );
INVx5_ASAP7_75t_SL g295 ( .A(n_137), .Y(n_295) );
AND2x2_ASAP7_75t_L g331 ( .A(n_137), .B(n_316), .Y(n_331) );
OR2x2_ASAP7_75t_L g370 ( .A(n_137), .B(n_172), .Y(n_370) );
OR2x2_ASAP7_75t_L g401 ( .A(n_137), .B(n_292), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_137), .B(n_305), .Y(n_437) );
AND2x2_ASAP7_75t_L g449 ( .A(n_137), .B(n_292), .Y(n_449) );
OR2x6_ASAP7_75t_L g137 ( .A(n_138), .B(n_170), .Y(n_137) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_147), .B(n_165), .Y(n_138) );
BUFx2_ASAP7_75t_L g218 ( .A(n_140), .Y(n_218) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_145), .Y(n_140) );
NAND2x1p5_ASAP7_75t_L g259 ( .A(n_141), .B(n_145), .Y(n_259) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
INVx1_ASAP7_75t_L g185 ( .A(n_142), .Y(n_185) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g151 ( .A(n_143), .Y(n_151) );
INVx1_ASAP7_75t_L g200 ( .A(n_143), .Y(n_200) );
INVx1_ASAP7_75t_L g152 ( .A(n_144), .Y(n_152) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_144), .Y(n_157) );
INVx3_ASAP7_75t_L g160 ( .A(n_144), .Y(n_160) );
INVx1_ASAP7_75t_L g196 ( .A(n_144), .Y(n_196) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_144), .Y(n_250) );
INVx4_ASAP7_75t_SL g164 ( .A(n_145), .Y(n_164) );
BUFx3_ASAP7_75t_L g201 ( .A(n_145), .Y(n_201) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
O2A1O1Ixp33_ASAP7_75t_L g178 ( .A1(n_149), .A2(n_164), .B(n_179), .C(n_180), .Y(n_178) );
O2A1O1Ixp33_ASAP7_75t_SL g243 ( .A1(n_149), .A2(n_164), .B(n_244), .C(n_245), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_SL g493 ( .A1(n_149), .A2(n_164), .B(n_494), .C(n_495), .Y(n_493) );
O2A1O1Ixp33_ASAP7_75t_SL g503 ( .A1(n_149), .A2(n_164), .B(n_504), .C(n_505), .Y(n_503) );
O2A1O1Ixp33_ASAP7_75t_SL g525 ( .A1(n_149), .A2(n_164), .B(n_526), .C(n_527), .Y(n_525) );
O2A1O1Ixp33_ASAP7_75t_L g554 ( .A1(n_149), .A2(n_164), .B(n_555), .C(n_556), .Y(n_554) );
O2A1O1Ixp33_ASAP7_75t_SL g590 ( .A1(n_149), .A2(n_164), .B(n_591), .C(n_592), .Y(n_590) );
INVx5_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x6_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
BUFx3_ASAP7_75t_L g162 ( .A(n_151), .Y(n_162) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_151), .Y(n_237) );
O2A1O1Ixp33_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_155), .B(n_158), .C(n_161), .Y(n_153) );
O2A1O1Ixp33_ASAP7_75t_L g209 ( .A1(n_155), .A2(n_161), .B(n_210), .C(n_211), .Y(n_209) );
O2A1O1Ixp5_ASAP7_75t_L g516 ( .A1(n_155), .A2(n_517), .B(n_518), .C(n_519), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_L g547 ( .A1(n_155), .A2(n_519), .B(n_548), .C(n_549), .Y(n_547) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx4_ASAP7_75t_L g182 ( .A(n_157), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_159), .B(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g246 ( .A(n_159), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_L g536 ( .A1(n_159), .A2(n_223), .B(n_537), .C(n_538), .Y(n_536) );
OAI22xp33_ASAP7_75t_L g593 ( .A1(n_159), .A2(n_182), .B1(n_594), .B2(n_595), .Y(n_593) );
INVx5_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_160), .B(n_498), .Y(n_497) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g251 ( .A(n_162), .Y(n_251) );
INVx1_ASAP7_75t_L g508 ( .A(n_162), .Y(n_508) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_165), .A2(n_207), .B(n_208), .Y(n_206) );
INVx2_ASAP7_75t_L g225 ( .A(n_165), .Y(n_225) );
INVx1_ASAP7_75t_L g228 ( .A(n_165), .Y(n_228) );
OA21x2_ASAP7_75t_L g491 ( .A1(n_165), .A2(n_492), .B(n_499), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_L g533 ( .A1(n_165), .A2(n_259), .B(n_534), .C(n_535), .Y(n_533) );
AND2x2_ASAP7_75t_SL g165 ( .A(n_166), .B(n_167), .Y(n_165) );
AND2x2_ASAP7_75t_L g176 ( .A(n_166), .B(n_167), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
AND2x2_ASAP7_75t_L g448 ( .A(n_171), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_SL g171 ( .A(n_172), .Y(n_171) );
OR2x2_ASAP7_75t_L g311 ( .A(n_172), .B(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g172 ( .A(n_173), .B(n_189), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_173), .B(n_292), .Y(n_291) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_173), .Y(n_304) );
INVx3_ASAP7_75t_L g319 ( .A(n_173), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_173), .B(n_189), .Y(n_343) );
OR2x2_ASAP7_75t_L g352 ( .A(n_173), .B(n_295), .Y(n_352) );
AND2x2_ASAP7_75t_L g356 ( .A(n_173), .B(n_316), .Y(n_356) );
AND2x2_ASAP7_75t_L g362 ( .A(n_173), .B(n_363), .Y(n_362) );
INVxp67_ASAP7_75t_L g399 ( .A(n_173), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_173), .B(n_256), .Y(n_413) );
OA21x2_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_177), .B(n_186), .Y(n_173) );
OA21x2_ASAP7_75t_L g501 ( .A1(n_174), .A2(n_502), .B(n_509), .Y(n_501) );
OA21x2_ASAP7_75t_L g523 ( .A1(n_174), .A2(n_524), .B(n_530), .Y(n_523) );
OA21x2_ASAP7_75t_L g552 ( .A1(n_174), .A2(n_553), .B(n_560), .Y(n_552) );
HB1xp67_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx4_ASAP7_75t_L g188 ( .A(n_175), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_175), .A2(n_192), .B(n_193), .Y(n_191) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g266 ( .A(n_176), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_L g233 ( .A1(n_181), .A2(n_234), .B(n_235), .C(n_236), .Y(n_233) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_182), .B(n_507), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_182), .B(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g223 ( .A(n_185), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_185), .B(n_593), .Y(n_592) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_187), .A2(n_242), .B(n_252), .Y(n_241) );
INVx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_188), .B(n_213), .Y(n_212) );
AO21x2_ASAP7_75t_L g230 ( .A1(n_188), .A2(n_231), .B(n_239), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_188), .B(n_240), .Y(n_239) );
AO21x2_ASAP7_75t_L g256 ( .A1(n_188), .A2(n_257), .B(n_264), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_188), .B(n_521), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_188), .B(n_540), .Y(n_539) );
AO21x2_ASAP7_75t_L g543 ( .A1(n_188), .A2(n_544), .B(n_550), .Y(n_543) );
OR2x2_ASAP7_75t_L g305 ( .A(n_189), .B(n_256), .Y(n_305) );
AND2x2_ASAP7_75t_L g316 ( .A(n_189), .B(n_292), .Y(n_316) );
AND2x2_ASAP7_75t_L g328 ( .A(n_189), .B(n_319), .Y(n_328) );
NAND2xp5_ASAP7_75t_SL g351 ( .A(n_189), .B(n_256), .Y(n_351) );
INVx1_ASAP7_75t_SL g363 ( .A(n_189), .Y(n_363) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AND2x2_ASAP7_75t_L g255 ( .A(n_190), .B(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_190), .B(n_295), .Y(n_294) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_197), .B(n_198), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_198), .A2(n_262), .B(n_263), .Y(n_261) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx3_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_214), .Y(n_203) );
AND2x2_ASAP7_75t_L g276 ( .A(n_204), .B(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_204), .B(n_229), .Y(n_280) );
AND2x2_ASAP7_75t_L g283 ( .A(n_204), .B(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_204), .B(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g308 ( .A(n_204), .B(n_299), .Y(n_308) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_204), .Y(n_327) );
AND2x2_ASAP7_75t_L g348 ( .A(n_204), .B(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g358 ( .A(n_204), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g404 ( .A(n_204), .B(n_287), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_204), .B(n_310), .Y(n_431) );
INVx5_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
BUFx2_ASAP7_75t_L g301 ( .A(n_205), .Y(n_301) );
AND2x2_ASAP7_75t_L g367 ( .A(n_205), .B(n_299), .Y(n_367) );
AND2x2_ASAP7_75t_L g451 ( .A(n_205), .B(n_319), .Y(n_451) );
OR2x6_ASAP7_75t_L g205 ( .A(n_206), .B(n_212), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_214), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g440 ( .A(n_214), .Y(n_440) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_229), .Y(n_214) );
AND2x2_ASAP7_75t_L g270 ( .A(n_215), .B(n_271), .Y(n_270) );
AND2x4_ASAP7_75t_L g279 ( .A(n_215), .B(n_277), .Y(n_279) );
INVx5_ASAP7_75t_L g287 ( .A(n_215), .Y(n_287) );
AND2x2_ASAP7_75t_L g310 ( .A(n_215), .B(n_241), .Y(n_310) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_215), .Y(n_347) );
OR2x6_ASAP7_75t_L g215 ( .A(n_216), .B(n_226), .Y(n_215) );
AOI21xp5_ASAP7_75t_SL g216 ( .A1(n_217), .A2(n_219), .B(n_224), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_223), .Y(n_220) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_225), .B(n_551), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_227), .B(n_228), .Y(n_226) );
AO21x2_ASAP7_75t_L g512 ( .A1(n_228), .A2(n_513), .B(n_520), .Y(n_512) );
INVx1_ASAP7_75t_L g388 ( .A(n_229), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_229), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g421 ( .A(n_229), .B(n_287), .Y(n_421) );
A2O1A1Ixp33_ASAP7_75t_L g450 ( .A1(n_229), .A2(n_344), .B(n_451), .C(n_452), .Y(n_450) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_241), .Y(n_229) );
BUFx2_ASAP7_75t_L g271 ( .A(n_230), .Y(n_271) );
INVx2_ASAP7_75t_L g275 ( .A(n_230), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_232), .B(n_238), .Y(n_231) );
HB1xp67_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx3_ASAP7_75t_L g559 ( .A(n_237), .Y(n_559) );
INVx2_ASAP7_75t_L g277 ( .A(n_241), .Y(n_277) );
AND2x2_ASAP7_75t_L g284 ( .A(n_241), .B(n_275), .Y(n_284) );
AND2x2_ASAP7_75t_L g375 ( .A(n_241), .B(n_287), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_249), .B(n_558), .Y(n_557) );
INVx4_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g496 ( .A(n_250), .Y(n_496) );
INVx2_ASAP7_75t_L g519 ( .A(n_251), .Y(n_519) );
AOI211x1_ASAP7_75t_SL g253 ( .A1(n_254), .A2(n_268), .B(n_281), .C(n_306), .Y(n_253) );
INVx1_ASAP7_75t_L g372 ( .A(n_254), .Y(n_372) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_267), .Y(n_254) );
INVx5_ASAP7_75t_SL g292 ( .A(n_256), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_256), .B(n_362), .Y(n_361) );
AOI311xp33_ASAP7_75t_L g380 ( .A1(n_256), .A2(n_381), .A3(n_383), .B(n_384), .C(n_390), .Y(n_380) );
A2O1A1Ixp33_ASAP7_75t_L g415 ( .A1(n_256), .A2(n_328), .B(n_416), .C(n_419), .Y(n_415) );
OAI21xp5_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_259), .B(n_260), .Y(n_257) );
OAI21xp5_ASAP7_75t_L g513 ( .A1(n_259), .A2(n_514), .B(n_515), .Y(n_513) );
OAI21xp5_ASAP7_75t_L g544 ( .A1(n_259), .A2(n_545), .B(n_546), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g587 ( .A(n_266), .Y(n_587) );
INVxp67_ASAP7_75t_L g335 ( .A(n_267), .Y(n_335) );
NAND4xp25_ASAP7_75t_SL g268 ( .A(n_269), .B(n_272), .C(n_278), .D(n_280), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_269), .B(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g326 ( .A(n_270), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_276), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_273), .B(n_279), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_273), .B(n_286), .Y(n_406) );
BUFx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_274), .B(n_287), .Y(n_424) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g299 ( .A(n_275), .Y(n_299) );
INVxp67_ASAP7_75t_L g334 ( .A(n_276), .Y(n_334) );
AND2x4_ASAP7_75t_L g286 ( .A(n_277), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g360 ( .A(n_277), .B(n_299), .Y(n_360) );
INVx1_ASAP7_75t_L g387 ( .A(n_277), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_277), .B(n_374), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_278), .B(n_348), .Y(n_368) );
INVx1_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_279), .B(n_301), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_279), .B(n_348), .Y(n_447) );
INVx1_ASAP7_75t_L g458 ( .A(n_280), .Y(n_458) );
A2O1A1Ixp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_285), .B(n_288), .C(n_296), .Y(n_281) );
INVx1_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g300 ( .A(n_284), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g338 ( .A(n_284), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g320 ( .A(n_285), .Y(n_320) );
AND2x2_ASAP7_75t_L g297 ( .A(n_286), .B(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_286), .B(n_348), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_286), .B(n_367), .Y(n_391) );
OR2x2_ASAP7_75t_L g307 ( .A(n_287), .B(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g339 ( .A(n_287), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_287), .B(n_299), .Y(n_354) );
AND2x2_ASAP7_75t_L g411 ( .A(n_287), .B(n_367), .Y(n_411) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_287), .Y(n_418) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AOI221xp5_ASAP7_75t_L g422 ( .A1(n_289), .A2(n_301), .B1(n_423), .B2(n_425), .C(n_428), .Y(n_422) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_293), .Y(n_289) );
INVx1_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g312 ( .A(n_292), .B(n_295), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_292), .B(n_362), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_292), .B(n_319), .Y(n_427) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g412 ( .A(n_294), .B(n_413), .Y(n_412) );
OR2x2_ASAP7_75t_L g426 ( .A(n_294), .B(n_427), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_295), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g323 ( .A(n_295), .B(n_316), .Y(n_323) );
AND2x2_ASAP7_75t_L g393 ( .A(n_295), .B(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_295), .B(n_342), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_295), .B(n_443), .Y(n_442) );
OAI21xp5_ASAP7_75t_SL g296 ( .A1(n_297), .A2(n_300), .B(n_302), .Y(n_296) );
INVx2_ASAP7_75t_L g329 ( .A(n_297), .Y(n_329) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g349 ( .A(n_299), .Y(n_349) );
OR2x2_ASAP7_75t_L g353 ( .A(n_301), .B(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g456 ( .A(n_301), .B(n_424), .Y(n_456) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
AOI21xp33_ASAP7_75t_SL g306 ( .A1(n_307), .A2(n_309), .B(n_311), .Y(n_306) );
INVx1_ASAP7_75t_L g460 ( .A(n_307), .Y(n_460) );
INVx2_ASAP7_75t_SL g374 ( .A(n_308), .Y(n_374) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
A2O1A1Ixp33_ASAP7_75t_L g455 ( .A1(n_311), .A2(n_392), .B(n_456), .C(n_457), .Y(n_455) );
OAI322xp33_ASAP7_75t_SL g324 ( .A1(n_312), .A2(n_325), .A3(n_328), .B1(n_329), .B2(n_330), .C1(n_332), .C2(n_335), .Y(n_324) );
INVx2_ASAP7_75t_L g344 ( .A(n_312), .Y(n_344) );
AOI221xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_320), .B1(n_321), .B2(n_323), .C(n_324), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OAI22xp33_ASAP7_75t_SL g390 ( .A1(n_315), .A2(n_391), .B1(n_392), .B2(n_395), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_316), .B(n_319), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_316), .B(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g389 ( .A(n_318), .B(n_351), .Y(n_389) );
INVx1_ASAP7_75t_L g379 ( .A(n_319), .Y(n_379) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g432 ( .A1(n_323), .A2(n_433), .B(n_435), .Y(n_432) );
AOI21xp33_ASAP7_75t_L g357 ( .A1(n_325), .A2(n_358), .B(n_361), .Y(n_357) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NOR2xp67_ASAP7_75t_SL g386 ( .A(n_327), .B(n_387), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_327), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_SL g443 ( .A(n_328), .Y(n_443) );
INVx1_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND4xp25_ASAP7_75t_L g336 ( .A(n_337), .B(n_364), .C(n_380), .D(n_396), .Y(n_336) );
AOI211xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_340), .B(n_345), .C(n_357), .Y(n_337) );
INVx1_ASAP7_75t_L g429 ( .A(n_338), .Y(n_429) );
AND2x2_ASAP7_75t_L g377 ( .A(n_339), .B(n_360), .Y(n_377) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_342), .B(n_344), .Y(n_341) );
INVx1_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_344), .B(n_379), .Y(n_378) );
OAI22xp33_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_350), .B1(n_353), .B2(n_355), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_347), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g395 ( .A(n_348), .Y(n_395) );
O2A1O1Ixp33_ASAP7_75t_L g409 ( .A1(n_348), .A2(n_387), .B(n_410), .C(n_412), .Y(n_409) );
OR2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
INVx1_ASAP7_75t_L g394 ( .A(n_351), .Y(n_394) );
INVx1_ASAP7_75t_L g454 ( .A(n_352), .Y(n_454) );
NAND2xp33_ASAP7_75t_SL g444 ( .A(n_353), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g383 ( .A(n_362), .Y(n_383) );
O2A1O1Ixp33_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_368), .B(n_369), .C(n_371), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OAI22xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_373), .B1(n_376), .B2(n_378), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_374), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_379), .B(n_400), .Y(n_462) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AOI21xp33_ASAP7_75t_SL g384 ( .A1(n_385), .A2(n_388), .B(n_389), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_402), .B1(n_405), .B2(n_407), .C(n_409), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
INVx1_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVxp67_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_412), .A2(n_429), .B1(n_430), .B2(n_431), .Y(n_428) );
NAND3xp33_ASAP7_75t_SL g414 ( .A(n_415), .B(n_422), .C(n_432), .Y(n_414) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_SL g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
CKINVDCx16_ASAP7_75t_R g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVxp67_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OAI211xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_440), .B(n_441), .C(n_450), .Y(n_438) );
INVx1_ASAP7_75t_L g459 ( .A(n_439), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_444), .B1(n_446), .B2(n_448), .Y(n_441) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_459), .B1(n_460), .B2(n_461), .Y(n_457) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g471 ( .A(n_466), .Y(n_471) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NAND3xp33_ASAP7_75t_L g472 ( .A(n_470), .B(n_473), .C(n_758), .Y(n_472) );
XNOR2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_484), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_477), .Y(n_476) );
CKINVDCx16_ASAP7_75t_R g479 ( .A(n_480), .Y(n_479) );
OR2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_683), .Y(n_486) );
NAND5xp2_ASAP7_75t_L g487 ( .A(n_488), .B(n_598), .C(n_630), .D(n_647), .E(n_670), .Y(n_487) );
AOI221xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_531), .B1(n_561), .B2(n_565), .C(n_569), .Y(n_488) );
INVx1_ASAP7_75t_L g710 ( .A(n_489), .Y(n_710) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_510), .Y(n_489) );
AND3x2_ASAP7_75t_L g685 ( .A(n_490), .B(n_512), .C(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_500), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_491), .B(n_567), .Y(n_566) );
BUFx3_ASAP7_75t_L g576 ( .A(n_491), .Y(n_576) );
AND2x2_ASAP7_75t_L g580 ( .A(n_491), .B(n_522), .Y(n_580) );
INVx2_ASAP7_75t_L g607 ( .A(n_491), .Y(n_607) );
OR2x2_ASAP7_75t_L g618 ( .A(n_491), .B(n_523), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_491), .B(n_511), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_491), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g697 ( .A(n_491), .B(n_523), .Y(n_697) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_500), .Y(n_579) );
AND2x2_ASAP7_75t_L g638 ( .A(n_500), .B(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_500), .B(n_511), .Y(n_657) );
INVx1_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
OR2x2_ASAP7_75t_L g568 ( .A(n_501), .B(n_511), .Y(n_568) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_501), .Y(n_575) );
AND2x2_ASAP7_75t_L g624 ( .A(n_501), .B(n_523), .Y(n_624) );
NAND3xp33_ASAP7_75t_L g649 ( .A(n_501), .B(n_510), .C(n_607), .Y(n_649) );
AND2x2_ASAP7_75t_L g714 ( .A(n_501), .B(n_512), .Y(n_714) );
AND2x2_ASAP7_75t_L g748 ( .A(n_501), .B(n_511), .Y(n_748) );
INVxp67_ASAP7_75t_L g577 ( .A(n_510), .Y(n_577) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_522), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_511), .B(n_607), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_511), .B(n_638), .Y(n_646) );
AND2x2_ASAP7_75t_L g696 ( .A(n_511), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g724 ( .A(n_511), .Y(n_724) );
INVx4_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g631 ( .A(n_512), .B(n_624), .Y(n_631) );
BUFx3_ASAP7_75t_L g663 ( .A(n_512), .Y(n_663) );
INVx2_ASAP7_75t_L g639 ( .A(n_522), .Y(n_639) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_523), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_531), .A2(n_699), .B1(n_701), .B2(n_702), .Y(n_698) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_541), .Y(n_531) );
AND2x2_ASAP7_75t_L g561 ( .A(n_532), .B(n_562), .Y(n_561) );
INVx3_ASAP7_75t_SL g572 ( .A(n_532), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_532), .B(n_602), .Y(n_634) );
OR2x2_ASAP7_75t_L g653 ( .A(n_532), .B(n_542), .Y(n_653) );
AND2x2_ASAP7_75t_L g658 ( .A(n_532), .B(n_610), .Y(n_658) );
AND2x2_ASAP7_75t_L g661 ( .A(n_532), .B(n_603), .Y(n_661) );
AND2x2_ASAP7_75t_L g673 ( .A(n_532), .B(n_552), .Y(n_673) );
AND2x2_ASAP7_75t_L g689 ( .A(n_532), .B(n_543), .Y(n_689) );
AND2x4_ASAP7_75t_L g692 ( .A(n_532), .B(n_563), .Y(n_692) );
OR2x2_ASAP7_75t_L g709 ( .A(n_532), .B(n_645), .Y(n_709) );
OR2x2_ASAP7_75t_L g740 ( .A(n_532), .B(n_585), .Y(n_740) );
NAND2xp5_ASAP7_75t_SL g742 ( .A(n_532), .B(n_668), .Y(n_742) );
OR2x6_ASAP7_75t_L g532 ( .A(n_533), .B(n_539), .Y(n_532) );
AND2x2_ASAP7_75t_L g616 ( .A(n_541), .B(n_583), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_541), .B(n_603), .Y(n_735) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_552), .Y(n_541) );
AND2x2_ASAP7_75t_L g571 ( .A(n_542), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g602 ( .A(n_542), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g610 ( .A(n_542), .B(n_585), .Y(n_610) );
AND2x2_ASAP7_75t_L g628 ( .A(n_542), .B(n_563), .Y(n_628) );
OR2x2_ASAP7_75t_L g645 ( .A(n_542), .B(n_603), .Y(n_645) );
INVx2_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
BUFx2_ASAP7_75t_L g564 ( .A(n_543), .Y(n_564) );
AND2x2_ASAP7_75t_L g668 ( .A(n_543), .B(n_552), .Y(n_668) );
INVx2_ASAP7_75t_L g563 ( .A(n_552), .Y(n_563) );
INVx1_ASAP7_75t_L g680 ( .A(n_552), .Y(n_680) );
AND2x2_ASAP7_75t_L g730 ( .A(n_552), .B(n_572), .Y(n_730) );
AND2x2_ASAP7_75t_L g582 ( .A(n_562), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g614 ( .A(n_562), .B(n_572), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_562), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
AND2x2_ASAP7_75t_L g601 ( .A(n_563), .B(n_572), .Y(n_601) );
OR2x2_ASAP7_75t_L g717 ( .A(n_564), .B(n_691), .Y(n_717) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_567), .B(n_697), .Y(n_703) );
INVx2_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
OAI32xp33_ASAP7_75t_L g659 ( .A1(n_568), .A2(n_660), .A3(n_662), .B1(n_664), .B2(n_665), .Y(n_659) );
OR2x2_ASAP7_75t_L g676 ( .A(n_568), .B(n_618), .Y(n_676) );
OAI21xp33_ASAP7_75t_SL g701 ( .A1(n_568), .A2(n_578), .B(n_606), .Y(n_701) );
OAI22xp33_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_573), .B1(n_578), .B2(n_581), .Y(n_569) );
INVxp33_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_571), .B(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_572), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g627 ( .A(n_572), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g727 ( .A(n_572), .B(n_668), .Y(n_727) );
OR2x2_ASAP7_75t_L g751 ( .A(n_572), .B(n_645), .Y(n_751) );
AOI21xp33_ASAP7_75t_L g734 ( .A1(n_573), .A2(n_633), .B(n_735), .Y(n_734) );
OR2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_577), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
INVx1_ASAP7_75t_L g611 ( .A(n_575), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_575), .B(n_580), .Y(n_629) );
AND2x2_ASAP7_75t_L g651 ( .A(n_576), .B(n_624), .Y(n_651) );
INVx1_ASAP7_75t_L g664 ( .A(n_576), .Y(n_664) );
OR2x2_ASAP7_75t_L g669 ( .A(n_576), .B(n_603), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_579), .B(n_618), .Y(n_617) );
OAI22xp33_ASAP7_75t_L g599 ( .A1(n_580), .A2(n_600), .B1(n_605), .B2(n_609), .Y(n_599) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_583), .A2(n_642), .B1(n_649), .B2(n_650), .Y(n_648) );
AND2x2_ASAP7_75t_L g726 ( .A(n_583), .B(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_585), .B(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g745 ( .A(n_585), .B(n_628), .Y(n_745) );
AO21x2_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_588), .B(n_596), .Y(n_585) );
INVx1_ASAP7_75t_L g604 ( .A(n_586), .Y(n_604) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OA21x2_ASAP7_75t_L g603 ( .A1(n_589), .A2(n_597), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AOI221xp5_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_611), .B1(n_612), .B2(n_617), .C(n_619), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_601), .B(n_603), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_601), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g620 ( .A(n_602), .Y(n_620) );
O2A1O1Ixp33_ASAP7_75t_L g707 ( .A1(n_602), .A2(n_708), .B(n_709), .C(n_710), .Y(n_707) );
AND2x2_ASAP7_75t_L g712 ( .A(n_602), .B(n_692), .Y(n_712) );
O2A1O1Ixp33_ASAP7_75t_SL g750 ( .A1(n_602), .A2(n_691), .B(n_751), .C(n_752), .Y(n_750) );
BUFx3_ASAP7_75t_L g642 ( .A(n_603), .Y(n_642) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_606), .B(n_663), .Y(n_706) );
AOI211xp5_ASAP7_75t_L g725 ( .A1(n_606), .A2(n_726), .B(n_728), .C(n_734), .Y(n_725) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
INVxp67_ASAP7_75t_L g686 ( .A(n_608), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_610), .B(n_730), .Y(n_729) );
NAND2xp5_ASAP7_75t_SL g612 ( .A(n_613), .B(n_615), .Y(n_612) );
INVx1_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
AOI211xp5_ASAP7_75t_L g630 ( .A1(n_614), .A2(n_631), .B(n_632), .C(n_640), .Y(n_630) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g715 ( .A(n_618), .Y(n_715) );
OR2x2_ASAP7_75t_L g732 ( .A(n_618), .B(n_662), .Y(n_732) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_621), .B1(n_626), .B2(n_629), .Y(n_619) );
OAI22xp33_ASAP7_75t_L g632 ( .A1(n_621), .A2(n_633), .B1(n_634), .B2(n_635), .Y(n_632) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_625), .Y(n_622) );
OR2x2_ASAP7_75t_L g719 ( .A(n_623), .B(n_663), .Y(n_719) );
INVx1_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g674 ( .A(n_624), .B(n_664), .Y(n_674) );
INVx1_ASAP7_75t_L g682 ( .A(n_625), .Y(n_682) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_628), .B(n_642), .Y(n_690) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g681 ( .A(n_638), .B(n_682), .Y(n_681) );
INVx2_ASAP7_75t_L g747 ( .A(n_639), .Y(n_747) );
AOI21xp33_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_643), .B(n_646), .Y(n_640) );
INVx1_ASAP7_75t_L g677 ( .A(n_641), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g652 ( .A(n_642), .B(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_642), .B(n_673), .Y(n_672) );
NAND2x1p5_ASAP7_75t_L g693 ( .A(n_642), .B(n_668), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g700 ( .A(n_642), .B(n_689), .Y(n_700) );
OAI211xp5_ASAP7_75t_L g704 ( .A1(n_642), .A2(n_652), .B(n_692), .C(n_705), .Y(n_704) );
INVx1_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
AOI221xp5_ASAP7_75t_SL g647 ( .A1(n_648), .A2(n_652), .B1(n_654), .B2(n_658), .C(n_659), .Y(n_647) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVxp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_656), .B(n_664), .Y(n_738) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
O2A1O1Ixp33_ASAP7_75t_L g749 ( .A1(n_658), .A2(n_673), .B(n_675), .C(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_661), .B(n_668), .Y(n_733) );
NAND2xp5_ASAP7_75t_SL g752 ( .A(n_662), .B(n_715), .Y(n_752) );
CKINVDCx16_ASAP7_75t_R g662 ( .A(n_663), .Y(n_662) );
INVxp33_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_669), .Y(n_666) );
AOI21xp33_ASAP7_75t_SL g678 ( .A1(n_667), .A2(n_679), .B(n_681), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_667), .B(n_740), .Y(n_739) );
INVx2_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_668), .B(n_722), .Y(n_721) );
AOI221xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_674), .B1(n_675), .B2(n_677), .C(n_678), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_674), .B(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g708 ( .A(n_680), .Y(n_708) );
NAND5xp2_ASAP7_75t_L g683 ( .A(n_684), .B(n_711), .C(n_725), .D(n_736), .E(n_749), .Y(n_683) );
AOI211xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_687), .B(n_694), .C(n_707), .Y(n_684) );
INVx2_ASAP7_75t_SL g731 ( .A(n_685), .Y(n_731) );
NAND4xp25_ASAP7_75t_SL g687 ( .A(n_688), .B(n_690), .C(n_691), .D(n_693), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx3_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OAI211xp5_ASAP7_75t_SL g694 ( .A1(n_693), .A2(n_695), .B(n_698), .C(n_704), .Y(n_694) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_696), .Y(n_695) );
AOI221xp5_ASAP7_75t_L g736 ( .A1(n_696), .A2(n_737), .B1(n_739), .B2(n_741), .C(n_743), .Y(n_736) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AOI221xp5_ASAP7_75t_SL g711 ( .A1(n_712), .A2(n_713), .B1(n_716), .B2(n_718), .C(n_720), .Y(n_711) );
AND2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_719), .A2(n_742), .B1(n_744), .B2(n_746), .Y(n_743) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_731), .B1(n_732), .B2(n_733), .Y(n_728) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
endmodule