module fake_netlist_6_3931_n_3520 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_695, n_507, n_580, n_762, n_209, n_367, n_465, n_680, n_741, n_760, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_726, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_740, n_578, n_703, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_106, n_725, n_358, n_160, n_751, n_449, n_131, n_749, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_396, n_495, n_350, n_78, n_84, n_585, n_732, n_568, n_392, n_442, n_480, n_142, n_724, n_143, n_382, n_673, n_180, n_62, n_628, n_557, n_349, n_643, n_233, n_617, n_698, n_255, n_739, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_768, n_38, n_471, n_289, n_421, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_769, n_202, n_320, n_108, n_639, n_676, n_327, n_727, n_369, n_597, n_685, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_669, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_718, n_747, n_667, n_71, n_74, n_229, n_542, n_644, n_682, n_621, n_305, n_72, n_721, n_750, n_532, n_742, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_704, n_748, n_506, n_56, n_763, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_710, n_387, n_452, n_616, n_658, n_744, n_39, n_344, n_73, n_581, n_428, n_761, n_746, n_609, n_765, n_432, n_641, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_720, n_525, n_758, n_611, n_156, n_491, n_145, n_42, n_133, n_656, n_772, n_96, n_8, n_666, n_371, n_770, n_567, n_189, n_738, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_653, n_752, n_112, n_172, n_713, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_734, n_708, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_709, n_366, n_777, n_407, n_450, n_103, n_272, n_526, n_185, n_712, n_348, n_711, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_717, n_46, n_330, n_771, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_686, n_252, n_757, n_228, n_565, n_594, n_719, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_745, n_654, n_323, n_606, n_393, n_411, n_503, n_716, n_152, n_623, n_92, n_599, n_513, n_776, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_731, n_406, n_483, n_735, n_102, n_204, n_482, n_755, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_714, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_767, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_345, n_409, n_231, n_354, n_689, n_40, n_505, n_240, n_756, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_635, n_95, n_311, n_10, n_403, n_723, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_764, n_556, n_159, n_157, n_162, n_692, n_733, n_754, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_560, n_753, n_642, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_737, n_318, n_303, n_511, n_715, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_582, n_4, n_199, n_138, n_266, n_296, n_674, n_775, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_759, n_355, n_426, n_317, n_149, n_632, n_702, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_773, n_675, n_85, n_99, n_257, n_730, n_655, n_13, n_706, n_670, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_690, n_29, n_75, n_401, n_324, n_743, n_766, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_728, n_681, n_729, n_110, n_151, n_774, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_688, n_722, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_637, n_295, n_385, n_701, n_629, n_388, n_190, n_262, n_484, n_613, n_736, n_187, n_501, n_531, n_60, n_361, n_508, n_663, n_379, n_170, n_778, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_3520);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_695;
input n_507;
input n_580;
input n_762;
input n_209;
input n_367;
input n_465;
input n_680;
input n_741;
input n_760;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_726;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_740;
input n_578;
input n_703;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_106;
input n_725;
input n_358;
input n_160;
input n_751;
input n_449;
input n_131;
input n_749;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_732;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_724;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_255;
input n_739;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_768;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_769;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_727;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_669;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_718;
input n_747;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_644;
input n_682;
input n_621;
input n_305;
input n_72;
input n_721;
input n_750;
input n_532;
input n_742;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_704;
input n_748;
input n_506;
input n_56;
input n_763;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_710;
input n_387;
input n_452;
input n_616;
input n_658;
input n_744;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_761;
input n_746;
input n_609;
input n_765;
input n_432;
input n_641;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_720;
input n_525;
input n_758;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_656;
input n_772;
input n_96;
input n_8;
input n_666;
input n_371;
input n_770;
input n_567;
input n_189;
input n_738;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_752;
input n_112;
input n_172;
input n_713;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_734;
input n_708;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_709;
input n_366;
input n_777;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_712;
input n_348;
input n_711;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_717;
input n_46;
input n_330;
input n_771;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_686;
input n_252;
input n_757;
input n_228;
input n_565;
input n_594;
input n_719;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_745;
input n_654;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_716;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_776;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_731;
input n_406;
input n_483;
input n_735;
input n_102;
input n_204;
input n_482;
input n_755;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_714;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_767;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_505;
input n_240;
input n_756;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_635;
input n_95;
input n_311;
input n_10;
input n_403;
input n_723;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_764;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_733;
input n_754;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_560;
input n_753;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_737;
input n_318;
input n_303;
input n_511;
input n_715;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_674;
input n_775;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_759;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_773;
input n_675;
input n_85;
input n_99;
input n_257;
input n_730;
input n_655;
input n_13;
input n_706;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_690;
input n_29;
input n_75;
input n_401;
input n_324;
input n_743;
input n_766;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_728;
input n_681;
input n_729;
input n_110;
input n_151;
input n_774;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_688;
input n_722;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_637;
input n_295;
input n_385;
input n_701;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_736;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_663;
input n_379;
input n_170;
input n_778;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_3520;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_1613;
wire n_1458;
wire n_2576;
wire n_1234;
wire n_3254;
wire n_1199;
wire n_1674;
wire n_3392;
wire n_1027;
wire n_1351;
wire n_3266;
wire n_1189;
wire n_3152;
wire n_1212;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_3301;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_3088;
wire n_3443;
wire n_1923;
wire n_3257;
wire n_1342;
wire n_1348;
wire n_1209;
wire n_1387;
wire n_2260;
wire n_3222;
wire n_1708;
wire n_805;
wire n_1151;
wire n_2977;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_3332;
wire n_3465;
wire n_1975;
wire n_1930;
wire n_1743;
wire n_1009;
wire n_2405;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_2382;
wire n_2672;
wire n_3030;
wire n_2291;
wire n_830;
wire n_2299;
wire n_3340;
wire n_1371;
wire n_873;
wire n_1285;
wire n_2886;
wire n_2974;
wire n_1985;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_2247;
wire n_1711;
wire n_1078;
wire n_3106;
wire n_2630;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_836;
wire n_3345;
wire n_2074;
wire n_2447;
wire n_2919;
wire n_3440;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1772;
wire n_1232;
wire n_1572;
wire n_1874;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_2480;
wire n_2739;
wire n_3023;
wire n_822;
wire n_3232;
wire n_1313;
wire n_2791;
wire n_3251;
wire n_1056;
wire n_3316;
wire n_2212;
wire n_3494;
wire n_3048;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3063;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_1798;
wire n_943;
wire n_1550;
wire n_2703;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_940;
wire n_1971;
wire n_1781;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_3028;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_3077;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3452;
wire n_3107;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_1421;
wire n_2836;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_3047;
wire n_1280;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_1467;
wire n_3297;
wire n_976;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_1088;
wire n_1894;
wire n_2996;
wire n_1231;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_2085;
wire n_3368;
wire n_917;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_3507;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_3506;
wire n_3269;
wire n_1230;
wire n_3413;
wire n_1967;
wire n_1193;
wire n_1054;
wire n_3412;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_1986;
wire n_2300;
wire n_2397;
wire n_824;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_2907;
wire n_3438;
wire n_2735;
wire n_1843;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_2850;
wire n_1909;
wire n_2080;
wire n_813;
wire n_1481;
wire n_1441;
wire n_818;
wire n_3373;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_1381;
wire n_2961;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_2059;
wire n_2198;
wire n_3319;
wire n_2669;
wire n_2925;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_792;
wire n_2522;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_2616;
wire n_3118;
wire n_3315;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_3488;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1599;
wire n_1068;
wire n_982;
wire n_2674;
wire n_2832;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_2831;
wire n_2998;
wire n_3446;
wire n_3317;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_3518;
wire n_1866;
wire n_1680;
wire n_2692;
wire n_993;
wire n_3248;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_3514;
wire n_2228;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_2455;
wire n_2876;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_2355;
wire n_966;
wire n_2908;
wire n_3168;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_2895;
wire n_2009;
wire n_3403;
wire n_1793;
wire n_2922;
wire n_1233;
wire n_2714;
wire n_1289;
wire n_2245;
wire n_3092;
wire n_3055;
wire n_3492;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_3294;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_1265;
wire n_2711;
wire n_3490;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_3369;
wire n_3419;
wire n_1982;
wire n_2878;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3247;
wire n_871;
wire n_3069;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_2641;
wire n_1664;
wire n_1722;
wire n_3022;
wire n_3052;
wire n_1165;
wire n_2008;
wire n_2749;
wire n_3298;
wire n_2192;
wire n_3281;
wire n_2254;
wire n_2345;
wire n_3346;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_780;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_928;
wire n_1801;
wire n_835;
wire n_2347;
wire n_850;
wire n_1886;
wire n_1214;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_3453;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3410;
wire n_3153;
wire n_3428;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_825;
wire n_2916;
wire n_3415;
wire n_1063;
wire n_1588;
wire n_2963;
wire n_2947;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_1624;
wire n_1124;
wire n_2096;
wire n_2980;
wire n_1965;
wire n_2476;
wire n_3280;
wire n_3434;
wire n_1515;
wire n_961;
wire n_3510;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_890;
wire n_2377;
wire n_2178;
wire n_3271;
wire n_950;
wire n_2812;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_3460;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_3237;
wire n_949;
wire n_1630;
wire n_2887;
wire n_3500;
wire n_2075;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_3192;
wire n_1546;
wire n_2583;
wire n_2606;
wire n_2279;
wire n_1052;
wire n_1033;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_3073;
wire n_2431;
wire n_2987;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_3252;
wire n_2932;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_3253;
wire n_3337;
wire n_3431;
wire n_3209;
wire n_3450;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2893;
wire n_2775;
wire n_1208;
wire n_1627;
wire n_1164;
wire n_1295;
wire n_2954;
wire n_3477;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_1487;
wire n_2691;
wire n_3421;
wire n_840;
wire n_2913;
wire n_874;
wire n_1756;
wire n_3183;
wire n_2493;
wire n_1128;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1565;
wire n_1067;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_3436;
wire n_1932;
wire n_925;
wire n_1101;
wire n_2535;
wire n_1026;
wire n_1880;
wire n_3366;
wire n_3442;
wire n_2631;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_963;
wire n_2767;
wire n_794;
wire n_894;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_2707;
wire n_3240;
wire n_1514;
wire n_1863;
wire n_826;
wire n_3385;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_1714;
wire n_872;
wire n_1139;
wire n_3179;
wire n_1018;
wire n_3400;
wire n_1521;
wire n_1366;
wire n_847;
wire n_851;
wire n_2537;
wire n_2897;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_2747;
wire n_3171;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_3491;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_3158;
wire n_1788;
wire n_3426;
wire n_1999;
wire n_2731;
wire n_2590;
wire n_2643;
wire n_3150;
wire n_3018;
wire n_3353;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_3470;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_1492;
wire n_987;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_3104;
wire n_3435;
wire n_842;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_1432;
wire n_2208;
wire n_843;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_2012;
wire n_3497;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_1809;
wire n_3119;
wire n_2948;
wire n_1577;
wire n_2958;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_2936;
wire n_3224;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_3173;
wire n_1992;
wire n_1049;
wire n_3223;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_1717;
wire n_1817;
wire n_926;
wire n_2449;
wire n_927;
wire n_2610;
wire n_3129;
wire n_1849;
wire n_2848;
wire n_919;
wire n_2868;
wire n_1698;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_2857;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_1299;
wire n_2896;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_3325;
wire n_2238;
wire n_2368;
wire n_2403;
wire n_1070;
wire n_3342;
wire n_2837;
wire n_998;
wire n_3200;
wire n_1665;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_3390;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_3324;
wire n_3341;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_1507;
wire n_2482;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3006;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_3201;
wire n_3447;
wire n_1142;
wire n_2849;
wire n_1475;
wire n_1774;
wire n_1398;
wire n_1201;
wire n_884;
wire n_1048;
wire n_2354;
wire n_2682;
wire n_3103;
wire n_3032;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_931;
wire n_1021;
wire n_3393;
wire n_811;
wire n_2442;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_3451;
wire n_3480;
wire n_1418;
wire n_958;
wire n_1250;
wire n_3331;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_889;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_1310;
wire n_3142;
wire n_819;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_1314;
wire n_1837;
wire n_831;
wire n_2218;
wire n_964;
wire n_2788;
wire n_3196;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2860;
wire n_2292;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2511;
wire n_2475;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_1877;
wire n_3144;
wire n_3211;
wire n_3244;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_3287;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_970;
wire n_3306;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_2329;
wire n_1092;
wire n_3481;
wire n_2237;
wire n_3026;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_3033;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_1223;
wire n_2990;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3226;
wire n_3323;
wire n_3364;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_1153;
wire n_1618;
wire n_3407;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_3425;
wire n_2384;
wire n_1745;
wire n_914;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_2801;
wire n_2920;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_2306;
wire n_1892;
wire n_1459;
wire n_1614;
wire n_3188;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_2889;
wire n_1169;
wire n_3243;
wire n_1617;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_1470;
wire n_2550;
wire n_3093;
wire n_3175;
wire n_3214;
wire n_1243;
wire n_848;
wire n_2732;
wire n_2928;
wire n_2249;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_3284;
wire n_983;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_1390;
wire n_906;
wire n_2289;
wire n_1733;
wire n_1077;
wire n_2315;
wire n_1419;
wire n_2863;
wire n_3299;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_3360;
wire n_2135;
wire n_3367;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_2627;
wire n_3234;
wire n_2276;
wire n_960;
wire n_956;
wire n_856;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_2993;
wire n_3016;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_1129;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_1869;
wire n_2911;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_1889;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_793;
wire n_3466;
wire n_1593;
wire n_1202;
wire n_1030;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_2942;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_2555;
wire n_3338;
wire n_3462;
wire n_2219;
wire n_1203;
wire n_2851;
wire n_3406;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_999;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_2984;
wire n_2263;
wire n_994;
wire n_3291;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_3194;
wire n_3250;
wire n_1934;
wire n_3276;
wire n_1020;
wire n_1042;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_2756;
wire n_1871;
wire n_3448;
wire n_845;
wire n_807;
wire n_2924;
wire n_1036;
wire n_1138;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_1510;
wire n_892;
wire n_3120;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_2052;
wire n_1847;
wire n_2302;
wire n_1667;
wire n_1206;
wire n_3230;
wire n_1397;
wire n_1037;
wire n_3236;
wire n_1279;
wire n_1115;
wire n_901;
wire n_1499;
wire n_2755;
wire n_3141;
wire n_923;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_3195;
wire n_2526;
wire n_3041;
wire n_2423;
wire n_1057;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_991;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_2439;
wire n_1818;
wire n_1108;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_3399;
wire n_2088;
wire n_1611;
wire n_785;
wire n_2740;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_3416;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_3042;
wire n_3213;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1943;
wire n_1216;
wire n_3228;
wire n_1320;
wire n_2716;
wire n_3249;
wire n_3081;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3010;
wire n_2499;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_3382;
wire n_2486;
wire n_3132;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3238;
wire n_2235;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_3424;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_809;
wire n_1043;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_2964;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_3485;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3475;
wire n_3501;
wire n_1840;
wire n_1152;
wire n_1705;
wire n_3262;
wire n_2904;
wire n_2244;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_3029;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_962;
wire n_1041;
wire n_2346;
wire n_3134;
wire n_1569;
wire n_936;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_1288;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_2882;
wire n_3320;
wire n_2541;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_934;
wire n_1637;
wire n_2635;
wire n_3307;
wire n_3439;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_2871;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_3502;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_3184;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_2390;
wire n_806;
wire n_879;
wire n_2310;
wire n_959;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_2986;
wire n_1900;
wire n_3246;
wire n_799;
wire n_1548;
wire n_3381;
wire n_3044;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_787;
wire n_2172;
wire n_3489;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2962;
wire n_2154;
wire n_2727;
wire n_3377;
wire n_2939;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_2533;
wire n_3157;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_3457;
wire n_2759;
wire n_1229;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_3469;
wire n_2266;
wire n_2960;
wire n_3005;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_1706;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_3375;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3379;
wire n_3156;
wire n_1931;
wire n_2083;
wire n_1269;
wire n_2834;
wire n_3207;
wire n_2668;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_1375;
wire n_1941;
wire n_3483;
wire n_2128;
wire n_1650;
wire n_1794;
wire n_786;
wire n_1962;
wire n_1045;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_3091;
wire n_834;
wire n_2695;
wire n_3124;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_3398;
wire n_2671;
wire n_2888;
wire n_2761;
wire n_2885;
wire n_2793;
wire n_2715;
wire n_2923;
wire n_1804;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_3511;
wire n_2054;
wire n_876;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_3308;
wire n_1600;
wire n_1113;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_1098;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_841;
wire n_1476;
wire n_2516;
wire n_3391;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_3458;
wire n_3515;
wire n_1150;
wire n_3190;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1882;
wire n_1023;
wire n_2951;
wire n_1076;
wire n_1118;
wire n_2949;
wire n_1807;
wire n_1929;
wire n_1007;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_1879;
wire n_853;
wire n_1542;
wire n_2587;
wire n_3199;
wire n_2931;
wire n_875;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_1953;
wire n_933;
wire n_3343;
wire n_3303;
wire n_978;
wire n_2752;
wire n_3135;
wire n_1976;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_2140;
wire n_988;
wire n_3503;
wire n_3160;
wire n_2796;
wire n_1065;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2186;
wire n_2163;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3034;
wire n_823;
wire n_1132;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_2969;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_3027;
wire n_781;
wire n_789;
wire n_1554;
wire n_3231;
wire n_1130;
wire n_3083;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_2380;
wire n_1120;
wire n_832;
wire n_1583;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_814;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_1461;
wire n_3432;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_3493;
wire n_2935;
wire n_863;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_2910;
wire n_2385;
wire n_1283;
wire n_918;
wire n_1848;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_3268;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3154;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_1994;
wire n_957;
wire n_3473;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_971;
wire n_2702;
wire n_3241;
wire n_946;
wire n_2906;
wire n_1303;
wire n_2769;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_2180;
wire n_1689;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_3334;
wire n_1245;
wire n_838;
wire n_3215;
wire n_3336;
wire n_844;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_1083;
wire n_1561;
wire n_2741;
wire n_3114;
wire n_930;
wire n_888;
wire n_2275;
wire n_2465;
wire n_1112;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_3486;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_2034;
wire n_1028;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_2444;
wire n_2437;
wire n_1215;
wire n_839;
wire n_2743;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_3204;
wire n_1104;
wire n_854;
wire n_1058;
wire n_3378;
wire n_2312;
wire n_3404;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_2242;
wire n_1266;
wire n_3362;
wire n_1509;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3290;
wire n_1109;
wire n_2222;
wire n_3256;
wire n_1276;
wire n_3176;
wire n_3309;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2505;
wire n_2188;
wire n_1989;
wire n_2609;
wire n_1161;
wire n_1085;
wire n_2802;
wire n_2999;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_1584;
wire n_2425;
wire n_924;
wire n_3461;
wire n_3408;
wire n_1582;
wire n_2318;
wire n_3286;
wire n_2408;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_1184;
wire n_2483;
wire n_2950;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_2592;
wire n_1525;
wire n_3098;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_1362;
wire n_1156;
wire n_829;
wire n_3123;
wire n_2600;
wire n_984;
wire n_3380;
wire n_1829;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_868;
wire n_3038;
wire n_859;
wire n_2033;
wire n_3086;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_3285;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_3361;
wire n_981;
wire n_3478;
wire n_1349;
wire n_2071;
wire n_1144;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_3233;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_3496;
wire n_1301;
wire n_2805;
wire n_802;
wire n_3310;
wire n_980;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_3344;
wire n_2334;
wire n_3295;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_1194;
wire n_3374;
wire n_2742;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_1996;
wire n_2367;
wire n_2867;
wire n_3198;
wire n_1039;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_941;
wire n_975;
wire n_3206;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_849;
wire n_2662;
wire n_3116;
wire n_3147;
wire n_3383;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_3187;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3330;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_2065;
wire n_2879;
wire n_861;
wire n_857;
wire n_967;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_2968;
wire n_1629;
wire n_2221;
wire n_1170;
wire n_1819;
wire n_2055;
wire n_1260;
wire n_1010;
wire n_3444;
wire n_2553;
wire n_1040;
wire n_915;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3467;
wire n_3001;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_3433;
wire n_1365;
wire n_1417;
wire n_2185;
wire n_2086;
wire n_1242;
wire n_2927;
wire n_1836;
wire n_2774;
wire n_3039;
wire n_1226;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3274;
wire n_3333;
wire n_3186;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_2579;
wire n_862;
wire n_2105;
wire n_3079;
wire n_2098;
wire n_3085;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_3387;
wire n_2027;
wire n_3070;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_3504;
wire n_1449;
wire n_827;
wire n_2912;
wire n_2659;
wire n_2930;
wire n_1025;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_1742;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g779 ( 
.A(n_527),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_663),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_490),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_61),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_158),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_671),
.Y(n_784)
);

INVx1_ASAP7_75t_SL g785 ( 
.A(n_402),
.Y(n_785)
);

INVx1_ASAP7_75t_SL g786 ( 
.A(n_768),
.Y(n_786)
);

BUFx10_ASAP7_75t_L g787 ( 
.A(n_756),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_675),
.Y(n_788)
);

CKINVDCx16_ASAP7_75t_R g789 ( 
.A(n_354),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_687),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_565),
.Y(n_791)
);

BUFx3_ASAP7_75t_L g792 ( 
.A(n_398),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_185),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_746),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_628),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_738),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_472),
.Y(n_797)
);

INVx1_ASAP7_75t_SL g798 ( 
.A(n_284),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_652),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_121),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_464),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_749),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_573),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_558),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_152),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_438),
.Y(n_806)
);

CKINVDCx14_ASAP7_75t_R g807 ( 
.A(n_362),
.Y(n_807)
);

CKINVDCx20_ASAP7_75t_R g808 ( 
.A(n_715),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_383),
.Y(n_809)
);

INVx1_ASAP7_75t_SL g810 ( 
.A(n_568),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_547),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_725),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_597),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_230),
.Y(n_814)
);

BUFx5_ASAP7_75t_L g815 ( 
.A(n_694),
.Y(n_815)
);

CKINVDCx20_ASAP7_75t_R g816 ( 
.A(n_357),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_631),
.Y(n_817)
);

INVx2_ASAP7_75t_SL g818 ( 
.A(n_610),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_717),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_741),
.Y(n_820)
);

BUFx5_ASAP7_75t_L g821 ( 
.A(n_386),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_634),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_656),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_706),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_550),
.Y(n_825)
);

BUFx3_ASAP7_75t_L g826 ( 
.A(n_724),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_740),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_342),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_100),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_403),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_676),
.Y(n_831)
);

CKINVDCx20_ASAP7_75t_R g832 ( 
.A(n_769),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_462),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_33),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_572),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_762),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_701),
.Y(n_837)
);

BUFx3_ASAP7_75t_L g838 ( 
.A(n_583),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_734),
.Y(n_839)
);

INVx2_ASAP7_75t_SL g840 ( 
.A(n_526),
.Y(n_840)
);

BUFx10_ASAP7_75t_L g841 ( 
.A(n_743),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_733),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_523),
.Y(n_843)
);

INVx1_ASAP7_75t_SL g844 ( 
.A(n_569),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_129),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_81),
.Y(n_846)
);

BUFx3_ASAP7_75t_L g847 ( 
.A(n_287),
.Y(n_847)
);

INVx1_ASAP7_75t_SL g848 ( 
.A(n_33),
.Y(n_848)
);

CKINVDCx20_ASAP7_75t_R g849 ( 
.A(n_739),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_125),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_392),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_337),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_552),
.Y(n_853)
);

CKINVDCx20_ASAP7_75t_R g854 ( 
.A(n_592),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_645),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_574),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_594),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_771),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_536),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_657),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_580),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_736),
.Y(n_862)
);

CKINVDCx20_ASAP7_75t_R g863 ( 
.A(n_325),
.Y(n_863)
);

CKINVDCx20_ASAP7_75t_R g864 ( 
.A(n_686),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_674),
.Y(n_865)
);

BUFx3_ASAP7_75t_L g866 ( 
.A(n_589),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_608),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_176),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_638),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_765),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_653),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_28),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_100),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_487),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_368),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_763),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_402),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_582),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_351),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_661),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_707),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_551),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_723),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_212),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_745),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_632),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_535),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_648),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_642),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_180),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_578),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_533),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_757),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_297),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_309),
.Y(n_895)
);

BUFx10_ASAP7_75t_L g896 ( 
.A(n_384),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_668),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_700),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_479),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_679),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_630),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_538),
.Y(n_902)
);

CKINVDCx20_ASAP7_75t_R g903 ( 
.A(n_629),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_264),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_655),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_772),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_627),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_68),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_525),
.Y(n_909)
);

CKINVDCx20_ASAP7_75t_R g910 ( 
.A(n_159),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_662),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_0),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_639),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_682),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_464),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_325),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_759),
.Y(n_917)
);

CKINVDCx20_ASAP7_75t_R g918 ( 
.A(n_542),
.Y(n_918)
);

INVx3_ASAP7_75t_L g919 ( 
.A(n_532),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_421),
.Y(n_920)
);

CKINVDCx20_ASAP7_75t_R g921 ( 
.A(n_534),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_117),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_358),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_252),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_425),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_584),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_48),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_263),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_773),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_716),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_305),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_315),
.Y(n_932)
);

BUFx10_ASAP7_75t_L g933 ( 
.A(n_714),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_683),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_195),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_590),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_670),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_431),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_327),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_684),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_262),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_195),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_74),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_316),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_98),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_123),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_549),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_555),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_338),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_484),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_767),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_444),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_651),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_774),
.Y(n_954)
);

CKINVDCx14_ASAP7_75t_R g955 ( 
.A(n_18),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_332),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_171),
.Y(n_957)
);

CKINVDCx16_ASAP7_75t_R g958 ( 
.A(n_228),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_224),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_690),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_465),
.Y(n_961)
);

HB1xp67_ASAP7_75t_L g962 ( 
.A(n_777),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_114),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_531),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_504),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_90),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_563),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_75),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_537),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_279),
.Y(n_970)
);

INVx2_ASAP7_75t_SL g971 ( 
.A(n_350),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_143),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_737),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_471),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_660),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_166),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_264),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_617),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_233),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_457),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_7),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_515),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_424),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_97),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_107),
.Y(n_985)
);

INVx2_ASAP7_75t_SL g986 ( 
.A(n_556),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_421),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_57),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_49),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_596),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_308),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_649),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_560),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_274),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_368),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_562),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_742),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_593),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_541),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_336),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_623),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_600),
.Y(n_1002)
);

CKINVDCx16_ASAP7_75t_R g1003 ( 
.A(n_761),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_776),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_728),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_727),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_514),
.Y(n_1007)
);

CKINVDCx16_ASAP7_75t_R g1008 ( 
.A(n_174),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_159),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_664),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_451),
.Y(n_1011)
);

BUFx3_ASAP7_75t_L g1012 ( 
.A(n_41),
.Y(n_1012)
);

CKINVDCx14_ASAP7_75t_R g1013 ( 
.A(n_555),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_260),
.Y(n_1014)
);

CKINVDCx20_ASAP7_75t_R g1015 ( 
.A(n_386),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_681),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_10),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_303),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_215),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_635),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_371),
.Y(n_1021)
);

CKINVDCx20_ASAP7_75t_R g1022 ( 
.A(n_541),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_329),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_722),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_297),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_281),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_551),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_747),
.Y(n_1028)
);

CKINVDCx20_ASAP7_75t_R g1029 ( 
.A(n_640),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_591),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_647),
.Y(n_1031)
);

BUFx10_ASAP7_75t_L g1032 ( 
.A(n_406),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_123),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_680),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_90),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_528),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_522),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_571),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_601),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_666),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_633),
.Y(n_1041)
);

INVx1_ASAP7_75t_SL g1042 ( 
.A(n_704),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_570),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_84),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_718),
.Y(n_1045)
);

BUFx5_ASAP7_75t_L g1046 ( 
.A(n_711),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_172),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_207),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_521),
.Y(n_1049)
);

CKINVDCx20_ASAP7_75t_R g1050 ( 
.A(n_708),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_382),
.Y(n_1051)
);

CKINVDCx20_ASAP7_75t_R g1052 ( 
.A(n_703),
.Y(n_1052)
);

CKINVDCx20_ASAP7_75t_R g1053 ( 
.A(n_702),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_699),
.Y(n_1054)
);

CKINVDCx20_ASAP7_75t_R g1055 ( 
.A(n_778),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_366),
.Y(n_1056)
);

CKINVDCx20_ASAP7_75t_R g1057 ( 
.A(n_587),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_430),
.Y(n_1058)
);

BUFx8_ASAP7_75t_SL g1059 ( 
.A(n_581),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_220),
.Y(n_1060)
);

CKINVDCx20_ASAP7_75t_R g1061 ( 
.A(n_542),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_592),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_554),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_443),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_473),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_347),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_197),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_301),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_454),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_248),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_41),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_117),
.Y(n_1072)
);

INVx1_ASAP7_75t_SL g1073 ( 
.A(n_528),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_245),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_389),
.Y(n_1075)
);

CKINVDCx20_ASAP7_75t_R g1076 ( 
.A(n_513),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_726),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_442),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_97),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_513),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_744),
.Y(n_1081)
);

BUFx8_ASAP7_75t_SL g1082 ( 
.A(n_677),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_465),
.Y(n_1083)
);

CKINVDCx20_ASAP7_75t_R g1084 ( 
.A(n_217),
.Y(n_1084)
);

CKINVDCx20_ASAP7_75t_R g1085 ( 
.A(n_665),
.Y(n_1085)
);

INVx1_ASAP7_75t_SL g1086 ( 
.A(n_685),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_263),
.Y(n_1087)
);

CKINVDCx20_ASAP7_75t_R g1088 ( 
.A(n_242),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_557),
.Y(n_1089)
);

BUFx2_ASAP7_75t_L g1090 ( 
.A(n_25),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_389),
.Y(n_1091)
);

INVx1_ASAP7_75t_SL g1092 ( 
.A(n_691),
.Y(n_1092)
);

CKINVDCx20_ASAP7_75t_R g1093 ( 
.A(n_92),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_543),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_468),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_221),
.Y(n_1096)
);

BUFx3_ASAP7_75t_L g1097 ( 
.A(n_345),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_579),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_383),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_70),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_593),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_74),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_561),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_644),
.Y(n_1104)
);

BUFx3_ASAP7_75t_L g1105 ( 
.A(n_315),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_167),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_278),
.Y(n_1107)
);

CKINVDCx20_ASAP7_75t_R g1108 ( 
.A(n_88),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_147),
.Y(n_1109)
);

BUFx3_ASAP7_75t_L g1110 ( 
.A(n_408),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_646),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_559),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_719),
.Y(n_1113)
);

BUFx2_ASAP7_75t_L g1114 ( 
.A(n_296),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_735),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_650),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_178),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_271),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_110),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_57),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_393),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_269),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_111),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_342),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_257),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_753),
.Y(n_1126)
);

CKINVDCx20_ASAP7_75t_R g1127 ( 
.A(n_546),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_112),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_556),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_364),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_176),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_673),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_299),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_536),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_140),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_42),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_689),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_564),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_4),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_294),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_211),
.Y(n_1142)
);

CKINVDCx11_ASAP7_75t_R g1143 ( 
.A(n_193),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_8),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_732),
.Y(n_1145)
);

INVx2_ASAP7_75t_SL g1146 ( 
.A(n_101),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_135),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_266),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_419),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_539),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_624),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_731),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_108),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_232),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_567),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_606),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_710),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_597),
.Y(n_1158)
);

BUFx10_ASAP7_75t_L g1159 ( 
.A(n_602),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_696),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_544),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_173),
.Y(n_1162)
);

CKINVDCx20_ASAP7_75t_R g1163 ( 
.A(n_119),
.Y(n_1163)
);

INVx2_ASAP7_75t_R g1164 ( 
.A(n_192),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_210),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_270),
.Y(n_1166)
);

BUFx10_ASAP7_75t_L g1167 ( 
.A(n_391),
.Y(n_1167)
);

BUFx3_ASAP7_75t_L g1168 ( 
.A(n_487),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_300),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_692),
.Y(n_1170)
);

INVxp67_ASAP7_75t_SL g1171 ( 
.A(n_238),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_253),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_190),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_729),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_571),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_626),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_522),
.Y(n_1177)
);

BUFx2_ASAP7_75t_L g1178 ( 
.A(n_538),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_524),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_130),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_328),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_512),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_529),
.Y(n_1183)
);

CKINVDCx16_ASAP7_75t_R g1184 ( 
.A(n_122),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_414),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_385),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_637),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_730),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_755),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_568),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_621),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_429),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_751),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_175),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_202),
.Y(n_1195)
);

INVx2_ASAP7_75t_SL g1196 ( 
.A(n_335),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_697),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_658),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_518),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_80),
.Y(n_1200)
);

CKINVDCx20_ASAP7_75t_R g1201 ( 
.A(n_575),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_709),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_486),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_441),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_174),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_292),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_449),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_3),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_586),
.Y(n_1209)
);

CKINVDCx20_ASAP7_75t_R g1210 ( 
.A(n_698),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_461),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_21),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_318),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_286),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_492),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_27),
.Y(n_1216)
);

CKINVDCx16_ASAP7_75t_R g1217 ( 
.A(n_688),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_576),
.Y(n_1218)
);

INVx1_ASAP7_75t_SL g1219 ( 
.A(n_764),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_748),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_43),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_387),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_625),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_659),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_108),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_484),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_288),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_760),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_179),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_299),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_588),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_306),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_382),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_583),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_219),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_326),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_643),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_252),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_566),
.Y(n_1239)
);

CKINVDCx16_ASAP7_75t_R g1240 ( 
.A(n_540),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_356),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_125),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_693),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_436),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_750),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_775),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_548),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_26),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_32),
.Y(n_1249)
);

CKINVDCx20_ASAP7_75t_R g1250 ( 
.A(n_287),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_358),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_61),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_585),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_495),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_232),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_530),
.Y(n_1256)
);

CKINVDCx16_ASAP7_75t_R g1257 ( 
.A(n_183),
.Y(n_1257)
);

BUFx8_ASAP7_75t_SL g1258 ( 
.A(n_221),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_534),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_488),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_261),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_641),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_69),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_236),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_705),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_669),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_463),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_244),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_329),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_766),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_180),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_280),
.Y(n_1272)
);

BUFx10_ASAP7_75t_L g1273 ( 
.A(n_667),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_201),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_553),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_29),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_96),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_378),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_154),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_133),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_713),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_239),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_84),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_712),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_247),
.Y(n_1285)
);

BUFx3_ASAP7_75t_L g1286 ( 
.A(n_288),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_262),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_577),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_66),
.Y(n_1289)
);

CKINVDCx14_ASAP7_75t_R g1290 ( 
.A(n_118),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_508),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_303),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_758),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_654),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_413),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_770),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_678),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_695),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_326),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_474),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_672),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_545),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_721),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_595),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_268),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_720),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_395),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_446),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_412),
.Y(n_1309)
);

CKINVDCx20_ASAP7_75t_R g1310 ( 
.A(n_754),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_752),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_636),
.Y(n_1312)
);

BUFx6f_ASAP7_75t_L g1313 ( 
.A(n_163),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_498),
.Y(n_1314)
);

INVxp33_ASAP7_75t_L g1315 ( 
.A(n_928),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_821),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_1143),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_821),
.Y(n_1318)
);

INVxp67_ASAP7_75t_SL g1319 ( 
.A(n_962),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_955),
.B(n_0),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_821),
.Y(n_1321)
);

INVxp67_ASAP7_75t_SL g1322 ( 
.A(n_1005),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_1059),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_821),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_821),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_792),
.Y(n_1326)
);

CKINVDCx16_ASAP7_75t_R g1327 ( 
.A(n_789),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_792),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_806),
.Y(n_1329)
);

CKINVDCx20_ASAP7_75t_R g1330 ( 
.A(n_1310),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1313),
.Y(n_1331)
);

INVxp67_ASAP7_75t_SL g1332 ( 
.A(n_919),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_806),
.Y(n_1333)
);

CKINVDCx14_ASAP7_75t_R g1334 ( 
.A(n_807),
.Y(n_1334)
);

INVxp67_ASAP7_75t_SL g1335 ( 
.A(n_999),
.Y(n_1335)
);

INVxp67_ASAP7_75t_SL g1336 ( 
.A(n_999),
.Y(n_1336)
);

CKINVDCx14_ASAP7_75t_R g1337 ( 
.A(n_807),
.Y(n_1337)
);

BUFx10_ASAP7_75t_L g1338 ( 
.A(n_1314),
.Y(n_1338)
);

CKINVDCx20_ASAP7_75t_R g1339 ( 
.A(n_808),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_834),
.Y(n_1340)
);

CKINVDCx20_ASAP7_75t_R g1341 ( 
.A(n_832),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_838),
.Y(n_1342)
);

CKINVDCx20_ASAP7_75t_R g1343 ( 
.A(n_849),
.Y(n_1343)
);

INVx1_ASAP7_75t_SL g1344 ( 
.A(n_1062),
.Y(n_1344)
);

INVxp67_ASAP7_75t_SL g1345 ( 
.A(n_826),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_847),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_847),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1313),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_861),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_861),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_866),
.Y(n_1351)
);

CKINVDCx20_ASAP7_75t_R g1352 ( 
.A(n_864),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_866),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_991),
.Y(n_1354)
);

CKINVDCx20_ASAP7_75t_R g1355 ( 
.A(n_903),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1012),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1012),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1089),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1089),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1097),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1258),
.Y(n_1361)
);

CKINVDCx16_ASAP7_75t_R g1362 ( 
.A(n_958),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1101),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1105),
.Y(n_1364)
);

INVxp67_ASAP7_75t_L g1365 ( 
.A(n_1087),
.Y(n_1365)
);

BUFx6f_ASAP7_75t_L g1366 ( 
.A(n_788),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1105),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1110),
.Y(n_1368)
);

INVxp67_ASAP7_75t_L g1369 ( 
.A(n_1090),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1110),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1168),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1168),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1286),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1008),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_805),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1184),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_805),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_805),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_780),
.Y(n_1379)
);

CKINVDCx20_ASAP7_75t_R g1380 ( 
.A(n_1029),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_805),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1313),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_809),
.Y(n_1383)
);

INVxp67_ASAP7_75t_L g1384 ( 
.A(n_1114),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_809),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_809),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_809),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1240),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_784),
.Y(n_1389)
);

BUFx8_ASAP7_75t_SL g1390 ( 
.A(n_1178),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_859),
.Y(n_1391)
);

CKINVDCx16_ASAP7_75t_R g1392 ( 
.A(n_1257),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_859),
.Y(n_1393)
);

CKINVDCx16_ASAP7_75t_R g1394 ( 
.A(n_1003),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_859),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_931),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_931),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_931),
.Y(n_1398)
);

BUFx3_ASAP7_75t_L g1399 ( 
.A(n_787),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_931),
.Y(n_1400)
);

CKINVDCx20_ASAP7_75t_R g1401 ( 
.A(n_1050),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_939),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_939),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_939),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_939),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_972),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_972),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_972),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_972),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_989),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_989),
.Y(n_1411)
);

INVxp33_ASAP7_75t_SL g1412 ( 
.A(n_781),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_794),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_989),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_989),
.Y(n_1415)
);

INVxp33_ASAP7_75t_L g1416 ( 
.A(n_779),
.Y(n_1416)
);

INVxp33_ASAP7_75t_L g1417 ( 
.A(n_783),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1021),
.Y(n_1418)
);

INVxp67_ASAP7_75t_SL g1419 ( 
.A(n_898),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1021),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1021),
.Y(n_1421)
);

INVxp67_ASAP7_75t_SL g1422 ( 
.A(n_929),
.Y(n_1422)
);

CKINVDCx20_ASAP7_75t_R g1423 ( 
.A(n_1052),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1021),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_795),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1094),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1094),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_799),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1117),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1304),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1117),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1199),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1199),
.Y(n_1433)
);

CKINVDCx20_ASAP7_75t_R g1434 ( 
.A(n_1053),
.Y(n_1434)
);

INVxp33_ASAP7_75t_SL g1435 ( 
.A(n_782),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1199),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1199),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_802),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1222),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1222),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1222),
.Y(n_1441)
);

INVxp67_ASAP7_75t_L g1442 ( 
.A(n_896),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1222),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1279),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1279),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1279),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1279),
.Y(n_1447)
);

CKINVDCx14_ASAP7_75t_R g1448 ( 
.A(n_955),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1300),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1305),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_788),
.Y(n_1451)
);

INVxp67_ASAP7_75t_SL g1452 ( 
.A(n_1115),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_812),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_817),
.Y(n_1454)
);

BUFx6f_ASAP7_75t_L g1455 ( 
.A(n_1366),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1348),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1382),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1405),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1445),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1375),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1334),
.B(n_1013),
.Y(n_1461)
);

BUFx6f_ASAP7_75t_L g1462 ( 
.A(n_1366),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1377),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1376),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1378),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1381),
.Y(n_1466)
);

BUFx6f_ASAP7_75t_L g1467 ( 
.A(n_1366),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1383),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1385),
.Y(n_1469)
);

BUFx8_ASAP7_75t_L g1470 ( 
.A(n_1399),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1389),
.B(n_818),
.Y(n_1471)
);

CKINVDCx11_ASAP7_75t_R g1472 ( 
.A(n_1338),
.Y(n_1472)
);

BUFx6f_ASAP7_75t_L g1473 ( 
.A(n_1451),
.Y(n_1473)
);

AND2x2_ASAP7_75t_SL g1474 ( 
.A(n_1394),
.B(n_1217),
.Y(n_1474)
);

INVx5_ASAP7_75t_L g1475 ( 
.A(n_1390),
.Y(n_1475)
);

AND2x4_ASAP7_75t_L g1476 ( 
.A(n_1322),
.B(n_1284),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_L g1477 ( 
.A(n_1451),
.Y(n_1477)
);

BUFx8_ASAP7_75t_L g1478 ( 
.A(n_1326),
.Y(n_1478)
);

AOI22x1_ASAP7_75t_R g1479 ( 
.A1(n_1330),
.A2(n_854),
.B1(n_863),
.B2(n_816),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1386),
.Y(n_1480)
);

INVx6_ASAP7_75t_L g1481 ( 
.A(n_1338),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_1412),
.B(n_1013),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1387),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1391),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1393),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1395),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1396),
.Y(n_1487)
);

BUFx6f_ASAP7_75t_L g1488 ( 
.A(n_1397),
.Y(n_1488)
);

BUFx6f_ASAP7_75t_L g1489 ( 
.A(n_1398),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1400),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1413),
.B(n_790),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1318),
.A2(n_886),
.B(n_824),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1402),
.Y(n_1493)
);

INVx3_ASAP7_75t_L g1494 ( 
.A(n_1403),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1388),
.Y(n_1495)
);

AOI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1344),
.A2(n_1290),
.B1(n_1055),
.B2(n_1210),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1337),
.B(n_1290),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1404),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1406),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1362),
.Y(n_1500)
);

INVx3_ASAP7_75t_L g1501 ( 
.A(n_1407),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_1425),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1345),
.B(n_786),
.Y(n_1503)
);

INVxp67_ASAP7_75t_L g1504 ( 
.A(n_1430),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1408),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1409),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1410),
.Y(n_1507)
);

BUFx6f_ASAP7_75t_L g1508 ( 
.A(n_1411),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1414),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1428),
.B(n_824),
.Y(n_1510)
);

BUFx6f_ASAP7_75t_L g1511 ( 
.A(n_1415),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1418),
.Y(n_1512)
);

BUFx6f_ASAP7_75t_L g1513 ( 
.A(n_1420),
.Y(n_1513)
);

BUFx6f_ASAP7_75t_L g1514 ( 
.A(n_1421),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1424),
.Y(n_1515)
);

INVx3_ASAP7_75t_L g1516 ( 
.A(n_1426),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1392),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1427),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1438),
.B(n_886),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1429),
.Y(n_1520)
);

AOI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1319),
.A2(n_1085),
.B1(n_1301),
.B2(n_1171),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1431),
.Y(n_1522)
);

INVx5_ASAP7_75t_L g1523 ( 
.A(n_1448),
.Y(n_1523)
);

AND2x6_ASAP7_75t_L g1524 ( 
.A(n_1320),
.B(n_785),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1432),
.Y(n_1525)
);

INVx3_ASAP7_75t_L g1526 ( 
.A(n_1433),
.Y(n_1526)
);

INVx3_ASAP7_75t_L g1527 ( 
.A(n_1436),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1437),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1439),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1440),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1441),
.Y(n_1531)
);

BUFx3_ASAP7_75t_L g1532 ( 
.A(n_1328),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1443),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1444),
.Y(n_1534)
);

CKINVDCx20_ASAP7_75t_R g1535 ( 
.A(n_1339),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1446),
.Y(n_1536)
);

BUFx6f_ASAP7_75t_L g1537 ( 
.A(n_1447),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_SL g1538 ( 
.A(n_1323),
.B(n_1082),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1321),
.Y(n_1539)
);

INVx3_ASAP7_75t_L g1540 ( 
.A(n_1329),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_1453),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1454),
.B(n_917),
.Y(n_1542)
);

INVx3_ASAP7_75t_L g1543 ( 
.A(n_1333),
.Y(n_1543)
);

CKINVDCx16_ASAP7_75t_R g1544 ( 
.A(n_1341),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1332),
.Y(n_1545)
);

BUFx6f_ASAP7_75t_L g1546 ( 
.A(n_1449),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1335),
.Y(n_1547)
);

AND2x6_ASAP7_75t_L g1548 ( 
.A(n_1340),
.B(n_798),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1324),
.Y(n_1549)
);

INVx3_ASAP7_75t_L g1550 ( 
.A(n_1342),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1325),
.Y(n_1551)
);

BUFx6f_ASAP7_75t_L g1552 ( 
.A(n_1450),
.Y(n_1552)
);

INVx5_ASAP7_75t_L g1553 ( 
.A(n_1435),
.Y(n_1553)
);

INVx3_ASAP7_75t_L g1554 ( 
.A(n_1346),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1336),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1419),
.B(n_787),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1422),
.B(n_973),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1347),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1349),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1350),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1452),
.B(n_841),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1351),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1353),
.Y(n_1563)
);

NAND2x1_ASAP7_75t_L g1564 ( 
.A(n_1354),
.B(n_788),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1356),
.Y(n_1565)
);

INVx3_ASAP7_75t_L g1566 ( 
.A(n_1357),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1358),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1359),
.Y(n_1568)
);

NOR2xp33_ASAP7_75t_L g1569 ( 
.A(n_1365),
.B(n_1042),
.Y(n_1569)
);

BUFx6f_ASAP7_75t_L g1570 ( 
.A(n_1360),
.Y(n_1570)
);

INVx3_ASAP7_75t_L g1571 ( 
.A(n_1363),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1364),
.Y(n_1572)
);

INVx5_ASAP7_75t_L g1573 ( 
.A(n_1416),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1367),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1368),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_L g1576 ( 
.A(n_1369),
.B(n_1086),
.Y(n_1576)
);

BUFx6f_ASAP7_75t_L g1577 ( 
.A(n_1370),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1315),
.B(n_841),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1384),
.B(n_1092),
.Y(n_1579)
);

BUFx6f_ASAP7_75t_L g1580 ( 
.A(n_1371),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1372),
.B(n_973),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1373),
.Y(n_1582)
);

BUFx6f_ASAP7_75t_L g1583 ( 
.A(n_1361),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1417),
.B(n_933),
.Y(n_1584)
);

BUFx6f_ASAP7_75t_L g1585 ( 
.A(n_1442),
.Y(n_1585)
);

AND2x4_ASAP7_75t_L g1586 ( 
.A(n_1343),
.B(n_1219),
.Y(n_1586)
);

BUFx2_ASAP7_75t_L g1587 ( 
.A(n_1352),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1355),
.Y(n_1588)
);

BUFx3_ASAP7_75t_L g1589 ( 
.A(n_1380),
.Y(n_1589)
);

AND2x6_ASAP7_75t_L g1590 ( 
.A(n_1401),
.B(n_810),
.Y(n_1590)
);

INVx5_ASAP7_75t_L g1591 ( 
.A(n_1423),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1434),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1334),
.B(n_933),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1331),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1331),
.Y(n_1595)
);

INVx3_ASAP7_75t_L g1596 ( 
.A(n_1331),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1379),
.B(n_1001),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1331),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_L g1599 ( 
.A(n_1412),
.B(n_1306),
.Y(n_1599)
);

BUFx2_ASAP7_75t_L g1600 ( 
.A(n_1317),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1331),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1331),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1331),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1331),
.Y(n_1604)
);

BUFx12f_ASAP7_75t_L g1605 ( 
.A(n_1323),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1331),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1331),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1331),
.Y(n_1608)
);

BUFx3_ASAP7_75t_L g1609 ( 
.A(n_1326),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1331),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1399),
.B(n_820),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1331),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1331),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1331),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_1379),
.Y(n_1615)
);

NOR2x1_ASAP7_75t_L g1616 ( 
.A(n_1399),
.B(n_822),
.Y(n_1616)
);

HB1xp67_ASAP7_75t_L g1617 ( 
.A(n_1374),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1331),
.Y(n_1618)
);

BUFx6f_ASAP7_75t_L g1619 ( 
.A(n_1366),
.Y(n_1619)
);

BUFx2_ASAP7_75t_L g1620 ( 
.A(n_1317),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1331),
.Y(n_1621)
);

BUFx6f_ASAP7_75t_L g1622 ( 
.A(n_1366),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1374),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1331),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1331),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1331),
.Y(n_1626)
);

NOR2xp33_ASAP7_75t_L g1627 ( 
.A(n_1412),
.B(n_1016),
.Y(n_1627)
);

BUFx12f_ASAP7_75t_L g1628 ( 
.A(n_1323),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1331),
.Y(n_1629)
);

BUFx2_ASAP7_75t_L g1630 ( 
.A(n_1317),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1331),
.Y(n_1631)
);

BUFx8_ASAP7_75t_L g1632 ( 
.A(n_1399),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1331),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1331),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1331),
.Y(n_1635)
);

NOR2x1_ASAP7_75t_L g1636 ( 
.A(n_1399),
.B(n_823),
.Y(n_1636)
);

BUFx3_ASAP7_75t_L g1637 ( 
.A(n_1326),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1331),
.Y(n_1638)
);

BUFx3_ASAP7_75t_L g1639 ( 
.A(n_1326),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1399),
.B(n_827),
.Y(n_1640)
);

OAI21x1_ASAP7_75t_L g1641 ( 
.A1(n_1316),
.A2(n_1224),
.B(n_1016),
.Y(n_1641)
);

BUFx6f_ASAP7_75t_L g1642 ( 
.A(n_1366),
.Y(n_1642)
);

BUFx6f_ASAP7_75t_L g1643 ( 
.A(n_1366),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1331),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1379),
.B(n_1224),
.Y(n_1645)
);

INVx4_ASAP7_75t_L g1646 ( 
.A(n_1379),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1344),
.B(n_844),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1331),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1399),
.B(n_836),
.Y(n_1649)
);

BUFx2_ASAP7_75t_L g1650 ( 
.A(n_1317),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1331),
.Y(n_1651)
);

CKINVDCx6p67_ASAP7_75t_R g1652 ( 
.A(n_1327),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1379),
.B(n_1270),
.Y(n_1653)
);

NAND2xp33_ASAP7_75t_L g1654 ( 
.A(n_1320),
.B(n_1302),
.Y(n_1654)
);

AOI22xp33_ASAP7_75t_SL g1655 ( 
.A1(n_1334),
.A2(n_918),
.B1(n_921),
.B2(n_910),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1412),
.B(n_1293),
.Y(n_1656)
);

BUFx3_ASAP7_75t_L g1657 ( 
.A(n_1326),
.Y(n_1657)
);

INVxp67_ASAP7_75t_L g1658 ( 
.A(n_1374),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1331),
.Y(n_1659)
);

AND2x4_ASAP7_75t_L g1660 ( 
.A(n_1399),
.B(n_865),
.Y(n_1660)
);

BUFx6f_ASAP7_75t_L g1661 ( 
.A(n_1366),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1379),
.B(n_1293),
.Y(n_1662)
);

AND2x6_ASAP7_75t_L g1663 ( 
.A(n_1399),
.B(n_848),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1379),
.B(n_1298),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1379),
.B(n_867),
.Y(n_1665)
);

INVx3_ASAP7_75t_L g1666 ( 
.A(n_1331),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1331),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1412),
.B(n_869),
.Y(n_1668)
);

BUFx3_ASAP7_75t_L g1669 ( 
.A(n_1326),
.Y(n_1669)
);

BUFx6f_ASAP7_75t_L g1670 ( 
.A(n_1366),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1331),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1331),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1379),
.B(n_876),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1331),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1379),
.B(n_883),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1331),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1331),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1331),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1331),
.Y(n_1679)
);

BUFx3_ASAP7_75t_L g1680 ( 
.A(n_1326),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1379),
.B(n_888),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1334),
.B(n_1159),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1331),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1331),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1331),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1379),
.B(n_906),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1331),
.Y(n_1687)
);

INVx4_ASAP7_75t_L g1688 ( 
.A(n_1379),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1331),
.Y(n_1689)
);

BUFx6f_ASAP7_75t_L g1690 ( 
.A(n_1366),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1331),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1399),
.B(n_914),
.Y(n_1692)
);

AND2x2_ASAP7_75t_SL g1693 ( 
.A(n_1394),
.B(n_853),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1379),
.B(n_930),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1374),
.Y(n_1695)
);

INVx3_ASAP7_75t_L g1696 ( 
.A(n_1331),
.Y(n_1696)
);

INVxp67_ASAP7_75t_L g1697 ( 
.A(n_1374),
.Y(n_1697)
);

OA21x2_ASAP7_75t_L g1698 ( 
.A1(n_1316),
.A2(n_951),
.B(n_940),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1331),
.Y(n_1699)
);

INVx5_ASAP7_75t_L g1700 ( 
.A(n_1390),
.Y(n_1700)
);

AND2x4_ASAP7_75t_L g1701 ( 
.A(n_1399),
.B(n_975),
.Y(n_1701)
);

INVx3_ASAP7_75t_L g1702 ( 
.A(n_1331),
.Y(n_1702)
);

INVx3_ASAP7_75t_L g1703 ( 
.A(n_1331),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1331),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_1502),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_1541),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1558),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1559),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_1615),
.Y(n_1709)
);

BUFx10_ASAP7_75t_L g1710 ( 
.A(n_1481),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1488),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_1535),
.Y(n_1712)
);

CKINVDCx5p33_ASAP7_75t_R g1713 ( 
.A(n_1544),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_1591),
.Y(n_1714)
);

CKINVDCx20_ASAP7_75t_R g1715 ( 
.A(n_1652),
.Y(n_1715)
);

CKINVDCx5p33_ASAP7_75t_R g1716 ( 
.A(n_1591),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_1589),
.Y(n_1717)
);

CKINVDCx5p33_ASAP7_75t_R g1718 ( 
.A(n_1605),
.Y(n_1718)
);

NOR2xp33_ASAP7_75t_R g1719 ( 
.A(n_1523),
.B(n_819),
.Y(n_1719)
);

INVx1_ASAP7_75t_SL g1720 ( 
.A(n_1573),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1488),
.Y(n_1721)
);

INVx3_ASAP7_75t_L g1722 ( 
.A(n_1455),
.Y(n_1722)
);

CKINVDCx5p33_ASAP7_75t_R g1723 ( 
.A(n_1628),
.Y(n_1723)
);

INVx5_ASAP7_75t_L g1724 ( 
.A(n_1523),
.Y(n_1724)
);

CKINVDCx20_ASAP7_75t_R g1725 ( 
.A(n_1587),
.Y(n_1725)
);

BUFx3_ASAP7_75t_L g1726 ( 
.A(n_1532),
.Y(n_1726)
);

NOR2x1p5_ASAP7_75t_L g1727 ( 
.A(n_1593),
.B(n_791),
.Y(n_1727)
);

NOR2xp67_ASAP7_75t_L g1728 ( 
.A(n_1646),
.B(n_1688),
.Y(n_1728)
);

CKINVDCx5p33_ASAP7_75t_R g1729 ( 
.A(n_1553),
.Y(n_1729)
);

CKINVDCx5p33_ASAP7_75t_R g1730 ( 
.A(n_1553),
.Y(n_1730)
);

CKINVDCx20_ASAP7_75t_R g1731 ( 
.A(n_1500),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1489),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1560),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1647),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_1475),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1562),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1489),
.Y(n_1737)
);

CKINVDCx20_ASAP7_75t_R g1738 ( 
.A(n_1517),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_1700),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1508),
.Y(n_1740)
);

NAND2xp33_ASAP7_75t_SL g1741 ( 
.A(n_1585),
.B(n_1015),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_1583),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_1472),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1565),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1508),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1511),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1567),
.Y(n_1747)
);

BUFx6f_ASAP7_75t_L g1748 ( 
.A(n_1455),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1568),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1511),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_1600),
.Y(n_1751)
);

BUFx6f_ASAP7_75t_L g1752 ( 
.A(n_1462),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_1620),
.Y(n_1753)
);

CKINVDCx20_ASAP7_75t_R g1754 ( 
.A(n_1630),
.Y(n_1754)
);

BUFx10_ASAP7_75t_L g1755 ( 
.A(n_1569),
.Y(n_1755)
);

CKINVDCx20_ASAP7_75t_R g1756 ( 
.A(n_1650),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1572),
.Y(n_1757)
);

NAND2xp33_ASAP7_75t_R g1758 ( 
.A(n_1586),
.B(n_793),
.Y(n_1758)
);

INVx3_ASAP7_75t_L g1759 ( 
.A(n_1462),
.Y(n_1759)
);

BUFx6f_ASAP7_75t_L g1760 ( 
.A(n_1467),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_R g1761 ( 
.A(n_1654),
.B(n_837),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1574),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1582),
.Y(n_1763)
);

CKINVDCx5p33_ASAP7_75t_R g1764 ( 
.A(n_1479),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1513),
.Y(n_1765)
);

AND3x1_ASAP7_75t_L g1766 ( 
.A(n_1496),
.B(n_840),
.C(n_825),
.Y(n_1766)
);

NOR2xp33_ASAP7_75t_R g1767 ( 
.A(n_1538),
.B(n_839),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_1588),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1513),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_1592),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1570),
.Y(n_1771)
);

CKINVDCx5p33_ASAP7_75t_R g1772 ( 
.A(n_1474),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1577),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_1590),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1491),
.B(n_842),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1580),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1580),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1563),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1514),
.Y(n_1779)
);

CKINVDCx20_ASAP7_75t_R g1780 ( 
.A(n_1464),
.Y(n_1780)
);

CKINVDCx5p33_ASAP7_75t_R g1781 ( 
.A(n_1590),
.Y(n_1781)
);

CKINVDCx20_ASAP7_75t_R g1782 ( 
.A(n_1495),
.Y(n_1782)
);

CKINVDCx5p33_ASAP7_75t_R g1783 ( 
.A(n_1470),
.Y(n_1783)
);

CKINVDCx20_ASAP7_75t_R g1784 ( 
.A(n_1617),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_1632),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1575),
.Y(n_1786)
);

INVx3_ASAP7_75t_L g1787 ( 
.A(n_1467),
.Y(n_1787)
);

INVx1_ASAP7_75t_SL g1788 ( 
.A(n_1584),
.Y(n_1788)
);

CKINVDCx5p33_ASAP7_75t_R g1789 ( 
.A(n_1482),
.Y(n_1789)
);

CKINVDCx5p33_ASAP7_75t_R g1790 ( 
.A(n_1471),
.Y(n_1790)
);

NOR2xp67_ASAP7_75t_L g1791 ( 
.A(n_1504),
.B(n_855),
.Y(n_1791)
);

NOR2xp33_ASAP7_75t_L g1792 ( 
.A(n_1665),
.B(n_971),
.Y(n_1792)
);

CKINVDCx5p33_ASAP7_75t_R g1793 ( 
.A(n_1668),
.Y(n_1793)
);

BUFx8_ASAP7_75t_L g1794 ( 
.A(n_1663),
.Y(n_1794)
);

INVx3_ASAP7_75t_L g1795 ( 
.A(n_1473),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1539),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_R g1797 ( 
.A(n_1545),
.B(n_858),
.Y(n_1797)
);

CKINVDCx5p33_ASAP7_75t_R g1798 ( 
.A(n_1510),
.Y(n_1798)
);

CKINVDCx5p33_ASAP7_75t_R g1799 ( 
.A(n_1519),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1531),
.Y(n_1800)
);

CKINVDCx20_ASAP7_75t_R g1801 ( 
.A(n_1623),
.Y(n_1801)
);

CKINVDCx5p33_ASAP7_75t_R g1802 ( 
.A(n_1542),
.Y(n_1802)
);

CKINVDCx5p33_ASAP7_75t_R g1803 ( 
.A(n_1597),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1549),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1551),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1609),
.Y(n_1806)
);

NOR2xp33_ASAP7_75t_R g1807 ( 
.A(n_1547),
.B(n_860),
.Y(n_1807)
);

CKINVDCx20_ASAP7_75t_R g1808 ( 
.A(n_1695),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1637),
.Y(n_1809)
);

CKINVDCx5p33_ASAP7_75t_R g1810 ( 
.A(n_1645),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1537),
.Y(n_1811)
);

BUFx2_ASAP7_75t_L g1812 ( 
.A(n_1663),
.Y(n_1812)
);

BUFx10_ASAP7_75t_L g1813 ( 
.A(n_1576),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_SL g1814 ( 
.A(n_1503),
.B(n_1273),
.Y(n_1814)
);

CKINVDCx5p33_ASAP7_75t_R g1815 ( 
.A(n_1653),
.Y(n_1815)
);

CKINVDCx5p33_ASAP7_75t_R g1816 ( 
.A(n_1662),
.Y(n_1816)
);

CKINVDCx5p33_ASAP7_75t_R g1817 ( 
.A(n_1664),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_1524),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1639),
.Y(n_1819)
);

CKINVDCx5p33_ASAP7_75t_R g1820 ( 
.A(n_1524),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1537),
.Y(n_1821)
);

CKINVDCx5p33_ASAP7_75t_R g1822 ( 
.A(n_1693),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1657),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1669),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1673),
.B(n_986),
.Y(n_1825)
);

INVx3_ASAP7_75t_L g1826 ( 
.A(n_1473),
.Y(n_1826)
);

CKINVDCx5p33_ASAP7_75t_R g1827 ( 
.A(n_1675),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1680),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1681),
.B(n_870),
.Y(n_1829)
);

CKINVDCx5p33_ASAP7_75t_R g1830 ( 
.A(n_1686),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1694),
.B(n_871),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1456),
.Y(n_1832)
);

INVxp67_ASAP7_75t_L g1833 ( 
.A(n_1578),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1546),
.Y(n_1834)
);

NOR2xp33_ASAP7_75t_L g1835 ( 
.A(n_1555),
.B(n_1146),
.Y(n_1835)
);

CKINVDCx20_ASAP7_75t_R g1836 ( 
.A(n_1521),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1552),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1552),
.Y(n_1838)
);

CKINVDCx5p33_ASAP7_75t_R g1839 ( 
.A(n_1599),
.Y(n_1839)
);

CKINVDCx5p33_ASAP7_75t_R g1840 ( 
.A(n_1627),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1458),
.Y(n_1841)
);

CKINVDCx5p33_ASAP7_75t_R g1842 ( 
.A(n_1656),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1594),
.Y(n_1843)
);

NOR2xp67_ASAP7_75t_L g1844 ( 
.A(n_1658),
.B(n_880),
.Y(n_1844)
);

CKINVDCx5p33_ASAP7_75t_R g1845 ( 
.A(n_1579),
.Y(n_1845)
);

CKINVDCx20_ASAP7_75t_R g1846 ( 
.A(n_1697),
.Y(n_1846)
);

CKINVDCx5p33_ASAP7_75t_R g1847 ( 
.A(n_1655),
.Y(n_1847)
);

CKINVDCx5p33_ASAP7_75t_R g1848 ( 
.A(n_1476),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_R g1849 ( 
.A(n_1461),
.B(n_881),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1556),
.B(n_885),
.Y(n_1850)
);

CKINVDCx20_ASAP7_75t_R g1851 ( 
.A(n_1497),
.Y(n_1851)
);

OAI21x1_ASAP7_75t_L g1852 ( 
.A1(n_1492),
.A2(n_1002),
.B(n_978),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1460),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1469),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1595),
.Y(n_1855)
);

NOR2xp33_ASAP7_75t_R g1856 ( 
.A(n_1682),
.B(n_889),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1480),
.Y(n_1857)
);

CKINVDCx5p33_ASAP7_75t_R g1858 ( 
.A(n_1561),
.Y(n_1858)
);

INVx8_ASAP7_75t_L g1859 ( 
.A(n_1548),
.Y(n_1859)
);

NOR2xp33_ASAP7_75t_L g1860 ( 
.A(n_1557),
.B(n_1611),
.Y(n_1860)
);

NOR2xp33_ASAP7_75t_R g1861 ( 
.A(n_1540),
.B(n_893),
.Y(n_1861)
);

CKINVDCx5p33_ASAP7_75t_R g1862 ( 
.A(n_1548),
.Y(n_1862)
);

HB1xp67_ASAP7_75t_L g1863 ( 
.A(n_1640),
.Y(n_1863)
);

CKINVDCx5p33_ASAP7_75t_R g1864 ( 
.A(n_1478),
.Y(n_1864)
);

NOR2xp33_ASAP7_75t_R g1865 ( 
.A(n_1543),
.B(n_897),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1649),
.B(n_1196),
.Y(n_1866)
);

CKINVDCx5p33_ASAP7_75t_R g1867 ( 
.A(n_1660),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1483),
.Y(n_1868)
);

INVx3_ASAP7_75t_L g1869 ( 
.A(n_1477),
.Y(n_1869)
);

INVx1_ASAP7_75t_SL g1870 ( 
.A(n_1692),
.Y(n_1870)
);

CKINVDCx5p33_ASAP7_75t_R g1871 ( 
.A(n_1701),
.Y(n_1871)
);

BUFx2_ASAP7_75t_L g1872 ( 
.A(n_1616),
.Y(n_1872)
);

NOR2xp33_ASAP7_75t_R g1873 ( 
.A(n_1550),
.B(n_901),
.Y(n_1873)
);

CKINVDCx5p33_ASAP7_75t_R g1874 ( 
.A(n_1554),
.Y(n_1874)
);

CKINVDCx20_ASAP7_75t_R g1875 ( 
.A(n_1581),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1487),
.Y(n_1876)
);

CKINVDCx5p33_ASAP7_75t_R g1877 ( 
.A(n_1566),
.Y(n_1877)
);

CKINVDCx5p33_ASAP7_75t_R g1878 ( 
.A(n_1571),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1493),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1499),
.Y(n_1880)
);

AND3x2_ASAP7_75t_L g1881 ( 
.A(n_1507),
.B(n_902),
.C(n_875),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1601),
.Y(n_1882)
);

CKINVDCx5p33_ASAP7_75t_R g1883 ( 
.A(n_1477),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1509),
.Y(n_1884)
);

INVx2_ASAP7_75t_SL g1885 ( 
.A(n_1636),
.Y(n_1885)
);

AO21x2_ASAP7_75t_L g1886 ( 
.A1(n_1641),
.A2(n_1010),
.B(n_1006),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1604),
.Y(n_1887)
);

BUFx6f_ASAP7_75t_L g1888 ( 
.A(n_1619),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_1622),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1606),
.B(n_905),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1607),
.Y(n_1891)
);

CKINVDCx5p33_ASAP7_75t_R g1892 ( 
.A(n_1642),
.Y(n_1892)
);

CKINVDCx5p33_ASAP7_75t_R g1893 ( 
.A(n_1642),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1512),
.Y(n_1894)
);

NOR2xp33_ASAP7_75t_R g1895 ( 
.A(n_1494),
.B(n_907),
.Y(n_1895)
);

CKINVDCx5p33_ASAP7_75t_R g1896 ( 
.A(n_1643),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1608),
.Y(n_1897)
);

BUFx3_ASAP7_75t_L g1898 ( 
.A(n_1564),
.Y(n_1898)
);

CKINVDCx5p33_ASAP7_75t_R g1899 ( 
.A(n_1643),
.Y(n_1899)
);

CKINVDCx5p33_ASAP7_75t_R g1900 ( 
.A(n_1661),
.Y(n_1900)
);

CKINVDCx5p33_ASAP7_75t_R g1901 ( 
.A(n_1661),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1596),
.B(n_1167),
.Y(n_1902)
);

BUFx3_ASAP7_75t_L g1903 ( 
.A(n_1670),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1612),
.Y(n_1904)
);

NAND2xp33_ASAP7_75t_SL g1905 ( 
.A(n_1670),
.B(n_1022),
.Y(n_1905)
);

CKINVDCx5p33_ASAP7_75t_R g1906 ( 
.A(n_1690),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1621),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1629),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1634),
.Y(n_1909)
);

BUFx3_ASAP7_75t_L g1910 ( 
.A(n_1690),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1518),
.Y(n_1911)
);

NOR2xp33_ASAP7_75t_R g1912 ( 
.A(n_1501),
.B(n_911),
.Y(n_1912)
);

CKINVDCx20_ASAP7_75t_R g1913 ( 
.A(n_1698),
.Y(n_1913)
);

AND3x2_ASAP7_75t_L g1914 ( 
.A(n_1520),
.B(n_902),
.C(n_875),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1827),
.B(n_1667),
.Y(n_1915)
);

INVx1_ASAP7_75t_SL g1916 ( 
.A(n_1734),
.Y(n_1916)
);

CKINVDCx5p33_ASAP7_75t_R g1917 ( 
.A(n_1705),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1707),
.Y(n_1918)
);

NAND2xp33_ASAP7_75t_R g1919 ( 
.A(n_1822),
.B(n_913),
.Y(n_1919)
);

AND2x6_ASAP7_75t_L g1920 ( 
.A(n_1788),
.B(n_788),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1830),
.B(n_1671),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1708),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1832),
.Y(n_1923)
);

BUFx2_ASAP7_75t_L g1924 ( 
.A(n_1845),
.Y(n_1924)
);

INVx4_ASAP7_75t_L g1925 ( 
.A(n_1742),
.Y(n_1925)
);

AOI22xp5_ASAP7_75t_SL g1926 ( 
.A1(n_1836),
.A2(n_1061),
.B1(n_1066),
.B2(n_1057),
.Y(n_1926)
);

OR2x6_ASAP7_75t_L g1927 ( 
.A(n_1859),
.B(n_1812),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1733),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1841),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1798),
.B(n_1674),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1799),
.B(n_1676),
.Y(n_1931)
);

BUFx6f_ASAP7_75t_L g1932 ( 
.A(n_1748),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1802),
.B(n_1683),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1736),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1744),
.Y(n_1935)
);

BUFx3_ASAP7_75t_L g1936 ( 
.A(n_1726),
.Y(n_1936)
);

BUFx6f_ASAP7_75t_L g1937 ( 
.A(n_1748),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1843),
.Y(n_1938)
);

AND2x2_ASAP7_75t_SL g1939 ( 
.A(n_1766),
.B(n_923),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1839),
.B(n_1032),
.Y(n_1940)
);

BUFx6f_ASAP7_75t_L g1941 ( 
.A(n_1748),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1803),
.B(n_1810),
.Y(n_1942)
);

INVxp67_ASAP7_75t_L g1943 ( 
.A(n_1758),
.Y(n_1943)
);

INVxp67_ASAP7_75t_SL g1944 ( 
.A(n_1752),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1747),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1749),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1840),
.B(n_1666),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1855),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1882),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1887),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1891),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1757),
.Y(n_1952)
);

INVx2_ASAP7_75t_SL g1953 ( 
.A(n_1902),
.Y(n_1953)
);

AND2x4_ASAP7_75t_L g1954 ( 
.A(n_1903),
.B(n_1529),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1897),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1762),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1763),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1842),
.B(n_1696),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1853),
.Y(n_1959)
);

AOI22xp33_ASAP7_75t_L g1960 ( 
.A1(n_1913),
.A2(n_1164),
.B1(n_1031),
.B2(n_1034),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1854),
.Y(n_1961)
);

INVx3_ASAP7_75t_L g1962 ( 
.A(n_1910),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1857),
.Y(n_1963)
);

CKINVDCx5p33_ASAP7_75t_R g1964 ( 
.A(n_1706),
.Y(n_1964)
);

NOR2xp33_ASAP7_75t_L g1965 ( 
.A(n_1793),
.B(n_1073),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1868),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1904),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1907),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1876),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_SL g1970 ( 
.A(n_1815),
.B(n_934),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1908),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1909),
.Y(n_1972)
);

CKINVDCx5p33_ASAP7_75t_R g1973 ( 
.A(n_1709),
.Y(n_1973)
);

BUFx6f_ASAP7_75t_L g1974 ( 
.A(n_1752),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_SL g1975 ( 
.A(n_1816),
.B(n_937),
.Y(n_1975)
);

INVx8_ASAP7_75t_L g1976 ( 
.A(n_1724),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_SL g1977 ( 
.A(n_1817),
.B(n_953),
.Y(n_1977)
);

INVx4_ASAP7_75t_L g1978 ( 
.A(n_1883),
.Y(n_1978)
);

AND2x6_ASAP7_75t_L g1979 ( 
.A(n_1860),
.B(n_796),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1796),
.Y(n_1980)
);

AND2x6_ASAP7_75t_L g1981 ( 
.A(n_1806),
.B(n_1809),
.Y(n_1981)
);

NOR2x1p5_ASAP7_75t_L g1982 ( 
.A(n_1864),
.B(n_797),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1755),
.B(n_1702),
.Y(n_1983)
);

INVx5_ASAP7_75t_L g1984 ( 
.A(n_1710),
.Y(n_1984)
);

INVx2_ASAP7_75t_SL g1985 ( 
.A(n_1710),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1804),
.Y(n_1986)
);

BUFx2_ASAP7_75t_L g1987 ( 
.A(n_1731),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1879),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1880),
.Y(n_1989)
);

CKINVDCx5p33_ASAP7_75t_R g1990 ( 
.A(n_1712),
.Y(n_1990)
);

AND2x6_ASAP7_75t_L g1991 ( 
.A(n_1819),
.B(n_1823),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1805),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1884),
.Y(n_1993)
);

OR2x6_ASAP7_75t_L g1994 ( 
.A(n_1833),
.B(n_938),
.Y(n_1994)
);

INVx1_ASAP7_75t_SL g1995 ( 
.A(n_1780),
.Y(n_1995)
);

BUFx6f_ASAP7_75t_L g1996 ( 
.A(n_1752),
.Y(n_1996)
);

INVx1_ASAP7_75t_SL g1997 ( 
.A(n_1782),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1894),
.Y(n_1998)
);

INVx5_ASAP7_75t_L g1999 ( 
.A(n_1724),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1778),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_SL g2001 ( 
.A(n_1790),
.B(n_954),
.Y(n_2001)
);

INVx3_ASAP7_75t_L g2002 ( 
.A(n_1760),
.Y(n_2002)
);

BUFx6f_ASAP7_75t_L g2003 ( 
.A(n_1760),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1813),
.B(n_1703),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1786),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1792),
.B(n_1530),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_SL g2007 ( 
.A(n_1858),
.B(n_1728),
.Y(n_2007)
);

INVx3_ASAP7_75t_L g2008 ( 
.A(n_1760),
.Y(n_2008)
);

BUFx6f_ASAP7_75t_L g2009 ( 
.A(n_1888),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1911),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_SL g2011 ( 
.A(n_1874),
.B(n_992),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1825),
.B(n_1533),
.Y(n_2012)
);

INVx4_ASAP7_75t_L g2013 ( 
.A(n_1889),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1711),
.Y(n_2014)
);

AND2x6_ASAP7_75t_L g2015 ( 
.A(n_1824),
.B(n_796),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1829),
.B(n_1536),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1834),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1831),
.B(n_1463),
.Y(n_2018)
);

NOR2xp33_ASAP7_75t_L g2019 ( 
.A(n_1789),
.B(n_800),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1775),
.B(n_1465),
.Y(n_2020)
);

CKINVDCx20_ASAP7_75t_R g2021 ( 
.A(n_1725),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1721),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1850),
.B(n_1466),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_SL g2024 ( 
.A(n_1877),
.B(n_997),
.Y(n_2024)
);

AOI22xp33_ASAP7_75t_L g2025 ( 
.A1(n_1886),
.A2(n_1040),
.B1(n_1041),
.B2(n_1039),
.Y(n_2025)
);

INVx4_ASAP7_75t_SL g2026 ( 
.A(n_1888),
.Y(n_2026)
);

AND2x6_ASAP7_75t_L g2027 ( 
.A(n_1828),
.B(n_796),
.Y(n_2027)
);

AND2x2_ASAP7_75t_L g2028 ( 
.A(n_1878),
.B(n_1672),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1732),
.Y(n_2029)
);

NAND2xp33_ASAP7_75t_L g2030 ( 
.A(n_1885),
.B(n_815),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1837),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1835),
.B(n_1468),
.Y(n_2032)
);

AND2x4_ASAP7_75t_L g2033 ( 
.A(n_1838),
.B(n_1457),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1737),
.Y(n_2034)
);

INVx3_ASAP7_75t_L g2035 ( 
.A(n_1722),
.Y(n_2035)
);

AO22x2_ASAP7_75t_L g2036 ( 
.A1(n_1814),
.A2(n_944),
.B1(n_1019),
.B2(n_942),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1870),
.B(n_1685),
.Y(n_2037)
);

AND2x4_ASAP7_75t_L g2038 ( 
.A(n_1771),
.B(n_1459),
.Y(n_2038)
);

BUFx3_ASAP7_75t_L g2039 ( 
.A(n_1892),
.Y(n_2039)
);

BUFx6f_ASAP7_75t_L g2040 ( 
.A(n_1898),
.Y(n_2040)
);

NOR2xp33_ASAP7_75t_L g2041 ( 
.A(n_1875),
.B(n_801),
.Y(n_2041)
);

AND2x6_ASAP7_75t_L g2042 ( 
.A(n_1866),
.B(n_796),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1773),
.Y(n_2043)
);

INVx3_ASAP7_75t_L g2044 ( 
.A(n_1722),
.Y(n_2044)
);

INVxp67_ASAP7_75t_SL g2045 ( 
.A(n_1759),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_1740),
.Y(n_2046)
);

AO22x2_ASAP7_75t_L g2047 ( 
.A1(n_1847),
.A2(n_944),
.B1(n_1019),
.B2(n_942),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_SL g2048 ( 
.A(n_1797),
.B(n_1004),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1776),
.Y(n_2049)
);

CKINVDCx5p33_ASAP7_75t_R g2050 ( 
.A(n_1717),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1791),
.B(n_1648),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1777),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1759),
.Y(n_2053)
);

INVx3_ASAP7_75t_L g2054 ( 
.A(n_1787),
.Y(n_2054)
);

INVx1_ASAP7_75t_SL g2055 ( 
.A(n_1784),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1787),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1890),
.B(n_1484),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1745),
.Y(n_2058)
);

BUFx6f_ASAP7_75t_L g2059 ( 
.A(n_1893),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1795),
.Y(n_2060)
);

AND2x6_ASAP7_75t_L g2061 ( 
.A(n_1720),
.B(n_831),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1826),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1869),
.Y(n_2063)
);

AND2x4_ASAP7_75t_L g2064 ( 
.A(n_1746),
.B(n_1598),
.Y(n_2064)
);

INVx1_ASAP7_75t_SL g2065 ( 
.A(n_1801),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1750),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1869),
.Y(n_2067)
);

AND2x4_ASAP7_75t_L g2068 ( 
.A(n_1765),
.B(n_1602),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1769),
.Y(n_2069)
);

BUFx6f_ASAP7_75t_L g2070 ( 
.A(n_1896),
.Y(n_2070)
);

AND2x4_ASAP7_75t_L g2071 ( 
.A(n_1779),
.B(n_1603),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1800),
.Y(n_2072)
);

CKINVDCx5p33_ASAP7_75t_R g2073 ( 
.A(n_1714),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1811),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_1844),
.B(n_1485),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_1821),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1886),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_1872),
.B(n_1486),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_1852),
.Y(n_2079)
);

BUFx3_ASAP7_75t_L g2080 ( 
.A(n_1899),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_1863),
.B(n_1704),
.Y(n_2081)
);

INVx4_ASAP7_75t_L g2082 ( 
.A(n_1900),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_1807),
.B(n_1490),
.Y(n_2083)
);

AND2x4_ASAP7_75t_L g2084 ( 
.A(n_1901),
.B(n_1610),
.Y(n_2084)
);

INVx3_ASAP7_75t_L g2085 ( 
.A(n_1906),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1881),
.Y(n_2086)
);

AND2x4_ASAP7_75t_L g2087 ( 
.A(n_1727),
.B(n_1613),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1914),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1848),
.Y(n_2089)
);

AND2x4_ASAP7_75t_L g2090 ( 
.A(n_1738),
.B(n_1614),
.Y(n_2090)
);

BUFx2_ASAP7_75t_L g2091 ( 
.A(n_1808),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1918),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_SL g2093 ( 
.A(n_1942),
.B(n_1768),
.Y(n_2093)
);

NOR2xp33_ASAP7_75t_L g2094 ( 
.A(n_1965),
.B(n_1770),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1922),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_1923),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_SL g2097 ( 
.A(n_1953),
.B(n_1818),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_2016),
.B(n_1960),
.Y(n_2098)
);

INVx5_ASAP7_75t_L g2099 ( 
.A(n_2059),
.Y(n_2099)
);

CKINVDCx20_ASAP7_75t_R g2100 ( 
.A(n_2021),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1928),
.Y(n_2101)
);

AND2x4_ASAP7_75t_L g2102 ( 
.A(n_1984),
.B(n_1715),
.Y(n_2102)
);

NOR2xp67_ASAP7_75t_L g2103 ( 
.A(n_1984),
.B(n_1716),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1934),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1935),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1945),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1946),
.Y(n_2107)
);

INVx3_ASAP7_75t_L g2108 ( 
.A(n_1932),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1952),
.Y(n_2109)
);

BUFx6f_ASAP7_75t_L g2110 ( 
.A(n_1932),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1956),
.Y(n_2111)
);

AND2x4_ASAP7_75t_L g2112 ( 
.A(n_1936),
.B(n_1851),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_1929),
.Y(n_2113)
);

INVx1_ASAP7_75t_SL g2114 ( 
.A(n_1916),
.Y(n_2114)
);

INVxp67_ASAP7_75t_L g2115 ( 
.A(n_1947),
.Y(n_2115)
);

NAND2x1p5_ASAP7_75t_L g2116 ( 
.A(n_2040),
.B(n_1618),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_1938),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_1948),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1957),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_SL g2120 ( 
.A(n_1943),
.B(n_1820),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1959),
.Y(n_2121)
);

INVxp67_ASAP7_75t_L g2122 ( 
.A(n_1958),
.Y(n_2122)
);

NAND2x1p5_ASAP7_75t_L g2123 ( 
.A(n_2040),
.B(n_1624),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_2023),
.B(n_1856),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_1949),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1961),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_1950),
.Y(n_2127)
);

NAND2x1p5_ASAP7_75t_L g2128 ( 
.A(n_2085),
.B(n_1625),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_2018),
.B(n_1849),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_1951),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_2020),
.B(n_1861),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_1955),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1963),
.Y(n_2133)
);

INVx8_ASAP7_75t_L g2134 ( 
.A(n_1976),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_1930),
.B(n_1865),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_1967),
.Y(n_2136)
);

AO22x2_ASAP7_75t_L g2137 ( 
.A1(n_1940),
.A2(n_1063),
.B1(n_1072),
.B2(n_1051),
.Y(n_2137)
);

AO22x2_ASAP7_75t_L g2138 ( 
.A1(n_1995),
.A2(n_1063),
.B1(n_1072),
.B2(n_1051),
.Y(n_2138)
);

AO22x2_ASAP7_75t_L g2139 ( 
.A1(n_1997),
.A2(n_2065),
.B1(n_2055),
.B2(n_1926),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1966),
.Y(n_2140)
);

BUFx8_ASAP7_75t_L g2141 ( 
.A(n_2091),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_1931),
.B(n_1873),
.Y(n_2142)
);

AOI22xp33_ASAP7_75t_L g2143 ( 
.A1(n_1969),
.A2(n_1988),
.B1(n_1993),
.B2(n_1989),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_1968),
.Y(n_2144)
);

INVx3_ASAP7_75t_L g2145 ( 
.A(n_1937),
.Y(n_2145)
);

AND2x4_ASAP7_75t_L g2146 ( 
.A(n_2039),
.B(n_2080),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1998),
.Y(n_2147)
);

CKINVDCx5p33_ASAP7_75t_R g2148 ( 
.A(n_1917),
.Y(n_2148)
);

NAND2xp33_ASAP7_75t_L g2149 ( 
.A(n_1981),
.B(n_1729),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_1933),
.B(n_1761),
.Y(n_2150)
);

AOI22x1_ASAP7_75t_L g2151 ( 
.A1(n_2077),
.A2(n_1862),
.B1(n_1772),
.B2(n_1867),
.Y(n_2151)
);

BUFx2_ASAP7_75t_L g2152 ( 
.A(n_1987),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_1971),
.Y(n_2153)
);

AND2x4_ASAP7_75t_L g2154 ( 
.A(n_2059),
.B(n_1754),
.Y(n_2154)
);

AND2x4_ASAP7_75t_L g2155 ( 
.A(n_2070),
.B(n_1756),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2010),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1972),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1980),
.Y(n_2158)
);

BUFx10_ASAP7_75t_L g2159 ( 
.A(n_2041),
.Y(n_2159)
);

AOI22xp33_ASAP7_75t_L g2160 ( 
.A1(n_2025),
.A2(n_1077),
.B1(n_1081),
.B2(n_1054),
.Y(n_2160)
);

NOR2x1_ASAP7_75t_L g2161 ( 
.A(n_1925),
.B(n_1846),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1986),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1992),
.Y(n_2163)
);

BUFx6f_ASAP7_75t_L g2164 ( 
.A(n_1937),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2000),
.Y(n_2165)
);

BUFx6f_ASAP7_75t_L g2166 ( 
.A(n_1941),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_1915),
.B(n_1871),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_2005),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_2064),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2081),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_1921),
.B(n_1895),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2068),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2071),
.Y(n_2173)
);

INVx2_ASAP7_75t_SL g2174 ( 
.A(n_1983),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_2019),
.B(n_1751),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_2006),
.B(n_1912),
.Y(n_2176)
);

OAI22x1_ASAP7_75t_R g2177 ( 
.A1(n_1990),
.A2(n_1743),
.B1(n_1785),
.B2(n_1783),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_2014),
.Y(n_2178)
);

BUFx6f_ASAP7_75t_L g2179 ( 
.A(n_1941),
.Y(n_2179)
);

OR2x2_ASAP7_75t_L g2180 ( 
.A(n_1994),
.B(n_1753),
.Y(n_2180)
);

AO22x2_ASAP7_75t_L g2181 ( 
.A1(n_2089),
.A2(n_1267),
.B1(n_1272),
.B2(n_1239),
.Y(n_2181)
);

AND2x4_ASAP7_75t_L g2182 ( 
.A(n_2070),
.B(n_1713),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_2022),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_2012),
.B(n_1156),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_2029),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2051),
.B(n_1157),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2017),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2031),
.Y(n_2188)
);

BUFx8_ASAP7_75t_L g2189 ( 
.A(n_1924),
.Y(n_2189)
);

AOI22x1_ASAP7_75t_L g2190 ( 
.A1(n_2036),
.A2(n_1764),
.B1(n_1781),
.B2(n_1774),
.Y(n_2190)
);

NOR2x1_ASAP7_75t_L g2191 ( 
.A(n_1978),
.B(n_1076),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_2034),
.Y(n_2192)
);

BUFx6f_ASAP7_75t_L g2193 ( 
.A(n_1974),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_2046),
.Y(n_2194)
);

AND2x6_ASAP7_75t_L g2195 ( 
.A(n_2087),
.B(n_1174),
.Y(n_2195)
);

A2O1A1Ixp33_ASAP7_75t_L g2196 ( 
.A1(n_2057),
.A2(n_1741),
.B(n_1187),
.C(n_1220),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2043),
.Y(n_2197)
);

NOR2xp33_ASAP7_75t_L g2198 ( 
.A(n_1970),
.B(n_1730),
.Y(n_2198)
);

AND2x4_ASAP7_75t_L g2199 ( 
.A(n_2026),
.B(n_1718),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_2032),
.B(n_1176),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2049),
.Y(n_2201)
);

NOR2xp33_ASAP7_75t_L g2202 ( 
.A(n_1975),
.B(n_1905),
.Y(n_2202)
);

BUFx6f_ASAP7_75t_L g2203 ( 
.A(n_1974),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2052),
.Y(n_2204)
);

OAI221xp5_ASAP7_75t_L g2205 ( 
.A1(n_2078),
.A2(n_1977),
.B1(n_2088),
.B2(n_2086),
.C(n_2001),
.Y(n_2205)
);

OR2x2_ASAP7_75t_L g2206 ( 
.A(n_2050),
.B(n_1723),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2033),
.Y(n_2207)
);

OAI22xp5_ASAP7_75t_L g2208 ( 
.A1(n_2007),
.A2(n_1237),
.B1(n_1243),
.B2(n_1228),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2038),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2069),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_SL g2211 ( 
.A(n_2083),
.B(n_1767),
.Y(n_2211)
);

BUFx3_ASAP7_75t_L g2212 ( 
.A(n_1964),
.Y(n_2212)
);

AOI22xp5_ASAP7_75t_SL g2213 ( 
.A1(n_1973),
.A2(n_1088),
.B1(n_1093),
.B2(n_1084),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_2004),
.B(n_1735),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_SL g2215 ( 
.A(n_2028),
.B(n_1719),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_2058),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_2037),
.B(n_1739),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_2066),
.Y(n_2218)
);

INVx2_ASAP7_75t_L g2219 ( 
.A(n_2076),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_SL g2220 ( 
.A(n_2013),
.B(n_1794),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_1920),
.B(n_1498),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2072),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_1920),
.B(n_1505),
.Y(n_2223)
);

INVx3_ASAP7_75t_R g2224 ( 
.A(n_2090),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2074),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_1920),
.B(n_1515),
.Y(n_2226)
);

NOR2xp33_ASAP7_75t_L g2227 ( 
.A(n_2082),
.B(n_1108),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2053),
.Y(n_2228)
);

NAND3xp33_ASAP7_75t_L g2229 ( 
.A(n_1919),
.B(n_804),
.C(n_803),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2056),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_2075),
.B(n_1522),
.Y(n_2231)
);

CKINVDCx11_ASAP7_75t_R g2232 ( 
.A(n_1927),
.Y(n_2232)
);

CKINVDCx5p33_ASAP7_75t_R g2233 ( 
.A(n_2073),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_2060),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_2062),
.Y(n_2235)
);

BUFx3_ASAP7_75t_L g2236 ( 
.A(n_1985),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_2063),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2067),
.Y(n_2238)
);

INVx2_ASAP7_75t_SL g2239 ( 
.A(n_1954),
.Y(n_2239)
);

INVxp67_ASAP7_75t_L g2240 ( 
.A(n_2047),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_2035),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2045),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_2044),
.Y(n_2243)
);

AOI21xp5_ASAP7_75t_L g2244 ( 
.A1(n_2150),
.A2(n_2079),
.B(n_1944),
.Y(n_2244)
);

A2O1A1Ixp33_ASAP7_75t_L g2245 ( 
.A1(n_2094),
.A2(n_2030),
.B(n_2011),
.C(n_2024),
.Y(n_2245)
);

INVxp67_ASAP7_75t_L g2246 ( 
.A(n_2114),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_2176),
.B(n_1981),
.Y(n_2247)
);

AOI21xp5_ASAP7_75t_L g2248 ( 
.A1(n_2098),
.A2(n_2048),
.B(n_1962),
.Y(n_2248)
);

AOI21xp5_ASAP7_75t_L g2249 ( 
.A1(n_2131),
.A2(n_2084),
.B(n_2009),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2092),
.Y(n_2250)
);

AOI21xp5_ASAP7_75t_L g2251 ( 
.A1(n_2129),
.A2(n_2009),
.B(n_2003),
.Y(n_2251)
);

BUFx2_ASAP7_75t_L g2252 ( 
.A(n_2152),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2095),
.Y(n_2253)
);

A2O1A1Ixp33_ASAP7_75t_L g2254 ( 
.A1(n_2202),
.A2(n_1939),
.B(n_2054),
.C(n_2008),
.Y(n_2254)
);

BUFx6f_ASAP7_75t_L g2255 ( 
.A(n_2110),
.Y(n_2255)
);

AOI21xp5_ASAP7_75t_L g2256 ( 
.A1(n_2124),
.A2(n_2003),
.B(n_1996),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_2135),
.B(n_1981),
.Y(n_2257)
);

AOI21xp5_ASAP7_75t_L g2258 ( 
.A1(n_2142),
.A2(n_1996),
.B(n_2002),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2171),
.B(n_1991),
.Y(n_2259)
);

NOR2x1_ASAP7_75t_R g2260 ( 
.A(n_2099),
.B(n_1999),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2101),
.Y(n_2261)
);

AOI21x1_ASAP7_75t_L g2262 ( 
.A1(n_2186),
.A2(n_1631),
.B(n_1626),
.Y(n_2262)
);

OAI21xp5_ASAP7_75t_L g2263 ( 
.A1(n_2200),
.A2(n_1979),
.B(n_1991),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2104),
.Y(n_2264)
);

BUFx4f_ASAP7_75t_L g2265 ( 
.A(n_2199),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_2184),
.B(n_1991),
.Y(n_2266)
);

CKINVDCx5p33_ASAP7_75t_R g2267 ( 
.A(n_2148),
.Y(n_2267)
);

BUFx2_ASAP7_75t_L g2268 ( 
.A(n_2154),
.Y(n_2268)
);

BUFx6f_ASAP7_75t_L g2269 ( 
.A(n_2110),
.Y(n_2269)
);

O2A1O1Ixp5_ASAP7_75t_L g2270 ( 
.A1(n_2211),
.A2(n_2196),
.B(n_2231),
.C(n_2208),
.Y(n_2270)
);

INVx2_ASAP7_75t_L g2271 ( 
.A(n_2096),
.Y(n_2271)
);

AND2x4_ASAP7_75t_L g2272 ( 
.A(n_2099),
.B(n_1982),
.Y(n_2272)
);

OAI21xp33_ASAP7_75t_SL g2273 ( 
.A1(n_2143),
.A2(n_835),
.B(n_830),
.Y(n_2273)
);

AOI21xp5_ASAP7_75t_L g2274 ( 
.A1(n_2167),
.A2(n_862),
.B(n_831),
.Y(n_2274)
);

HB1xp67_ASAP7_75t_L g2275 ( 
.A(n_2146),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2170),
.B(n_1979),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_2105),
.B(n_1979),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_2106),
.B(n_2107),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_2109),
.B(n_2061),
.Y(n_2279)
);

AOI21xp5_ASAP7_75t_L g2280 ( 
.A1(n_2205),
.A2(n_862),
.B(n_831),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2111),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_2119),
.B(n_2061),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2121),
.B(n_2042),
.Y(n_2283)
);

AOI21xp5_ASAP7_75t_L g2284 ( 
.A1(n_2242),
.A2(n_862),
.B(n_831),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2126),
.Y(n_2285)
);

NOR2xp33_ASAP7_75t_L g2286 ( 
.A(n_2175),
.B(n_2115),
.Y(n_2286)
);

AOI21xp5_ASAP7_75t_L g2287 ( 
.A1(n_2093),
.A2(n_900),
.B(n_862),
.Y(n_2287)
);

AOI22xp5_ASAP7_75t_L g2288 ( 
.A1(n_2122),
.A2(n_2042),
.B1(n_1020),
.B2(n_1028),
.Y(n_2288)
);

AND2x4_ASAP7_75t_L g2289 ( 
.A(n_2174),
.B(n_1633),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_2217),
.B(n_1127),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2133),
.Y(n_2291)
);

OAI22xp5_ASAP7_75t_L g2292 ( 
.A1(n_2140),
.A2(n_1201),
.B1(n_1250),
.B2(n_1163),
.Y(n_2292)
);

AND2x2_ASAP7_75t_L g2293 ( 
.A(n_2214),
.B(n_1635),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2147),
.Y(n_2294)
);

OR2x6_ASAP7_75t_SL g2295 ( 
.A(n_2233),
.B(n_811),
.Y(n_2295)
);

AND2x2_ASAP7_75t_L g2296 ( 
.A(n_2227),
.B(n_1638),
.Y(n_2296)
);

AOI21xp5_ASAP7_75t_L g2297 ( 
.A1(n_2156),
.A2(n_960),
.B(n_900),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2187),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2158),
.B(n_1525),
.Y(n_2299)
);

BUFx2_ASAP7_75t_L g2300 ( 
.A(n_2155),
.Y(n_2300)
);

BUFx2_ASAP7_75t_L g2301 ( 
.A(n_2100),
.Y(n_2301)
);

NOR2xp33_ASAP7_75t_R g2302 ( 
.A(n_2134),
.B(n_2212),
.Y(n_2302)
);

NOR2xp33_ASAP7_75t_R g2303 ( 
.A(n_2134),
.B(n_1024),
.Y(n_2303)
);

AOI21xp5_ASAP7_75t_L g2304 ( 
.A1(n_2215),
.A2(n_960),
.B(n_900),
.Y(n_2304)
);

AOI21xp5_ASAP7_75t_L g2305 ( 
.A1(n_2113),
.A2(n_960),
.B(n_900),
.Y(n_2305)
);

NAND3xp33_ASAP7_75t_L g2306 ( 
.A(n_2229),
.B(n_814),
.C(n_813),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2188),
.Y(n_2307)
);

INVxp67_ASAP7_75t_L g2308 ( 
.A(n_2180),
.Y(n_2308)
);

AOI21xp5_ASAP7_75t_L g2309 ( 
.A1(n_2117),
.A2(n_2125),
.B(n_2118),
.Y(n_2309)
);

BUFx6f_ASAP7_75t_L g2310 ( 
.A(n_2164),
.Y(n_2310)
);

BUFx4f_ASAP7_75t_L g2311 ( 
.A(n_2182),
.Y(n_2311)
);

INVxp67_ASAP7_75t_SL g2312 ( 
.A(n_2164),
.Y(n_2312)
);

OAI21xp5_ASAP7_75t_L g2313 ( 
.A1(n_2162),
.A2(n_2015),
.B(n_2027),
.Y(n_2313)
);

AOI21xp5_ASAP7_75t_L g2314 ( 
.A1(n_2127),
.A2(n_1202),
.B(n_960),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2163),
.B(n_1528),
.Y(n_2315)
);

AOI21x1_ASAP7_75t_L g2316 ( 
.A1(n_2228),
.A2(n_1651),
.B(n_1644),
.Y(n_2316)
);

AOI21xp5_ASAP7_75t_L g2317 ( 
.A1(n_2130),
.A2(n_1265),
.B(n_1202),
.Y(n_2317)
);

AO21x1_ASAP7_75t_L g2318 ( 
.A1(n_2221),
.A2(n_2226),
.B(n_2223),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_SL g2319 ( 
.A(n_2159),
.B(n_1045),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_2165),
.B(n_1534),
.Y(n_2320)
);

OAI21xp5_ASAP7_75t_L g2321 ( 
.A1(n_2157),
.A2(n_2027),
.B(n_2015),
.Y(n_2321)
);

AOI21x1_ASAP7_75t_L g2322 ( 
.A1(n_2230),
.A2(n_1677),
.B(n_1659),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2197),
.Y(n_2323)
);

AOI21xp5_ASAP7_75t_L g2324 ( 
.A1(n_2132),
.A2(n_1265),
.B(n_1202),
.Y(n_2324)
);

AOI21xp5_ASAP7_75t_L g2325 ( 
.A1(n_2136),
.A2(n_2153),
.B(n_2144),
.Y(n_2325)
);

BUFx4f_ASAP7_75t_L g2326 ( 
.A(n_2102),
.Y(n_2326)
);

OAI22xp5_ASAP7_75t_L g2327 ( 
.A1(n_2201),
.A2(n_1111),
.B1(n_1113),
.B2(n_1104),
.Y(n_2327)
);

AOI21xp5_ASAP7_75t_L g2328 ( 
.A1(n_2168),
.A2(n_1265),
.B(n_1202),
.Y(n_2328)
);

OAI21xp5_ASAP7_75t_L g2329 ( 
.A1(n_2204),
.A2(n_2027),
.B(n_2015),
.Y(n_2329)
);

OR2x6_ASAP7_75t_SL g2330 ( 
.A(n_2206),
.B(n_828),
.Y(n_2330)
);

CKINVDCx8_ASAP7_75t_R g2331 ( 
.A(n_2112),
.Y(n_2331)
);

AOI21xp5_ASAP7_75t_L g2332 ( 
.A1(n_2149),
.A2(n_2097),
.B(n_2169),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_2178),
.Y(n_2333)
);

AOI21xp5_ASAP7_75t_L g2334 ( 
.A1(n_2120),
.A2(n_1265),
.B(n_1126),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_SL g2335 ( 
.A(n_2198),
.B(n_1116),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2210),
.Y(n_2336)
);

OAI22xp5_ASAP7_75t_L g2337 ( 
.A1(n_2160),
.A2(n_1138),
.B1(n_1145),
.B2(n_1133),
.Y(n_2337)
);

NOR2xp33_ASAP7_75t_L g2338 ( 
.A(n_2240),
.B(n_829),
.Y(n_2338)
);

AND2x4_ASAP7_75t_L g2339 ( 
.A(n_2241),
.B(n_1678),
.Y(n_2339)
);

CKINVDCx20_ASAP7_75t_R g2340 ( 
.A(n_2141),
.Y(n_2340)
);

AOI21xp5_ASAP7_75t_L g2341 ( 
.A1(n_2183),
.A2(n_1152),
.B(n_1151),
.Y(n_2341)
);

AOI21xp5_ASAP7_75t_L g2342 ( 
.A1(n_2185),
.A2(n_1170),
.B(n_1160),
.Y(n_2342)
);

OAI21xp33_ASAP7_75t_L g2343 ( 
.A1(n_2191),
.A2(n_2138),
.B(n_2137),
.Y(n_2343)
);

AOI21x1_ASAP7_75t_L g2344 ( 
.A1(n_2238),
.A2(n_1684),
.B(n_1679),
.Y(n_2344)
);

AOI21xp5_ASAP7_75t_L g2345 ( 
.A1(n_2192),
.A2(n_1312),
.B(n_1311),
.Y(n_2345)
);

OAI22xp5_ASAP7_75t_L g2346 ( 
.A1(n_2234),
.A2(n_1189),
.B1(n_1191),
.B2(n_1188),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2194),
.B(n_1687),
.Y(n_2347)
);

AOI21xp5_ASAP7_75t_L g2348 ( 
.A1(n_2216),
.A2(n_2219),
.B(n_2218),
.Y(n_2348)
);

AND2x4_ASAP7_75t_L g2349 ( 
.A(n_2243),
.B(n_1689),
.Y(n_2349)
);

HB1xp67_ASAP7_75t_L g2350 ( 
.A(n_2166),
.Y(n_2350)
);

AO21x1_ASAP7_75t_L g2351 ( 
.A1(n_2222),
.A2(n_884),
.B(n_879),
.Y(n_2351)
);

OAI22xp5_ASAP7_75t_L g2352 ( 
.A1(n_2235),
.A2(n_2237),
.B1(n_2225),
.B2(n_2151),
.Y(n_2352)
);

OR2x2_ASAP7_75t_L g2353 ( 
.A(n_2239),
.B(n_1691),
.Y(n_2353)
);

AOI22xp5_ASAP7_75t_L g2354 ( 
.A1(n_2195),
.A2(n_1197),
.B1(n_1198),
.B2(n_1193),
.Y(n_2354)
);

AOI21x1_ASAP7_75t_L g2355 ( 
.A1(n_2181),
.A2(n_1699),
.B(n_908),
.Y(n_2355)
);

AOI21xp5_ASAP7_75t_L g2356 ( 
.A1(n_2172),
.A2(n_1303),
.B(n_1297),
.Y(n_2356)
);

INVx3_ASAP7_75t_L g2357 ( 
.A(n_2179),
.Y(n_2357)
);

AND2x2_ASAP7_75t_L g2358 ( 
.A(n_2290),
.B(n_2139),
.Y(n_2358)
);

NOR2xp67_ASAP7_75t_SL g2359 ( 
.A(n_2267),
.B(n_2236),
.Y(n_2359)
);

INVx2_ASAP7_75t_L g2360 ( 
.A(n_2250),
.Y(n_2360)
);

INVxp67_ASAP7_75t_L g2361 ( 
.A(n_2252),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_SL g2362 ( 
.A(n_2286),
.B(n_2161),
.Y(n_2362)
);

CKINVDCx5p33_ASAP7_75t_R g2363 ( 
.A(n_2302),
.Y(n_2363)
);

OAI22xp5_ASAP7_75t_L g2364 ( 
.A1(n_2278),
.A2(n_2173),
.B1(n_2190),
.B2(n_2207),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_2296),
.B(n_2195),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_2253),
.B(n_2195),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_SL g2367 ( 
.A(n_2246),
.B(n_2213),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_SL g2368 ( 
.A(n_2311),
.B(n_2179),
.Y(n_2368)
);

OAI22xp5_ASAP7_75t_L g2369 ( 
.A1(n_2245),
.A2(n_2209),
.B1(n_2108),
.B2(n_2145),
.Y(n_2369)
);

O2A1O1Ixp33_ASAP7_75t_SL g2370 ( 
.A1(n_2254),
.A2(n_2220),
.B(n_912),
.C(n_920),
.Y(n_2370)
);

BUFx2_ASAP7_75t_L g2371 ( 
.A(n_2275),
.Y(n_2371)
);

OAI21xp5_ASAP7_75t_L g2372 ( 
.A1(n_2270),
.A2(n_2128),
.B(n_2103),
.Y(n_2372)
);

CKINVDCx14_ASAP7_75t_R g2373 ( 
.A(n_2340),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2261),
.Y(n_2374)
);

OAI21xp5_ASAP7_75t_L g2375 ( 
.A1(n_2248),
.A2(n_2123),
.B(n_2116),
.Y(n_2375)
);

CKINVDCx5p33_ASAP7_75t_R g2376 ( 
.A(n_2301),
.Y(n_2376)
);

AOI21xp5_ASAP7_75t_L g2377 ( 
.A1(n_2244),
.A2(n_2203),
.B(n_2193),
.Y(n_2377)
);

A2O1A1Ixp33_ASAP7_75t_SL g2378 ( 
.A1(n_2263),
.A2(n_1516),
.B(n_1526),
.C(n_1506),
.Y(n_2378)
);

NAND2x1p5_ASAP7_75t_L g2379 ( 
.A(n_2265),
.B(n_2193),
.Y(n_2379)
);

NOR2xp67_ASAP7_75t_L g2380 ( 
.A(n_2306),
.B(n_2224),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2264),
.Y(n_2381)
);

BUFx4f_ASAP7_75t_L g2382 ( 
.A(n_2255),
.Y(n_2382)
);

AOI21xp5_ASAP7_75t_L g2383 ( 
.A1(n_2266),
.A2(n_1246),
.B(n_1223),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_2281),
.B(n_2189),
.Y(n_2384)
);

NOR2xp33_ASAP7_75t_L g2385 ( 
.A(n_2292),
.B(n_2232),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2285),
.Y(n_2386)
);

BUFx2_ASAP7_75t_L g2387 ( 
.A(n_2255),
.Y(n_2387)
);

BUFx6f_ASAP7_75t_L g2388 ( 
.A(n_2269),
.Y(n_2388)
);

A2O1A1Ixp33_ASAP7_75t_SL g2389 ( 
.A1(n_2338),
.A2(n_1527),
.B(n_922),
.C(n_927),
.Y(n_2389)
);

AOI21xp5_ASAP7_75t_L g2390 ( 
.A1(n_2257),
.A2(n_1262),
.B(n_1245),
.Y(n_2390)
);

NOR2xp33_ASAP7_75t_L g2391 ( 
.A(n_2343),
.B(n_833),
.Y(n_2391)
);

AOI22xp5_ASAP7_75t_L g2392 ( 
.A1(n_2308),
.A2(n_1281),
.B1(n_1294),
.B2(n_1266),
.Y(n_2392)
);

AOI21xp5_ASAP7_75t_L g2393 ( 
.A1(n_2259),
.A2(n_1296),
.B(n_936),
.Y(n_2393)
);

A2O1A1Ixp33_ASAP7_75t_L g2394 ( 
.A1(n_2332),
.A2(n_941),
.B(n_943),
.C(n_915),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_2291),
.B(n_948),
.Y(n_2395)
);

NAND2x1p5_ASAP7_75t_L g2396 ( 
.A(n_2269),
.B(n_2177),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_2294),
.B(n_950),
.Y(n_2397)
);

BUFx12f_ASAP7_75t_L g2398 ( 
.A(n_2272),
.Y(n_2398)
);

AOI21xp5_ASAP7_75t_L g2399 ( 
.A1(n_2247),
.A2(n_961),
.B(n_957),
.Y(n_2399)
);

AOI21xp5_ASAP7_75t_L g2400 ( 
.A1(n_2249),
.A2(n_966),
.B(n_963),
.Y(n_2400)
);

OR2x6_ASAP7_75t_L g2401 ( 
.A(n_2272),
.B(n_2268),
.Y(n_2401)
);

INVx2_ASAP7_75t_SL g2402 ( 
.A(n_2269),
.Y(n_2402)
);

OAI22xp5_ASAP7_75t_L g2403 ( 
.A1(n_2298),
.A2(n_2323),
.B1(n_2307),
.B2(n_2336),
.Y(n_2403)
);

CKINVDCx5p33_ASAP7_75t_R g2404 ( 
.A(n_2331),
.Y(n_2404)
);

AOI21x1_ASAP7_75t_L g2405 ( 
.A1(n_2262),
.A2(n_2318),
.B(n_2280),
.Y(n_2405)
);

INVx2_ASAP7_75t_L g2406 ( 
.A(n_2271),
.Y(n_2406)
);

AOI21x1_ASAP7_75t_L g2407 ( 
.A1(n_2316),
.A2(n_988),
.B(n_985),
.Y(n_2407)
);

AOI21xp5_ASAP7_75t_L g2408 ( 
.A1(n_2251),
.A2(n_994),
.B(n_990),
.Y(n_2408)
);

INVx3_ASAP7_75t_L g2409 ( 
.A(n_2310),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2333),
.Y(n_2410)
);

OAI22xp5_ASAP7_75t_SL g2411 ( 
.A1(n_2300),
.A2(n_845),
.B1(n_846),
.B2(n_843),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2293),
.B(n_995),
.Y(n_2412)
);

O2A1O1Ixp33_ASAP7_75t_SL g2413 ( 
.A1(n_2277),
.A2(n_996),
.B(n_1000),
.C(n_998),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_L g2414 ( 
.A(n_2335),
.B(n_1007),
.Y(n_2414)
);

CKINVDCx6p67_ASAP7_75t_R g2415 ( 
.A(n_2310),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2347),
.Y(n_2416)
);

HB1xp67_ASAP7_75t_L g2417 ( 
.A(n_2350),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2299),
.Y(n_2418)
);

INVx4_ASAP7_75t_L g2419 ( 
.A(n_2310),
.Y(n_2419)
);

OAI22xp5_ASAP7_75t_L g2420 ( 
.A1(n_2276),
.A2(n_851),
.B1(n_852),
.B2(n_850),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_2256),
.B(n_1014),
.Y(n_2421)
);

BUFx2_ASAP7_75t_L g2422 ( 
.A(n_2357),
.Y(n_2422)
);

AO21x1_ASAP7_75t_L g2423 ( 
.A1(n_2352),
.A2(n_1027),
.B(n_1018),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_2258),
.B(n_1035),
.Y(n_2424)
);

INVx5_ASAP7_75t_L g2425 ( 
.A(n_2289),
.Y(n_2425)
);

AOI21xp5_ASAP7_75t_L g2426 ( 
.A1(n_2309),
.A2(n_1048),
.B(n_1043),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2315),
.Y(n_2427)
);

AOI21xp5_ASAP7_75t_L g2428 ( 
.A1(n_2325),
.A2(n_1080),
.B(n_1058),
.Y(n_2428)
);

INVx3_ASAP7_75t_L g2429 ( 
.A(n_2326),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_2273),
.B(n_2279),
.Y(n_2430)
);

A2O1A1Ixp33_ASAP7_75t_L g2431 ( 
.A1(n_2348),
.A2(n_1096),
.B(n_1098),
.C(n_1091),
.Y(n_2431)
);

OR2x2_ASAP7_75t_L g2432 ( 
.A(n_2353),
.B(n_856),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2320),
.Y(n_2433)
);

NOR2xp33_ASAP7_75t_L g2434 ( 
.A(n_2319),
.B(n_857),
.Y(n_2434)
);

BUFx12f_ASAP7_75t_L g2435 ( 
.A(n_2339),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2339),
.Y(n_2436)
);

INVx3_ASAP7_75t_L g2437 ( 
.A(n_2349),
.Y(n_2437)
);

OAI21xp33_ASAP7_75t_SL g2438 ( 
.A1(n_2282),
.A2(n_2283),
.B(n_2329),
.Y(n_2438)
);

O2A1O1Ixp33_ASAP7_75t_SL g2439 ( 
.A1(n_2313),
.A2(n_1121),
.B(n_1122),
.C(n_1120),
.Y(n_2439)
);

CKINVDCx5p33_ASAP7_75t_R g2440 ( 
.A(n_2303),
.Y(n_2440)
);

OAI21x1_ASAP7_75t_L g2441 ( 
.A1(n_2322),
.A2(n_1295),
.B(n_1130),
.Y(n_2441)
);

CKINVDCx5p33_ASAP7_75t_R g2442 ( 
.A(n_2330),
.Y(n_2442)
);

INVx3_ASAP7_75t_L g2443 ( 
.A(n_2349),
.Y(n_2443)
);

BUFx12f_ASAP7_75t_L g2444 ( 
.A(n_2260),
.Y(n_2444)
);

BUFx3_ASAP7_75t_L g2445 ( 
.A(n_2295),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2344),
.Y(n_2446)
);

OAI21x1_ASAP7_75t_L g2447 ( 
.A1(n_2284),
.A2(n_1135),
.B(n_1129),
.Y(n_2447)
);

OR2x2_ASAP7_75t_L g2448 ( 
.A(n_2312),
.B(n_868),
.Y(n_2448)
);

OAI21x1_ASAP7_75t_L g2449 ( 
.A1(n_2304),
.A2(n_1166),
.B(n_1162),
.Y(n_2449)
);

AOI21xp5_ASAP7_75t_L g2450 ( 
.A1(n_2274),
.A2(n_1179),
.B(n_1177),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2351),
.Y(n_2451)
);

BUFx2_ASAP7_75t_L g2452 ( 
.A(n_2354),
.Y(n_2452)
);

INVx4_ASAP7_75t_L g2453 ( 
.A(n_2355),
.Y(n_2453)
);

O2A1O1Ixp33_ASAP7_75t_L g2454 ( 
.A1(n_2327),
.A2(n_1181),
.B(n_1203),
.C(n_1180),
.Y(n_2454)
);

AOI21xp5_ASAP7_75t_L g2455 ( 
.A1(n_2287),
.A2(n_1225),
.B(n_1214),
.Y(n_2455)
);

INVx3_ASAP7_75t_L g2456 ( 
.A(n_2356),
.Y(n_2456)
);

INVx2_ASAP7_75t_L g2457 ( 
.A(n_2321),
.Y(n_2457)
);

AOI22xp5_ASAP7_75t_L g2458 ( 
.A1(n_2346),
.A2(n_2337),
.B1(n_2288),
.B2(n_2341),
.Y(n_2458)
);

AND2x2_ASAP7_75t_L g2459 ( 
.A(n_2334),
.B(n_872),
.Y(n_2459)
);

OAI22xp5_ASAP7_75t_L g2460 ( 
.A1(n_2342),
.A2(n_874),
.B1(n_877),
.B2(n_873),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_L g2461 ( 
.A(n_2345),
.B(n_1226),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_L g2462 ( 
.A(n_2416),
.B(n_878),
.Y(n_2462)
);

INVx4_ASAP7_75t_L g2463 ( 
.A(n_2382),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2360),
.Y(n_2464)
);

INVx8_ASAP7_75t_L g2465 ( 
.A(n_2398),
.Y(n_2465)
);

BUFx12f_ASAP7_75t_L g2466 ( 
.A(n_2404),
.Y(n_2466)
);

BUFx12f_ASAP7_75t_L g2467 ( 
.A(n_2363),
.Y(n_2467)
);

INVx6_ASAP7_75t_SL g2468 ( 
.A(n_2401),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2374),
.Y(n_2469)
);

INVx3_ASAP7_75t_L g2470 ( 
.A(n_2379),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2381),
.Y(n_2471)
);

BUFx6f_ASAP7_75t_L g2472 ( 
.A(n_2388),
.Y(n_2472)
);

BUFx2_ASAP7_75t_R g2473 ( 
.A(n_2440),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2386),
.Y(n_2474)
);

OR2x6_ASAP7_75t_L g2475 ( 
.A(n_2401),
.B(n_2297),
.Y(n_2475)
);

CKINVDCx14_ASAP7_75t_R g2476 ( 
.A(n_2373),
.Y(n_2476)
);

NAND2x1p5_ASAP7_75t_L g2477 ( 
.A(n_2425),
.B(n_2328),
.Y(n_2477)
);

INVx2_ASAP7_75t_L g2478 ( 
.A(n_2406),
.Y(n_2478)
);

BUFx6f_ASAP7_75t_L g2479 ( 
.A(n_2388),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2403),
.Y(n_2480)
);

CKINVDCx11_ASAP7_75t_R g2481 ( 
.A(n_2444),
.Y(n_2481)
);

BUFx2_ASAP7_75t_SL g2482 ( 
.A(n_2425),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2410),
.Y(n_2483)
);

INVx1_ASAP7_75t_SL g2484 ( 
.A(n_2371),
.Y(n_2484)
);

CKINVDCx11_ASAP7_75t_R g2485 ( 
.A(n_2445),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2436),
.Y(n_2486)
);

BUFx4_ASAP7_75t_SL g2487 ( 
.A(n_2376),
.Y(n_2487)
);

BUFx4f_ASAP7_75t_L g2488 ( 
.A(n_2415),
.Y(n_2488)
);

CKINVDCx16_ASAP7_75t_R g2489 ( 
.A(n_2435),
.Y(n_2489)
);

INVx1_ASAP7_75t_SL g2490 ( 
.A(n_2417),
.Y(n_2490)
);

INVx3_ASAP7_75t_L g2491 ( 
.A(n_2429),
.Y(n_2491)
);

BUFx2_ASAP7_75t_L g2492 ( 
.A(n_2361),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2395),
.Y(n_2493)
);

INVx5_ASAP7_75t_L g2494 ( 
.A(n_2388),
.Y(n_2494)
);

BUFx3_ASAP7_75t_L g2495 ( 
.A(n_2387),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_L g2496 ( 
.A(n_2418),
.B(n_882),
.Y(n_2496)
);

INVx3_ASAP7_75t_L g2497 ( 
.A(n_2419),
.Y(n_2497)
);

INVx8_ASAP7_75t_L g2498 ( 
.A(n_2425),
.Y(n_2498)
);

NAND2x1p5_ASAP7_75t_L g2499 ( 
.A(n_2359),
.B(n_2305),
.Y(n_2499)
);

BUFx2_ASAP7_75t_SL g2500 ( 
.A(n_2402),
.Y(n_2500)
);

BUFx6f_ASAP7_75t_L g2501 ( 
.A(n_2422),
.Y(n_2501)
);

BUFx2_ASAP7_75t_R g2502 ( 
.A(n_2367),
.Y(n_2502)
);

INVxp67_ASAP7_75t_SL g2503 ( 
.A(n_2437),
.Y(n_2503)
);

INVx8_ASAP7_75t_L g2504 ( 
.A(n_2409),
.Y(n_2504)
);

INVx3_ASAP7_75t_L g2505 ( 
.A(n_2443),
.Y(n_2505)
);

BUFx2_ASAP7_75t_SL g2506 ( 
.A(n_2380),
.Y(n_2506)
);

CKINVDCx14_ASAP7_75t_R g2507 ( 
.A(n_2442),
.Y(n_2507)
);

INVx3_ASAP7_75t_L g2508 ( 
.A(n_2396),
.Y(n_2508)
);

INVx2_ASAP7_75t_L g2509 ( 
.A(n_2427),
.Y(n_2509)
);

INVx4_ASAP7_75t_L g2510 ( 
.A(n_2448),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_2433),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2397),
.Y(n_2512)
);

BUFx4f_ASAP7_75t_L g2513 ( 
.A(n_2358),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2421),
.Y(n_2514)
);

BUFx2_ASAP7_75t_SL g2515 ( 
.A(n_2368),
.Y(n_2515)
);

BUFx3_ASAP7_75t_L g2516 ( 
.A(n_2384),
.Y(n_2516)
);

NAND2x1p5_ASAP7_75t_L g2517 ( 
.A(n_2362),
.B(n_2314),
.Y(n_2517)
);

CKINVDCx11_ASAP7_75t_R g2518 ( 
.A(n_2452),
.Y(n_2518)
);

NAND2x1_ASAP7_75t_L g2519 ( 
.A(n_2456),
.B(n_2317),
.Y(n_2519)
);

BUFx6f_ASAP7_75t_L g2520 ( 
.A(n_2366),
.Y(n_2520)
);

BUFx3_ASAP7_75t_L g2521 ( 
.A(n_2385),
.Y(n_2521)
);

INVx2_ASAP7_75t_SL g2522 ( 
.A(n_2432),
.Y(n_2522)
);

BUFx12f_ASAP7_75t_L g2523 ( 
.A(n_2453),
.Y(n_2523)
);

BUFx2_ASAP7_75t_L g2524 ( 
.A(n_2365),
.Y(n_2524)
);

BUFx3_ASAP7_75t_L g2525 ( 
.A(n_2412),
.Y(n_2525)
);

INVx3_ASAP7_75t_L g2526 ( 
.A(n_2459),
.Y(n_2526)
);

INVx5_ASAP7_75t_L g2527 ( 
.A(n_2453),
.Y(n_2527)
);

INVx2_ASAP7_75t_L g2528 ( 
.A(n_2446),
.Y(n_2528)
);

INVx5_ASAP7_75t_L g2529 ( 
.A(n_2457),
.Y(n_2529)
);

INVx1_ASAP7_75t_SL g2530 ( 
.A(n_2411),
.Y(n_2530)
);

INVx2_ASAP7_75t_SL g2531 ( 
.A(n_2414),
.Y(n_2531)
);

BUFx3_ASAP7_75t_L g2532 ( 
.A(n_2434),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2424),
.Y(n_2533)
);

INVx2_ASAP7_75t_SL g2534 ( 
.A(n_2369),
.Y(n_2534)
);

INVx3_ASAP7_75t_L g2535 ( 
.A(n_2451),
.Y(n_2535)
);

BUFx6f_ASAP7_75t_L g2536 ( 
.A(n_2461),
.Y(n_2536)
);

NAND2x1p5_ASAP7_75t_L g2537 ( 
.A(n_2377),
.B(n_2324),
.Y(n_2537)
);

BUFx6f_ASAP7_75t_SL g2538 ( 
.A(n_2370),
.Y(n_2538)
);

BUFx3_ASAP7_75t_L g2539 ( 
.A(n_2391),
.Y(n_2539)
);

NOR2xp67_ASAP7_75t_SL g2540 ( 
.A(n_2372),
.B(n_887),
.Y(n_2540)
);

INVx4_ASAP7_75t_L g2541 ( 
.A(n_2364),
.Y(n_2541)
);

BUFx3_ASAP7_75t_L g2542 ( 
.A(n_2392),
.Y(n_2542)
);

NAND2x1p5_ASAP7_75t_L g2543 ( 
.A(n_2458),
.B(n_1238),
.Y(n_2543)
);

INVx3_ASAP7_75t_L g2544 ( 
.A(n_2449),
.Y(n_2544)
);

INVx5_ASAP7_75t_L g2545 ( 
.A(n_2389),
.Y(n_2545)
);

OR2x6_ASAP7_75t_L g2546 ( 
.A(n_2375),
.B(n_1249),
.Y(n_2546)
);

BUFx6f_ASAP7_75t_L g2547 ( 
.A(n_2430),
.Y(n_2547)
);

NOR2xp33_ASAP7_75t_L g2548 ( 
.A(n_2539),
.B(n_2532),
.Y(n_2548)
);

BUFx2_ASAP7_75t_SL g2549 ( 
.A(n_2529),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2478),
.Y(n_2550)
);

AO21x2_ASAP7_75t_L g2551 ( 
.A1(n_2528),
.A2(n_2405),
.B(n_2423),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2469),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2493),
.B(n_2399),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_2512),
.B(n_2394),
.Y(n_2554)
);

AO32x2_ASAP7_75t_L g2555 ( 
.A1(n_2541),
.A2(n_2420),
.A3(n_2460),
.B1(n_2438),
.B2(n_2454),
.Y(n_2555)
);

OA21x2_ASAP7_75t_L g2556 ( 
.A1(n_2480),
.A2(n_2441),
.B(n_2447),
.Y(n_2556)
);

OAI21x1_ASAP7_75t_L g2557 ( 
.A1(n_2519),
.A2(n_2407),
.B(n_2426),
.Y(n_2557)
);

NAND2xp5_ASAP7_75t_L g2558 ( 
.A(n_2509),
.B(n_2400),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_L g2559 ( 
.A(n_2511),
.B(n_2431),
.Y(n_2559)
);

INVxp67_ASAP7_75t_SL g2560 ( 
.A(n_2547),
.Y(n_2560)
);

INVx1_ASAP7_75t_SL g2561 ( 
.A(n_2484),
.Y(n_2561)
);

OAI21x1_ASAP7_75t_L g2562 ( 
.A1(n_2537),
.A2(n_2428),
.B(n_2408),
.Y(n_2562)
);

NAND2x1p5_ASAP7_75t_L g2563 ( 
.A(n_2529),
.B(n_2393),
.Y(n_2563)
);

BUFx12f_ASAP7_75t_L g2564 ( 
.A(n_2481),
.Y(n_2564)
);

INVx1_ASAP7_75t_SL g2565 ( 
.A(n_2518),
.Y(n_2565)
);

OAI21x1_ASAP7_75t_L g2566 ( 
.A1(n_2544),
.A2(n_2450),
.B(n_2455),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2471),
.Y(n_2567)
);

OAI21x1_ASAP7_75t_L g2568 ( 
.A1(n_2517),
.A2(n_2390),
.B(n_2383),
.Y(n_2568)
);

OR2x2_ASAP7_75t_L g2569 ( 
.A(n_2524),
.B(n_2378),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2474),
.Y(n_2570)
);

OAI21x1_ASAP7_75t_L g2571 ( 
.A1(n_2535),
.A2(n_2439),
.B(n_2413),
.Y(n_2571)
);

AO31x2_ASAP7_75t_L g2572 ( 
.A1(n_2533),
.A2(n_1255),
.A3(n_1285),
.B(n_1256),
.Y(n_2572)
);

NOR2xp33_ASAP7_75t_L g2573 ( 
.A(n_2542),
.B(n_2530),
.Y(n_2573)
);

OAI21x1_ASAP7_75t_L g2574 ( 
.A1(n_2499),
.A2(n_1046),
.B(n_815),
.Y(n_2574)
);

OAI21x1_ASAP7_75t_L g2575 ( 
.A1(n_2477),
.A2(n_1046),
.B(n_815),
.Y(n_2575)
);

OAI21x1_ASAP7_75t_L g2576 ( 
.A1(n_2483),
.A2(n_1046),
.B(n_815),
.Y(n_2576)
);

BUFx2_ASAP7_75t_L g2577 ( 
.A(n_2468),
.Y(n_2577)
);

OAI21x1_ASAP7_75t_L g2578 ( 
.A1(n_2526),
.A2(n_1046),
.B(n_815),
.Y(n_2578)
);

INVx5_ASAP7_75t_L g2579 ( 
.A(n_2463),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2464),
.Y(n_2580)
);

NAND2x1_ASAP7_75t_L g2581 ( 
.A(n_2547),
.B(n_598),
.Y(n_2581)
);

OAI21x1_ASAP7_75t_L g2582 ( 
.A1(n_2543),
.A2(n_603),
.B(n_599),
.Y(n_2582)
);

OAI21x1_ASAP7_75t_L g2583 ( 
.A1(n_2514),
.A2(n_605),
.B(n_604),
.Y(n_2583)
);

OAI221xp5_ASAP7_75t_L g2584 ( 
.A1(n_2525),
.A2(n_892),
.B1(n_894),
.B2(n_891),
.C(n_890),
.Y(n_2584)
);

INVx1_ASAP7_75t_SL g2585 ( 
.A(n_2490),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2486),
.Y(n_2586)
);

BUFx6f_ASAP7_75t_L g2587 ( 
.A(n_2488),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2503),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2520),
.Y(n_2589)
);

OA21x2_ASAP7_75t_L g2590 ( 
.A1(n_2534),
.A2(n_899),
.B(n_895),
.Y(n_2590)
);

OAI21x1_ASAP7_75t_L g2591 ( 
.A1(n_2505),
.A2(n_609),
.B(n_607),
.Y(n_2591)
);

NOR2x1_ASAP7_75t_SL g2592 ( 
.A(n_2546),
.B(n_611),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2520),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2527),
.Y(n_2594)
);

OAI21x1_ASAP7_75t_L g2595 ( 
.A1(n_2540),
.A2(n_613),
.B(n_612),
.Y(n_2595)
);

HB1xp67_ASAP7_75t_L g2596 ( 
.A(n_2536),
.Y(n_2596)
);

OAI21x1_ASAP7_75t_L g2597 ( 
.A1(n_2527),
.A2(n_615),
.B(n_614),
.Y(n_2597)
);

HB1xp67_ASAP7_75t_L g2598 ( 
.A(n_2536),
.Y(n_2598)
);

AO21x2_ASAP7_75t_L g2599 ( 
.A1(n_2496),
.A2(n_909),
.B(n_904),
.Y(n_2599)
);

INVx2_ASAP7_75t_SL g2600 ( 
.A(n_2487),
.Y(n_2600)
);

OR2x2_ASAP7_75t_L g2601 ( 
.A(n_2492),
.B(n_2),
.Y(n_2601)
);

OAI21x1_ASAP7_75t_L g2602 ( 
.A1(n_2508),
.A2(n_618),
.B(n_616),
.Y(n_2602)
);

OA21x2_ASAP7_75t_L g2603 ( 
.A1(n_2462),
.A2(n_924),
.B(n_916),
.Y(n_2603)
);

OAI21x1_ASAP7_75t_L g2604 ( 
.A1(n_2523),
.A2(n_620),
.B(n_619),
.Y(n_2604)
);

AND2x2_ASAP7_75t_L g2605 ( 
.A(n_2513),
.B(n_622),
.Y(n_2605)
);

AO21x2_ASAP7_75t_L g2606 ( 
.A1(n_2545),
.A2(n_926),
.B(n_925),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2515),
.Y(n_2607)
);

CKINVDCx16_ASAP7_75t_R g2608 ( 
.A(n_2489),
.Y(n_2608)
);

AO21x2_ASAP7_75t_L g2609 ( 
.A1(n_2576),
.A2(n_2538),
.B(n_2545),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2552),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2567),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2570),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_2580),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2586),
.Y(n_2614)
);

INVx2_ASAP7_75t_L g2615 ( 
.A(n_2550),
.Y(n_2615)
);

CKINVDCx5p33_ASAP7_75t_R g2616 ( 
.A(n_2564),
.Y(n_2616)
);

BUFx2_ASAP7_75t_L g2617 ( 
.A(n_2569),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2588),
.Y(n_2618)
);

INVx2_ASAP7_75t_L g2619 ( 
.A(n_2589),
.Y(n_2619)
);

OAI21x1_ASAP7_75t_L g2620 ( 
.A1(n_2557),
.A2(n_2497),
.B(n_2470),
.Y(n_2620)
);

INVx2_ASAP7_75t_L g2621 ( 
.A(n_2593),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_L g2622 ( 
.A(n_2560),
.B(n_2531),
.Y(n_2622)
);

NAND2x1p5_ASAP7_75t_L g2623 ( 
.A(n_2579),
.B(n_2494),
.Y(n_2623)
);

AND2x4_ASAP7_75t_L g2624 ( 
.A(n_2607),
.B(n_2495),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2572),
.Y(n_2625)
);

AOI21x1_ASAP7_75t_L g2626 ( 
.A1(n_2553),
.A2(n_2475),
.B(n_2522),
.Y(n_2626)
);

HB1xp67_ASAP7_75t_L g2627 ( 
.A(n_2596),
.Y(n_2627)
);

BUFx6f_ASAP7_75t_L g2628 ( 
.A(n_2587),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2594),
.Y(n_2629)
);

INVxp67_ASAP7_75t_L g2630 ( 
.A(n_2585),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2551),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_L g2632 ( 
.A(n_2598),
.B(n_2510),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2558),
.Y(n_2633)
);

BUFx2_ASAP7_75t_L g2634 ( 
.A(n_2574),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2549),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2559),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_2578),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2554),
.Y(n_2638)
);

BUFx3_ASAP7_75t_L g2639 ( 
.A(n_2577),
.Y(n_2639)
);

INVx2_ASAP7_75t_L g2640 ( 
.A(n_2575),
.Y(n_2640)
);

BUFx8_ASAP7_75t_SL g2641 ( 
.A(n_2587),
.Y(n_2641)
);

INVx3_ASAP7_75t_L g2642 ( 
.A(n_2600),
.Y(n_2642)
);

NOR2xp33_ASAP7_75t_L g2643 ( 
.A(n_2573),
.B(n_2502),
.Y(n_2643)
);

INVxp67_ASAP7_75t_L g2644 ( 
.A(n_2561),
.Y(n_2644)
);

INVx1_ASAP7_75t_SL g2645 ( 
.A(n_2548),
.Y(n_2645)
);

HB1xp67_ASAP7_75t_L g2646 ( 
.A(n_2563),
.Y(n_2646)
);

CKINVDCx5p33_ASAP7_75t_R g2647 ( 
.A(n_2608),
.Y(n_2647)
);

AND2x4_ASAP7_75t_L g2648 ( 
.A(n_2605),
.B(n_2501),
.Y(n_2648)
);

CKINVDCx14_ASAP7_75t_R g2649 ( 
.A(n_2601),
.Y(n_2649)
);

INVx2_ASAP7_75t_SL g2650 ( 
.A(n_2565),
.Y(n_2650)
);

BUFx6f_ASAP7_75t_L g2651 ( 
.A(n_2581),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2556),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2555),
.Y(n_2653)
);

OAI21x1_ASAP7_75t_L g2654 ( 
.A1(n_2562),
.A2(n_2491),
.B(n_2482),
.Y(n_2654)
);

OAI21x1_ASAP7_75t_L g2655 ( 
.A1(n_2566),
.A2(n_2498),
.B(n_2506),
.Y(n_2655)
);

BUFx4f_ASAP7_75t_SL g2656 ( 
.A(n_2628),
.Y(n_2656)
);

AND2x2_ASAP7_75t_L g2657 ( 
.A(n_2617),
.B(n_2521),
.Y(n_2657)
);

NOR2xp33_ASAP7_75t_R g2658 ( 
.A(n_2647),
.B(n_2476),
.Y(n_2658)
);

INVxp67_ASAP7_75t_L g2659 ( 
.A(n_2627),
.Y(n_2659)
);

AND2x2_ASAP7_75t_L g2660 ( 
.A(n_2617),
.B(n_2516),
.Y(n_2660)
);

CKINVDCx16_ASAP7_75t_R g2661 ( 
.A(n_2639),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2610),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2613),
.Y(n_2663)
);

NOR2xp33_ASAP7_75t_R g2664 ( 
.A(n_2616),
.B(n_2507),
.Y(n_2664)
);

INVx2_ASAP7_75t_L g2665 ( 
.A(n_2629),
.Y(n_2665)
);

AO21x2_ASAP7_75t_L g2666 ( 
.A1(n_2631),
.A2(n_2568),
.B(n_2606),
.Y(n_2666)
);

INVx2_ASAP7_75t_L g2667 ( 
.A(n_2611),
.Y(n_2667)
);

CKINVDCx16_ASAP7_75t_R g2668 ( 
.A(n_2649),
.Y(n_2668)
);

BUFx6f_ASAP7_75t_L g2669 ( 
.A(n_2628),
.Y(n_2669)
);

INVx4_ASAP7_75t_SL g2670 ( 
.A(n_2651),
.Y(n_2670)
);

BUFx3_ASAP7_75t_L g2671 ( 
.A(n_2641),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2612),
.Y(n_2672)
);

INVx3_ASAP7_75t_L g2673 ( 
.A(n_2624),
.Y(n_2673)
);

NOR2xp33_ASAP7_75t_R g2674 ( 
.A(n_2642),
.B(n_2466),
.Y(n_2674)
);

NOR2xp33_ASAP7_75t_R g2675 ( 
.A(n_2650),
.B(n_2485),
.Y(n_2675)
);

CKINVDCx5p33_ASAP7_75t_R g2676 ( 
.A(n_2645),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2614),
.Y(n_2677)
);

AND2x4_ASAP7_75t_L g2678 ( 
.A(n_2624),
.B(n_2604),
.Y(n_2678)
);

OR2x2_ASAP7_75t_L g2679 ( 
.A(n_2618),
.B(n_2590),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_L g2680 ( 
.A(n_2633),
.B(n_2638),
.Y(n_2680)
);

NAND2xp33_ASAP7_75t_R g2681 ( 
.A(n_2635),
.B(n_2603),
.Y(n_2681)
);

BUFx6f_ASAP7_75t_L g2682 ( 
.A(n_2648),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_L g2683 ( 
.A(n_2636),
.B(n_2599),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2615),
.Y(n_2684)
);

AND2x2_ASAP7_75t_L g2685 ( 
.A(n_2619),
.B(n_2592),
.Y(n_2685)
);

OR2x6_ASAP7_75t_L g2686 ( 
.A(n_2626),
.B(n_2597),
.Y(n_2686)
);

INVx2_ASAP7_75t_L g2687 ( 
.A(n_2621),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2625),
.Y(n_2688)
);

NAND2xp33_ASAP7_75t_R g2689 ( 
.A(n_2643),
.B(n_4),
.Y(n_2689)
);

AND2x2_ASAP7_75t_L g2690 ( 
.A(n_2630),
.B(n_2602),
.Y(n_2690)
);

CKINVDCx5p33_ASAP7_75t_R g2691 ( 
.A(n_2644),
.Y(n_2691)
);

INVx2_ASAP7_75t_L g2692 ( 
.A(n_2622),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2646),
.Y(n_2693)
);

OAI22xp33_ASAP7_75t_SL g2694 ( 
.A1(n_2653),
.A2(n_2584),
.B1(n_932),
.B2(n_935),
.Y(n_2694)
);

OR2x2_ASAP7_75t_L g2695 ( 
.A(n_2632),
.B(n_2571),
.Y(n_2695)
);

AND2x2_ASAP7_75t_L g2696 ( 
.A(n_2634),
.B(n_2591),
.Y(n_2696)
);

AND2x2_ASAP7_75t_SL g2697 ( 
.A(n_2634),
.B(n_2473),
.Y(n_2697)
);

INVx4_ASAP7_75t_L g2698 ( 
.A(n_2623),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2652),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2637),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2654),
.Y(n_2701)
);

OR2x6_ASAP7_75t_L g2702 ( 
.A(n_2655),
.B(n_2595),
.Y(n_2702)
);

HB1xp67_ASAP7_75t_L g2703 ( 
.A(n_2620),
.Y(n_2703)
);

CKINVDCx5p33_ASAP7_75t_R g2704 ( 
.A(n_2640),
.Y(n_2704)
);

NAND2x1_ASAP7_75t_L g2705 ( 
.A(n_2609),
.B(n_2472),
.Y(n_2705)
);

AND2x2_ASAP7_75t_L g2706 ( 
.A(n_2673),
.B(n_2657),
.Y(n_2706)
);

AND2x2_ASAP7_75t_L g2707 ( 
.A(n_2660),
.B(n_2467),
.Y(n_2707)
);

INVx2_ASAP7_75t_L g2708 ( 
.A(n_2693),
.Y(n_2708)
);

OR2x2_ASAP7_75t_L g2709 ( 
.A(n_2659),
.B(n_2583),
.Y(n_2709)
);

AND2x2_ASAP7_75t_L g2710 ( 
.A(n_2692),
.B(n_2582),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2662),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2672),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2677),
.Y(n_2713)
);

INVx3_ASAP7_75t_L g2714 ( 
.A(n_2682),
.Y(n_2714)
);

OR2x2_ASAP7_75t_L g2715 ( 
.A(n_2699),
.B(n_2500),
.Y(n_2715)
);

AND2x2_ASAP7_75t_L g2716 ( 
.A(n_2661),
.B(n_2472),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_2665),
.Y(n_2717)
);

HB1xp67_ASAP7_75t_L g2718 ( 
.A(n_2679),
.Y(n_2718)
);

OA21x2_ASAP7_75t_L g2719 ( 
.A1(n_2701),
.A2(n_946),
.B(n_945),
.Y(n_2719)
);

BUFx2_ASAP7_75t_L g2720 ( 
.A(n_2678),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2667),
.Y(n_2721)
);

AOI22xp33_ASAP7_75t_SL g2722 ( 
.A1(n_2668),
.A2(n_2465),
.B1(n_949),
.B2(n_952),
.Y(n_2722)
);

INVxp67_ASAP7_75t_L g2723 ( 
.A(n_2683),
.Y(n_2723)
);

OAI22xp33_ASAP7_75t_L g2724 ( 
.A1(n_2689),
.A2(n_2479),
.B1(n_956),
.B2(n_959),
.Y(n_2724)
);

AND2x2_ASAP7_75t_L g2725 ( 
.A(n_2687),
.B(n_5),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2688),
.Y(n_2726)
);

AND2x4_ASAP7_75t_L g2727 ( 
.A(n_2690),
.B(n_6),
.Y(n_2727)
);

BUFx2_ASAP7_75t_L g2728 ( 
.A(n_2704),
.Y(n_2728)
);

AND2x2_ASAP7_75t_L g2729 ( 
.A(n_2663),
.B(n_6),
.Y(n_2729)
);

BUFx3_ASAP7_75t_L g2730 ( 
.A(n_2671),
.Y(n_2730)
);

OR2x2_ASAP7_75t_L g2731 ( 
.A(n_2684),
.B(n_9),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2680),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2700),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2703),
.Y(n_2734)
);

OR2x2_ASAP7_75t_L g2735 ( 
.A(n_2695),
.B(n_10),
.Y(n_2735)
);

INVxp67_ASAP7_75t_SL g2736 ( 
.A(n_2718),
.Y(n_2736)
);

OR2x2_ASAP7_75t_L g2737 ( 
.A(n_2723),
.B(n_2696),
.Y(n_2737)
);

BUFx6f_ASAP7_75t_L g2738 ( 
.A(n_2730),
.Y(n_2738)
);

INVx4_ASAP7_75t_L g2739 ( 
.A(n_2716),
.Y(n_2739)
);

OA21x2_ASAP7_75t_L g2740 ( 
.A1(n_2734),
.A2(n_2691),
.B(n_2676),
.Y(n_2740)
);

AO31x2_ASAP7_75t_L g2741 ( 
.A1(n_2726),
.A2(n_2698),
.A3(n_2681),
.B(n_2666),
.Y(n_2741)
);

AND2x2_ASAP7_75t_L g2742 ( 
.A(n_2720),
.B(n_2682),
.Y(n_2742)
);

AOI21x1_ASAP7_75t_L g2743 ( 
.A1(n_2728),
.A2(n_2705),
.B(n_2686),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2711),
.Y(n_2744)
);

AOI22xp33_ASAP7_75t_L g2745 ( 
.A1(n_2719),
.A2(n_2694),
.B1(n_2697),
.B2(n_2686),
.Y(n_2745)
);

AND2x2_ASAP7_75t_L g2746 ( 
.A(n_2706),
.B(n_2685),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2712),
.Y(n_2747)
);

AND2x2_ASAP7_75t_L g2748 ( 
.A(n_2728),
.B(n_2702),
.Y(n_2748)
);

A2O1A1Ixp33_ASAP7_75t_L g2749 ( 
.A1(n_2722),
.A2(n_964),
.B(n_993),
.C(n_977),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2713),
.Y(n_2750)
);

CKINVDCx20_ASAP7_75t_R g2751 ( 
.A(n_2707),
.Y(n_2751)
);

OAI221xp5_ASAP7_75t_L g2752 ( 
.A1(n_2735),
.A2(n_2702),
.B1(n_967),
.B2(n_968),
.C(n_965),
.Y(n_2752)
);

INVx2_ASAP7_75t_L g2753 ( 
.A(n_2715),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2733),
.Y(n_2754)
);

INVx2_ASAP7_75t_L g2755 ( 
.A(n_2717),
.Y(n_2755)
);

OAI211xp5_ASAP7_75t_L g2756 ( 
.A1(n_2731),
.A2(n_2675),
.B(n_969),
.C(n_970),
.Y(n_2756)
);

BUFx6f_ASAP7_75t_L g2757 ( 
.A(n_2725),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_2721),
.Y(n_2758)
);

INVx2_ASAP7_75t_L g2759 ( 
.A(n_2708),
.Y(n_2759)
);

OAI21xp33_ASAP7_75t_L g2760 ( 
.A1(n_2709),
.A2(n_976),
.B(n_947),
.Y(n_2760)
);

BUFx3_ASAP7_75t_L g2761 ( 
.A(n_2714),
.Y(n_2761)
);

INVx2_ASAP7_75t_L g2762 ( 
.A(n_2732),
.Y(n_2762)
);

AO21x1_ASAP7_75t_L g2763 ( 
.A1(n_2724),
.A2(n_2658),
.B(n_2670),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2729),
.Y(n_2764)
);

OAI21xp33_ASAP7_75t_L g2765 ( 
.A1(n_2710),
.A2(n_980),
.B(n_974),
.Y(n_2765)
);

INVx2_ASAP7_75t_L g2766 ( 
.A(n_2759),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_L g2767 ( 
.A(n_2753),
.B(n_2727),
.Y(n_2767)
);

INVx5_ASAP7_75t_SL g2768 ( 
.A(n_2738),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2754),
.Y(n_2769)
);

INVx2_ASAP7_75t_L g2770 ( 
.A(n_2755),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2744),
.Y(n_2771)
);

NAND2xp33_ASAP7_75t_R g2772 ( 
.A(n_2740),
.B(n_2664),
.Y(n_2772)
);

NOR2xp33_ASAP7_75t_L g2773 ( 
.A(n_2763),
.B(n_2656),
.Y(n_2773)
);

AND2x2_ASAP7_75t_L g2774 ( 
.A(n_2748),
.B(n_2669),
.Y(n_2774)
);

BUFx2_ASAP7_75t_L g2775 ( 
.A(n_2739),
.Y(n_2775)
);

HB1xp67_ASAP7_75t_L g2776 ( 
.A(n_2762),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_L g2777 ( 
.A(n_2764),
.B(n_2669),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2747),
.Y(n_2778)
);

NAND2xp5_ASAP7_75t_L g2779 ( 
.A(n_2750),
.B(n_2670),
.Y(n_2779)
);

OR2x2_ASAP7_75t_L g2780 ( 
.A(n_2737),
.B(n_11),
.Y(n_2780)
);

INVx2_ASAP7_75t_L g2781 ( 
.A(n_2758),
.Y(n_2781)
);

AND2x2_ASAP7_75t_L g2782 ( 
.A(n_2742),
.B(n_2674),
.Y(n_2782)
);

OR2x2_ASAP7_75t_L g2783 ( 
.A(n_2736),
.B(n_11),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2757),
.Y(n_2784)
);

AND2x4_ASAP7_75t_L g2785 ( 
.A(n_2761),
.B(n_13),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_L g2786 ( 
.A(n_2760),
.B(n_979),
.Y(n_2786)
);

OAI211xp5_ASAP7_75t_L g2787 ( 
.A1(n_2745),
.A2(n_2752),
.B(n_2756),
.C(n_2765),
.Y(n_2787)
);

INVx2_ASAP7_75t_L g2788 ( 
.A(n_2746),
.Y(n_2788)
);

AOI222xp33_ASAP7_75t_L g2789 ( 
.A1(n_2749),
.A2(n_984),
.B1(n_982),
.B2(n_987),
.C1(n_983),
.C2(n_981),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2757),
.Y(n_2790)
);

HB1xp67_ASAP7_75t_L g2791 ( 
.A(n_2741),
.Y(n_2791)
);

AND2x2_ASAP7_75t_L g2792 ( 
.A(n_2743),
.B(n_2741),
.Y(n_2792)
);

AOI22xp5_ASAP7_75t_L g2793 ( 
.A1(n_2751),
.A2(n_1011),
.B1(n_1017),
.B2(n_1009),
.Y(n_2793)
);

BUFx2_ASAP7_75t_SL g2794 ( 
.A(n_2763),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2754),
.Y(n_2795)
);

AND2x4_ASAP7_75t_SL g2796 ( 
.A(n_2782),
.B(n_2504),
.Y(n_2796)
);

INVx2_ASAP7_75t_L g2797 ( 
.A(n_2775),
.Y(n_2797)
);

AOI22xp33_ASAP7_75t_L g2798 ( 
.A1(n_2794),
.A2(n_1025),
.B1(n_1026),
.B2(n_1023),
.Y(n_2798)
);

OR2x2_ASAP7_75t_L g2799 ( 
.A(n_2780),
.B(n_12),
.Y(n_2799)
);

OR2x2_ASAP7_75t_L g2800 ( 
.A(n_2766),
.B(n_12),
.Y(n_2800)
);

INVx2_ASAP7_75t_SL g2801 ( 
.A(n_2785),
.Y(n_2801)
);

OR2x2_ASAP7_75t_L g2802 ( 
.A(n_2770),
.B(n_13),
.Y(n_2802)
);

AND2x2_ASAP7_75t_L g2803 ( 
.A(n_2788),
.B(n_14),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2769),
.Y(n_2804)
);

AND2x4_ASAP7_75t_L g2805 ( 
.A(n_2784),
.B(n_14),
.Y(n_2805)
);

INVx2_ASAP7_75t_L g2806 ( 
.A(n_2774),
.Y(n_2806)
);

INVx6_ASAP7_75t_L g2807 ( 
.A(n_2783),
.Y(n_2807)
);

AND2x2_ASAP7_75t_L g2808 ( 
.A(n_2790),
.B(n_15),
.Y(n_2808)
);

AND2x2_ASAP7_75t_L g2809 ( 
.A(n_2773),
.B(n_2776),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2771),
.Y(n_2810)
);

AND2x2_ASAP7_75t_L g2811 ( 
.A(n_2767),
.B(n_15),
.Y(n_2811)
);

AND2x2_ASAP7_75t_L g2812 ( 
.A(n_2768),
.B(n_16),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2778),
.Y(n_2813)
);

AND2x4_ASAP7_75t_L g2814 ( 
.A(n_2779),
.B(n_16),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2795),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2781),
.Y(n_2816)
);

INVx2_ASAP7_75t_L g2817 ( 
.A(n_2768),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2777),
.Y(n_2818)
);

AND2x2_ASAP7_75t_L g2819 ( 
.A(n_2792),
.B(n_17),
.Y(n_2819)
);

OR2x6_ASAP7_75t_L g2820 ( 
.A(n_2787),
.B(n_17),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2791),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_2793),
.B(n_1030),
.Y(n_2822)
);

OR2x2_ASAP7_75t_L g2823 ( 
.A(n_2786),
.B(n_19),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_2789),
.B(n_2772),
.Y(n_2824)
);

INVxp67_ASAP7_75t_L g2825 ( 
.A(n_2801),
.Y(n_2825)
);

INVx2_ASAP7_75t_L g2826 ( 
.A(n_2817),
.Y(n_2826)
);

HB1xp67_ASAP7_75t_L g2827 ( 
.A(n_2807),
.Y(n_2827)
);

AOI21xp5_ASAP7_75t_L g2828 ( 
.A1(n_2824),
.A2(n_1036),
.B(n_1033),
.Y(n_2828)
);

AND2x4_ASAP7_75t_SL g2829 ( 
.A(n_2812),
.B(n_20),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2804),
.Y(n_2830)
);

AND2x2_ASAP7_75t_L g2831 ( 
.A(n_2809),
.B(n_20),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_L g2832 ( 
.A(n_2819),
.B(n_1037),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_L g2833 ( 
.A(n_2797),
.B(n_1038),
.Y(n_2833)
);

INVx2_ASAP7_75t_L g2834 ( 
.A(n_2806),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2810),
.Y(n_2835)
);

INVxp67_ASAP7_75t_L g2836 ( 
.A(n_2820),
.Y(n_2836)
);

INVxp67_ASAP7_75t_SL g2837 ( 
.A(n_2800),
.Y(n_2837)
);

NOR2x1_ASAP7_75t_L g2838 ( 
.A(n_2820),
.B(n_22),
.Y(n_2838)
);

AND2x2_ASAP7_75t_L g2839 ( 
.A(n_2818),
.B(n_22),
.Y(n_2839)
);

OR2x2_ASAP7_75t_L g2840 ( 
.A(n_2816),
.B(n_23),
.Y(n_2840)
);

OAI21xp33_ASAP7_75t_L g2841 ( 
.A1(n_2798),
.A2(n_2815),
.B(n_2813),
.Y(n_2841)
);

INVx2_ASAP7_75t_L g2842 ( 
.A(n_2802),
.Y(n_2842)
);

INVx2_ASAP7_75t_L g2843 ( 
.A(n_2807),
.Y(n_2843)
);

AND2x2_ASAP7_75t_L g2844 ( 
.A(n_2796),
.B(n_23),
.Y(n_2844)
);

INVx2_ASAP7_75t_SL g2845 ( 
.A(n_2805),
.Y(n_2845)
);

OR2x2_ASAP7_75t_L g2846 ( 
.A(n_2799),
.B(n_24),
.Y(n_2846)
);

OR2x2_ASAP7_75t_L g2847 ( 
.A(n_2823),
.B(n_24),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2821),
.Y(n_2848)
);

AND2x2_ASAP7_75t_L g2849 ( 
.A(n_2814),
.B(n_2811),
.Y(n_2849)
);

INVx2_ASAP7_75t_L g2850 ( 
.A(n_2803),
.Y(n_2850)
);

AND2x4_ASAP7_75t_L g2851 ( 
.A(n_2808),
.B(n_2822),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2804),
.Y(n_2852)
);

INVx2_ASAP7_75t_L g2853 ( 
.A(n_2817),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2804),
.Y(n_2854)
);

NAND2xp5_ASAP7_75t_L g2855 ( 
.A(n_2819),
.B(n_1044),
.Y(n_2855)
);

INVx2_ASAP7_75t_L g2856 ( 
.A(n_2817),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2804),
.Y(n_2857)
);

INVx1_ASAP7_75t_SL g2858 ( 
.A(n_2812),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2804),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2817),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2804),
.Y(n_2861)
);

INVxp67_ASAP7_75t_L g2862 ( 
.A(n_2801),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_L g2863 ( 
.A(n_2819),
.B(n_1047),
.Y(n_2863)
);

INVx2_ASAP7_75t_SL g2864 ( 
.A(n_2817),
.Y(n_2864)
);

INVx1_ASAP7_75t_SL g2865 ( 
.A(n_2829),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_L g2866 ( 
.A(n_2858),
.B(n_1049),
.Y(n_2866)
);

INVx1_ASAP7_75t_SL g2867 ( 
.A(n_2827),
.Y(n_2867)
);

INVx3_ASAP7_75t_L g2868 ( 
.A(n_2843),
.Y(n_2868)
);

AND2x2_ASAP7_75t_L g2869 ( 
.A(n_2849),
.B(n_26),
.Y(n_2869)
);

AND2x4_ASAP7_75t_L g2870 ( 
.A(n_2826),
.B(n_27),
.Y(n_2870)
);

AND2x2_ASAP7_75t_L g2871 ( 
.A(n_2845),
.B(n_30),
.Y(n_2871)
);

OR2x2_ASAP7_75t_L g2872 ( 
.A(n_2836),
.B(n_30),
.Y(n_2872)
);

INVx2_ASAP7_75t_L g2873 ( 
.A(n_2853),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_L g2874 ( 
.A(n_2838),
.B(n_1056),
.Y(n_2874)
);

AND2x2_ASAP7_75t_L g2875 ( 
.A(n_2856),
.B(n_31),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_L g2876 ( 
.A(n_2860),
.B(n_2825),
.Y(n_2876)
);

INVxp67_ASAP7_75t_SL g2877 ( 
.A(n_2862),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_SL g2878 ( 
.A(n_2851),
.B(n_1060),
.Y(n_2878)
);

NAND2x1p5_ASAP7_75t_L g2879 ( 
.A(n_2844),
.B(n_32),
.Y(n_2879)
);

AND2x2_ASAP7_75t_L g2880 ( 
.A(n_2851),
.B(n_31),
.Y(n_2880)
);

OR2x2_ASAP7_75t_L g2881 ( 
.A(n_2850),
.B(n_34),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_2837),
.B(n_1064),
.Y(n_2882)
);

INVx2_ASAP7_75t_L g2883 ( 
.A(n_2842),
.Y(n_2883)
);

INVx2_ASAP7_75t_L g2884 ( 
.A(n_2840),
.Y(n_2884)
);

INVx1_ASAP7_75t_SL g2885 ( 
.A(n_2831),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2830),
.Y(n_2886)
);

OR2x2_ASAP7_75t_L g2887 ( 
.A(n_2834),
.B(n_35),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2830),
.Y(n_2888)
);

AND2x2_ASAP7_75t_L g2889 ( 
.A(n_2839),
.B(n_36),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2848),
.Y(n_2890)
);

INVx2_ASAP7_75t_L g2891 ( 
.A(n_2846),
.Y(n_2891)
);

OR2x2_ASAP7_75t_L g2892 ( 
.A(n_2847),
.B(n_36),
.Y(n_2892)
);

NOR2xp33_ASAP7_75t_L g2893 ( 
.A(n_2832),
.B(n_1065),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2835),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2852),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2854),
.Y(n_2896)
);

NAND2xp5_ASAP7_75t_L g2897 ( 
.A(n_2841),
.B(n_1067),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_L g2898 ( 
.A(n_2833),
.B(n_1068),
.Y(n_2898)
);

AOI22xp5_ASAP7_75t_SL g2899 ( 
.A1(n_2828),
.A2(n_1070),
.B1(n_1071),
.B2(n_1069),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2857),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2859),
.Y(n_2901)
);

AND2x2_ASAP7_75t_L g2902 ( 
.A(n_2861),
.B(n_37),
.Y(n_2902)
);

HB1xp67_ASAP7_75t_L g2903 ( 
.A(n_2855),
.Y(n_2903)
);

BUFx2_ASAP7_75t_L g2904 ( 
.A(n_2863),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2827),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_L g2906 ( 
.A(n_2858),
.B(n_1074),
.Y(n_2906)
);

INVx1_ASAP7_75t_SL g2907 ( 
.A(n_2829),
.Y(n_2907)
);

OR2x2_ASAP7_75t_L g2908 ( 
.A(n_2858),
.B(n_37),
.Y(n_2908)
);

NAND4xp75_ASAP7_75t_L g2909 ( 
.A(n_2838),
.B(n_40),
.C(n_38),
.D(n_39),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2827),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_L g2911 ( 
.A(n_2858),
.B(n_1075),
.Y(n_2911)
);

INVx2_ASAP7_75t_L g2912 ( 
.A(n_2864),
.Y(n_2912)
);

INVx2_ASAP7_75t_L g2913 ( 
.A(n_2864),
.Y(n_2913)
);

BUFx2_ASAP7_75t_L g2914 ( 
.A(n_2827),
.Y(n_2914)
);

INVx1_ASAP7_75t_SL g2915 ( 
.A(n_2829),
.Y(n_2915)
);

NAND2xp5_ASAP7_75t_L g2916 ( 
.A(n_2858),
.B(n_1078),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2827),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2827),
.Y(n_2918)
);

OR2x2_ASAP7_75t_L g2919 ( 
.A(n_2858),
.B(n_39),
.Y(n_2919)
);

AND2x2_ASAP7_75t_L g2920 ( 
.A(n_2864),
.B(n_44),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_L g2921 ( 
.A(n_2914),
.B(n_1079),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2872),
.Y(n_2922)
);

INVx2_ASAP7_75t_L g2923 ( 
.A(n_2879),
.Y(n_2923)
);

OR2x2_ASAP7_75t_L g2924 ( 
.A(n_2905),
.B(n_45),
.Y(n_2924)
);

NAND2x1p5_ASAP7_75t_L g2925 ( 
.A(n_2865),
.B(n_46),
.Y(n_2925)
);

AND2x2_ASAP7_75t_L g2926 ( 
.A(n_2907),
.B(n_1083),
.Y(n_2926)
);

HB1xp67_ASAP7_75t_L g2927 ( 
.A(n_2915),
.Y(n_2927)
);

INVx2_ASAP7_75t_L g2928 ( 
.A(n_2868),
.Y(n_2928)
);

AND2x2_ASAP7_75t_L g2929 ( 
.A(n_2877),
.B(n_1095),
.Y(n_2929)
);

NOR2xp33_ASAP7_75t_SL g2930 ( 
.A(n_2909),
.B(n_1100),
.Y(n_2930)
);

AND2x2_ASAP7_75t_L g2931 ( 
.A(n_2912),
.B(n_1099),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2881),
.Y(n_2932)
);

AND2x2_ASAP7_75t_L g2933 ( 
.A(n_2913),
.B(n_1102),
.Y(n_2933)
);

OR2x6_ASAP7_75t_L g2934 ( 
.A(n_2910),
.B(n_46),
.Y(n_2934)
);

INVx2_ASAP7_75t_L g2935 ( 
.A(n_2920),
.Y(n_2935)
);

INVx2_ASAP7_75t_L g2936 ( 
.A(n_2917),
.Y(n_2936)
);

AND2x2_ASAP7_75t_L g2937 ( 
.A(n_2918),
.B(n_1103),
.Y(n_2937)
);

INVx2_ASAP7_75t_L g2938 ( 
.A(n_2871),
.Y(n_2938)
);

HB1xp67_ASAP7_75t_L g2939 ( 
.A(n_2885),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2880),
.Y(n_2940)
);

AOI22xp33_ASAP7_75t_L g2941 ( 
.A1(n_2904),
.A2(n_2903),
.B1(n_2891),
.B2(n_2884),
.Y(n_2941)
);

AND2x4_ASAP7_75t_L g2942 ( 
.A(n_2873),
.B(n_48),
.Y(n_2942)
);

INVx2_ASAP7_75t_SL g2943 ( 
.A(n_2870),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2887),
.Y(n_2944)
);

INVx2_ASAP7_75t_L g2945 ( 
.A(n_2870),
.Y(n_2945)
);

OR2x2_ASAP7_75t_L g2946 ( 
.A(n_2876),
.B(n_47),
.Y(n_2946)
);

AOI22xp33_ASAP7_75t_L g2947 ( 
.A1(n_2883),
.A2(n_1107),
.B1(n_1109),
.B2(n_1106),
.Y(n_2947)
);

AND2x4_ASAP7_75t_L g2948 ( 
.A(n_2875),
.B(n_47),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2892),
.Y(n_2949)
);

AND2x2_ASAP7_75t_L g2950 ( 
.A(n_2869),
.B(n_1112),
.Y(n_2950)
);

AND2x2_ASAP7_75t_L g2951 ( 
.A(n_2889),
.B(n_1118),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2902),
.Y(n_2952)
);

INVx1_ASAP7_75t_SL g2953 ( 
.A(n_2908),
.Y(n_2953)
);

INVx2_ASAP7_75t_L g2954 ( 
.A(n_2919),
.Y(n_2954)
);

HB1xp67_ASAP7_75t_L g2955 ( 
.A(n_2909),
.Y(n_2955)
);

OR2x2_ASAP7_75t_L g2956 ( 
.A(n_2882),
.B(n_50),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_L g2957 ( 
.A(n_2899),
.B(n_1119),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2886),
.Y(n_2958)
);

NAND2xp5_ASAP7_75t_L g2959 ( 
.A(n_2893),
.B(n_1123),
.Y(n_2959)
);

AND2x2_ASAP7_75t_L g2960 ( 
.A(n_2878),
.B(n_1124),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2888),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_L g2962 ( 
.A(n_2866),
.B(n_1125),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2890),
.Y(n_2963)
);

INVx4_ASAP7_75t_L g2964 ( 
.A(n_2901),
.Y(n_2964)
);

AND2x2_ASAP7_75t_L g2965 ( 
.A(n_2894),
.B(n_2895),
.Y(n_2965)
);

INVx2_ASAP7_75t_SL g2966 ( 
.A(n_2896),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2900),
.Y(n_2967)
);

AOI22xp5_ASAP7_75t_L g2968 ( 
.A1(n_2897),
.A2(n_1131),
.B1(n_1132),
.B2(n_1128),
.Y(n_2968)
);

INVx1_ASAP7_75t_SL g2969 ( 
.A(n_2874),
.Y(n_2969)
);

INVx2_ASAP7_75t_SL g2970 ( 
.A(n_2906),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2916),
.Y(n_2971)
);

OR2x2_ASAP7_75t_L g2972 ( 
.A(n_2911),
.B(n_51),
.Y(n_2972)
);

NAND2x1_ASAP7_75t_L g2973 ( 
.A(n_2898),
.B(n_52),
.Y(n_2973)
);

BUFx2_ASAP7_75t_L g2974 ( 
.A(n_2914),
.Y(n_2974)
);

NOR2xp33_ASAP7_75t_L g2975 ( 
.A(n_2865),
.B(n_1134),
.Y(n_2975)
);

NAND2xp5_ASAP7_75t_L g2976 ( 
.A(n_2914),
.B(n_1136),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2914),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2914),
.Y(n_2978)
);

NAND2xp5_ASAP7_75t_L g2979 ( 
.A(n_2914),
.B(n_1137),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_L g2980 ( 
.A(n_2914),
.B(n_1139),
.Y(n_2980)
);

INVx2_ASAP7_75t_L g2981 ( 
.A(n_2914),
.Y(n_2981)
);

AND2x2_ASAP7_75t_L g2982 ( 
.A(n_2914),
.B(n_1140),
.Y(n_2982)
);

NAND3xp33_ASAP7_75t_L g2983 ( 
.A(n_2914),
.B(n_1142),
.C(n_1141),
.Y(n_2983)
);

NOR2xp33_ASAP7_75t_L g2984 ( 
.A(n_2865),
.B(n_1144),
.Y(n_2984)
);

AND2x2_ASAP7_75t_L g2985 ( 
.A(n_2914),
.B(n_1147),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_L g2986 ( 
.A(n_2914),
.B(n_1148),
.Y(n_2986)
);

AOI22xp33_ASAP7_75t_L g2987 ( 
.A1(n_2867),
.A2(n_1150),
.B1(n_1153),
.B2(n_1149),
.Y(n_2987)
);

INVx1_ASAP7_75t_SL g2988 ( 
.A(n_2914),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2914),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_L g2990 ( 
.A(n_2914),
.B(n_1154),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2914),
.Y(n_2991)
);

OAI21xp33_ASAP7_75t_L g2992 ( 
.A1(n_2867),
.A2(n_1158),
.B(n_1155),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_L g2993 ( 
.A(n_2914),
.B(n_1161),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_2914),
.B(n_1165),
.Y(n_2994)
);

INVx2_ASAP7_75t_L g2995 ( 
.A(n_2914),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2914),
.Y(n_2996)
);

OAI21xp33_ASAP7_75t_L g2997 ( 
.A1(n_2927),
.A2(n_1172),
.B(n_1169),
.Y(n_2997)
);

NAND2x1_ASAP7_75t_SL g2998 ( 
.A(n_2955),
.B(n_52),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2974),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2939),
.Y(n_3000)
);

OAI21xp5_ASAP7_75t_L g3001 ( 
.A1(n_2988),
.A2(n_1175),
.B(n_1173),
.Y(n_3001)
);

NAND2x1_ASAP7_75t_L g3002 ( 
.A(n_2943),
.B(n_2981),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2995),
.B(n_1182),
.Y(n_3003)
);

OAI22xp5_ASAP7_75t_L g3004 ( 
.A1(n_2925),
.A2(n_2978),
.B1(n_2989),
.B2(n_2977),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_L g3005 ( 
.A(n_2991),
.B(n_1183),
.Y(n_3005)
);

AOI22xp33_ASAP7_75t_L g3006 ( 
.A1(n_2996),
.A2(n_1186),
.B1(n_1190),
.B2(n_1185),
.Y(n_3006)
);

INVxp67_ASAP7_75t_L g3007 ( 
.A(n_2930),
.Y(n_3007)
);

AOI221xp5_ASAP7_75t_L g3008 ( 
.A1(n_2936),
.A2(n_1195),
.B1(n_1200),
.B2(n_1194),
.C(n_1192),
.Y(n_3008)
);

INVx2_ASAP7_75t_L g3009 ( 
.A(n_2923),
.Y(n_3009)
);

OR2x2_ASAP7_75t_L g3010 ( 
.A(n_2945),
.B(n_2953),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2924),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2934),
.Y(n_3012)
);

NAND2xp5_ASAP7_75t_R g3013 ( 
.A(n_2970),
.B(n_53),
.Y(n_3013)
);

INVx2_ASAP7_75t_L g3014 ( 
.A(n_2928),
.Y(n_3014)
);

AND2x4_ASAP7_75t_L g3015 ( 
.A(n_2938),
.B(n_53),
.Y(n_3015)
);

A2O1A1O1Ixp25_ASAP7_75t_L g3016 ( 
.A1(n_2952),
.A2(n_56),
.B(n_54),
.C(n_55),
.D(n_58),
.Y(n_3016)
);

INVx2_ASAP7_75t_L g3017 ( 
.A(n_2948),
.Y(n_3017)
);

AOI22xp5_ASAP7_75t_L g3018 ( 
.A1(n_2940),
.A2(n_1205),
.B1(n_1206),
.B2(n_1204),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2942),
.Y(n_3019)
);

OAI22xp5_ASAP7_75t_L g3020 ( 
.A1(n_2935),
.A2(n_2954),
.B1(n_2987),
.B2(n_2969),
.Y(n_3020)
);

OAI22xp33_ASAP7_75t_L g3021 ( 
.A1(n_2964),
.A2(n_1208),
.B1(n_1209),
.B2(n_1207),
.Y(n_3021)
);

INVxp67_ASAP7_75t_L g3022 ( 
.A(n_2975),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2942),
.Y(n_3023)
);

OAI21xp33_ASAP7_75t_L g3024 ( 
.A1(n_2922),
.A2(n_1212),
.B(n_1211),
.Y(n_3024)
);

AND2x2_ASAP7_75t_L g3025 ( 
.A(n_2926),
.B(n_1213),
.Y(n_3025)
);

AOI221xp5_ASAP7_75t_L g3026 ( 
.A1(n_2966),
.A2(n_1218),
.B1(n_1221),
.B2(n_1216),
.C(n_1215),
.Y(n_3026)
);

AOI322xp5_ASAP7_75t_L g3027 ( 
.A1(n_2963),
.A2(n_1231),
.A3(n_1229),
.B1(n_1232),
.B2(n_1233),
.C1(n_1230),
.C2(n_1227),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2949),
.Y(n_3028)
);

AND2x2_ASAP7_75t_L g3029 ( 
.A(n_2932),
.B(n_1234),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2946),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_SL g3031 ( 
.A(n_2982),
.B(n_1235),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_2950),
.B(n_1236),
.Y(n_3032)
);

AOI221xp5_ASAP7_75t_L g3033 ( 
.A1(n_2967),
.A2(n_1244),
.B1(n_1247),
.B2(n_1242),
.C(n_1241),
.Y(n_3033)
);

NAND2xp5_ASAP7_75t_L g3034 ( 
.A(n_2951),
.B(n_1248),
.Y(n_3034)
);

AND2x2_ASAP7_75t_L g3035 ( 
.A(n_2944),
.B(n_1251),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2965),
.Y(n_3036)
);

OAI21xp5_ASAP7_75t_L g3037 ( 
.A1(n_2983),
.A2(n_1253),
.B(n_1252),
.Y(n_3037)
);

AOI21xp5_ASAP7_75t_L g3038 ( 
.A1(n_2973),
.A2(n_1259),
.B(n_1254),
.Y(n_3038)
);

OR2x2_ASAP7_75t_L g3039 ( 
.A(n_2971),
.B(n_2994),
.Y(n_3039)
);

INVx2_ASAP7_75t_L g3040 ( 
.A(n_2972),
.Y(n_3040)
);

NAND3xp33_ASAP7_75t_L g3041 ( 
.A(n_2958),
.B(n_1261),
.C(n_1260),
.Y(n_3041)
);

AOI22xp5_ASAP7_75t_L g3042 ( 
.A1(n_2984),
.A2(n_1264),
.B1(n_1268),
.B2(n_1263),
.Y(n_3042)
);

AOI21xp33_ASAP7_75t_L g3043 ( 
.A1(n_2921),
.A2(n_1271),
.B(n_1269),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_2956),
.Y(n_3044)
);

NOR2x1_ASAP7_75t_L g3045 ( 
.A(n_2985),
.B(n_54),
.Y(n_3045)
);

INVx1_ASAP7_75t_SL g3046 ( 
.A(n_2929),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_L g3047 ( 
.A(n_2931),
.B(n_1274),
.Y(n_3047)
);

NOR2xp67_ASAP7_75t_L g3048 ( 
.A(n_2961),
.B(n_56),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2933),
.B(n_1275),
.Y(n_3049)
);

NOR2xp33_ASAP7_75t_L g3050 ( 
.A(n_2992),
.B(n_1276),
.Y(n_3050)
);

INVx1_ASAP7_75t_SL g3051 ( 
.A(n_2960),
.Y(n_3051)
);

AOI21xp5_ASAP7_75t_L g3052 ( 
.A1(n_2957),
.A2(n_1278),
.B(n_1277),
.Y(n_3052)
);

AOI22xp5_ASAP7_75t_L g3053 ( 
.A1(n_2937),
.A2(n_1282),
.B1(n_1283),
.B2(n_1280),
.Y(n_3053)
);

NAND2xp5_ASAP7_75t_L g3054 ( 
.A(n_2968),
.B(n_2947),
.Y(n_3054)
);

AOI222xp33_ASAP7_75t_L g3055 ( 
.A1(n_2976),
.A2(n_1291),
.B1(n_1288),
.B2(n_1292),
.C1(n_1289),
.C2(n_1287),
.Y(n_3055)
);

NOR2xp33_ASAP7_75t_L g3056 ( 
.A(n_2962),
.B(n_1299),
.Y(n_3056)
);

OAI322xp33_ASAP7_75t_L g3057 ( 
.A1(n_2979),
.A2(n_1308),
.A3(n_1309),
.B1(n_1307),
.B2(n_59),
.C1(n_63),
.C2(n_62),
.Y(n_3057)
);

AND2x4_ASAP7_75t_L g3058 ( 
.A(n_2980),
.B(n_55),
.Y(n_3058)
);

OR2x2_ASAP7_75t_L g3059 ( 
.A(n_2986),
.B(n_58),
.Y(n_3059)
);

OAI22xp33_ASAP7_75t_L g3060 ( 
.A1(n_2990),
.A2(n_62),
.B1(n_59),
.B2(n_60),
.Y(n_3060)
);

AOI22xp5_ASAP7_75t_L g3061 ( 
.A1(n_2993),
.A2(n_64),
.B1(n_60),
.B2(n_63),
.Y(n_3061)
);

AOI211xp5_ASAP7_75t_L g3062 ( 
.A1(n_2959),
.A2(n_69),
.B(n_65),
.C(n_67),
.Y(n_3062)
);

AOI22xp5_ASAP7_75t_L g3063 ( 
.A1(n_2988),
.A2(n_70),
.B1(n_65),
.B2(n_67),
.Y(n_3063)
);

AOI22xp5_ASAP7_75t_L g3064 ( 
.A1(n_2988),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_3064)
);

AOI21xp5_ASAP7_75t_L g3065 ( 
.A1(n_2955),
.A2(n_73),
.B(n_75),
.Y(n_3065)
);

AND2x2_ASAP7_75t_L g3066 ( 
.A(n_2927),
.B(n_76),
.Y(n_3066)
);

NAND3xp33_ASAP7_75t_L g3067 ( 
.A(n_2955),
.B(n_76),
.C(n_77),
.Y(n_3067)
);

O2A1O1Ixp33_ASAP7_75t_L g3068 ( 
.A1(n_2955),
.A2(n_80),
.B(n_78),
.C(n_79),
.Y(n_3068)
);

NAND2x1_ASAP7_75t_L g3069 ( 
.A(n_2974),
.B(n_78),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_L g3070 ( 
.A(n_2927),
.B(n_79),
.Y(n_3070)
);

HB1xp67_ASAP7_75t_L g3071 ( 
.A(n_2974),
.Y(n_3071)
);

INVx2_ASAP7_75t_L g3072 ( 
.A(n_2974),
.Y(n_3072)
);

OAI32xp33_ASAP7_75t_L g3073 ( 
.A1(n_2955),
.A2(n_83),
.A3(n_86),
.B1(n_82),
.B2(n_85),
.Y(n_3073)
);

OAI22xp33_ASAP7_75t_L g3074 ( 
.A1(n_2988),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_3074)
);

HB1xp67_ASAP7_75t_L g3075 ( 
.A(n_2974),
.Y(n_3075)
);

OAI211xp5_ASAP7_75t_L g3076 ( 
.A1(n_2955),
.A2(n_89),
.B(n_86),
.C(n_87),
.Y(n_3076)
);

OAI31xp33_ASAP7_75t_L g3077 ( 
.A1(n_2955),
.A2(n_93),
.A3(n_89),
.B(n_91),
.Y(n_3077)
);

O2A1O1Ixp33_ASAP7_75t_L g3078 ( 
.A1(n_2955),
.A2(n_95),
.B(n_93),
.C(n_94),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2974),
.Y(n_3079)
);

AOI221xp5_ASAP7_75t_L g3080 ( 
.A1(n_2955),
.A2(n_116),
.B1(n_126),
.B2(n_105),
.C(n_94),
.Y(n_3080)
);

OAI22xp5_ASAP7_75t_L g3081 ( 
.A1(n_2988),
.A2(n_99),
.B1(n_95),
.B2(n_96),
.Y(n_3081)
);

OAI21xp5_ASAP7_75t_SL g3082 ( 
.A1(n_2955),
.A2(n_102),
.B(n_103),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_2927),
.B(n_104),
.Y(n_3083)
);

INVx1_ASAP7_75t_SL g3084 ( 
.A(n_2974),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_2974),
.Y(n_3085)
);

AOI21xp33_ASAP7_75t_SL g3086 ( 
.A1(n_2925),
.A2(n_104),
.B(n_106),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2974),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2974),
.Y(n_3088)
);

OAI33xp33_ASAP7_75t_L g3089 ( 
.A1(n_2977),
.A2(n_109),
.A3(n_113),
.B1(n_106),
.B2(n_107),
.B3(n_112),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_2927),
.B(n_114),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_2974),
.Y(n_3091)
);

INVx2_ASAP7_75t_L g3092 ( 
.A(n_2974),
.Y(n_3092)
);

INVxp67_ASAP7_75t_SL g3093 ( 
.A(n_2925),
.Y(n_3093)
);

NAND2xp33_ASAP7_75t_L g3094 ( 
.A(n_2925),
.B(n_115),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2974),
.Y(n_3095)
);

OAI211xp5_ASAP7_75t_SL g3096 ( 
.A1(n_2941),
.A2(n_124),
.B(n_120),
.C(n_122),
.Y(n_3096)
);

NAND2xp5_ASAP7_75t_L g3097 ( 
.A(n_2927),
.B(n_126),
.Y(n_3097)
);

AOI221xp5_ASAP7_75t_L g3098 ( 
.A1(n_2955),
.A2(n_148),
.B1(n_156),
.B2(n_138),
.C(n_127),
.Y(n_3098)
);

INVxp67_ASAP7_75t_L g3099 ( 
.A(n_2974),
.Y(n_3099)
);

OAI21xp5_ASAP7_75t_L g3100 ( 
.A1(n_2955),
.A2(n_127),
.B(n_128),
.Y(n_3100)
);

AOI22xp5_ASAP7_75t_L g3101 ( 
.A1(n_2988),
.A2(n_132),
.B1(n_128),
.B2(n_131),
.Y(n_3101)
);

OAI322xp33_ASAP7_75t_L g3102 ( 
.A1(n_2988),
.A2(n_139),
.A3(n_137),
.B1(n_135),
.B2(n_132),
.C1(n_134),
.C2(n_136),
.Y(n_3102)
);

AND2x2_ASAP7_75t_L g3103 ( 
.A(n_2927),
.B(n_134),
.Y(n_3103)
);

OAI22xp5_ASAP7_75t_L g3104 ( 
.A1(n_2988),
.A2(n_139),
.B1(n_136),
.B2(n_137),
.Y(n_3104)
);

OAI211xp5_ASAP7_75t_SL g3105 ( 
.A1(n_2941),
.A2(n_143),
.B(n_141),
.C(n_142),
.Y(n_3105)
);

OAI21xp33_ASAP7_75t_SL g3106 ( 
.A1(n_2988),
.A2(n_141),
.B(n_144),
.Y(n_3106)
);

OAI322xp33_ASAP7_75t_L g3107 ( 
.A1(n_2988),
.A2(n_150),
.A3(n_149),
.B1(n_146),
.B2(n_144),
.C1(n_145),
.C2(n_148),
.Y(n_3107)
);

OAI21xp33_ASAP7_75t_L g3108 ( 
.A1(n_2927),
.A2(n_149),
.B(n_151),
.Y(n_3108)
);

OR2x6_ASAP7_75t_L g3109 ( 
.A(n_2925),
.B(n_152),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_L g3110 ( 
.A(n_2927),
.B(n_153),
.Y(n_3110)
);

OR2x2_ASAP7_75t_L g3111 ( 
.A(n_2974),
.B(n_153),
.Y(n_3111)
);

AOI221xp5_ASAP7_75t_L g3112 ( 
.A1(n_2955),
.A2(n_168),
.B1(n_183),
.B2(n_161),
.C(n_154),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_2974),
.Y(n_3113)
);

AND2x2_ASAP7_75t_L g3114 ( 
.A(n_2927),
.B(n_155),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_3071),
.Y(n_3115)
);

NOR2xp33_ASAP7_75t_L g3116 ( 
.A(n_3109),
.B(n_157),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_3075),
.Y(n_3117)
);

OR2x2_ASAP7_75t_L g3118 ( 
.A(n_3084),
.B(n_158),
.Y(n_3118)
);

INVxp67_ASAP7_75t_L g3119 ( 
.A(n_3109),
.Y(n_3119)
);

HB1xp67_ASAP7_75t_L g3120 ( 
.A(n_3069),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_3066),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_L g3122 ( 
.A(n_3093),
.B(n_160),
.Y(n_3122)
);

AND2x2_ASAP7_75t_L g3123 ( 
.A(n_3072),
.B(n_161),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_3103),
.B(n_162),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_3114),
.Y(n_3125)
);

AOI21xp33_ASAP7_75t_L g3126 ( 
.A1(n_3002),
.A2(n_162),
.B(n_163),
.Y(n_3126)
);

NOR2xp33_ASAP7_75t_L g3127 ( 
.A(n_3106),
.B(n_164),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_3010),
.Y(n_3128)
);

INVx1_ASAP7_75t_L g3129 ( 
.A(n_3111),
.Y(n_3129)
);

INVxp67_ASAP7_75t_L g3130 ( 
.A(n_3094),
.Y(n_3130)
);

INVx1_ASAP7_75t_L g3131 ( 
.A(n_3048),
.Y(n_3131)
);

NAND2xp5_ASAP7_75t_L g3132 ( 
.A(n_2998),
.B(n_164),
.Y(n_3132)
);

INVx1_ASAP7_75t_SL g3133 ( 
.A(n_3045),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_SL g3134 ( 
.A(n_3004),
.B(n_3086),
.Y(n_3134)
);

NAND2xp5_ASAP7_75t_L g3135 ( 
.A(n_3092),
.B(n_165),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_2999),
.Y(n_3136)
);

NAND2x1p5_ASAP7_75t_L g3137 ( 
.A(n_3046),
.B(n_167),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_3079),
.Y(n_3138)
);

AND2x2_ASAP7_75t_L g3139 ( 
.A(n_3085),
.B(n_166),
.Y(n_3139)
);

AND2x2_ASAP7_75t_L g3140 ( 
.A(n_3087),
.B(n_168),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_3088),
.Y(n_3141)
);

INVxp67_ASAP7_75t_SL g3142 ( 
.A(n_3099),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_L g3143 ( 
.A(n_3091),
.B(n_3095),
.Y(n_3143)
);

OAI33xp33_ASAP7_75t_L g3144 ( 
.A1(n_3020),
.A2(n_172),
.A3(n_179),
.B1(n_169),
.B2(n_170),
.B3(n_177),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_3113),
.Y(n_3145)
);

OAI221xp5_ASAP7_75t_L g3146 ( 
.A1(n_3000),
.A2(n_184),
.B1(n_181),
.B2(n_182),
.C(n_185),
.Y(n_3146)
);

OAI21xp33_ASAP7_75t_L g3147 ( 
.A1(n_3009),
.A2(n_181),
.B(n_182),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_L g3148 ( 
.A(n_3019),
.B(n_186),
.Y(n_3148)
);

INVx2_ASAP7_75t_L g3149 ( 
.A(n_3023),
.Y(n_3149)
);

NOR2x1_ASAP7_75t_L g3150 ( 
.A(n_3076),
.B(n_186),
.Y(n_3150)
);

NOR3xp33_ASAP7_75t_SL g3151 ( 
.A(n_3012),
.B(n_187),
.C(n_188),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_3070),
.Y(n_3152)
);

NAND2xp33_ASAP7_75t_SL g3153 ( 
.A(n_3083),
.B(n_187),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_3090),
.Y(n_3154)
);

INVx2_ASAP7_75t_L g3155 ( 
.A(n_3015),
.Y(n_3155)
);

AOI22xp33_ASAP7_75t_L g3156 ( 
.A1(n_3017),
.A2(n_192),
.B1(n_189),
.B2(n_191),
.Y(n_3156)
);

OR2x2_ASAP7_75t_L g3157 ( 
.A(n_3097),
.B(n_193),
.Y(n_3157)
);

NAND2xp5_ASAP7_75t_L g3158 ( 
.A(n_3015),
.B(n_194),
.Y(n_3158)
);

INVx1_ASAP7_75t_L g3159 ( 
.A(n_3110),
.Y(n_3159)
);

NOR2xp33_ASAP7_75t_L g3160 ( 
.A(n_3108),
.B(n_196),
.Y(n_3160)
);

NOR2xp33_ASAP7_75t_L g3161 ( 
.A(n_3007),
.B(n_196),
.Y(n_3161)
);

NAND2xp33_ASAP7_75t_L g3162 ( 
.A(n_3011),
.B(n_3036),
.Y(n_3162)
);

AND2x2_ASAP7_75t_L g3163 ( 
.A(n_3014),
.B(n_197),
.Y(n_3163)
);

AND2x2_ASAP7_75t_L g3164 ( 
.A(n_3040),
.B(n_198),
.Y(n_3164)
);

NAND2x1p5_ASAP7_75t_L g3165 ( 
.A(n_3051),
.B(n_200),
.Y(n_3165)
);

HB1xp67_ASAP7_75t_L g3166 ( 
.A(n_3028),
.Y(n_3166)
);

NAND2xp5_ASAP7_75t_L g3167 ( 
.A(n_3065),
.B(n_199),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_3058),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_3058),
.Y(n_3169)
);

AND2x2_ASAP7_75t_L g3170 ( 
.A(n_3030),
.B(n_200),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_L g3171 ( 
.A(n_3025),
.B(n_201),
.Y(n_3171)
);

OR2x2_ASAP7_75t_L g3172 ( 
.A(n_3082),
.B(n_203),
.Y(n_3172)
);

NAND2xp33_ASAP7_75t_L g3173 ( 
.A(n_2997),
.B(n_203),
.Y(n_3173)
);

XOR2x2_ASAP7_75t_L g3174 ( 
.A(n_3067),
.B(n_204),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_3059),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_3044),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_L g3177 ( 
.A(n_3077),
.B(n_204),
.Y(n_3177)
);

INVxp67_ASAP7_75t_L g3178 ( 
.A(n_3050),
.Y(n_3178)
);

INVx2_ASAP7_75t_L g3179 ( 
.A(n_3039),
.Y(n_3179)
);

NAND2xp5_ASAP7_75t_L g3180 ( 
.A(n_3074),
.B(n_205),
.Y(n_3180)
);

INVx4_ASAP7_75t_L g3181 ( 
.A(n_3029),
.Y(n_3181)
);

NOR2xp67_ASAP7_75t_SL g3182 ( 
.A(n_3100),
.B(n_205),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_3035),
.Y(n_3183)
);

OR2x2_ASAP7_75t_L g3184 ( 
.A(n_3022),
.B(n_206),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_3013),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_3003),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_L g3187 ( 
.A(n_3062),
.B(n_207),
.Y(n_3187)
);

NOR2xp33_ASAP7_75t_L g3188 ( 
.A(n_3089),
.B(n_208),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_3005),
.Y(n_3189)
);

INVx2_ASAP7_75t_SL g3190 ( 
.A(n_3081),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_3104),
.Y(n_3191)
);

NAND2x1_ASAP7_75t_L g3192 ( 
.A(n_3001),
.B(n_208),
.Y(n_3192)
);

INVx2_ASAP7_75t_SL g3193 ( 
.A(n_3031),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_3073),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_L g3195 ( 
.A(n_3063),
.B(n_209),
.Y(n_3195)
);

INVx2_ASAP7_75t_L g3196 ( 
.A(n_3032),
.Y(n_3196)
);

NOR2xp33_ASAP7_75t_L g3197 ( 
.A(n_3096),
.B(n_3105),
.Y(n_3197)
);

INVxp33_ASAP7_75t_L g3198 ( 
.A(n_3056),
.Y(n_3198)
);

OR4x1_ASAP7_75t_L g3199 ( 
.A(n_3016),
.B(n_214),
.C(n_212),
.D(n_213),
.Y(n_3199)
);

INVx2_ASAP7_75t_SL g3200 ( 
.A(n_3064),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_3034),
.Y(n_3201)
);

NOR2x1_ASAP7_75t_L g3202 ( 
.A(n_3102),
.B(n_213),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_L g3203 ( 
.A(n_3101),
.B(n_214),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_L g3204 ( 
.A(n_3080),
.B(n_215),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_L g3205 ( 
.A(n_3098),
.B(n_216),
.Y(n_3205)
);

AND2x2_ASAP7_75t_L g3206 ( 
.A(n_3119),
.B(n_3054),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_3120),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_L g3208 ( 
.A(n_3131),
.B(n_3112),
.Y(n_3208)
);

NAND2xp5_ASAP7_75t_L g3209 ( 
.A(n_3133),
.B(n_3068),
.Y(n_3209)
);

AND2x2_ASAP7_75t_L g3210 ( 
.A(n_3142),
.B(n_3006),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_3137),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_L g3212 ( 
.A(n_3127),
.B(n_3078),
.Y(n_3212)
);

INVxp67_ASAP7_75t_L g3213 ( 
.A(n_3116),
.Y(n_3213)
);

AND2x2_ASAP7_75t_L g3214 ( 
.A(n_3128),
.B(n_3018),
.Y(n_3214)
);

OR2x2_ASAP7_75t_L g3215 ( 
.A(n_3165),
.B(n_3155),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_3115),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_3117),
.Y(n_3217)
);

INVx1_ASAP7_75t_L g3218 ( 
.A(n_3132),
.Y(n_3218)
);

NAND2xp5_ASAP7_75t_L g3219 ( 
.A(n_3185),
.B(n_3055),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_3118),
.Y(n_3220)
);

NAND2xp5_ASAP7_75t_L g3221 ( 
.A(n_3149),
.B(n_3053),
.Y(n_3221)
);

OAI31xp33_ASAP7_75t_SL g3222 ( 
.A1(n_3202),
.A2(n_3060),
.A3(n_3021),
.B(n_3041),
.Y(n_3222)
);

INVx1_ASAP7_75t_L g3223 ( 
.A(n_3139),
.Y(n_3223)
);

AND2x2_ASAP7_75t_L g3224 ( 
.A(n_3121),
.B(n_3125),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_3140),
.Y(n_3225)
);

AND2x2_ASAP7_75t_L g3226 ( 
.A(n_3130),
.B(n_3047),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_3143),
.Y(n_3227)
);

INVx3_ASAP7_75t_L g3228 ( 
.A(n_3181),
.Y(n_3228)
);

AND2x2_ASAP7_75t_L g3229 ( 
.A(n_3194),
.B(n_3049),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_L g3230 ( 
.A(n_3168),
.B(n_3042),
.Y(n_3230)
);

NAND3xp33_ASAP7_75t_L g3231 ( 
.A(n_3162),
.B(n_3026),
.C(n_3008),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_3123),
.Y(n_3232)
);

INVx2_ASAP7_75t_L g3233 ( 
.A(n_3169),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_3166),
.Y(n_3234)
);

NAND3xp33_ASAP7_75t_L g3235 ( 
.A(n_3150),
.B(n_3033),
.C(n_3024),
.Y(n_3235)
);

NOR2xp33_ASAP7_75t_L g3236 ( 
.A(n_3134),
.B(n_3057),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_L g3237 ( 
.A(n_3197),
.B(n_3027),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_3158),
.Y(n_3238)
);

AND2x2_ASAP7_75t_L g3239 ( 
.A(n_3190),
.B(n_3061),
.Y(n_3239)
);

NAND2xp5_ASAP7_75t_L g3240 ( 
.A(n_3200),
.B(n_3038),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_3124),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_L g3242 ( 
.A(n_3129),
.B(n_3052),
.Y(n_3242)
);

A2O1A1Ixp33_ASAP7_75t_L g3243 ( 
.A1(n_3188),
.A2(n_3037),
.B(n_3043),
.C(n_3107),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_L g3244 ( 
.A(n_3136),
.B(n_217),
.Y(n_3244)
);

NAND2x2_ASAP7_75t_L g3245 ( 
.A(n_3193),
.B(n_3192),
.Y(n_3245)
);

INVx2_ASAP7_75t_L g3246 ( 
.A(n_3184),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_3122),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_3170),
.Y(n_3248)
);

NOR2xp33_ASAP7_75t_L g3249 ( 
.A(n_3181),
.B(n_218),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_L g3250 ( 
.A(n_3138),
.B(n_218),
.Y(n_3250)
);

AND2x2_ASAP7_75t_L g3251 ( 
.A(n_3151),
.B(n_222),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_L g3252 ( 
.A(n_3141),
.B(n_223),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_3148),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_3163),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_3164),
.Y(n_3255)
);

AOI22x1_ASAP7_75t_SL g3256 ( 
.A1(n_3145),
.A2(n_226),
.B1(n_224),
.B2(n_225),
.Y(n_3256)
);

INVxp67_ASAP7_75t_L g3257 ( 
.A(n_3182),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_3135),
.Y(n_3258)
);

AOI22xp33_ASAP7_75t_L g3259 ( 
.A1(n_3191),
.A2(n_229),
.B1(n_226),
.B2(n_227),
.Y(n_3259)
);

AND2x2_ASAP7_75t_L g3260 ( 
.A(n_3179),
.B(n_227),
.Y(n_3260)
);

NOR2x1_ASAP7_75t_L g3261 ( 
.A(n_3172),
.B(n_229),
.Y(n_3261)
);

NOR2xp33_ASAP7_75t_L g3262 ( 
.A(n_3126),
.B(n_231),
.Y(n_3262)
);

INVx1_ASAP7_75t_SL g3263 ( 
.A(n_3153),
.Y(n_3263)
);

NAND2xp5_ASAP7_75t_L g3264 ( 
.A(n_3183),
.B(n_231),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_3171),
.Y(n_3265)
);

NAND2xp5_ASAP7_75t_L g3266 ( 
.A(n_3160),
.B(n_233),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_L g3267 ( 
.A(n_3175),
.B(n_234),
.Y(n_3267)
);

INVx2_ASAP7_75t_L g3268 ( 
.A(n_3157),
.Y(n_3268)
);

INVx2_ASAP7_75t_SL g3269 ( 
.A(n_3176),
.Y(n_3269)
);

HB1xp67_ASAP7_75t_L g3270 ( 
.A(n_3167),
.Y(n_3270)
);

NOR2x1_ASAP7_75t_L g3271 ( 
.A(n_3180),
.B(n_235),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_3161),
.Y(n_3272)
);

OR2x2_ASAP7_75t_L g3273 ( 
.A(n_3177),
.B(n_3204),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_3174),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_3147),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_L g3276 ( 
.A(n_3152),
.B(n_237),
.Y(n_3276)
);

INVx1_ASAP7_75t_L g3277 ( 
.A(n_3154),
.Y(n_3277)
);

AND2x2_ASAP7_75t_L g3278 ( 
.A(n_3159),
.B(n_240),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_L g3279 ( 
.A(n_3196),
.B(n_241),
.Y(n_3279)
);

AND2x2_ASAP7_75t_L g3280 ( 
.A(n_3198),
.B(n_241),
.Y(n_3280)
);

INVx3_ASAP7_75t_L g3281 ( 
.A(n_3201),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_3187),
.Y(n_3282)
);

AOI22xp33_ASAP7_75t_SL g3283 ( 
.A1(n_3205),
.A2(n_244),
.B1(n_242),
.B2(n_243),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_SL g3284 ( 
.A(n_3195),
.B(n_243),
.Y(n_3284)
);

AND2x2_ASAP7_75t_L g3285 ( 
.A(n_3186),
.B(n_245),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_3203),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_3156),
.B(n_246),
.Y(n_3287)
);

OR2x2_ASAP7_75t_L g3288 ( 
.A(n_3189),
.B(n_246),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_3146),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_3178),
.B(n_248),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_L g3291 ( 
.A(n_3173),
.B(n_3199),
.Y(n_3291)
);

AOI22xp33_ASAP7_75t_L g3292 ( 
.A1(n_3144),
.A2(n_251),
.B1(n_249),
.B2(n_250),
.Y(n_3292)
);

INVx1_ASAP7_75t_SL g3293 ( 
.A(n_3133),
.Y(n_3293)
);

INVxp33_ASAP7_75t_L g3294 ( 
.A(n_3120),
.Y(n_3294)
);

AND2x2_ASAP7_75t_L g3295 ( 
.A(n_3119),
.B(n_254),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_3120),
.Y(n_3296)
);

INVx2_ASAP7_75t_L g3297 ( 
.A(n_3120),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_3120),
.Y(n_3298)
);

AOI21xp33_ASAP7_75t_L g3299 ( 
.A1(n_3131),
.A2(n_255),
.B(n_256),
.Y(n_3299)
);

INVx1_ASAP7_75t_SL g3300 ( 
.A(n_3133),
.Y(n_3300)
);

BUFx2_ASAP7_75t_L g3301 ( 
.A(n_3120),
.Y(n_3301)
);

AND2x4_ASAP7_75t_SL g3302 ( 
.A(n_3120),
.B(n_255),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_SL g3303 ( 
.A(n_3133),
.B(n_256),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_3120),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_3120),
.Y(n_3305)
);

NOR2xp33_ASAP7_75t_L g3306 ( 
.A(n_3120),
.B(n_257),
.Y(n_3306)
);

OAI21xp5_ASAP7_75t_L g3307 ( 
.A1(n_3120),
.A2(n_258),
.B(n_259),
.Y(n_3307)
);

OAI21xp33_ASAP7_75t_L g3308 ( 
.A1(n_3194),
.A2(n_258),
.B(n_259),
.Y(n_3308)
);

AND2x4_ASAP7_75t_L g3309 ( 
.A(n_3120),
.B(n_261),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_3120),
.Y(n_3310)
);

OAI21xp33_ASAP7_75t_L g3311 ( 
.A1(n_3194),
.A2(n_265),
.B(n_267),
.Y(n_3311)
);

INVx1_ASAP7_75t_L g3312 ( 
.A(n_3120),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_3120),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_L g3314 ( 
.A(n_3120),
.B(n_265),
.Y(n_3314)
);

INVx1_ASAP7_75t_SL g3315 ( 
.A(n_3133),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_L g3316 ( 
.A(n_3120),
.B(n_269),
.Y(n_3316)
);

INVx2_ASAP7_75t_L g3317 ( 
.A(n_3120),
.Y(n_3317)
);

OR2x2_ASAP7_75t_L g3318 ( 
.A(n_3133),
.B(n_271),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_L g3319 ( 
.A(n_3120),
.B(n_272),
.Y(n_3319)
);

XNOR2xp5_ASAP7_75t_L g3320 ( 
.A(n_3174),
.B(n_273),
.Y(n_3320)
);

NAND2xp5_ASAP7_75t_L g3321 ( 
.A(n_3120),
.B(n_273),
.Y(n_3321)
);

NAND2xp5_ASAP7_75t_L g3322 ( 
.A(n_3120),
.B(n_274),
.Y(n_3322)
);

NOR3xp33_ASAP7_75t_SL g3323 ( 
.A(n_3236),
.B(n_3209),
.C(n_3231),
.Y(n_3323)
);

INVxp67_ASAP7_75t_L g3324 ( 
.A(n_3301),
.Y(n_3324)
);

AOI221xp5_ASAP7_75t_L g3325 ( 
.A1(n_3294),
.A2(n_277),
.B1(n_279),
.B2(n_276),
.C(n_278),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_3228),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_3228),
.Y(n_3327)
);

AOI21xp5_ASAP7_75t_L g3328 ( 
.A1(n_3212),
.A2(n_275),
.B(n_280),
.Y(n_3328)
);

NOR3xp33_ASAP7_75t_SL g3329 ( 
.A(n_3208),
.B(n_281),
.C(n_282),
.Y(n_3329)
);

INVx1_ASAP7_75t_L g3330 ( 
.A(n_3215),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3302),
.Y(n_3331)
);

NOR2xp67_ASAP7_75t_L g3332 ( 
.A(n_3211),
.B(n_282),
.Y(n_3332)
);

NOR3xp33_ASAP7_75t_L g3333 ( 
.A(n_3235),
.B(n_294),
.C(n_283),
.Y(n_3333)
);

AOI21xp5_ASAP7_75t_L g3334 ( 
.A1(n_3291),
.A2(n_283),
.B(n_284),
.Y(n_3334)
);

NAND2xp5_ASAP7_75t_L g3335 ( 
.A(n_3309),
.B(n_285),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_L g3336 ( 
.A(n_3309),
.B(n_3293),
.Y(n_3336)
);

O2A1O1Ixp33_ASAP7_75t_L g3337 ( 
.A1(n_3243),
.A2(n_290),
.B(n_286),
.C(n_289),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_L g3338 ( 
.A(n_3300),
.B(n_289),
.Y(n_3338)
);

INVx1_ASAP7_75t_L g3339 ( 
.A(n_3297),
.Y(n_3339)
);

OAI21xp33_ASAP7_75t_L g3340 ( 
.A1(n_3315),
.A2(n_290),
.B(n_291),
.Y(n_3340)
);

NAND3xp33_ASAP7_75t_L g3341 ( 
.A(n_3222),
.B(n_291),
.C(n_293),
.Y(n_3341)
);

INVx2_ASAP7_75t_L g3342 ( 
.A(n_3317),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_3207),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_3296),
.Y(n_3344)
);

OAI21xp5_ASAP7_75t_SL g3345 ( 
.A1(n_3292),
.A2(n_293),
.B(n_295),
.Y(n_3345)
);

A2O1A1Ixp33_ASAP7_75t_L g3346 ( 
.A1(n_3306),
.A2(n_301),
.B(n_295),
.C(n_298),
.Y(n_3346)
);

NOR2x1_ASAP7_75t_L g3347 ( 
.A(n_3261),
.B(n_302),
.Y(n_3347)
);

AND4x1_ASAP7_75t_L g3348 ( 
.A(n_3271),
.B(n_305),
.C(n_302),
.D(n_304),
.Y(n_3348)
);

INVx1_ASAP7_75t_L g3349 ( 
.A(n_3298),
.Y(n_3349)
);

NAND3xp33_ASAP7_75t_L g3350 ( 
.A(n_3304),
.B(n_3310),
.C(n_3305),
.Y(n_3350)
);

INVx2_ASAP7_75t_SL g3351 ( 
.A(n_3312),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_3313),
.Y(n_3352)
);

OR2x2_ASAP7_75t_L g3353 ( 
.A(n_3233),
.B(n_306),
.Y(n_3353)
);

OAI22xp33_ASAP7_75t_L g3354 ( 
.A1(n_3245),
.A2(n_311),
.B1(n_307),
.B2(n_310),
.Y(n_3354)
);

NOR4xp25_ASAP7_75t_SL g3355 ( 
.A(n_3234),
.B(n_311),
.C(n_307),
.D(n_310),
.Y(n_3355)
);

XNOR2xp5_ASAP7_75t_L g3356 ( 
.A(n_3320),
.B(n_3256),
.Y(n_3356)
);

AOI211x1_ASAP7_75t_L g3357 ( 
.A1(n_3308),
.A2(n_314),
.B(n_312),
.C(n_313),
.Y(n_3357)
);

NOR3xp33_ASAP7_75t_L g3358 ( 
.A(n_3257),
.B(n_312),
.C(n_313),
.Y(n_3358)
);

AOI21xp5_ASAP7_75t_L g3359 ( 
.A1(n_3303),
.A2(n_314),
.B(n_316),
.Y(n_3359)
);

NOR2xp33_ASAP7_75t_L g3360 ( 
.A(n_3311),
.B(n_317),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_SL g3361 ( 
.A(n_3263),
.B(n_317),
.Y(n_3361)
);

AOI21xp33_ASAP7_75t_L g3362 ( 
.A1(n_3274),
.A2(n_318),
.B(n_319),
.Y(n_3362)
);

INVx2_ASAP7_75t_L g3363 ( 
.A(n_3318),
.Y(n_3363)
);

INVx2_ASAP7_75t_L g3364 ( 
.A(n_3295),
.Y(n_3364)
);

NAND2xp5_ASAP7_75t_SL g3365 ( 
.A(n_3269),
.B(n_320),
.Y(n_3365)
);

INVx2_ASAP7_75t_L g3366 ( 
.A(n_3288),
.Y(n_3366)
);

NOR3xp33_ASAP7_75t_L g3367 ( 
.A(n_3240),
.B(n_321),
.C(n_322),
.Y(n_3367)
);

OAI211xp5_ASAP7_75t_SL g3368 ( 
.A1(n_3213),
.A2(n_323),
.B(n_321),
.C(n_322),
.Y(n_3368)
);

OR2x2_ASAP7_75t_L g3369 ( 
.A(n_3314),
.B(n_323),
.Y(n_3369)
);

INVx2_ASAP7_75t_L g3370 ( 
.A(n_3224),
.Y(n_3370)
);

NOR2xp33_ASAP7_75t_L g3371 ( 
.A(n_3223),
.B(n_324),
.Y(n_3371)
);

AOI211xp5_ASAP7_75t_L g3372 ( 
.A1(n_3216),
.A2(n_3217),
.B(n_3275),
.C(n_3289),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_L g3373 ( 
.A(n_3251),
.B(n_330),
.Y(n_3373)
);

AO21x1_ASAP7_75t_L g3374 ( 
.A1(n_3316),
.A2(n_330),
.B(n_331),
.Y(n_3374)
);

NOR2x1_ASAP7_75t_L g3375 ( 
.A(n_3319),
.B(n_331),
.Y(n_3375)
);

NOR3xp33_ASAP7_75t_L g3376 ( 
.A(n_3237),
.B(n_332),
.C(n_333),
.Y(n_3376)
);

O2A1O1Ixp33_ASAP7_75t_L g3377 ( 
.A1(n_3321),
.A2(n_335),
.B(n_333),
.C(n_334),
.Y(n_3377)
);

HB1xp67_ASAP7_75t_L g3378 ( 
.A(n_3322),
.Y(n_3378)
);

AND2x2_ASAP7_75t_L g3379 ( 
.A(n_3206),
.B(n_339),
.Y(n_3379)
);

AND2x2_ASAP7_75t_L g3380 ( 
.A(n_3225),
.B(n_340),
.Y(n_3380)
);

AOI211xp5_ASAP7_75t_L g3381 ( 
.A1(n_3227),
.A2(n_343),
.B(n_340),
.C(n_341),
.Y(n_3381)
);

NAND2x1_ASAP7_75t_L g3382 ( 
.A(n_3281),
.B(n_341),
.Y(n_3382)
);

AOI22xp5_ASAP7_75t_L g3383 ( 
.A1(n_3239),
.A2(n_345),
.B1(n_343),
.B2(n_344),
.Y(n_3383)
);

XOR2x2_ASAP7_75t_L g3384 ( 
.A(n_3229),
.B(n_346),
.Y(n_3384)
);

NAND3xp33_ASAP7_75t_L g3385 ( 
.A(n_3283),
.B(n_346),
.C(n_347),
.Y(n_3385)
);

NAND4xp25_ASAP7_75t_L g3386 ( 
.A(n_3219),
.B(n_350),
.C(n_348),
.D(n_349),
.Y(n_3386)
);

NAND5xp2_ASAP7_75t_L g3387 ( 
.A(n_3232),
.B(n_353),
.C(n_349),
.D(n_352),
.E(n_355),
.Y(n_3387)
);

NAND4xp25_ASAP7_75t_L g3388 ( 
.A(n_3273),
.B(n_359),
.C(n_355),
.D(n_357),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_SL g3389 ( 
.A(n_3220),
.B(n_359),
.Y(n_3389)
);

OAI22x1_ASAP7_75t_L g3390 ( 
.A1(n_3248),
.A2(n_3255),
.B1(n_3254),
.B2(n_3246),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_SL g3391 ( 
.A(n_3307),
.B(n_360),
.Y(n_3391)
);

OAI21xp5_ASAP7_75t_L g3392 ( 
.A1(n_3324),
.A2(n_3260),
.B(n_3218),
.Y(n_3392)
);

XNOR2xp5_ASAP7_75t_L g3393 ( 
.A(n_3356),
.B(n_3226),
.Y(n_3393)
);

AOI221xp5_ASAP7_75t_L g3394 ( 
.A1(n_3341),
.A2(n_3277),
.B1(n_3272),
.B2(n_3282),
.C(n_3286),
.Y(n_3394)
);

AOI221xp5_ASAP7_75t_L g3395 ( 
.A1(n_3354),
.A2(n_3247),
.B1(n_3210),
.B2(n_3238),
.C(n_3253),
.Y(n_3395)
);

XNOR2xp5_ASAP7_75t_L g3396 ( 
.A(n_3384),
.B(n_3270),
.Y(n_3396)
);

AOI221xp5_ASAP7_75t_L g3397 ( 
.A1(n_3350),
.A2(n_3241),
.B1(n_3258),
.B2(n_3265),
.C(n_3299),
.Y(n_3397)
);

NOR3xp33_ASAP7_75t_L g3398 ( 
.A(n_3330),
.B(n_3221),
.C(n_3230),
.Y(n_3398)
);

AOI221x1_ASAP7_75t_L g3399 ( 
.A1(n_3333),
.A2(n_3250),
.B1(n_3252),
.B2(n_3244),
.C(n_3267),
.Y(n_3399)
);

NOR4xp25_ASAP7_75t_L g3400 ( 
.A(n_3336),
.B(n_3242),
.C(n_3214),
.D(n_3268),
.Y(n_3400)
);

OAI211xp5_ASAP7_75t_SL g3401 ( 
.A1(n_3323),
.A2(n_3284),
.B(n_3259),
.C(n_3266),
.Y(n_3401)
);

NOR2xp33_ASAP7_75t_L g3402 ( 
.A(n_3348),
.B(n_3262),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_3332),
.B(n_3249),
.Y(n_3403)
);

AOI211xp5_ASAP7_75t_L g3404 ( 
.A1(n_3345),
.A2(n_3276),
.B(n_3278),
.C(n_3287),
.Y(n_3404)
);

AOI22xp33_ASAP7_75t_L g3405 ( 
.A1(n_3342),
.A2(n_3370),
.B1(n_3351),
.B2(n_3339),
.Y(n_3405)
);

AOI22x1_ASAP7_75t_SL g3406 ( 
.A1(n_3331),
.A2(n_3280),
.B1(n_3264),
.B2(n_3290),
.Y(n_3406)
);

NAND2xp5_ASAP7_75t_SL g3407 ( 
.A(n_3347),
.B(n_3279),
.Y(n_3407)
);

AOI222xp33_ASAP7_75t_L g3408 ( 
.A1(n_3326),
.A2(n_3285),
.B1(n_363),
.B2(n_365),
.C1(n_361),
.C2(n_362),
.Y(n_3408)
);

A2O1A1Ixp33_ASAP7_75t_L g3409 ( 
.A1(n_3337),
.A2(n_366),
.B(n_364),
.C(n_365),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_3382),
.Y(n_3410)
);

NOR2xp33_ASAP7_75t_L g3411 ( 
.A(n_3388),
.B(n_367),
.Y(n_3411)
);

AOI222xp33_ASAP7_75t_L g3412 ( 
.A1(n_3327),
.A2(n_3349),
.B1(n_3344),
.B2(n_3352),
.C1(n_3343),
.C2(n_3390),
.Y(n_3412)
);

AOI221xp5_ASAP7_75t_L g3413 ( 
.A1(n_3376),
.A2(n_371),
.B1(n_369),
.B2(n_370),
.C(n_372),
.Y(n_3413)
);

AOI221xp5_ASAP7_75t_L g3414 ( 
.A1(n_3372),
.A2(n_372),
.B1(n_369),
.B2(n_370),
.C(n_373),
.Y(n_3414)
);

AOI21xp33_ASAP7_75t_L g3415 ( 
.A1(n_3363),
.A2(n_374),
.B(n_375),
.Y(n_3415)
);

NOR4xp25_ASAP7_75t_L g3416 ( 
.A(n_3364),
.B(n_377),
.C(n_375),
.D(n_376),
.Y(n_3416)
);

NAND4xp75_ASAP7_75t_L g3417 ( 
.A(n_3375),
.B(n_379),
.C(n_376),
.D(n_377),
.Y(n_3417)
);

NAND4xp25_ASAP7_75t_SL g3418 ( 
.A(n_3338),
.B(n_385),
.C(n_380),
.D(n_381),
.Y(n_3418)
);

OAI21xp5_ASAP7_75t_L g3419 ( 
.A1(n_3385),
.A2(n_3334),
.B(n_3329),
.Y(n_3419)
);

NOR2xp67_ASAP7_75t_L g3420 ( 
.A(n_3387),
.B(n_380),
.Y(n_3420)
);

AOI21xp5_ASAP7_75t_L g3421 ( 
.A1(n_3391),
.A2(n_381),
.B(n_387),
.Y(n_3421)
);

AOI211xp5_ASAP7_75t_L g3422 ( 
.A1(n_3374),
.A2(n_392),
.B(n_388),
.C(n_390),
.Y(n_3422)
);

A2O1A1Ixp33_ASAP7_75t_L g3423 ( 
.A1(n_3377),
.A2(n_397),
.B(n_394),
.C(n_396),
.Y(n_3423)
);

NAND4xp75_ASAP7_75t_L g3424 ( 
.A(n_3379),
.B(n_399),
.C(n_397),
.D(n_398),
.Y(n_3424)
);

NAND4xp25_ASAP7_75t_SL g3425 ( 
.A(n_3366),
.B(n_401),
.C(n_399),
.D(n_400),
.Y(n_3425)
);

OAI21xp5_ASAP7_75t_L g3426 ( 
.A1(n_3328),
.A2(n_403),
.B(n_404),
.Y(n_3426)
);

AOI21xp5_ASAP7_75t_L g3427 ( 
.A1(n_3361),
.A2(n_404),
.B(n_405),
.Y(n_3427)
);

AOI211xp5_ASAP7_75t_L g3428 ( 
.A1(n_3362),
.A2(n_408),
.B(n_406),
.C(n_407),
.Y(n_3428)
);

AOI221xp5_ASAP7_75t_L g3429 ( 
.A1(n_3357),
.A2(n_410),
.B1(n_407),
.B2(n_409),
.C(n_411),
.Y(n_3429)
);

AOI221xp5_ASAP7_75t_L g3430 ( 
.A1(n_3367),
.A2(n_411),
.B1(n_409),
.B2(n_410),
.C(n_414),
.Y(n_3430)
);

AOI211xp5_ASAP7_75t_L g3431 ( 
.A1(n_3340),
.A2(n_417),
.B(n_415),
.C(n_416),
.Y(n_3431)
);

OAI21xp33_ASAP7_75t_L g3432 ( 
.A1(n_3378),
.A2(n_416),
.B(n_417),
.Y(n_3432)
);

AOI211xp5_ASAP7_75t_L g3433 ( 
.A1(n_3368),
.A2(n_420),
.B(n_418),
.C(n_419),
.Y(n_3433)
);

OAI221xp5_ASAP7_75t_L g3434 ( 
.A1(n_3358),
.A2(n_422),
.B1(n_418),
.B2(n_420),
.C(n_423),
.Y(n_3434)
);

AOI211xp5_ASAP7_75t_L g3435 ( 
.A1(n_3359),
.A2(n_425),
.B(n_422),
.C(n_423),
.Y(n_3435)
);

OAI222xp33_ASAP7_75t_L g3436 ( 
.A1(n_3373),
.A2(n_428),
.B1(n_432),
.B2(n_426),
.C1(n_427),
.C2(n_430),
.Y(n_3436)
);

AOI21xp5_ASAP7_75t_L g3437 ( 
.A1(n_3389),
.A2(n_433),
.B(n_434),
.Y(n_3437)
);

OAI21xp33_ASAP7_75t_L g3438 ( 
.A1(n_3386),
.A2(n_3360),
.B(n_3380),
.Y(n_3438)
);

OAI22x1_ASAP7_75t_L g3439 ( 
.A1(n_3383),
.A2(n_438),
.B1(n_435),
.B2(n_437),
.Y(n_3439)
);

NAND4xp25_ASAP7_75t_L g3440 ( 
.A(n_3405),
.B(n_3381),
.C(n_3325),
.D(n_3371),
.Y(n_3440)
);

A2O1A1Ixp33_ASAP7_75t_L g3441 ( 
.A1(n_3420),
.A2(n_3346),
.B(n_3365),
.C(n_3369),
.Y(n_3441)
);

OAI211xp5_ASAP7_75t_L g3442 ( 
.A1(n_3412),
.A2(n_3355),
.B(n_3335),
.C(n_3353),
.Y(n_3442)
);

AOI211xp5_ASAP7_75t_L g3443 ( 
.A1(n_3400),
.A2(n_440),
.B(n_437),
.C(n_439),
.Y(n_3443)
);

AOI222xp33_ASAP7_75t_L g3444 ( 
.A1(n_3419),
.A2(n_442),
.B1(n_444),
.B2(n_440),
.C1(n_441),
.C2(n_443),
.Y(n_3444)
);

OAI21xp5_ASAP7_75t_L g3445 ( 
.A1(n_3393),
.A2(n_445),
.B(n_447),
.Y(n_3445)
);

AOI221xp5_ASAP7_75t_L g3446 ( 
.A1(n_3416),
.A2(n_448),
.B1(n_445),
.B2(n_447),
.C(n_449),
.Y(n_3446)
);

AOI211xp5_ASAP7_75t_SL g3447 ( 
.A1(n_3410),
.A2(n_452),
.B(n_450),
.C(n_451),
.Y(n_3447)
);

OAI221xp5_ASAP7_75t_SL g3448 ( 
.A1(n_3397),
.A2(n_453),
.B1(n_450),
.B2(n_452),
.C(n_454),
.Y(n_3448)
);

INVx1_ASAP7_75t_L g3449 ( 
.A(n_3396),
.Y(n_3449)
);

OAI22xp33_ASAP7_75t_SL g3450 ( 
.A1(n_3403),
.A2(n_456),
.B1(n_453),
.B2(n_455),
.Y(n_3450)
);

OAI221xp5_ASAP7_75t_L g3451 ( 
.A1(n_3394),
.A2(n_458),
.B1(n_455),
.B2(n_456),
.C(n_459),
.Y(n_3451)
);

A2O1A1Ixp33_ASAP7_75t_L g3452 ( 
.A1(n_3411),
.A2(n_461),
.B(n_459),
.C(n_460),
.Y(n_3452)
);

OAI221xp5_ASAP7_75t_L g3453 ( 
.A1(n_3392),
.A2(n_466),
.B1(n_462),
.B2(n_463),
.C(n_467),
.Y(n_3453)
);

AOI221xp5_ASAP7_75t_L g3454 ( 
.A1(n_3401),
.A2(n_468),
.B1(n_466),
.B2(n_467),
.C(n_469),
.Y(n_3454)
);

AOI211xp5_ASAP7_75t_SL g3455 ( 
.A1(n_3402),
.A2(n_472),
.B(n_469),
.C(n_470),
.Y(n_3455)
);

OAI311xp33_ASAP7_75t_L g3456 ( 
.A1(n_3395),
.A2(n_474),
.A3(n_470),
.B1(n_473),
.C1(n_475),
.Y(n_3456)
);

AOI22xp5_ASAP7_75t_L g3457 ( 
.A1(n_3398),
.A2(n_477),
.B1(n_475),
.B2(n_476),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3417),
.Y(n_3458)
);

AOI21xp5_ASAP7_75t_L g3459 ( 
.A1(n_3407),
.A2(n_3421),
.B(n_3437),
.Y(n_3459)
);

XNOR2x1_ASAP7_75t_L g3460 ( 
.A(n_3424),
.B(n_476),
.Y(n_3460)
);

XNOR2xp5_ASAP7_75t_L g3461 ( 
.A(n_3406),
.B(n_477),
.Y(n_3461)
);

NAND3xp33_ASAP7_75t_SL g3462 ( 
.A(n_3422),
.B(n_478),
.C(n_479),
.Y(n_3462)
);

OAI321xp33_ASAP7_75t_L g3463 ( 
.A1(n_3438),
.A2(n_481),
.A3(n_483),
.B1(n_478),
.B2(n_480),
.C(n_482),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_3439),
.Y(n_3464)
);

HB1xp67_ASAP7_75t_L g3465 ( 
.A(n_3425),
.Y(n_3465)
);

AOI211x1_ASAP7_75t_L g3466 ( 
.A1(n_3426),
.A2(n_488),
.B(n_485),
.C(n_486),
.Y(n_3466)
);

AO22x2_ASAP7_75t_L g3467 ( 
.A1(n_3399),
.A2(n_490),
.B1(n_485),
.B2(n_489),
.Y(n_3467)
);

OAI211xp5_ASAP7_75t_L g3468 ( 
.A1(n_3404),
.A2(n_492),
.B(n_489),
.C(n_491),
.Y(n_3468)
);

OAI21xp5_ASAP7_75t_L g3469 ( 
.A1(n_3461),
.A2(n_3423),
.B(n_3409),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_3467),
.Y(n_3470)
);

OAI321xp33_ASAP7_75t_L g3471 ( 
.A1(n_3440),
.A2(n_3429),
.A3(n_3433),
.B1(n_3414),
.B2(n_3434),
.C(n_3435),
.Y(n_3471)
);

OAI221xp5_ASAP7_75t_L g3472 ( 
.A1(n_3443),
.A2(n_3413),
.B1(n_3430),
.B2(n_3428),
.C(n_3431),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_3467),
.Y(n_3473)
);

OAI322xp33_ASAP7_75t_SL g3474 ( 
.A1(n_3458),
.A2(n_3418),
.A3(n_3427),
.B1(n_3408),
.B2(n_3432),
.C1(n_3415),
.C2(n_3436),
.Y(n_3474)
);

NAND2xp5_ASAP7_75t_L g3475 ( 
.A(n_3447),
.B(n_493),
.Y(n_3475)
);

OAI22xp5_ASAP7_75t_L g3476 ( 
.A1(n_3464),
.A2(n_495),
.B1(n_493),
.B2(n_494),
.Y(n_3476)
);

INVx1_ASAP7_75t_SL g3477 ( 
.A(n_3460),
.Y(n_3477)
);

OAI211xp5_ASAP7_75t_SL g3478 ( 
.A1(n_3441),
.A2(n_498),
.B(n_496),
.C(n_497),
.Y(n_3478)
);

NAND3xp33_ASAP7_75t_L g3479 ( 
.A(n_3446),
.B(n_497),
.C(n_499),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_L g3480 ( 
.A(n_3455),
.B(n_499),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3465),
.Y(n_3481)
);

NOR2xp67_ASAP7_75t_L g3482 ( 
.A(n_3442),
.B(n_500),
.Y(n_3482)
);

AOI21xp33_ASAP7_75t_SL g3483 ( 
.A1(n_3449),
.A2(n_501),
.B(n_502),
.Y(n_3483)
);

AOI21xp5_ASAP7_75t_L g3484 ( 
.A1(n_3459),
.A2(n_502),
.B(n_503),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_L g3485 ( 
.A(n_3470),
.B(n_3466),
.Y(n_3485)
);

OAI22xp33_ASAP7_75t_L g3486 ( 
.A1(n_3481),
.A2(n_3451),
.B1(n_3457),
.B2(n_3453),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3473),
.Y(n_3487)
);

HB1xp67_ASAP7_75t_L g3488 ( 
.A(n_3482),
.Y(n_3488)
);

OA21x2_ASAP7_75t_L g3489 ( 
.A1(n_3469),
.A2(n_3445),
.B(n_3454),
.Y(n_3489)
);

OAI22xp5_ASAP7_75t_L g3490 ( 
.A1(n_3479),
.A2(n_3448),
.B1(n_3452),
.B2(n_3468),
.Y(n_3490)
);

OR2x2_ASAP7_75t_L g3491 ( 
.A(n_3475),
.B(n_3462),
.Y(n_3491)
);

AND2x4_ASAP7_75t_L g3492 ( 
.A(n_3477),
.B(n_3456),
.Y(n_3492)
);

AND2x4_ASAP7_75t_L g3493 ( 
.A(n_3480),
.B(n_3450),
.Y(n_3493)
);

INVx5_ASAP7_75t_L g3494 ( 
.A(n_3483),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_L g3495 ( 
.A(n_3476),
.B(n_3444),
.Y(n_3495)
);

BUFx2_ASAP7_75t_L g3496 ( 
.A(n_3488),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_3492),
.B(n_3484),
.Y(n_3497)
);

CKINVDCx20_ASAP7_75t_R g3498 ( 
.A(n_3489),
.Y(n_3498)
);

INVx1_ASAP7_75t_SL g3499 ( 
.A(n_3494),
.Y(n_3499)
);

AO22x2_ASAP7_75t_L g3500 ( 
.A1(n_3487),
.A2(n_3474),
.B1(n_3471),
.B2(n_3478),
.Y(n_3500)
);

CKINVDCx5p33_ASAP7_75t_R g3501 ( 
.A(n_3485),
.Y(n_3501)
);

INVx1_ASAP7_75t_L g3502 ( 
.A(n_3491),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_SL g3503 ( 
.A(n_3486),
.B(n_3463),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3493),
.Y(n_3504)
);

INVx1_ASAP7_75t_L g3505 ( 
.A(n_3496),
.Y(n_3505)
);

XNOR2x1_ASAP7_75t_L g3506 ( 
.A(n_3500),
.B(n_3490),
.Y(n_3506)
);

INVxp67_ASAP7_75t_SL g3507 ( 
.A(n_3497),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_3500),
.Y(n_3508)
);

INVxp33_ASAP7_75t_L g3509 ( 
.A(n_3506),
.Y(n_3509)
);

AND2x4_ASAP7_75t_L g3510 ( 
.A(n_3505),
.B(n_3504),
.Y(n_3510)
);

INVx1_ASAP7_75t_L g3511 ( 
.A(n_3508),
.Y(n_3511)
);

INVx2_ASAP7_75t_L g3512 ( 
.A(n_3510),
.Y(n_3512)
);

AND2x2_ASAP7_75t_L g3513 ( 
.A(n_3512),
.B(n_3499),
.Y(n_3513)
);

AOI22x1_ASAP7_75t_L g3514 ( 
.A1(n_3513),
.A2(n_3501),
.B1(n_3511),
.B2(n_3507),
.Y(n_3514)
);

OAI22xp5_ASAP7_75t_L g3515 ( 
.A1(n_3514),
.A2(n_3498),
.B1(n_3509),
.B2(n_3495),
.Y(n_3515)
);

AOI22xp5_ASAP7_75t_L g3516 ( 
.A1(n_3515),
.A2(n_3503),
.B1(n_3502),
.B2(n_3472),
.Y(n_3516)
);

AOI22xp5_ASAP7_75t_L g3517 ( 
.A1(n_3516),
.A2(n_507),
.B1(n_505),
.B2(n_506),
.Y(n_3517)
);

OA21x2_ASAP7_75t_L g3518 ( 
.A1(n_3517),
.A2(n_508),
.B(n_509),
.Y(n_3518)
);

AOI221xp5_ASAP7_75t_SL g3519 ( 
.A1(n_3518),
.A2(n_516),
.B1(n_510),
.B2(n_511),
.C(n_517),
.Y(n_3519)
);

AOI211xp5_ASAP7_75t_L g3520 ( 
.A1(n_3519),
.A2(n_520),
.B(n_517),
.C(n_519),
.Y(n_3520)
);


endmodule