module fake_netlist_1_10246_n_39 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_39);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_39;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
NAND2xp5_ASAP7_75t_L g11 ( .A(n_1), .B(n_3), .Y(n_11) );
AND2x4_ASAP7_75t_L g12 ( .A(n_0), .B(n_7), .Y(n_12) );
OAI22xp5_ASAP7_75t_SL g13 ( .A1(n_3), .A2(n_9), .B1(n_6), .B2(n_7), .Y(n_13) );
NAND2xp5_ASAP7_75t_SL g14 ( .A(n_6), .B(n_0), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
AND2x4_ASAP7_75t_L g16 ( .A(n_2), .B(n_5), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_15), .Y(n_17) );
AOI22xp33_ASAP7_75t_L g18 ( .A1(n_15), .A2(n_2), .B1(n_4), .B2(n_5), .Y(n_18) );
AND2x4_ASAP7_75t_L g19 ( .A(n_12), .B(n_4), .Y(n_19) );
BUFx6f_ASAP7_75t_L g20 ( .A(n_12), .Y(n_20) );
OAI21x1_ASAP7_75t_L g21 ( .A1(n_17), .A2(n_11), .B(n_14), .Y(n_21) );
AO21x2_ASAP7_75t_L g22 ( .A1(n_19), .A2(n_14), .B(n_12), .Y(n_22) );
OAI21x1_ASAP7_75t_L g23 ( .A1(n_17), .A2(n_8), .B(n_10), .Y(n_23) );
OR2x6_ASAP7_75t_L g24 ( .A(n_21), .B(n_13), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_22), .B(n_19), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
NAND2xp5_ASAP7_75t_SL g27 ( .A(n_25), .B(n_19), .Y(n_27) );
AOI22xp5_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_24), .B1(n_22), .B2(n_19), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_26), .Y(n_29) );
NOR2xp33_ASAP7_75t_L g30 ( .A(n_29), .B(n_24), .Y(n_30) );
AOI211xp5_ASAP7_75t_L g31 ( .A1(n_28), .A2(n_16), .B(n_27), .C(n_19), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_29), .Y(n_32) );
XNOR2x1_ASAP7_75t_L g33 ( .A(n_32), .B(n_24), .Y(n_33) );
NOR2x1_ASAP7_75t_L g34 ( .A(n_30), .B(n_16), .Y(n_34) );
OAI221xp5_ASAP7_75t_L g35 ( .A1(n_31), .A2(n_18), .B1(n_20), .B2(n_22), .C(n_21), .Y(n_35) );
OAI22xp5_ASAP7_75t_L g36 ( .A1(n_33), .A2(n_20), .B1(n_23), .B2(n_34), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_35), .Y(n_37) );
OAI22xp5_ASAP7_75t_SL g38 ( .A1(n_36), .A2(n_20), .B1(n_23), .B2(n_37), .Y(n_38) );
AOI22xp33_ASAP7_75t_L g39 ( .A1(n_38), .A2(n_20), .B1(n_37), .B2(n_36), .Y(n_39) );
endmodule