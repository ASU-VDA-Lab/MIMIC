module fake_jpeg_21978_n_78 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_78);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_78;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_13),
.B(n_32),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_31),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_28),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_47),
.Y(n_52)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_0),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_50),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_46),
.A2(n_36),
.B1(n_42),
.B2(n_33),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_49),
.A2(n_54),
.B1(n_0),
.B2(n_1),
.Y(n_56)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_51),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_39),
.B1(n_38),
.B2(n_37),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_52),
.A2(n_35),
.B(n_34),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_2),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_57),
.B(n_52),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_59),
.B(n_60),
.Y(n_68)
);

NOR2x1_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_49),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_55),
.B(n_1),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_61),
.A2(n_62),
.B(n_63),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_2),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_63),
.A2(n_53),
.B1(n_7),
.B2(n_8),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_3),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_65),
.A2(n_4),
.B(n_9),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_66),
.B(n_67),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_68),
.C(n_12),
.Y(n_71)
);

OAI321xp33_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_69),
.A3(n_14),
.B1(n_15),
.B2(n_16),
.C(n_17),
.Y(n_72)
);

NOR3xp33_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_10),
.C(n_19),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_20),
.C(n_22),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_23),
.C(n_24),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_30),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_26),
.Y(n_78)
);


endmodule