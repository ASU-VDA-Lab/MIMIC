module fake_netlist_6_2086_n_1067 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1067);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1067;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_367;
wire n_465;
wire n_680;
wire n_760;
wire n_741;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_222;
wire n_300;
wire n_248;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_989;
wire n_843;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_886;
wire n_448;
wire n_844;
wire n_953;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_947;
wire n_381;
wire n_911;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_964;
wire n_802;
wire n_982;
wire n_831;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_1055;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1063;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_127),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_190),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_120),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_46),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_209),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_146),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_92),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_114),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_134),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_16),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_69),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_136),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_150),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_30),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_111),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_147),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_152),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_144),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_151),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_174),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_19),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_96),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_198),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_186),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_80),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_7),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_195),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_43),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_132),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_176),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_53),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_101),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_8),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_107),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_157),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_52),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_197),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_47),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_48),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_29),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_166),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_131),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_24),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_70),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_148),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_84),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_105),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_189),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_182),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_141),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_155),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_37),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_63),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_109),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_59),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_170),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_99),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_102),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_17),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_104),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_26),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_72),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_126),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_129),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_158),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_61),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_192),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_173),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_219),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_268),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_211),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_274),
.Y(n_281)
);

BUFx10_ASAP7_75t_L g282 ( 
.A(n_237),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_230),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_235),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_242),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_244),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_212),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_217),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_262),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_213),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_214),
.Y(n_292)
);

INVxp67_ASAP7_75t_SL g293 ( 
.A(n_225),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_218),
.Y(n_294)
);

INVxp67_ASAP7_75t_SL g295 ( 
.A(n_275),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_244),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_220),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_262),
.B(n_0),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_221),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_227),
.Y(n_300)
);

INVxp33_ASAP7_75t_SL g301 ( 
.A(n_252),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_258),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_228),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g304 ( 
.A(n_270),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_223),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_224),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_226),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_229),
.Y(n_308)
);

INVxp67_ASAP7_75t_SL g309 ( 
.A(n_262),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_246),
.Y(n_310)
);

INVxp33_ASAP7_75t_SL g311 ( 
.A(n_210),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_231),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_247),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_258),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_232),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_260),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_233),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_264),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_266),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_272),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_271),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_273),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_222),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_234),
.Y(n_324)
);

INVxp33_ASAP7_75t_SL g325 ( 
.A(n_210),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_222),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_272),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_290),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_290),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_291),
.Y(n_330)
);

BUFx8_ASAP7_75t_L g331 ( 
.A(n_320),
.Y(n_331)
);

AND2x4_ASAP7_75t_L g332 ( 
.A(n_309),
.B(n_251),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_316),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_293),
.A2(n_241),
.B1(n_253),
.B2(n_215),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_280),
.B(n_251),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_316),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_290),
.Y(n_337)
);

INVxp33_ASAP7_75t_SL g338 ( 
.A(n_288),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_290),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_278),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_323),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_279),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_326),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_292),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_294),
.Y(n_345)
);

INVx5_ASAP7_75t_L g346 ( 
.A(n_282),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_289),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_295),
.A2(n_215),
.B1(n_276),
.B2(n_216),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_297),
.Y(n_349)
);

AND2x4_ASAP7_75t_L g350 ( 
.A(n_284),
.B(n_257),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_299),
.Y(n_351)
);

INVx2_ASAP7_75t_SL g352 ( 
.A(n_282),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_305),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_301),
.A2(n_216),
.B1(n_276),
.B2(n_277),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_311),
.B(n_257),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_306),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_311),
.B(n_277),
.Y(n_357)
);

AND2x6_ASAP7_75t_L g358 ( 
.A(n_298),
.B(n_27),
.Y(n_358)
);

CKINVDCx6p67_ASAP7_75t_R g359 ( 
.A(n_286),
.Y(n_359)
);

INVx5_ASAP7_75t_L g360 ( 
.A(n_282),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_307),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_283),
.B(n_236),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_308),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_310),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_313),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_318),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_319),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_281),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_321),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_300),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_301),
.A2(n_254),
.B1(n_267),
.B2(n_265),
.Y(n_371)
);

OA21x2_ASAP7_75t_L g372 ( 
.A1(n_322),
.A2(n_239),
.B(n_238),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_287),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_303),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_312),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_304),
.Y(n_376)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_285),
.B(n_315),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_317),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_324),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_325),
.B(n_240),
.Y(n_380)
);

AND2x4_ASAP7_75t_L g381 ( 
.A(n_325),
.B(n_243),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_330),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_359),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_331),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_329),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_375),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_329),
.Y(n_387)
);

BUFx10_ASAP7_75t_L g388 ( 
.A(n_377),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_328),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_344),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_337),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_331),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_375),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_333),
.Y(n_394)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_333),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_338),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_377),
.A2(n_261),
.B1(n_248),
.B2(n_249),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_334),
.A2(n_327),
.B1(n_314),
.B2(n_302),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_353),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_364),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_365),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_347),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_338),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_R g404 ( 
.A(n_374),
.B(n_286),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_370),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_369),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_378),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_378),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_378),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_378),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_337),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_339),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_336),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_328),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_374),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_379),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_380),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_339),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_336),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_376),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_346),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_346),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_346),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_346),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_362),
.Y(n_425)
);

BUFx10_ASAP7_75t_L g426 ( 
.A(n_352),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_360),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_373),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_360),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_376),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_360),
.Y(n_431)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_328),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_360),
.B(n_296),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_R g434 ( 
.A(n_355),
.B(n_296),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_335),
.B(n_245),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_362),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_371),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_348),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_328),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_351),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_332),
.B(n_250),
.Y(n_441)
);

NAND2xp33_ASAP7_75t_R g442 ( 
.A(n_372),
.B(n_0),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_356),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_368),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_R g445 ( 
.A(n_355),
.B(n_302),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_354),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_368),
.Y(n_447)
);

NOR2xp67_ASAP7_75t_L g448 ( 
.A(n_381),
.B(n_357),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_R g449 ( 
.A(n_357),
.B(n_314),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_332),
.B(n_255),
.Y(n_450)
);

NAND3xp33_ASAP7_75t_L g451 ( 
.A(n_442),
.B(n_372),
.C(n_350),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_420),
.B(n_350),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_430),
.B(n_381),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_382),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_390),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_399),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_435),
.B(n_446),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_391),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_448),
.B(n_381),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_400),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_416),
.B(n_327),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_401),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_391),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_419),
.B(n_345),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_441),
.B(n_372),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_406),
.Y(n_466)
);

NAND3xp33_ASAP7_75t_L g467 ( 
.A(n_442),
.B(n_450),
.C(n_428),
.Y(n_467)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_407),
.Y(n_468)
);

AND2x2_ASAP7_75t_SL g469 ( 
.A(n_433),
.B(n_345),
.Y(n_469)
);

OR2x2_ASAP7_75t_L g470 ( 
.A(n_394),
.B(n_349),
.Y(n_470)
);

AND3x1_ASAP7_75t_L g471 ( 
.A(n_397),
.B(n_361),
.C(n_349),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_438),
.B(n_356),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_411),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_411),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_408),
.B(n_410),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_415),
.B(n_356),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_418),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_395),
.B(n_361),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_444),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_447),
.B(n_363),
.Y(n_480)
);

OR2x6_ASAP7_75t_L g481 ( 
.A(n_398),
.B(n_366),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_385),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_386),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_387),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_440),
.B(n_358),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_412),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_389),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_437),
.B(n_363),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_393),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_419),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_396),
.Y(n_491)
);

AND2x6_ASAP7_75t_L g492 ( 
.A(n_443),
.B(n_358),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_388),
.B(n_366),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_413),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_426),
.B(n_363),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_439),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_389),
.Y(n_497)
);

INVx1_ASAP7_75t_SL g498 ( 
.A(n_404),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_389),
.Y(n_499)
);

NAND2x1p5_ASAP7_75t_L g500 ( 
.A(n_432),
.B(n_414),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_414),
.B(n_432),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_404),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_426),
.B(n_363),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_414),
.Y(n_504)
);

NAND3xp33_ASAP7_75t_SL g505 ( 
.A(n_434),
.B(n_259),
.C(n_256),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_388),
.B(n_367),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_421),
.B(n_340),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_422),
.B(n_343),
.Y(n_508)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_423),
.Y(n_509)
);

INVx8_ASAP7_75t_L g510 ( 
.A(n_409),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_403),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_424),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_405),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_434),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_427),
.B(n_367),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_429),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_425),
.B(n_340),
.Y(n_517)
);

INVx4_ASAP7_75t_L g518 ( 
.A(n_431),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_436),
.B(n_343),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_417),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_402),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_383),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g523 ( 
.A(n_384),
.B(n_263),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_449),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_445),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_449),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_445),
.B(n_340),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_392),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_451),
.A2(n_342),
.B1(n_340),
.B2(n_343),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_474),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_517),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_477),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_463),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_487),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_457),
.A2(n_269),
.B1(n_343),
.B2(n_342),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_454),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_463),
.Y(n_537)
);

OAI221xp5_ASAP7_75t_L g538 ( 
.A1(n_467),
.A2(n_342),
.B1(n_341),
.B2(n_3),
.C(n_4),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_459),
.A2(n_471),
.B1(n_467),
.B2(n_453),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_455),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_456),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g542 ( 
.A(n_472),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_460),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_462),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_458),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_466),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_471),
.A2(n_342),
.B1(n_341),
.B2(n_97),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_519),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_484),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_488),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_486),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g552 ( 
.A(n_470),
.Y(n_552)
);

AO22x2_ASAP7_75t_L g553 ( 
.A1(n_451),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_473),
.Y(n_554)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_452),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_461),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_482),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_464),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_480),
.B(n_5),
.Y(n_559)
);

NAND3xp33_ASAP7_75t_L g560 ( 
.A(n_479),
.B(n_5),
.C(n_6),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_490),
.B(n_464),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_490),
.B(n_28),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_482),
.Y(n_563)
);

NAND2xp33_ASAP7_75t_L g564 ( 
.A(n_524),
.B(n_31),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_510),
.Y(n_565)
);

INVx4_ASAP7_75t_SL g566 ( 
.A(n_524),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_504),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_496),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_478),
.Y(n_569)
);

INVx2_ASAP7_75t_SL g570 ( 
.A(n_510),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_499),
.Y(n_571)
);

O2A1O1Ixp33_ASAP7_75t_L g572 ( 
.A1(n_465),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_493),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_527),
.B(n_9),
.Y(n_574)
);

NAND2x1p5_ASAP7_75t_L g575 ( 
.A(n_468),
.B(n_32),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_475),
.B(n_468),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_490),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_494),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_506),
.B(n_9),
.Y(n_579)
);

INVxp67_ASAP7_75t_L g580 ( 
.A(n_521),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_514),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_509),
.B(n_33),
.Y(n_582)
);

NAND3xp33_ASAP7_75t_L g583 ( 
.A(n_526),
.B(n_10),
.C(n_11),
.Y(n_583)
);

OR2x2_ASAP7_75t_L g584 ( 
.A(n_498),
.B(n_10),
.Y(n_584)
);

INVx2_ASAP7_75t_SL g585 ( 
.A(n_510),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_497),
.Y(n_586)
);

INVxp67_ASAP7_75t_L g587 ( 
.A(n_502),
.Y(n_587)
);

AND2x2_ASAP7_75t_SL g588 ( 
.A(n_565),
.B(n_524),
.Y(n_588)
);

NAND3xp33_ASAP7_75t_L g589 ( 
.A(n_542),
.B(n_513),
.C(n_550),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_531),
.B(n_525),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_548),
.B(n_498),
.Y(n_591)
);

OAI21xp33_ASAP7_75t_L g592 ( 
.A1(n_573),
.A2(n_523),
.B(n_489),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_569),
.B(n_536),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_552),
.B(n_483),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_540),
.B(n_469),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_541),
.B(n_515),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_543),
.B(n_515),
.Y(n_597)
);

O2A1O1Ixp33_ASAP7_75t_L g598 ( 
.A1(n_579),
.A2(n_505),
.B(n_481),
.C(n_476),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_530),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_544),
.B(n_546),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_555),
.B(n_491),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_539),
.B(n_495),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_553),
.A2(n_481),
.B1(n_492),
.B2(n_485),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_532),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_561),
.B(n_508),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_578),
.B(n_511),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_L g607 ( 
.A1(n_547),
.A2(n_492),
.B(n_501),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_561),
.B(n_520),
.Y(n_608)
);

A2O1A1Ixp33_ASAP7_75t_L g609 ( 
.A1(n_576),
.A2(n_516),
.B(n_507),
.C(n_503),
.Y(n_609)
);

A2O1A1Ixp33_ASAP7_75t_L g610 ( 
.A1(n_574),
.A2(n_523),
.B(n_522),
.C(n_520),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_549),
.B(n_509),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_551),
.B(n_512),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_566),
.B(n_512),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_558),
.B(n_532),
.Y(n_614)
);

BUFx12f_ASAP7_75t_L g615 ( 
.A(n_570),
.Y(n_615)
);

AO21x1_ASAP7_75t_L g616 ( 
.A1(n_559),
.A2(n_572),
.B(n_564),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_581),
.B(n_587),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_L g618 ( 
.A1(n_553),
.A2(n_520),
.B1(n_518),
.B2(n_497),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_577),
.B(n_518),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_545),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_538),
.A2(n_492),
.B1(n_497),
.B2(n_500),
.Y(n_621)
);

AND2x4_ASAP7_75t_L g622 ( 
.A(n_566),
.B(n_528),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_529),
.A2(n_35),
.B(n_34),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_577),
.B(n_528),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_577),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_545),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_582),
.B(n_528),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_585),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_554),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_586),
.A2(n_38),
.B(n_36),
.Y(n_630)
);

O2A1O1Ixp33_ASAP7_75t_L g631 ( 
.A1(n_584),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_L g632 ( 
.A1(n_571),
.A2(n_208),
.B(n_40),
.Y(n_632)
);

O2A1O1Ixp33_ASAP7_75t_L g633 ( 
.A1(n_568),
.A2(n_583),
.B(n_580),
.C(n_560),
.Y(n_633)
);

BUFx12f_ASAP7_75t_L g634 ( 
.A(n_582),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_557),
.B(n_12),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_562),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_563),
.B(n_13),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_562),
.B(n_535),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_586),
.A2(n_115),
.B(n_206),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_533),
.B(n_537),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_534),
.B(n_567),
.Y(n_641)
);

A2O1A1Ixp33_ASAP7_75t_L g642 ( 
.A1(n_598),
.A2(n_567),
.B(n_534),
.C(n_556),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_596),
.B(n_575),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_625),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_594),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_645)
);

O2A1O1Ixp33_ASAP7_75t_L g646 ( 
.A1(n_610),
.A2(n_14),
.B(n_15),
.C(n_17),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_599),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_591),
.B(n_590),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_626),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_622),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_638),
.A2(n_117),
.B(n_205),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_604),
.Y(n_652)
);

O2A1O1Ixp33_ASAP7_75t_L g653 ( 
.A1(n_631),
.A2(n_18),
.B(n_19),
.C(n_20),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_597),
.B(n_18),
.Y(n_654)
);

AOI22x1_ASAP7_75t_L g655 ( 
.A1(n_623),
.A2(n_118),
.B1(n_204),
.B2(n_203),
.Y(n_655)
);

INVxp67_ASAP7_75t_SL g656 ( 
.A(n_636),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_636),
.B(n_39),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_607),
.A2(n_116),
.B(n_202),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_620),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_622),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_589),
.B(n_20),
.Y(n_661)
);

NOR2x1_ASAP7_75t_L g662 ( 
.A(n_602),
.B(n_41),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_600),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_593),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_629),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_614),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_636),
.B(n_21),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_606),
.B(n_21),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_588),
.B(n_22),
.Y(n_669)
);

NOR3xp33_ASAP7_75t_L g670 ( 
.A(n_592),
.B(n_22),
.C(n_23),
.Y(n_670)
);

INVx3_ASAP7_75t_SL g671 ( 
.A(n_628),
.Y(n_671)
);

INVxp67_ASAP7_75t_L g672 ( 
.A(n_617),
.Y(n_672)
);

BUFx2_ASAP7_75t_L g673 ( 
.A(n_601),
.Y(n_673)
);

O2A1O1Ixp33_ASAP7_75t_L g674 ( 
.A1(n_609),
.A2(n_23),
.B(n_24),
.C(n_25),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_640),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_605),
.B(n_595),
.Y(n_676)
);

O2A1O1Ixp33_ASAP7_75t_L g677 ( 
.A1(n_633),
.A2(n_25),
.B(n_26),
.C(n_42),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_611),
.B(n_44),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_612),
.B(n_608),
.Y(n_679)
);

OAI22xp5_ASAP7_75t_L g680 ( 
.A1(n_603),
.A2(n_45),
.B1(n_49),
.B2(n_50),
.Y(n_680)
);

AND2x4_ASAP7_75t_L g681 ( 
.A(n_613),
.B(n_51),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_627),
.B(n_54),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_635),
.B(n_613),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_634),
.B(n_55),
.Y(n_684)
);

NAND2x1p5_ASAP7_75t_L g685 ( 
.A(n_625),
.B(n_56),
.Y(n_685)
);

NOR2xp67_ASAP7_75t_SL g686 ( 
.A(n_615),
.B(n_57),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_641),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_618),
.A2(n_58),
.B1(n_60),
.B2(n_62),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_618),
.B(n_64),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_637),
.B(n_65),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_625),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_624),
.B(n_66),
.Y(n_692)
);

AND2x4_ASAP7_75t_L g693 ( 
.A(n_619),
.B(n_207),
.Y(n_693)
);

AND2x4_ASAP7_75t_SL g694 ( 
.A(n_621),
.B(n_616),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_632),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_632),
.A2(n_67),
.B1(n_68),
.B2(n_71),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_630),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_671),
.Y(n_698)
);

BUFx3_ASAP7_75t_L g699 ( 
.A(n_650),
.Y(n_699)
);

INVx8_ASAP7_75t_L g700 ( 
.A(n_644),
.Y(n_700)
);

INVx1_ASAP7_75t_SL g701 ( 
.A(n_673),
.Y(n_701)
);

INVx5_ASAP7_75t_L g702 ( 
.A(n_644),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_647),
.Y(n_703)
);

HB1xp67_ASAP7_75t_L g704 ( 
.A(n_652),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_665),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_670),
.A2(n_639),
.B1(n_74),
.B2(n_75),
.Y(n_706)
);

BUFx4_ASAP7_75t_SL g707 ( 
.A(n_660),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_659),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_644),
.Y(n_709)
);

BUFx2_ASAP7_75t_SL g710 ( 
.A(n_691),
.Y(n_710)
);

BUFx12f_ASAP7_75t_L g711 ( 
.A(n_691),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_691),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_672),
.B(n_73),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_681),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_681),
.Y(n_715)
);

BUFx3_ASAP7_75t_L g716 ( 
.A(n_657),
.Y(n_716)
);

CKINVDCx6p67_ASAP7_75t_R g717 ( 
.A(n_683),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_649),
.Y(n_718)
);

BUFx2_ASAP7_75t_SL g719 ( 
.A(n_656),
.Y(n_719)
);

INVxp67_ASAP7_75t_SL g720 ( 
.A(n_666),
.Y(n_720)
);

BUFx12f_ASAP7_75t_L g721 ( 
.A(n_657),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_675),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_667),
.Y(n_723)
);

BUFx12f_ASAP7_75t_L g724 ( 
.A(n_693),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_663),
.Y(n_725)
);

CKINVDCx11_ASAP7_75t_R g726 ( 
.A(n_693),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_687),
.Y(n_727)
);

INVx4_ASAP7_75t_L g728 ( 
.A(n_685),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_661),
.Y(n_729)
);

INVx4_ASAP7_75t_L g730 ( 
.A(n_682),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_664),
.Y(n_731)
);

INVx4_ASAP7_75t_L g732 ( 
.A(n_694),
.Y(n_732)
);

HB1xp67_ASAP7_75t_L g733 ( 
.A(n_695),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_SL g734 ( 
.A1(n_689),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_734)
);

BUFx12f_ASAP7_75t_L g735 ( 
.A(n_686),
.Y(n_735)
);

INVx4_ASAP7_75t_L g736 ( 
.A(n_697),
.Y(n_736)
);

INVxp67_ASAP7_75t_SL g737 ( 
.A(n_676),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_654),
.Y(n_738)
);

AND2x4_ASAP7_75t_L g739 ( 
.A(n_642),
.B(n_79),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_648),
.B(n_81),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_679),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_669),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_643),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_646),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_668),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_696),
.A2(n_82),
.B1(n_83),
.B2(n_85),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_684),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_655),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_674),
.Y(n_749)
);

BUFx6f_ASAP7_75t_SL g750 ( 
.A(n_688),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_692),
.Y(n_751)
);

BUFx2_ASAP7_75t_SL g752 ( 
.A(n_688),
.Y(n_752)
);

INVx3_ASAP7_75t_SL g753 ( 
.A(n_678),
.Y(n_753)
);

BUFx8_ASAP7_75t_L g754 ( 
.A(n_645),
.Y(n_754)
);

INVx8_ASAP7_75t_L g755 ( 
.A(n_651),
.Y(n_755)
);

INVx8_ASAP7_75t_L g756 ( 
.A(n_662),
.Y(n_756)
);

NAND2x1p5_ASAP7_75t_L g757 ( 
.A(n_662),
.B(n_86),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_690),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_696),
.Y(n_759)
);

BUFx12f_ASAP7_75t_L g760 ( 
.A(n_677),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_653),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_704),
.Y(n_762)
);

INVx1_ASAP7_75t_SL g763 ( 
.A(n_701),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_729),
.B(n_680),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_704),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_703),
.Y(n_766)
);

INVx3_ASAP7_75t_L g767 ( 
.A(n_731),
.Y(n_767)
);

NOR2x1_ASAP7_75t_R g768 ( 
.A(n_698),
.B(n_658),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_708),
.Y(n_769)
);

INVxp67_ASAP7_75t_SL g770 ( 
.A(n_720),
.Y(n_770)
);

OR2x2_ASAP7_75t_L g771 ( 
.A(n_701),
.B(n_87),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_698),
.Y(n_772)
);

OAI21x1_ASAP7_75t_L g773 ( 
.A1(n_748),
.A2(n_88),
.B(n_89),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_709),
.Y(n_774)
);

OAI222xp33_ASAP7_75t_L g775 ( 
.A1(n_759),
.A2(n_729),
.B1(n_746),
.B2(n_706),
.C1(n_749),
.C2(n_739),
.Y(n_775)
);

AO32x2_ASAP7_75t_L g776 ( 
.A1(n_736),
.A2(n_90),
.A3(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_776)
);

INVx2_ASAP7_75t_SL g777 ( 
.A(n_707),
.Y(n_777)
);

OA21x2_ASAP7_75t_L g778 ( 
.A1(n_748),
.A2(n_95),
.B(n_98),
.Y(n_778)
);

OAI21x1_ASAP7_75t_L g779 ( 
.A1(n_757),
.A2(n_100),
.B(n_103),
.Y(n_779)
);

AOI22x1_ASAP7_75t_L g780 ( 
.A1(n_760),
.A2(n_106),
.B1(n_108),
.B2(n_110),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_711),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_759),
.A2(n_112),
.B1(n_113),
.B2(n_119),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_750),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_723),
.B(n_124),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_720),
.Y(n_785)
);

OA21x2_ASAP7_75t_L g786 ( 
.A1(n_744),
.A2(n_125),
.B(n_128),
.Y(n_786)
);

INVx5_ASAP7_75t_L g787 ( 
.A(n_756),
.Y(n_787)
);

OR2x2_ASAP7_75t_L g788 ( 
.A(n_737),
.B(n_130),
.Y(n_788)
);

BUFx2_ASAP7_75t_SL g789 ( 
.A(n_699),
.Y(n_789)
);

OAI21x1_ASAP7_75t_L g790 ( 
.A1(n_757),
.A2(n_133),
.B(n_135),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_727),
.Y(n_791)
);

INVx6_ASAP7_75t_L g792 ( 
.A(n_702),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_727),
.Y(n_793)
);

XNOR2xp5_ASAP7_75t_L g794 ( 
.A(n_747),
.B(n_201),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_718),
.Y(n_795)
);

OAI21x1_ASAP7_75t_L g796 ( 
.A1(n_743),
.A2(n_137),
.B(n_138),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_L g797 ( 
.A1(n_750),
.A2(n_139),
.B1(n_140),
.B2(n_142),
.Y(n_797)
);

OAI21x1_ASAP7_75t_SL g798 ( 
.A1(n_732),
.A2(n_143),
.B(n_145),
.Y(n_798)
);

OA21x2_ASAP7_75t_L g799 ( 
.A1(n_706),
.A2(n_737),
.B(n_733),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_717),
.B(n_149),
.Y(n_800)
);

CKINVDCx20_ASAP7_75t_R g801 ( 
.A(n_726),
.Y(n_801)
);

BUFx2_ASAP7_75t_L g802 ( 
.A(n_699),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_742),
.B(n_153),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_754),
.A2(n_200),
.B1(n_156),
.B2(n_159),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_752),
.A2(n_154),
.B1(n_160),
.B2(n_161),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_705),
.Y(n_806)
);

OAI21x1_ASAP7_75t_L g807 ( 
.A1(n_733),
.A2(n_162),
.B(n_163),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_707),
.Y(n_808)
);

OAI21x1_ASAP7_75t_SL g809 ( 
.A1(n_732),
.A2(n_164),
.B(n_165),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_725),
.Y(n_810)
);

OA21x2_ASAP7_75t_L g811 ( 
.A1(n_738),
.A2(n_167),
.B(n_168),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_741),
.B(n_169),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_700),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_722),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_741),
.B(n_171),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_700),
.Y(n_816)
);

INVx8_ASAP7_75t_L g817 ( 
.A(n_700),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_763),
.B(n_810),
.Y(n_818)
);

OR2x2_ASAP7_75t_L g819 ( 
.A(n_762),
.B(n_731),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_791),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_766),
.B(n_739),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_769),
.B(n_758),
.Y(n_822)
);

INVxp67_ASAP7_75t_L g823 ( 
.A(n_763),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_765),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_793),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_770),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_764),
.A2(n_754),
.B1(n_761),
.B2(n_742),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_770),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_806),
.B(n_742),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_785),
.Y(n_830)
);

OAI21x1_ASAP7_75t_L g831 ( 
.A1(n_773),
.A2(n_740),
.B(n_755),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_795),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_802),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_814),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_767),
.Y(n_835)
);

AOI21x1_ASAP7_75t_L g836 ( 
.A1(n_786),
.A2(n_713),
.B(n_756),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_767),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_787),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_799),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_799),
.Y(n_840)
);

INVx4_ASAP7_75t_SL g841 ( 
.A(n_792),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_776),
.Y(n_842)
);

OAI21x1_ASAP7_75t_SL g843 ( 
.A1(n_798),
.A2(n_736),
.B(n_730),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_776),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_788),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_776),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_778),
.Y(n_847)
);

OAI21x1_ASAP7_75t_L g848 ( 
.A1(n_796),
.A2(n_755),
.B(n_756),
.Y(n_848)
);

INVxp67_ASAP7_75t_SL g849 ( 
.A(n_768),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_812),
.Y(n_850)
);

CKINVDCx20_ASAP7_75t_R g851 ( 
.A(n_801),
.Y(n_851)
);

BUFx4f_ASAP7_75t_SL g852 ( 
.A(n_801),
.Y(n_852)
);

NAND2x1_ASAP7_75t_L g853 ( 
.A(n_786),
.B(n_728),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_811),
.Y(n_854)
);

BUFx2_ASAP7_75t_R g855 ( 
.A(n_772),
.Y(n_855)
);

OR2x6_ASAP7_75t_L g856 ( 
.A(n_789),
.B(n_755),
.Y(n_856)
);

OR2x2_ASAP7_75t_L g857 ( 
.A(n_771),
.B(n_747),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_812),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_811),
.B(n_730),
.Y(n_859)
);

NAND2x1p5_ASAP7_75t_L g860 ( 
.A(n_853),
.B(n_787),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_851),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_SL g862 ( 
.A1(n_827),
.A2(n_775),
.B(n_764),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_830),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_830),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_819),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_835),
.Y(n_866)
);

OR2x6_ASAP7_75t_L g867 ( 
.A(n_856),
.B(n_792),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_835),
.Y(n_868)
);

NAND2xp33_ASAP7_75t_SL g869 ( 
.A(n_851),
.B(n_772),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_852),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_820),
.Y(n_871)
);

A2O1A1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_849),
.A2(n_783),
.B(n_804),
.C(n_803),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_820),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_837),
.B(n_787),
.Y(n_874)
);

INVx4_ASAP7_75t_L g875 ( 
.A(n_841),
.Y(n_875)
);

OR2x2_ASAP7_75t_L g876 ( 
.A(n_826),
.B(n_777),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_825),
.Y(n_877)
);

A2O1A1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_842),
.A2(n_783),
.B(n_804),
.C(n_803),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_825),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_855),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_824),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_828),
.Y(n_882)
);

INVx8_ASAP7_75t_L g883 ( 
.A(n_856),
.Y(n_883)
);

NAND2xp33_ASAP7_75t_R g884 ( 
.A(n_857),
.B(n_800),
.Y(n_884)
);

NOR2x1_ASAP7_75t_SL g885 ( 
.A(n_856),
.B(n_787),
.Y(n_885)
);

INVx2_ASAP7_75t_SL g886 ( 
.A(n_822),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_819),
.Y(n_887)
);

INVxp33_ASAP7_75t_L g888 ( 
.A(n_857),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_833),
.B(n_808),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_850),
.A2(n_775),
.B(n_797),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_823),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_818),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_822),
.B(n_781),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_838),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_858),
.B(n_761),
.Y(n_895)
);

OR2x2_ASAP7_75t_L g896 ( 
.A(n_865),
.B(n_839),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_894),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_863),
.Y(n_898)
);

INVx4_ASAP7_75t_L g899 ( 
.A(n_875),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_887),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_864),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_871),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_892),
.B(n_845),
.Y(n_903)
);

NAND4xp25_ASAP7_75t_L g904 ( 
.A(n_890),
.B(n_829),
.C(n_840),
.D(n_821),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_888),
.B(n_834),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_861),
.B(n_745),
.Y(n_906)
);

AND2x4_ASAP7_75t_SL g907 ( 
.A(n_875),
.B(n_856),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_886),
.B(n_866),
.Y(n_908)
);

INVxp67_ASAP7_75t_SL g909 ( 
.A(n_866),
.Y(n_909)
);

AOI211xp5_ASAP7_75t_L g910 ( 
.A1(n_862),
.A2(n_782),
.B(n_794),
.C(n_805),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_877),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_879),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_870),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_873),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_868),
.B(n_894),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_874),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_891),
.B(n_745),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_885),
.B(n_859),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_881),
.Y(n_919)
);

AO21x2_ASAP7_75t_L g920 ( 
.A1(n_918),
.A2(n_847),
.B(n_854),
.Y(n_920)
);

OAI22xp33_ASAP7_75t_L g921 ( 
.A1(n_904),
.A2(n_862),
.B1(n_884),
.B2(n_844),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_897),
.Y(n_922)
);

OAI221xp5_ASAP7_75t_L g923 ( 
.A1(n_910),
.A2(n_872),
.B1(n_878),
.B2(n_869),
.C(n_895),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_916),
.B(n_893),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_913),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_913),
.Y(n_926)
);

AOI211xp5_ASAP7_75t_L g927 ( 
.A1(n_918),
.A2(n_761),
.B(n_876),
.C(n_889),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_917),
.A2(n_842),
.B(n_844),
.C(n_846),
.Y(n_928)
);

BUFx2_ASAP7_75t_L g929 ( 
.A(n_899),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_898),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_903),
.B(n_880),
.Y(n_931)
);

OR2x6_ASAP7_75t_L g932 ( 
.A(n_899),
.B(n_883),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_916),
.B(n_874),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_896),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_933),
.B(n_916),
.Y(n_935)
);

OR2x2_ASAP7_75t_L g936 ( 
.A(n_934),
.B(n_900),
.Y(n_936)
);

OR2x2_ASAP7_75t_L g937 ( 
.A(n_934),
.B(n_905),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_930),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_929),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_924),
.B(n_918),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_932),
.B(n_908),
.Y(n_941)
);

BUFx2_ASAP7_75t_L g942 ( 
.A(n_932),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_920),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_926),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_920),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_939),
.B(n_921),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_944),
.Y(n_947)
);

INVx5_ASAP7_75t_SL g948 ( 
.A(n_944),
.Y(n_948)
);

OR2x2_ASAP7_75t_L g949 ( 
.A(n_936),
.B(n_937),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_938),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_941),
.B(n_932),
.Y(n_951)
);

OR2x2_ASAP7_75t_L g952 ( 
.A(n_942),
.B(n_921),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_944),
.B(n_927),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_951),
.B(n_944),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_950),
.Y(n_955)
);

INVxp67_ASAP7_75t_L g956 ( 
.A(n_952),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_948),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_948),
.Y(n_958)
);

OR2x2_ASAP7_75t_L g959 ( 
.A(n_949),
.B(n_946),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_947),
.B(n_935),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_956),
.B(n_953),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_954),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_955),
.Y(n_963)
);

OAI31xp33_ASAP7_75t_L g964 ( 
.A1(n_959),
.A2(n_923),
.A3(n_945),
.B(n_928),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_957),
.A2(n_935),
.B1(n_926),
.B2(n_925),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_958),
.B(n_926),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_954),
.Y(n_967)
);

OR2x6_ASAP7_75t_L g968 ( 
.A(n_960),
.B(n_926),
.Y(n_968)
);

AOI22xp5_ASAP7_75t_L g969 ( 
.A1(n_960),
.A2(n_925),
.B1(n_940),
.B2(n_931),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_954),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_957),
.B(n_931),
.Y(n_971)
);

OR2x2_ASAP7_75t_L g972 ( 
.A(n_961),
.B(n_945),
.Y(n_972)
);

NOR2x1_ASAP7_75t_L g973 ( 
.A(n_970),
.B(n_943),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_963),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_962),
.B(n_922),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_968),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_967),
.Y(n_977)
);

OR2x2_ASAP7_75t_L g978 ( 
.A(n_966),
.B(n_943),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_968),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_977),
.Y(n_980)
);

INVxp67_ASAP7_75t_L g981 ( 
.A(n_979),
.Y(n_981)
);

XOR2x2_ASAP7_75t_L g982 ( 
.A(n_975),
.B(n_971),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_973),
.A2(n_964),
.B(n_965),
.Y(n_983)
);

OR2x2_ASAP7_75t_L g984 ( 
.A(n_976),
.B(n_969),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_972),
.A2(n_906),
.B(n_928),
.Y(n_985)
);

INVxp67_ASAP7_75t_L g986 ( 
.A(n_978),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_981),
.B(n_974),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_980),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_983),
.B(n_919),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_984),
.B(n_899),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_986),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_991),
.B(n_982),
.Y(n_992)
);

INVx1_ASAP7_75t_SL g993 ( 
.A(n_987),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_988),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_989),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_990),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_991),
.Y(n_997)
);

O2A1O1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_992),
.A2(n_985),
.B(n_809),
.C(n_784),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_993),
.A2(n_780),
.B(n_745),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_997),
.B(n_898),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_994),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_996),
.B(n_908),
.Y(n_1002)
);

NOR5xp2_ASAP7_75t_L g1003 ( 
.A(n_995),
.B(n_909),
.C(n_901),
.D(n_914),
.E(n_735),
.Y(n_1003)
);

OAI322xp33_ASAP7_75t_L g1004 ( 
.A1(n_1001),
.A2(n_896),
.A3(n_897),
.B1(n_860),
.B2(n_901),
.C1(n_853),
.C2(n_914),
.Y(n_1004)
);

OAI21xp33_ASAP7_75t_L g1005 ( 
.A1(n_1002),
.A2(n_907),
.B(n_897),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_R g1006 ( 
.A(n_1000),
.B(n_726),
.Y(n_1006)
);

NOR2x1_ASAP7_75t_L g1007 ( 
.A(n_999),
.B(n_710),
.Y(n_1007)
);

AOI211xp5_ASAP7_75t_L g1008 ( 
.A1(n_1006),
.A2(n_998),
.B(n_1005),
.C(n_1004),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_1007),
.A2(n_1003),
.B1(n_907),
.B2(n_860),
.Y(n_1009)
);

NAND5xp2_ASAP7_75t_L g1010 ( 
.A(n_1005),
.B(n_734),
.C(n_815),
.D(n_859),
.E(n_836),
.Y(n_1010)
);

AOI311xp33_ASAP7_75t_L g1011 ( 
.A1(n_1007),
.A2(n_882),
.A3(n_847),
.B(n_832),
.C(n_734),
.Y(n_1011)
);

NOR2x1_ASAP7_75t_L g1012 ( 
.A(n_1007),
.B(n_712),
.Y(n_1012)
);

OA22x2_ASAP7_75t_L g1013 ( 
.A1(n_1005),
.A2(n_816),
.B1(n_813),
.B2(n_843),
.Y(n_1013)
);

AOI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_1005),
.A2(n_724),
.B1(n_721),
.B2(n_915),
.Y(n_1014)
);

NAND3xp33_ASAP7_75t_SL g1015 ( 
.A(n_1006),
.B(n_728),
.C(n_915),
.Y(n_1015)
);

NAND3x1_ASAP7_75t_SL g1016 ( 
.A(n_1012),
.B(n_817),
.C(n_702),
.Y(n_1016)
);

NAND4xp25_ASAP7_75t_SL g1017 ( 
.A(n_1008),
.B(n_1014),
.C(n_1011),
.D(n_1015),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_1009),
.A2(n_817),
.B(n_790),
.Y(n_1018)
);

AOI222xp33_ASAP7_75t_L g1019 ( 
.A1(n_1010),
.A2(n_753),
.B1(n_807),
.B2(n_779),
.C1(n_715),
.C2(n_912),
.Y(n_1019)
);

OAI321xp33_ASAP7_75t_L g1020 ( 
.A1(n_1013),
.A2(n_867),
.A3(n_709),
.B1(n_836),
.B2(n_774),
.C(n_714),
.Y(n_1020)
);

AOI21xp33_ASAP7_75t_L g1021 ( 
.A1(n_1008),
.A2(n_817),
.B(n_175),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_1012),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_1012),
.B(n_841),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1012),
.Y(n_1024)
);

NAND4xp75_ASAP7_75t_L g1025 ( 
.A(n_1021),
.B(n_172),
.C(n_177),
.D(n_178),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_1023),
.B(n_912),
.Y(n_1026)
);

NOR4xp75_ASAP7_75t_L g1027 ( 
.A(n_1017),
.B(n_843),
.C(n_838),
.D(n_868),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1022),
.Y(n_1028)
);

OAI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_1018),
.A2(n_774),
.B1(n_792),
.B2(n_753),
.Y(n_1029)
);

NAND2x1_ASAP7_75t_L g1030 ( 
.A(n_1024),
.B(n_709),
.Y(n_1030)
);

NAND4xp25_ASAP7_75t_L g1031 ( 
.A(n_1019),
.B(n_712),
.C(n_716),
.D(n_838),
.Y(n_1031)
);

OAI221xp5_ASAP7_75t_L g1032 ( 
.A1(n_1016),
.A2(n_867),
.B1(n_702),
.B2(n_719),
.C(n_716),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_1020),
.B(n_911),
.Y(n_1033)
);

NOR3xp33_ASAP7_75t_L g1034 ( 
.A(n_1021),
.B(n_848),
.C(n_831),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_1017),
.A2(n_774),
.B1(n_883),
.B2(n_751),
.Y(n_1035)
);

NOR2x1_ASAP7_75t_L g1036 ( 
.A(n_1022),
.B(n_867),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_1023),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_1028),
.Y(n_1038)
);

INVxp67_ASAP7_75t_L g1039 ( 
.A(n_1037),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_1035),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_1029),
.Y(n_1041)
);

HB1xp67_ASAP7_75t_L g1042 ( 
.A(n_1030),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_1036),
.A2(n_702),
.B1(n_902),
.B2(n_911),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1026),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1027),
.Y(n_1045)
);

INVx1_ASAP7_75t_SL g1046 ( 
.A(n_1025),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_1039),
.A2(n_1031),
.B(n_1032),
.Y(n_1047)
);

AOI21xp33_ASAP7_75t_L g1048 ( 
.A1(n_1038),
.A2(n_1033),
.B(n_1034),
.Y(n_1048)
);

XNOR2x1_ASAP7_75t_L g1049 ( 
.A(n_1040),
.B(n_1046),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1042),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_R g1051 ( 
.A1(n_1043),
.A2(n_902),
.B(n_180),
.C(n_181),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1045),
.Y(n_1052)
);

INVx3_ASAP7_75t_L g1053 ( 
.A(n_1050),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1049),
.Y(n_1054)
);

AO22x2_ASAP7_75t_L g1055 ( 
.A1(n_1052),
.A2(n_1044),
.B1(n_1041),
.B2(n_841),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1055),
.Y(n_1056)
);

INVxp67_ASAP7_75t_L g1057 ( 
.A(n_1056),
.Y(n_1057)
);

OAI22x1_ASAP7_75t_L g1058 ( 
.A1(n_1057),
.A2(n_1054),
.B1(n_1053),
.B2(n_1048),
.Y(n_1058)
);

O2A1O1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_1058),
.A2(n_1047),
.B(n_1051),
.C(n_184),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1058),
.Y(n_1060)
);

AOI222xp33_ASAP7_75t_SL g1061 ( 
.A1(n_1060),
.A2(n_179),
.B1(n_183),
.B2(n_185),
.C1(n_187),
.C2(n_188),
.Y(n_1061)
);

INVx2_ASAP7_75t_SL g1062 ( 
.A(n_1059),
.Y(n_1062)
);

AOI22xp5_ASAP7_75t_SL g1063 ( 
.A1(n_1062),
.A2(n_714),
.B1(n_193),
.B2(n_194),
.Y(n_1063)
);

AOI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_1061),
.A2(n_714),
.B1(n_883),
.B2(n_751),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_SL g1065 ( 
.A1(n_1063),
.A2(n_191),
.B1(n_196),
.B2(n_199),
.Y(n_1065)
);

OAI21xp5_ASAP7_75t_SL g1066 ( 
.A1(n_1065),
.A2(n_1064),
.B(n_751),
.Y(n_1066)
);

AOI211xp5_ASAP7_75t_L g1067 ( 
.A1(n_1066),
.A2(n_848),
.B(n_831),
.C(n_821),
.Y(n_1067)
);


endmodule