module real_aes_3587_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_87;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_393;
wire n_294;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_L g359 ( .A(n_0), .B(n_291), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g373 ( .A(n_1), .Y(n_373) );
O2A1O1Ixp33_ASAP7_75t_SL g295 ( .A1(n_2), .A2(n_257), .B(n_296), .C(n_298), .Y(n_295) );
AOI22xp33_ASAP7_75t_L g176 ( .A1(n_3), .A2(n_56), .B1(n_177), .B2(n_180), .Y(n_176) );
OAI22xp33_ASAP7_75t_L g364 ( .A1(n_4), .A2(n_63), .B1(n_256), .B2(n_262), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_5), .Y(n_391) );
OAI22xp5_ASAP7_75t_L g259 ( .A1(n_6), .A2(n_52), .B1(n_260), .B2(n_262), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g643 ( .A(n_6), .Y(n_643) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_7), .Y(n_283) );
INVx1_ASAP7_75t_L g134 ( .A(n_8), .Y(n_134) );
INVxp67_ASAP7_75t_L g148 ( .A(n_8), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_8), .B(n_54), .Y(n_157) );
AOI22xp5_ASAP7_75t_L g253 ( .A1(n_9), .A2(n_43), .B1(n_254), .B2(n_256), .Y(n_253) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_9), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g216 ( .A1(n_10), .A2(n_20), .B1(n_217), .B2(n_221), .Y(n_216) );
OA21x2_ASAP7_75t_L g269 ( .A1(n_11), .A2(n_51), .B(n_270), .Y(n_269) );
OA21x2_ASAP7_75t_L g272 ( .A1(n_11), .A2(n_51), .B(n_270), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g130 ( .A(n_12), .B(n_119), .Y(n_130) );
HB1xp67_ASAP7_75t_L g83 ( .A(n_13), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_14), .Y(n_104) );
BUFx3_ASAP7_75t_L g229 ( .A(n_15), .Y(n_229) );
O2A1O1Ixp33_ASAP7_75t_L g302 ( .A1(n_16), .A2(n_303), .B(n_304), .C(n_306), .Y(n_302) );
OAI22xp33_ASAP7_75t_SL g362 ( .A1(n_17), .A2(n_32), .B1(n_256), .B2(n_282), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_18), .A2(n_23), .B1(n_282), .B2(n_286), .Y(n_351) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_19), .Y(n_119) );
O2A1O1Ixp5_ASAP7_75t_L g318 ( .A1(n_21), .A2(n_257), .B(n_319), .C(n_321), .Y(n_318) );
INVx1_ASAP7_75t_L g120 ( .A(n_22), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_22), .B(n_53), .Y(n_145) );
HB1xp67_ASAP7_75t_L g86 ( .A(n_24), .Y(n_86) );
AOI22xp33_ASAP7_75t_L g184 ( .A1(n_25), .A2(n_73), .B1(n_185), .B2(n_193), .Y(n_184) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_26), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_27), .B(n_336), .Y(n_355) );
HB1xp67_ASAP7_75t_L g89 ( .A(n_28), .Y(n_89) );
AOI22xp33_ASAP7_75t_L g197 ( .A1(n_29), .A2(n_74), .B1(n_198), .B2(n_202), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_30), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g206 ( .A1(n_31), .A2(n_62), .B1(n_207), .B2(n_211), .Y(n_206) );
INVx1_ASAP7_75t_L g270 ( .A(n_33), .Y(n_270) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_34), .Y(n_240) );
AND2x4_ASAP7_75t_L g266 ( .A(n_34), .B(n_238), .Y(n_266) );
AND2x4_ASAP7_75t_L g309 ( .A(n_34), .B(n_238), .Y(n_309) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_35), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_36), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_37), .Y(n_328) );
INVx2_ASAP7_75t_L g287 ( .A(n_38), .Y(n_287) );
O2A1O1Ixp33_ASAP7_75t_L g388 ( .A1(n_39), .A2(n_257), .B(n_389), .C(n_390), .Y(n_388) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_40), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g165 ( .A1(n_41), .A2(n_50), .B1(n_166), .B2(n_171), .Y(n_165) );
AOI22xp33_ASAP7_75t_SL g635 ( .A1(n_42), .A2(n_106), .B1(n_107), .B2(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_42), .Y(n_636) );
AOI21xp5_ASAP7_75t_L g110 ( .A1(n_44), .A2(n_111), .B(n_137), .Y(n_110) );
AOI22xp5_ASAP7_75t_L g352 ( .A1(n_45), .A2(n_60), .B1(n_297), .B2(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_46), .B(n_267), .Y(n_375) );
OA22x2_ASAP7_75t_L g124 ( .A1(n_47), .A2(n_54), .B1(n_119), .B2(n_123), .Y(n_124) );
INVx1_ASAP7_75t_L g164 ( .A(n_47), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_48), .Y(n_374) );
NAND2xp33_ASAP7_75t_R g271 ( .A(n_49), .B(n_272), .Y(n_271) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_49), .A2(n_77), .B1(n_336), .B2(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g136 ( .A(n_53), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_53), .B(n_161), .Y(n_160) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_53), .Y(n_232) );
OAI21xp33_ASAP7_75t_L g175 ( .A1(n_54), .A2(n_61), .B(n_149), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_55), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_57), .Y(n_285) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_58), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_59), .Y(n_102) );
INVx1_ASAP7_75t_L g122 ( .A(n_61), .Y(n_122) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_61), .B(n_72), .Y(n_158) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_64), .Y(n_255) );
BUFx5_ASAP7_75t_L g256 ( .A(n_64), .Y(n_256) );
INVx1_ASAP7_75t_L g261 ( .A(n_64), .Y(n_261) );
INVx2_ASAP7_75t_L g311 ( .A(n_65), .Y(n_311) );
INVx2_ASAP7_75t_L g393 ( .A(n_66), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g305 ( .A(n_67), .Y(n_305) );
INVx1_ASAP7_75t_L g138 ( .A(n_68), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_69), .B(n_151), .Y(n_150) );
INVx2_ASAP7_75t_SL g238 ( .A(n_70), .Y(n_238) );
INVx1_ASAP7_75t_L g326 ( .A(n_71), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_72), .B(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g331 ( .A(n_75), .Y(n_331) );
OAI21xp33_ASAP7_75t_SL g386 ( .A1(n_76), .A2(n_256), .B(n_387), .Y(n_386) );
INVxp67_ASAP7_75t_SL g289 ( .A(n_77), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_77), .B(n_336), .Y(n_335) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_224), .B1(n_241), .B2(n_622), .C(n_629), .Y(n_78) );
XOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_98), .Y(n_79) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_81), .A2(n_82), .B1(n_96), .B2(n_97), .Y(n_80) );
CKINVDCx14_ASAP7_75t_R g96 ( .A(n_81), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_82), .Y(n_97) );
AOI22xp5_ASAP7_75t_L g82 ( .A1(n_83), .A2(n_84), .B1(n_94), .B2(n_95), .Y(n_82) );
INVx1_ASAP7_75t_L g94 ( .A(n_83), .Y(n_94) );
CKINVDCx20_ASAP7_75t_R g95 ( .A(n_84), .Y(n_95) );
AOI22xp5_ASAP7_75t_L g84 ( .A1(n_85), .A2(n_87), .B1(n_88), .B2(n_93), .Y(n_84) );
CKINVDCx20_ASAP7_75t_R g93 ( .A(n_85), .Y(n_93) );
BUFx2_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
INVx1_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
OAI22xp5_ASAP7_75t_L g88 ( .A1(n_89), .A2(n_90), .B1(n_91), .B2(n_92), .Y(n_88) );
INVx1_ASAP7_75t_L g91 ( .A(n_89), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_90), .Y(n_92) );
AOI22xp33_ASAP7_75t_SL g98 ( .A1(n_99), .A2(n_100), .B1(n_106), .B2(n_107), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
OAI22xp5_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_103), .B1(n_104), .B2(n_105), .Y(n_100) );
INVx1_ASAP7_75t_L g105 ( .A(n_101), .Y(n_105) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_102), .A2(n_256), .B1(n_282), .B2(n_283), .Y(n_281) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
NAND2xp5_ASAP7_75t_SL g387 ( .A(n_104), .B(n_256), .Y(n_387) );
AOI22xp33_ASAP7_75t_SL g630 ( .A1(n_106), .A2(n_107), .B1(n_631), .B2(n_632), .Y(n_630) );
INVxp67_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
NOR2x1_ASAP7_75t_L g108 ( .A(n_109), .B(n_183), .Y(n_108) );
NAND3xp33_ASAP7_75t_L g109 ( .A(n_110), .B(n_165), .C(n_176), .Y(n_109) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx3_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_125), .Y(n_115) );
AND2x2_ASAP7_75t_L g182 ( .A(n_116), .B(n_179), .Y(n_182) );
AND2x2_ASAP7_75t_L g199 ( .A(n_116), .B(n_200), .Y(n_199) );
AND2x4_ASAP7_75t_L g204 ( .A(n_116), .B(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_124), .Y(n_116) );
INVx1_ASAP7_75t_L g170 ( .A(n_117), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_121), .Y(n_117) );
NAND2xp33_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
INVx2_ASAP7_75t_L g123 ( .A(n_119), .Y(n_123) );
INVx3_ASAP7_75t_L g129 ( .A(n_119), .Y(n_129) );
NAND2xp33_ASAP7_75t_L g135 ( .A(n_119), .B(n_136), .Y(n_135) );
HB1xp67_ASAP7_75t_L g144 ( .A(n_119), .Y(n_144) );
INVx1_ASAP7_75t_L g149 ( .A(n_119), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_120), .B(n_164), .Y(n_163) );
INVxp67_ASAP7_75t_L g233 ( .A(n_120), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
OAI21xp5_ASAP7_75t_L g147 ( .A1(n_122), .A2(n_148), .B(n_149), .Y(n_147) );
AND2x2_ASAP7_75t_L g146 ( .A(n_124), .B(n_147), .Y(n_146) );
AND2x2_ASAP7_75t_L g169 ( .A(n_124), .B(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g189 ( .A(n_124), .Y(n_189) );
AND2x4_ASAP7_75t_L g168 ( .A(n_125), .B(n_169), .Y(n_168) );
AND2x4_ASAP7_75t_L g173 ( .A(n_125), .B(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g215 ( .A(n_125), .B(n_188), .Y(n_215) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_131), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g142 ( .A(n_127), .B(n_143), .Y(n_142) );
AND2x4_ASAP7_75t_L g179 ( .A(n_127), .B(n_131), .Y(n_179) );
OR2x2_ASAP7_75t_L g191 ( .A(n_127), .B(n_192), .Y(n_191) );
AND2x4_ASAP7_75t_L g200 ( .A(n_127), .B(n_201), .Y(n_200) );
AND2x4_ASAP7_75t_L g127 ( .A(n_128), .B(n_130), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_129), .B(n_134), .Y(n_133) );
INVxp67_ASAP7_75t_L g161 ( .A(n_129), .Y(n_161) );
NAND3xp33_ASAP7_75t_L g159 ( .A(n_130), .B(n_160), .C(n_162), .Y(n_159) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g192 ( .A(n_132), .Y(n_192) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_135), .Y(n_132) );
OAI21xp33_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_139), .B(n_150), .Y(n_137) );
INVx2_ASAP7_75t_SL g139 ( .A(n_140), .Y(n_139) );
BUFx4f_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_146), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
INVx1_ASAP7_75t_L g155 ( .A(n_144), .Y(n_155) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_145), .Y(n_230) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx4_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AO21x2_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_156), .B(n_159), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_161), .B(n_163), .Y(n_162) );
AND2x2_ASAP7_75t_L g174 ( .A(n_162), .B(n_175), .Y(n_174) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_164), .Y(n_234) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x4_ASAP7_75t_L g178 ( .A(n_169), .B(n_179), .Y(n_178) );
AND2x4_ASAP7_75t_L g188 ( .A(n_170), .B(n_189), .Y(n_188) );
BUFx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AND2x4_ASAP7_75t_L g196 ( .A(n_174), .B(n_190), .Y(n_196) );
AND2x4_ASAP7_75t_L g223 ( .A(n_174), .B(n_200), .Y(n_223) );
BUFx3_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AND2x4_ASAP7_75t_L g210 ( .A(n_179), .B(n_188), .Y(n_210) );
BUFx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
BUFx3_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NAND4xp25_ASAP7_75t_L g183 ( .A(n_184), .B(n_197), .C(n_206), .D(n_216), .Y(n_183) );
BUFx3_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AND2x4_ASAP7_75t_L g187 ( .A(n_188), .B(n_190), .Y(n_187) );
AND2x4_ASAP7_75t_L g220 ( .A(n_188), .B(n_200), .Y(n_220) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g205 ( .A(n_191), .Y(n_205) );
INVx1_ASAP7_75t_L g201 ( .A(n_192), .Y(n_201) );
BUFx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx6_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
BUFx8_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
BUFx3_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
BUFx4f_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx3_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
BUFx12f_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx4_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx8_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
BUFx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_227), .B(n_235), .Y(n_226) );
INVxp67_ASAP7_75t_SL g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g634 ( .A(n_228), .B(n_235), .Y(n_634) );
AOI211xp5_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_231), .C(n_234), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_232), .B(n_233), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_236), .B(n_239), .Y(n_235) );
OR2x2_ASAP7_75t_L g638 ( .A(n_236), .B(n_240), .Y(n_638) );
INVx1_ASAP7_75t_L g641 ( .A(n_236), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_236), .B(n_239), .Y(n_642) );
HB1xp67_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x4_ASAP7_75t_L g242 ( .A(n_243), .B(n_519), .Y(n_242) );
NOR3xp33_ASAP7_75t_L g243 ( .A(n_244), .B(n_430), .C(n_478), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_376), .Y(n_244) );
OAI21xp33_ASAP7_75t_SL g245 ( .A1(n_246), .A2(n_312), .B(n_343), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_246), .A2(n_590), .B(n_592), .Y(n_589) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
OR2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_273), .Y(n_247) );
OR2x2_ASAP7_75t_L g517 ( .A(n_248), .B(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_248), .B(n_550), .Y(n_549) );
INVx2_ASAP7_75t_SL g248 ( .A(n_249), .Y(n_248) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g398 ( .A(n_250), .Y(n_398) );
INVx2_ASAP7_75t_L g429 ( .A(n_250), .Y(n_429) );
AND2x2_ASAP7_75t_L g450 ( .A(n_250), .B(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g569 ( .A(n_250), .B(n_275), .Y(n_569) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_271), .Y(n_250) );
AND2x2_ASAP7_75t_L g470 ( .A(n_251), .B(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_264), .Y(n_251) );
AOI22xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_257), .B1(n_259), .B2(n_263), .Y(n_252) );
AOI22xp5_ASAP7_75t_L g284 ( .A1(n_254), .A2(n_285), .B1(n_286), .B2(n_287), .Y(n_284) );
INVx1_ASAP7_75t_L g303 ( .A(n_254), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_254), .A2(n_256), .B1(n_373), .B2(n_374), .Y(n_372) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g262 ( .A(n_255), .Y(n_262) );
INVx6_ASAP7_75t_L g282 ( .A(n_255), .Y(n_282) );
INVx3_ASAP7_75t_L g320 ( .A(n_255), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_256), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_256), .B(n_328), .Y(n_327) );
AOI22xp33_ASAP7_75t_SL g369 ( .A1(n_256), .A2(n_282), .B1(n_370), .B2(n_371), .Y(n_369) );
OAI22xp33_ASAP7_75t_L g280 ( .A1(n_257), .A2(n_263), .B1(n_281), .B2(n_284), .Y(n_280) );
INVx1_ASAP7_75t_L g342 ( .A(n_257), .Y(n_342) );
OAI221xp5_ASAP7_75t_L g368 ( .A1(n_257), .A2(n_266), .B1(n_306), .B2(n_369), .C(n_372), .Y(n_368) );
BUFx6f_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx4_ASAP7_75t_L g263 ( .A(n_258), .Y(n_263) );
INVx3_ASAP7_75t_L g306 ( .A(n_258), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_258), .B(n_326), .Y(n_325) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_258), .Y(n_350) );
INVx1_ASAP7_75t_L g354 ( .A(n_258), .Y(n_354) );
NAND2xp5_ASAP7_75t_SL g361 ( .A(n_258), .B(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g297 ( .A(n_260), .Y(n_297) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g286 ( .A(n_261), .Y(n_286) );
OAI22xp5_ASAP7_75t_L g323 ( .A1(n_263), .A2(n_324), .B1(n_325), .B2(n_327), .Y(n_323) );
INVx2_ASAP7_75t_L g339 ( .A(n_263), .Y(n_339) );
NOR2xp67_ASAP7_75t_L g264 ( .A(n_265), .B(n_267), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_266), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_266), .B(n_292), .Y(n_365) );
INVx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
BUFx3_ASAP7_75t_L g329 ( .A(n_268), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_268), .B(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx4_ASAP7_75t_L g292 ( .A(n_269), .Y(n_292) );
BUFx3_ASAP7_75t_L g416 ( .A(n_269), .Y(n_416) );
BUFx3_ASAP7_75t_L g279 ( .A(n_272), .Y(n_279) );
INVx1_ASAP7_75t_L g332 ( .A(n_272), .Y(n_332) );
INVx1_ASAP7_75t_L g384 ( .A(n_272), .Y(n_384) );
INVx2_ASAP7_75t_L g473 ( .A(n_272), .Y(n_473) );
INVx2_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_274), .B(n_402), .Y(n_522) );
AND2x2_ASAP7_75t_L g609 ( .A(n_274), .B(n_553), .Y(n_609) );
AND2x4_ASAP7_75t_L g274 ( .A(n_275), .B(n_293), .Y(n_274) );
INVx1_ASAP7_75t_L g426 ( .A(n_275), .Y(n_426) );
OAI21x1_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_280), .B(n_288), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
AND2x2_ASAP7_75t_SL g623 ( .A(n_277), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_278), .B(n_309), .Y(n_348) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g340 ( .A(n_281), .Y(n_340) );
INVx2_ASAP7_75t_L g299 ( .A(n_282), .Y(n_299) );
INVx2_ASAP7_75t_SL g353 ( .A(n_282), .Y(n_353) );
INVx1_ASAP7_75t_L g341 ( .A(n_284), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_286), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_SL g390 ( .A(n_286), .B(n_391), .Y(n_390) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
INVx2_ASAP7_75t_L g367 ( .A(n_290), .Y(n_367) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NOR2xp33_ASAP7_75t_SL g307 ( .A(n_291), .B(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_SL g310 ( .A(n_292), .B(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g336 ( .A(n_292), .Y(n_336) );
OR2x2_ASAP7_75t_L g333 ( .A(n_293), .B(n_334), .Y(n_333) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_293), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_293), .B(n_316), .Y(n_407) );
INVx2_ASAP7_75t_L g428 ( .A(n_293), .Y(n_428) );
INVx1_ASAP7_75t_L g467 ( .A(n_293), .Y(n_467) );
INVx1_ASAP7_75t_L g508 ( .A(n_293), .Y(n_508) );
AND2x2_ASAP7_75t_L g543 ( .A(n_293), .B(n_334), .Y(n_543) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_293), .Y(n_598) );
AO31x2_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_301), .A3(n_307), .B(n_310), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_303), .Y(n_625) );
AOI21xp5_ASAP7_75t_L g363 ( .A1(n_306), .A2(n_364), .B(n_365), .Y(n_363) );
NOR3xp33_ASAP7_75t_L g317 ( .A(n_308), .B(n_318), .C(n_323), .Y(n_317) );
AOI221xp5_ASAP7_75t_L g338 ( .A1(n_308), .A2(n_339), .B1(n_340), .B2(n_341), .C(n_342), .Y(n_338) );
INVx4_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g383 ( .A(n_309), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_333), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g397 ( .A(n_316), .B(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g436 ( .A(n_316), .B(n_428), .Y(n_436) );
INVx2_ASAP7_75t_L g451 ( .A(n_316), .Y(n_451) );
INVx2_ASAP7_75t_L g477 ( .A(n_316), .Y(n_477) );
AO21x2_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_329), .B(n_330), .Y(n_316) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g324 ( .A(n_320), .Y(n_324) );
INVx1_ASAP7_75t_L g389 ( .A(n_320), .Y(n_389) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_329), .B(n_338), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_333), .Y(n_433) );
OR2x2_ASAP7_75t_L g448 ( .A(n_333), .B(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g525 ( .A(n_333), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_334), .B(n_477), .Y(n_476) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_334), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_334), .B(n_533), .Y(n_559) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
AND2x2_ASAP7_75t_L g469 ( .A(n_337), .B(n_470), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g385 ( .A1(n_339), .A2(n_386), .B(n_388), .Y(n_385) );
AOI322xp5_ASAP7_75t_L g551 ( .A1(n_343), .A2(n_491), .A3(n_529), .B1(n_552), .B2(n_554), .C1(n_555), .C2(n_556), .Y(n_551) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_356), .Y(n_343) );
AND2x2_ASAP7_75t_L g556 ( .A(n_344), .B(n_536), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_344), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g607 ( .A(n_344), .B(n_499), .Y(n_607) );
INVx3_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_345), .B(n_404), .Y(n_422) );
AND2x2_ASAP7_75t_L g483 ( .A(n_345), .B(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_345), .B(n_445), .Y(n_527) );
AND2x4_ASAP7_75t_L g564 ( .A(n_345), .B(n_356), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_345), .B(n_486), .Y(n_605) );
INVx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g394 ( .A(n_346), .B(n_366), .Y(n_394) );
INVx1_ASAP7_75t_L g443 ( .A(n_346), .Y(n_443) );
AND2x2_ASAP7_75t_L g587 ( .A(n_346), .B(n_420), .Y(n_587) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g405 ( .A(n_347), .Y(n_405) );
OAI21x1_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_349), .B(n_355), .Y(n_347) );
INVx1_ASAP7_75t_L g414 ( .A(n_349), .Y(n_414) );
OA22x2_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_351), .B1(n_352), .B2(n_354), .Y(n_349) );
INVx4_ASAP7_75t_L g628 ( .A(n_350), .Y(n_628) );
INVx1_ASAP7_75t_L g417 ( .A(n_355), .Y(n_417) );
INVx1_ASAP7_75t_SL g512 ( .A(n_356), .Y(n_512) );
AND2x4_ASAP7_75t_L g356 ( .A(n_357), .B(n_366), .Y(n_356) );
AND2x2_ASAP7_75t_L g404 ( .A(n_357), .B(n_381), .Y(n_404) );
INVx1_ASAP7_75t_L g445 ( .A(n_357), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_357), .B(n_380), .Y(n_621) );
INVx3_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g420 ( .A(n_358), .Y(n_420) );
INVx1_ASAP7_75t_L g462 ( .A(n_358), .Y(n_462) );
AND2x2_ASAP7_75t_L g486 ( .A(n_358), .B(n_366), .Y(n_486) );
AND2x2_ASAP7_75t_L g536 ( .A(n_358), .B(n_381), .Y(n_536) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_358), .Y(n_540) );
AND2x4_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_363), .Y(n_360) );
OR2x2_ASAP7_75t_L g412 ( .A(n_366), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g442 ( .A(n_366), .B(n_443), .Y(n_442) );
OA21x2_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_368), .B(n_375), .Y(n_366) );
OA21x2_ASAP7_75t_L g457 ( .A1(n_367), .A2(n_368), .B(n_375), .Y(n_457) );
AOI221xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_395), .B1(n_402), .B2(n_406), .C(n_408), .Y(n_376) );
INVxp67_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_379), .B(n_394), .Y(n_378) );
AND2x2_ASAP7_75t_L g582 ( .A(n_379), .B(n_442), .Y(n_582) );
BUFx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OR2x2_ASAP7_75t_L g596 ( .A(n_380), .B(n_477), .Y(n_596) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OR2x2_ASAP7_75t_L g419 ( .A(n_381), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g440 ( .A(n_381), .Y(n_440) );
AND2x2_ASAP7_75t_L g463 ( .A(n_381), .B(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g485 ( .A(n_381), .Y(n_485) );
BUFx2_ASAP7_75t_L g573 ( .A(n_381), .Y(n_573) );
INVx3_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AOI21x1_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_385), .B(n_392), .Y(n_382) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_394), .A2(n_418), .B(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g585 ( .A(n_394), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_395), .A2(n_432), .B1(n_437), .B2(n_444), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_396), .B(n_399), .Y(n_395) );
OR2x2_ASAP7_75t_L g493 ( .A(n_396), .B(n_494), .Y(n_493) );
INVx2_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
AND2x4_ASAP7_75t_L g524 ( .A(n_397), .B(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g542 ( .A(n_397), .B(n_543), .Y(n_542) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g616 ( .A(n_401), .B(n_532), .Y(n_616) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NOR2xp33_ASAP7_75t_SL g528 ( .A(n_403), .B(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
AND2x2_ASAP7_75t_L g504 ( .A(n_405), .B(n_485), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_405), .B(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g591 ( .A(n_405), .Y(n_591) );
OR2x2_ASAP7_75t_L g620 ( .A(n_405), .B(n_621), .Y(n_620) );
AND2x4_ASAP7_75t_L g588 ( .A(n_406), .B(n_569), .Y(n_588) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AOI21xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_421), .B(n_423), .Y(n_408) );
INVx2_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_418), .Y(n_410) );
AND2x2_ASAP7_75t_L g444 ( .A(n_411), .B(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g546 ( .A(n_411), .B(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AND2x4_ASAP7_75t_L g455 ( .A(n_413), .B(n_456), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_415), .B(n_417), .Y(n_413) );
INVx3_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AND2x4_ASAP7_75t_L g499 ( .A(n_420), .B(n_456), .Y(n_499) );
OAI21xp33_ASAP7_75t_L g617 ( .A1(n_421), .A2(n_506), .B(n_618), .Y(n_617) );
BUFx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_424), .B(n_427), .Y(n_423) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OR2x2_ASAP7_75t_L g599 ( .A(n_425), .B(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g474 ( .A(n_427), .B(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g558 ( .A(n_427), .B(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
INVx1_ASAP7_75t_L g495 ( .A(n_428), .Y(n_495) );
INVx1_ASAP7_75t_L g534 ( .A(n_429), .Y(n_534) );
AND2x4_ASAP7_75t_L g553 ( .A(n_429), .B(n_477), .Y(n_553) );
INVx1_ASAP7_75t_SL g600 ( .A(n_429), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_431), .B(n_446), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g568 ( .A(n_436), .B(n_569), .Y(n_568) );
NOR2x1_ASAP7_75t_L g437 ( .A(n_438), .B(n_441), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OR2x2_ASAP7_75t_L g453 ( .A(n_439), .B(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g552 ( .A(n_439), .B(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_440), .B(n_464), .Y(n_614) );
INVx3_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_444), .B(n_465), .Y(n_500) );
AND2x2_ASAP7_75t_L g491 ( .A(n_445), .B(n_455), .Y(n_491) );
AOI222xp33_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_452), .B1(n_458), .B2(n_460), .C1(n_465), .C2(n_474), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OAI21xp33_ASAP7_75t_L g497 ( .A1(n_448), .A2(n_498), .B(n_500), .Y(n_497) );
OAI221xp5_ASAP7_75t_L g565 ( .A1(n_448), .A2(n_566), .B1(n_567), .B2(n_570), .C(n_574), .Y(n_565) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
BUFx2_ASAP7_75t_L g480 ( .A(n_450), .Y(n_480) );
AND2x2_ASAP7_75t_L g509 ( .A(n_451), .B(n_469), .Y(n_509) );
INVx1_ASAP7_75t_L g533 ( .A(n_451), .Y(n_533) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_451), .Y(n_562) );
OAI21xp5_ASAP7_75t_L g545 ( .A1(n_452), .A2(n_546), .B(n_548), .Y(n_545) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g576 ( .A(n_455), .B(n_547), .Y(n_576) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g464 ( .A(n_457), .Y(n_464) );
INVxp67_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
AND2x4_ASAP7_75t_L g460 ( .A(n_461), .B(n_463), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_463), .Y(n_490) );
INVx2_ASAP7_75t_L g541 ( .A(n_464), .Y(n_541) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
OR2x2_ASAP7_75t_L g597 ( .A(n_468), .B(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g563 ( .A(n_469), .Y(n_563) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_474), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
OR2x2_ASAP7_75t_L g518 ( .A(n_476), .B(n_495), .Y(n_518) );
NAND4xp25_ASAP7_75t_L g478 ( .A(n_479), .B(n_487), .C(n_496), .D(n_501), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
A2O1A1Ixp33_ASAP7_75t_L g574 ( .A1(n_480), .A2(n_575), .B(n_576), .C(n_577), .Y(n_574) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_486), .Y(n_484) );
INVx1_ASAP7_75t_L g515 ( .A(n_485), .Y(n_515) );
INVx1_ASAP7_75t_L g547 ( .A(n_485), .Y(n_547) );
OAI21xp5_ASAP7_75t_SL g487 ( .A1(n_488), .A2(n_491), .B(n_492), .Y(n_487) );
INVxp67_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVxp33_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
NAND2x1p5_ASAP7_75t_L g578 ( .A(n_499), .B(n_573), .Y(n_578) );
AND2x4_ASAP7_75t_L g590 ( .A(n_499), .B(n_591), .Y(n_590) );
NAND2x1p5_ASAP7_75t_L g601 ( .A(n_499), .B(n_514), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_505), .B1(n_510), .B2(n_516), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
NAND2x1p5_ASAP7_75t_SL g506 ( .A(n_507), .B(n_509), .Y(n_506) );
INVx2_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g575 ( .A(n_508), .Y(n_575) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_509), .Y(n_555) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_513), .Y(n_511) );
OR2x2_ASAP7_75t_L g566 ( .A(n_513), .B(n_539), .Y(n_566) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g554 ( .A(n_518), .Y(n_554) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_579), .Y(n_519) );
NOR3xp33_ASAP7_75t_L g520 ( .A(n_521), .B(n_544), .C(n_565), .Y(n_520) );
NAND3xp33_ASAP7_75t_L g521 ( .A(n_522), .B(n_523), .C(n_535), .Y(n_521) );
AOI22x1_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_526), .B1(n_528), .B2(n_530), .Y(n_523) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
OAI21xp33_ASAP7_75t_SL g535 ( .A1(n_536), .A2(n_537), .B(n_542), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_541), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVxp67_ASAP7_75t_L g613 ( .A(n_540), .Y(n_613) );
INVx1_ASAP7_75t_L g593 ( .A(n_541), .Y(n_593) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_543), .Y(n_550) );
NAND3xp33_ASAP7_75t_L g544 ( .A(n_545), .B(n_551), .C(n_557), .Y(n_544) );
INVx1_ASAP7_75t_L g586 ( .A(n_547), .Y(n_586) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
OAI21xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_560), .B(n_564), .Y(n_557) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_558), .A2(n_576), .B1(n_611), .B2(n_615), .Y(n_610) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVxp67_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NOR3xp33_ASAP7_75t_L g579 ( .A(n_580), .B(n_602), .C(n_617), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_589), .Y(n_580) );
OAI31xp33_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_583), .A3(n_587), .B(n_588), .Y(n_581) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_594), .B1(n_599), .B2(n_601), .Y(n_592) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NOR2x1_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
A2O1A1Ixp33_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_606), .B(n_608), .C(n_610), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
OR2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
BUFx3_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OA21x2_ASAP7_75t_L g640 ( .A1(n_624), .A2(n_641), .B(n_642), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
CKINVDCx20_ASAP7_75t_R g626 ( .A(n_627), .Y(n_626) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OAI222xp33_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_633), .B1(n_635), .B2(n_637), .C1(n_639), .C2(n_643), .Y(n_629) );
CKINVDCx5p33_ASAP7_75t_R g632 ( .A(n_631), .Y(n_632) );
INVx1_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
BUFx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
BUFx3_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
endmodule