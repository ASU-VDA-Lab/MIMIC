module fake_jpeg_26799_n_324 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_40),
.Y(n_50)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_24),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_39),
.C(n_40),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_46),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_19),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_21),
.Y(n_80)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_53),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_25),
.B1(n_31),
.B2(n_28),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_51),
.A2(n_58),
.B1(n_60),
.B2(n_36),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_39),
.A2(n_25),
.B1(n_29),
.B2(n_28),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_52),
.A2(n_23),
.B1(n_20),
.B2(n_32),
.Y(n_92)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_40),
.B(n_19),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_54),
.B(n_59),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_18),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_64),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_36),
.A2(n_25),
.B1(n_29),
.B2(n_26),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_36),
.A2(n_29),
.B1(n_26),
.B2(n_23),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_20),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_65),
.A2(n_69),
.B1(n_77),
.B2(n_92),
.Y(n_94)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_67),
.B(n_70),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_68),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_36),
.B1(n_34),
.B2(n_26),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_71),
.Y(n_99)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_48),
.A2(n_24),
.B1(n_21),
.B2(n_17),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_49),
.Y(n_76)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_45),
.A2(n_36),
.B1(n_34),
.B2(n_32),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_59),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_46),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_85),
.Y(n_101)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_90),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_55),
.A2(n_17),
.B1(n_16),
.B2(n_33),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_88),
.A2(n_91),
.B1(n_46),
.B2(n_52),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_57),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_89),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_43),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_55),
.A2(n_16),
.B1(n_33),
.B2(n_23),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_47),
.B(n_43),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_38),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_80),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_100),
.B1(n_113),
.B2(n_115),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_64),
.C(n_56),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_104),
.C(n_86),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_64),
.B1(n_51),
.B2(n_56),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_73),
.B(n_53),
.C(n_57),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_106),
.B(n_116),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_89),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_112),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_85),
.A2(n_55),
.B1(n_61),
.B2(n_49),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_82),
.A2(n_61),
.B1(n_62),
.B2(n_54),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_93),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_86),
.A2(n_0),
.B(n_1),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_68),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_119),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_84),
.A2(n_62),
.B1(n_43),
.B2(n_41),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_121),
.A2(n_65),
.B1(n_67),
.B2(n_75),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_87),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_123),
.B(n_129),
.C(n_130),
.Y(n_171)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_124),
.B(n_145),
.Y(n_154)
);

INVxp33_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_125),
.B(n_126),
.Y(n_168)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_102),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_77),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_83),
.Y(n_131)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_109),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_132),
.Y(n_176)
);

OAI32xp33_ASAP7_75t_L g133 ( 
.A1(n_101),
.A2(n_86),
.A3(n_92),
.B1(n_83),
.B2(n_69),
.Y(n_133)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_135),
.A2(n_140),
.B1(n_108),
.B2(n_110),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_96),
.A2(n_94),
.B1(n_120),
.B2(n_115),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_137),
.A2(n_128),
.B1(n_94),
.B2(n_149),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_78),
.C(n_79),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_138),
.B(n_142),
.C(n_151),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_120),
.A2(n_75),
.B1(n_71),
.B2(n_72),
.Y(n_140)
);

NAND2xp33_ASAP7_75t_SL g141 ( 
.A(n_118),
.B(n_33),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_141),
.A2(n_111),
.B1(n_76),
.B2(n_99),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_98),
.B(n_78),
.C(n_66),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_67),
.Y(n_143)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_62),
.Y(n_144)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_97),
.Y(n_145)
);

BUFx24_ASAP7_75t_SL g146 ( 
.A(n_95),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_146),
.B(n_148),
.Y(n_167)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_149),
.B(n_150),
.Y(n_174)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_98),
.B(n_35),
.C(n_38),
.Y(n_151)
);

OAI21xp33_ASAP7_75t_SL g208 ( 
.A1(n_152),
.A2(n_22),
.B(n_30),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_153),
.B(n_157),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_150),
.A2(n_117),
.B(n_102),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_155),
.A2(n_160),
.B(n_183),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_106),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_156),
.B(n_165),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_158),
.A2(n_159),
.B1(n_162),
.B2(n_164),
.Y(n_199)
);

NAND2x1_ASAP7_75t_L g160 ( 
.A(n_122),
.B(n_100),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_137),
.A2(n_95),
.B1(n_103),
.B2(n_110),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_161),
.A2(n_177),
.B1(n_182),
.B2(n_153),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_128),
.A2(n_105),
.B1(n_103),
.B2(n_71),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_148),
.A2(n_105),
.B1(n_108),
.B2(n_119),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_95),
.Y(n_165)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_173),
.Y(n_194)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_133),
.A2(n_107),
.B1(n_76),
.B2(n_68),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_130),
.A2(n_107),
.B1(n_43),
.B2(n_41),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_178),
.A2(n_181),
.B1(n_41),
.B2(n_23),
.Y(n_201)
);

MAJx2_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_22),
.C(n_38),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_1),
.C(n_2),
.Y(n_209)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_136),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_180),
.B(n_30),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_151),
.A2(n_142),
.B1(n_139),
.B2(n_147),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_147),
.A2(n_41),
.B1(n_38),
.B2(n_35),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_139),
.A2(n_22),
.B(n_30),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_124),
.A2(n_0),
.B(n_1),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_182),
.Y(n_193)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_186),
.B(n_188),
.Y(n_238)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_156),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_169),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_196),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_163),
.B(n_123),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_190),
.B(n_197),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_177),
.A2(n_145),
.B1(n_126),
.B2(n_20),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_192),
.A2(n_195),
.B1(n_202),
.B2(n_203),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_193),
.A2(n_208),
.B(n_211),
.Y(n_222)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_169),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_164),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_206),
.Y(n_233)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_200),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_178),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_160),
.A2(n_32),
.B1(n_22),
.B2(n_27),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_166),
.A2(n_27),
.B1(n_30),
.B2(n_22),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_27),
.Y(n_204)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_204),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_174),
.B(n_170),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_162),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_207),
.B(n_210),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_185),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_175),
.B(n_173),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_161),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_166),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_212),
.A2(n_214),
.B1(n_157),
.B2(n_4),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_172),
.B(n_13),
.Y(n_213)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_213),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_159),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_215),
.B(n_224),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_211),
.A2(n_160),
.B1(n_165),
.B2(n_184),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_216),
.A2(n_229),
.B1(n_220),
.B2(n_230),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_234),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_181),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_220),
.B(n_230),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_194),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_187),
.A2(n_152),
.B(n_157),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_226),
.A2(n_232),
.B(n_237),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_231),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_195),
.A2(n_184),
.B1(n_179),
.B2(n_171),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_171),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_194),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_197),
.A2(n_155),
.B(n_183),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_210),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_201),
.B(n_167),
.C(n_13),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_215),
.C(n_227),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_191),
.Y(n_236)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_236),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_207),
.A2(n_12),
.B(n_11),
.Y(n_237)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_228),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_241),
.Y(n_267)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_223),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_239),
.B(n_188),
.Y(n_244)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_244),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_206),
.Y(n_245)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_246),
.A2(n_257),
.B1(n_209),
.B2(n_237),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_186),
.Y(n_248)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_248),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_191),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_254),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_226),
.A2(n_198),
.B(n_199),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_253),
.A2(n_222),
.B(n_232),
.Y(n_261)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_233),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_256),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_203),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_3),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_221),
.A2(n_192),
.B1(n_214),
.B2(n_212),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_216),
.B(n_190),
.C(n_199),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_258),
.B(n_222),
.C(n_217),
.Y(n_260)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_218),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_259),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_249),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_261),
.A2(n_242),
.B(n_252),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_264),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_235),
.C(n_221),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_246),
.C(n_258),
.Y(n_277)
);

AO221x1_ASAP7_75t_L g266 ( 
.A1(n_241),
.A2(n_225),
.B1(n_196),
.B2(n_189),
.C(n_219),
.Y(n_266)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_266),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_243),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_245),
.Y(n_271)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_271),
.Y(n_282)
);

XOR2x1_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_12),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_272),
.A2(n_10),
.B(n_6),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_242),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_274)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_273),
.B(n_259),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_276),
.B(n_277),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_278),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_260),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_240),
.Y(n_283)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_283),
.Y(n_294)
);

A2O1A1Ixp33_ASAP7_75t_SL g284 ( 
.A1(n_272),
.A2(n_253),
.B(n_248),
.C(n_251),
.Y(n_284)
);

AO21x1_ASAP7_75t_L g292 ( 
.A1(n_284),
.A2(n_261),
.B(n_275),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_244),
.Y(n_285)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_285),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_286),
.A2(n_288),
.B1(n_265),
.B2(n_268),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_247),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_289),
.A2(n_270),
.B1(n_269),
.B2(n_250),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_296),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_292),
.A2(n_301),
.B1(n_284),
.B2(n_7),
.Y(n_307)
);

FAx1_ASAP7_75t_SL g293 ( 
.A(n_284),
.B(n_278),
.CI(n_279),
.CON(n_293),
.SN(n_293)
);

NOR2x1_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_10),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_263),
.C(n_262),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_299),
.C(n_294),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_298),
.B(n_282),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_287),
.A2(n_250),
.B1(n_10),
.B2(n_7),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_285),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_293),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_295),
.B(n_281),
.C(n_284),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_303),
.B(n_305),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_292),
.Y(n_306)
);

OAI21x1_ASAP7_75t_L g313 ( 
.A1(n_306),
.A2(n_293),
.B(n_291),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_308),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_297),
.A2(n_6),
.B(n_7),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_309),
.A2(n_291),
.B(n_9),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_300),
.B(n_8),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_310),
.B(n_301),
.Y(n_311)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_311),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_315),
.C(n_316),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_304),
.C(n_290),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_319),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_320),
.Y(n_321)
);

OAI321xp33_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_312),
.A3(n_318),
.B1(n_306),
.B2(n_307),
.C(n_317),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_8),
.C(n_9),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_8),
.Y(n_324)
);


endmodule