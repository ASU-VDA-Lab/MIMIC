module fake_jpeg_30850_n_508 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_508);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_508;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_6),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_53),
.Y(n_137)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_54),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_9),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_55),
.B(n_59),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_48),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_56),
.B(n_58),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_57),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_48),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_31),
.B(n_9),
.Y(n_59)
);

HAxp5_ASAP7_75t_SL g60 ( 
.A(n_28),
.B(n_16),
.CON(n_60),
.SN(n_60)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_60),
.B(n_71),
.Y(n_121)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_62),
.Y(n_117)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_64),
.Y(n_153)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_72),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_69),
.Y(n_156)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_70),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_17),
.B(n_7),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_42),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_18),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_74),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_17),
.B(n_7),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_75),
.B(n_87),
.Y(n_149)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_38),
.B(n_7),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_77),
.B(n_81),
.Y(n_125)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_78),
.Y(n_124)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_80),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_29),
.B(n_6),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_82),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_83),
.Y(n_151)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_19),
.B(n_10),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_33),
.Y(n_88)
);

INVx4_ASAP7_75t_SL g112 ( 
.A(n_88),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_90),
.Y(n_130)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_91),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_92),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_94),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_20),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_96),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_19),
.B(n_10),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_33),
.Y(n_97)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_97),
.Y(n_138)
);

INVx3_ASAP7_75t_SL g98 ( 
.A(n_43),
.Y(n_98)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_57),
.A2(n_100),
.B1(n_99),
.B2(n_93),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_103),
.A2(n_123),
.B1(n_146),
.B2(n_65),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_74),
.A2(n_51),
.B1(n_49),
.B2(n_39),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_104),
.A2(n_140),
.B1(n_154),
.B2(n_155),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_53),
.A2(n_51),
.B1(n_49),
.B2(n_27),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_108),
.A2(n_113),
.B1(n_133),
.B2(n_142),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_68),
.A2(n_49),
.B1(n_21),
.B2(n_47),
.Y(n_113)
);

HAxp5_ASAP7_75t_SL g119 ( 
.A(n_60),
.B(n_20),
.CON(n_119),
.SN(n_119)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_119),
.B(n_40),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_80),
.A2(n_50),
.B1(n_25),
.B2(n_24),
.Y(n_123)
);

AOI21xp33_ASAP7_75t_SL g131 ( 
.A1(n_77),
.A2(n_23),
.B(n_30),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_131),
.B(n_40),
.C(n_20),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_89),
.A2(n_26),
.B1(n_47),
.B2(n_44),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_90),
.A2(n_47),
.B1(n_44),
.B2(n_23),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_92),
.A2(n_44),
.B1(n_24),
.B2(n_50),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_54),
.A2(n_25),
.B1(n_36),
.B2(n_46),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_81),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_29),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_98),
.A2(n_30),
.B1(n_23),
.B2(n_36),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_94),
.A2(n_30),
.B1(n_23),
.B2(n_35),
.Y(n_155)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_115),
.Y(n_158)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_158),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_105),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_159),
.B(n_169),
.Y(n_213)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_160),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_161),
.Y(n_230)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_115),
.Y(n_162)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_162),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_106),
.B(n_59),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_163),
.B(n_164),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_55),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_101),
.Y(n_165)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_110),
.Y(n_166)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_166),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_78),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_167),
.B(n_173),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_168),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_121),
.A2(n_86),
.B1(n_88),
.B2(n_52),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_170),
.A2(n_204),
.B1(n_157),
.B2(n_108),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_149),
.B(n_61),
.Y(n_171)
);

AOI21xp33_ASAP7_75t_L g243 ( 
.A1(n_171),
.A2(n_192),
.B(n_197),
.Y(n_243)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_141),
.Y(n_172)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_172),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_121),
.B(n_69),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_122),
.Y(n_174)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_174),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_178),
.Y(n_214)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_177),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_119),
.A2(n_91),
.B1(n_64),
.B2(n_76),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_129),
.A2(n_142),
.B(n_102),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_207),
.C(n_114),
.Y(n_210)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_109),
.Y(n_180)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_180),
.Y(n_252)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_118),
.Y(n_181)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_181),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_129),
.B(n_63),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_182),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_117),
.B(n_147),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_183),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_73),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_184),
.Y(n_246)
);

INVx3_ASAP7_75t_SL g185 ( 
.A(n_137),
.Y(n_185)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_185),
.Y(n_248)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_107),
.Y(n_186)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_186),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_152),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_187),
.A2(n_198),
.B1(n_199),
.B2(n_201),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_188),
.A2(n_202),
.B1(n_208),
.B2(n_148),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_114),
.A2(n_70),
.B1(n_84),
.B2(n_79),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_189),
.A2(n_205),
.B1(n_206),
.B2(n_0),
.Y(n_240)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_193),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_156),
.B(n_46),
.Y(n_191)
);

OAI32xp33_ASAP7_75t_L g241 ( 
.A1(n_191),
.A2(n_200),
.A3(n_11),
.B1(n_1),
.B2(n_2),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_116),
.B(n_85),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_112),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_112),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_194),
.B(n_195),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_SL g245 ( 
.A(n_196),
.B(n_2),
.C(n_3),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_126),
.B(n_83),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_154),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_152),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_135),
.B(n_83),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_127),
.Y(n_201)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_143),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_203),
.A2(n_67),
.B1(n_13),
.B2(n_12),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_144),
.A2(n_12),
.B1(n_15),
.B2(n_14),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_127),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_139),
.B(n_82),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_113),
.B(n_40),
.Y(n_207)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_143),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_198),
.A2(n_148),
.B1(n_111),
.B2(n_137),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_209),
.A2(n_218),
.B1(n_224),
.B2(n_225),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_210),
.B(n_233),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_212),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_176),
.A2(n_130),
.B1(n_120),
.B2(n_134),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_220),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_207),
.A2(n_111),
.B1(n_145),
.B2(n_136),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_221),
.A2(n_222),
.B1(n_227),
.B2(n_228),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_207),
.A2(n_133),
.B1(n_107),
.B2(n_134),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_167),
.A2(n_104),
.B1(n_140),
.B2(n_155),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_157),
.A2(n_128),
.B1(n_132),
.B2(n_120),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_196),
.A2(n_128),
.B1(n_132),
.B2(n_139),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_196),
.A2(n_12),
.B1(n_15),
.B2(n_14),
.Y(n_228)
);

AOI32xp33_ASAP7_75t_L g233 ( 
.A1(n_195),
.A2(n_82),
.A3(n_67),
.B1(n_30),
.B2(n_40),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_234),
.A2(n_185),
.B1(n_205),
.B2(n_201),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_163),
.B(n_0),
.C(n_1),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_236),
.B(n_228),
.C(n_247),
.Y(n_269)
);

AOI22x1_ASAP7_75t_L g238 ( 
.A1(n_178),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_238),
.A2(n_194),
.B1(n_193),
.B2(n_185),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_240),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_204),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_160),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_242),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_245),
.B(n_3),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_173),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_247),
.A2(n_186),
.B1(n_188),
.B2(n_190),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_235),
.A2(n_214),
.B(n_250),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_254),
.A2(n_245),
.B(n_236),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_255),
.A2(n_293),
.B1(n_248),
.B2(n_251),
.Y(n_296)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_215),
.Y(n_256)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_256),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_232),
.B(n_164),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_258),
.B(n_262),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_259),
.A2(n_248),
.B1(n_237),
.B2(n_217),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_230),
.Y(n_261)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_261),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_230),
.Y(n_263)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_263),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_229),
.B(n_171),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_264),
.B(n_272),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_235),
.B(n_170),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_265),
.B(n_270),
.C(n_275),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_219),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_266),
.B(n_279),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_269),
.B(n_278),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_179),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_218),
.A2(n_166),
.B1(n_165),
.B2(n_177),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_271),
.A2(n_285),
.B1(n_286),
.B2(n_291),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_232),
.B(n_191),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_215),
.Y(n_273)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_273),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_224),
.A2(n_187),
.B1(n_199),
.B2(n_159),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_274),
.A2(n_217),
.B(n_221),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_200),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_211),
.Y(n_276)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_276),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_219),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_216),
.Y(n_280)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_280),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_219),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_282),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_229),
.B(n_181),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_283),
.B(n_287),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_225),
.A2(n_180),
.B1(n_174),
.B2(n_208),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_214),
.A2(n_246),
.B1(n_222),
.B2(n_210),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_246),
.B(n_168),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_213),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_289),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_244),
.B(n_188),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_216),
.Y(n_290)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_290),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_214),
.A2(n_202),
.B1(n_168),
.B2(n_186),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_227),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_294),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_244),
.B(n_172),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_296),
.A2(n_285),
.B1(n_259),
.B2(n_291),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_302),
.A2(n_284),
.B(n_287),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_304),
.A2(n_318),
.B1(n_319),
.B2(n_321),
.Y(n_348)
);

AO22x1_ASAP7_75t_SL g305 ( 
.A1(n_257),
.A2(n_241),
.B1(n_238),
.B2(n_223),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_305),
.B(n_329),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_306),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_254),
.B(n_233),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_312),
.B(n_324),
.C(n_325),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_260),
.A2(n_238),
.B(n_223),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_314),
.A2(n_327),
.B(n_255),
.Y(n_359)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_256),
.Y(n_316)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_316),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_264),
.B(n_237),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_317),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_257),
.A2(n_243),
.B1(n_251),
.B2(n_239),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_267),
.A2(n_271),
.B1(n_262),
.B2(n_286),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_273),
.Y(n_320)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_320),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_267),
.A2(n_239),
.B1(n_211),
.B2(n_249),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_280),
.Y(n_323)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_323),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_275),
.B(n_226),
.C(n_231),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_270),
.B(n_226),
.C(n_231),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_260),
.A2(n_253),
.B(n_169),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_258),
.B(n_252),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_328),
.B(n_330),
.C(n_331),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_292),
.A2(n_252),
.B1(n_249),
.B2(n_253),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_272),
.B(n_158),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_265),
.B(n_161),
.C(n_162),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_302),
.A2(n_274),
.B1(n_277),
.B2(n_268),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_333),
.A2(n_339),
.B1(n_300),
.B2(n_318),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_326),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_335),
.B(n_336),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_322),
.B(n_279),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_311),
.B(n_283),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_338),
.B(n_345),
.C(n_351),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_313),
.B(n_290),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_340),
.B(n_346),
.Y(n_382)
);

NAND2x1_ASAP7_75t_SL g384 ( 
.A(n_343),
.B(n_362),
.Y(n_384)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_295),
.Y(n_344)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_344),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_311),
.B(n_269),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_295),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_303),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_347),
.B(n_349),
.Y(n_389)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_303),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_301),
.B(n_294),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_313),
.B(n_266),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_352),
.Y(n_388)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_308),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_353),
.B(n_357),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_326),
.B(n_282),
.Y(n_355)
);

XNOR2x2_ASAP7_75t_SL g391 ( 
.A(n_355),
.B(n_359),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_310),
.B(n_289),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_308),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_358),
.B(n_361),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_301),
.B(n_278),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_360),
.B(n_324),
.C(n_327),
.Y(n_375)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_315),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_299),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_332),
.Y(n_363)
);

INVxp33_ASAP7_75t_SL g368 ( 
.A(n_363),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_298),
.B(n_281),
.Y(n_365)
);

FAx1_ASAP7_75t_SL g392 ( 
.A(n_365),
.B(n_281),
.CI(n_321),
.CON(n_392),
.SN(n_392)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_369),
.A2(n_394),
.B1(n_355),
.B2(n_361),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_345),
.B(n_312),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_371),
.B(n_376),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_354),
.A2(n_298),
.B1(n_296),
.B2(n_309),
.Y(n_372)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_372),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_359),
.A2(n_331),
.B(n_325),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_374),
.A2(n_371),
.B(n_385),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_375),
.B(n_337),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_360),
.B(n_328),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_351),
.B(n_338),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_377),
.B(n_352),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_350),
.A2(n_333),
.B(n_336),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_378),
.B(n_379),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_362),
.B(n_314),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_356),
.B(n_319),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_380),
.B(n_385),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_365),
.A2(n_305),
.B1(n_323),
.B2(n_315),
.Y(n_381)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_381),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_356),
.B(n_330),
.C(n_306),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_383),
.B(n_341),
.C(n_349),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_364),
.B(n_300),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_364),
.B(n_278),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_387),
.B(n_337),
.Y(n_419)
);

AOI22x1_ASAP7_75t_L g390 ( 
.A1(n_334),
.A2(n_305),
.B1(n_297),
.B2(n_332),
.Y(n_390)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_390),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_392),
.B(n_348),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_SL g393 ( 
.A(n_343),
.B(n_261),
.C(n_263),
.Y(n_393)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_393),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_339),
.A2(n_293),
.B1(n_316),
.B2(n_320),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_334),
.A2(n_297),
.B1(n_307),
.B2(n_261),
.Y(n_395)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_395),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_368),
.Y(n_396)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_396),
.Y(n_424)
);

XNOR2x1_ASAP7_75t_L g425 ( 
.A(n_397),
.B(n_416),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_386),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_399),
.B(n_373),
.Y(n_432)
);

NOR2x1_ASAP7_75t_L g401 ( 
.A(n_373),
.B(n_357),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_401),
.B(n_404),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_384),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_367),
.Y(n_405)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_405),
.Y(n_427)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_386),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g430 ( 
.A(n_408),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_409),
.B(n_415),
.Y(n_434)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_386),
.Y(n_410)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_410),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_412),
.B(n_418),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_369),
.A2(n_348),
.B1(n_335),
.B2(n_340),
.Y(n_413)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_413),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_376),
.B(n_357),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_388),
.A2(n_341),
.B1(n_358),
.B2(n_353),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_417),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_419),
.B(n_366),
.Y(n_438)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_389),
.Y(n_420)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_420),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_421),
.B(n_383),
.C(n_366),
.Y(n_431)
);

XOR2x2_ASAP7_75t_L g422 ( 
.A(n_418),
.B(n_391),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_422),
.B(n_416),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_398),
.A2(n_394),
.B1(n_374),
.B2(n_390),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_426),
.A2(n_428),
.B1(n_441),
.B2(n_400),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_402),
.A2(n_382),
.B1(n_391),
.B2(n_370),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_404),
.A2(n_384),
.B(n_373),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_429),
.B(n_437),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_431),
.B(n_406),
.C(n_407),
.Y(n_451)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_432),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_411),
.A2(n_390),
.B(n_392),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_438),
.B(n_442),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_405),
.A2(n_344),
.B1(n_347),
.B2(n_346),
.Y(n_441)
);

A2O1A1O1Ixp25_ASAP7_75t_L g442 ( 
.A1(n_403),
.A2(n_380),
.B(n_377),
.C(n_375),
.D(n_392),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_440),
.B(n_401),
.Y(n_443)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_443),
.Y(n_469)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_427),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_446),
.B(n_454),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_423),
.B(n_406),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_447),
.B(n_448),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_438),
.B(n_407),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_450),
.B(n_451),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_431),
.B(n_421),
.C(n_412),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_452),
.B(n_453),
.C(n_455),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_423),
.B(n_419),
.C(n_414),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_425),
.B(n_397),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_440),
.A2(n_403),
.B1(n_415),
.B2(n_410),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_456),
.B(n_458),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_422),
.B(n_387),
.C(n_408),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_457),
.B(n_459),
.Y(n_464)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_435),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_436),
.B(n_409),
.C(n_342),
.Y(n_459)
);

BUFx24_ASAP7_75t_SL g460 ( 
.A(n_444),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_460),
.B(n_466),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_449),
.A2(n_437),
.B(n_433),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_462),
.A2(n_470),
.B(n_472),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_452),
.A2(n_433),
.B(n_429),
.Y(n_465)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_465),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_451),
.B(n_424),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_457),
.A2(n_430),
.B1(n_426),
.B2(n_439),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_467),
.B(n_455),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_459),
.A2(n_430),
.B(n_439),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_453),
.A2(n_434),
.B(n_442),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_445),
.A2(n_434),
.B(n_425),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_474),
.B(n_307),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_462),
.B(n_445),
.Y(n_475)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_475),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_476),
.B(n_483),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_467),
.A2(n_342),
.B(n_447),
.Y(n_477)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_477),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_478),
.B(n_480),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_461),
.A2(n_464),
.B(n_468),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_479),
.B(n_473),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_468),
.B(n_363),
.C(n_263),
.Y(n_480)
);

OR2x2_ASAP7_75t_L g481 ( 
.A(n_469),
.B(n_363),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_481),
.A2(n_471),
.B1(n_463),
.B2(n_473),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_472),
.A2(n_276),
.B1(n_161),
.B2(n_5),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_470),
.B(n_161),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_486),
.B(n_5),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_488),
.A2(n_489),
.B(n_494),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_491),
.B(n_493),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_480),
.B(n_3),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_482),
.B(n_4),
.Y(n_494)
);

MAJx2_ASAP7_75t_L g496 ( 
.A(n_492),
.B(n_484),
.C(n_485),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_496),
.B(n_476),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_487),
.A2(n_485),
.B(n_481),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_497),
.A2(n_498),
.B(n_477),
.Y(n_502)
);

INVxp33_ASAP7_75t_L g498 ( 
.A(n_495),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g505 ( 
.A(n_501),
.B(n_503),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_502),
.A2(n_490),
.B1(n_494),
.B2(n_483),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_499),
.B(n_495),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_504),
.B(n_490),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_506),
.B(n_505),
.C(n_486),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_507),
.B(n_500),
.Y(n_508)
);


endmodule