module real_jpeg_25361_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_173;
wire n_40;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_0),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_0),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_0),
.B(n_46),
.Y(n_61)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_2),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_2),
.B(n_25),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_2),
.B(n_42),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_2),
.B(n_27),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_2),
.B(n_105),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_3),
.B(n_30),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_3),
.B(n_63),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_3),
.B(n_25),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_3),
.B(n_42),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_3),
.B(n_27),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_4),
.B(n_27),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_4),
.B(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_4),
.B(n_38),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_5),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_8),
.B(n_25),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_8),
.B(n_30),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_8),
.B(n_63),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_8),
.B(n_42),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_8),
.B(n_46),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_8),
.B(n_27),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_8),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_9),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_9),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_9),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_9),
.B(n_27),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_9),
.B(n_46),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_9),
.B(n_158),
.Y(n_157)
);

INVx8_ASAP7_75t_SL g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_12),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_13),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_13),
.B(n_63),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_13),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_13),
.B(n_25),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_13),
.B(n_42),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_13),
.B(n_46),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_13),
.B(n_27),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_13),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_14),
.B(n_80),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_14),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_16),
.Y(n_106)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_16),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_125),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_110),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_73),
.B2(n_109),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_48),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_32),
.C(n_40),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_23),
.B(n_123),
.Y(n_122)
);

BUFx24_ASAP7_75t_SL g202 ( 
.A(n_23),
.Y(n_202)
);

FAx1_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_26),
.CI(n_29),
.CON(n_23),
.SN(n_23)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_24),
.B(n_26),
.C(n_29),
.Y(n_96)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_27),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_32),
.A2(n_33),
.B1(n_40),
.B2(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_34),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_40),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_44),
.C(n_45),
.Y(n_40)
);

FAx1_ASAP7_75t_SL g115 ( 
.A(n_41),
.B(n_44),
.CI(n_45),
.CON(n_115),
.SN(n_115)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx13_ASAP7_75t_L g179 ( 
.A(n_46),
.Y(n_179)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_58),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_56),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_67),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_66),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_62),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_71),
.C(n_72),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_69),
.B(n_179),
.Y(n_178)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_72),
.Y(n_76)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_94),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_77),
.C(n_83),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_75),
.A2(n_77),
.B1(n_78),
.B2(n_113),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_75),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_81),
.B(n_82),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_81),
.Y(n_82)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_80),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_96),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_83),
.B(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_90),
.C(n_92),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_84),
.A2(n_85),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_86),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_147)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_90),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_107),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_114),
.C(n_121),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_111),
.B(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_114),
.A2(n_121),
.B1(n_122),
.B2(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_114),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.C(n_120),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_115),
.B(n_192),
.Y(n_191)
);

BUFx24_ASAP7_75t_SL g203 ( 
.A(n_115),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_116),
.B(n_120),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.C(n_119),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_119),
.Y(n_138)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_198),
.C(n_199),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_189),
.C(n_190),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_148),
.C(n_161),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_139),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_137),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_130),
.B(n_137),
.C(n_139),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.C(n_135),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_131),
.A2(n_132),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_133),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_145),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_140),
.B(n_146),
.C(n_147),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_143),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_160)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.C(n_160),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_149),
.B(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_152),
.A2(n_153),
.B1(n_160),
.B2(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_154),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_159),
.Y(n_173)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_185),
.C(n_186),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_170),
.C(n_176),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_168),
.C(n_169),
.Y(n_185)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_174),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_171),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.C(n_180),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_194),
.C(n_197),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);


endmodule