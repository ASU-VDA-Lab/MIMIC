module real_jpeg_6968_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g163 ( 
.A(n_0),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_0),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_0),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_0),
.Y(n_278)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_0),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_0),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_1),
.A2(n_197),
.B1(n_199),
.B2(n_200),
.Y(n_196)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_1),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_1),
.A2(n_122),
.B1(n_199),
.B2(n_269),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_SL g384 ( 
.A1(n_1),
.A2(n_199),
.B1(n_280),
.B2(n_385),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_SL g445 ( 
.A1(n_1),
.A2(n_199),
.B1(n_446),
.B2(n_448),
.Y(n_445)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_2),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_2),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_2),
.Y(n_185)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_2),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_2),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_3),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_3),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_3),
.A2(n_89),
.B1(n_116),
.B2(n_118),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_3),
.A2(n_89),
.B1(n_131),
.B2(n_133),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_3),
.A2(n_89),
.B1(n_280),
.B2(n_282),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_4),
.A2(n_33),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_4),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_4),
.A2(n_184),
.B1(n_253),
.B2(n_255),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g396 ( 
.A1(n_4),
.A2(n_184),
.B1(n_397),
.B2(n_398),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_4),
.A2(n_184),
.B1(n_419),
.B2(n_422),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_5),
.Y(n_526)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_7),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_8),
.Y(n_100)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_8),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_8),
.Y(n_379)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_9),
.Y(n_74)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_10),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_10),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_10),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_11),
.A2(n_212),
.B1(n_214),
.B2(n_217),
.Y(n_211)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_11),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_11),
.A2(n_217),
.B1(n_255),
.B2(n_266),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g299 ( 
.A1(n_11),
.A2(n_176),
.B1(n_217),
.B2(n_300),
.Y(n_299)
);

OAI22xp33_ASAP7_75t_L g359 ( 
.A1(n_11),
.A2(n_217),
.B1(n_360),
.B2(n_361),
.Y(n_359)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_13),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g372 ( 
.A1(n_13),
.A2(n_157),
.B1(n_214),
.B2(n_373),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_13),
.B(n_379),
.C(n_380),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_13),
.B(n_70),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_13),
.B(n_413),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_13),
.B(n_114),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_13),
.B(n_207),
.Y(n_453)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_14),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_52)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_14),
.A2(n_55),
.B1(n_175),
.B2(n_177),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_14),
.A2(n_55),
.B1(n_213),
.B2(n_221),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_14),
.A2(n_55),
.B1(n_343),
.B2(n_344),
.Y(n_342)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_16),
.A2(n_45),
.B1(n_47),
.B2(n_49),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_16),
.A2(n_49),
.B1(n_164),
.B2(n_169),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_16),
.A2(n_49),
.B1(n_220),
.B2(n_225),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_16),
.A2(n_49),
.B1(n_204),
.B2(n_317),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_17),
.A2(n_80),
.B1(n_82),
.B2(n_84),
.Y(n_79)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_17),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_17),
.A2(n_84),
.B1(n_121),
.B2(n_125),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_17),
.A2(n_84),
.B1(n_164),
.B2(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_17),
.A2(n_84),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_18),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_18),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_18),
.A2(n_188),
.B1(n_204),
.B2(n_206),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_18),
.A2(n_188),
.B1(n_240),
.B2(n_242),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g391 ( 
.A1(n_18),
.A2(n_188),
.B1(n_301),
.B2(n_392),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_522),
.B(n_524),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_136),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_134),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_129),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_23),
.B(n_129),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_119),
.C(n_126),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_24),
.A2(n_25),
.B1(n_518),
.B2(n_519),
.Y(n_517)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_56),
.C(n_90),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g509 ( 
.A(n_26),
.B(n_510),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_44),
.B1(n_50),
.B2(n_52),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_27),
.A2(n_50),
.B1(n_52),
.B2(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_27),
.A2(n_50),
.B1(n_120),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_27),
.A2(n_37),
.B1(n_183),
.B2(n_268),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_27),
.A2(n_250),
.B(n_268),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_27),
.A2(n_44),
.B1(n_50),
.B2(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_28),
.B(n_187),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_28),
.A2(n_245),
.B(n_249),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_37),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_32),
.Y(n_151)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_33),
.Y(n_133)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_33),
.Y(n_189)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_34),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_34),
.B(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_38),
.B1(n_39),
.B2(n_42),
.Y(n_37)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_37),
.B(n_157),
.Y(n_305)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_41),
.Y(n_147)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_41),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_43),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_43),
.Y(n_201)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_43),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_43),
.Y(n_319)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_50),
.A2(n_183),
.B(n_186),
.Y(n_182)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_51),
.B(n_187),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_51),
.B(n_359),
.Y(n_358)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_53),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_56),
.A2(n_90),
.B1(n_91),
.B2(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_56),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_79),
.B1(n_85),
.B2(n_86),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g127 ( 
.A(n_57),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_57),
.A2(n_85),
.B1(n_196),
.B2(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_57),
.A2(n_85),
.B1(n_265),
.B2(n_316),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_57),
.A2(n_79),
.B1(n_85),
.B2(n_499),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_70),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_62),
.Y(n_459)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_64),
.Y(n_207)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_65),
.Y(n_347)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_68),
.Y(n_343)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_69),
.Y(n_198)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_69),
.Y(n_254)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_70),
.A2(n_127),
.B(n_128),
.Y(n_126)
);

AOI22x1_ASAP7_75t_L g262 ( 
.A1(n_70),
.A2(n_127),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_70),
.A2(n_127),
.B1(n_341),
.B2(n_342),
.Y(n_340)
);

AO22x2_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_73),
.B1(n_75),
.B2(n_77),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_73),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_74),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_74),
.Y(n_241)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_74),
.Y(n_399)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_74),
.Y(n_462)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_95),
.B1(n_98),
.B2(n_101),
.Y(n_94)
);

INVx11_ASAP7_75t_L g397 ( 
.A(n_75),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_76),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_76),
.Y(n_228)
);

INVx4_ASAP7_75t_L g463 ( 
.A(n_77),
.Y(n_463)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_80),
.Y(n_255)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_85),
.B(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_85),
.A2(n_252),
.B(n_297),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_90),
.A2(n_91),
.B1(n_497),
.B2(n_498),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_90),
.B(n_494),
.C(n_497),
.Y(n_505)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_113),
.B(n_115),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_92),
.A2(n_113),
.B1(n_211),
.B2(n_218),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_92),
.A2(n_372),
.B(n_374),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_92),
.A2(n_113),
.B1(n_396),
.B2(n_445),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_92),
.A2(n_374),
.B(n_445),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_93),
.B(n_239),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_93),
.A2(n_114),
.B1(n_219),
.B2(n_274),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_93),
.A2(n_114),
.B1(n_274),
.B2(n_324),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_93),
.A2(n_114),
.B1(n_324),
.B2(n_350),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_104),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_104),
.A2(n_238),
.B(n_396),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_110),
.B2(n_112),
.Y(n_104)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_107),
.Y(n_176)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_108),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_109),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_109),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_111),
.Y(n_281)
);

BUFx5_ASAP7_75t_L g423 ( 
.A(n_111),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_113),
.A2(n_211),
.B(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_114),
.B(n_239),
.Y(n_374)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_115),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_117),
.Y(n_327)
);

INVx5_ASAP7_75t_L g447 ( 
.A(n_117),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_119),
.B(n_126),
.Y(n_519)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_124),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_127),
.A2(n_195),
.B(n_202),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_127),
.B(n_263),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_127),
.A2(n_202),
.B(n_451),
.Y(n_450)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_516),
.B(n_521),
.Y(n_136)
);

AOI21x1_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_488),
.B(n_513),
.Y(n_137)
);

OAI311xp33_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_309),
.A3(n_365),
.B1(n_482),
.C1(n_487),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_287),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_141),
.A2(n_484),
.B(n_485),
.Y(n_483)
);

NOR2x1_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_256),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_142),
.B(n_256),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_208),
.C(n_236),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_143),
.B(n_307),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_180),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_144),
.B(n_181),
.C(n_194),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_158),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_145),
.A2(n_158),
.B1(n_159),
.B2(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_145),
.Y(n_294)
);

OAI32xp33_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_148),
.A3(n_149),
.B1(n_152),
.B2(n_156),
.Y(n_145)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_150),
.B(n_153),
.Y(n_152)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_SL g245 ( 
.A1(n_156),
.A2(n_157),
.B(n_246),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_157),
.A2(n_160),
.B(n_388),
.Y(n_415)
);

OAI21xp33_ASAP7_75t_SL g451 ( 
.A1(n_157),
.A2(n_317),
.B(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_167),
.B1(n_170),
.B2(n_173),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_160),
.A2(n_231),
.B1(n_276),
.B2(n_279),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_160),
.A2(n_279),
.B(n_329),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_160),
.A2(n_384),
.B(n_388),
.Y(n_383)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_161),
.A2(n_174),
.B1(n_230),
.B2(n_234),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_161),
.A2(n_168),
.B1(n_299),
.B2(n_304),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_161),
.B(n_391),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_161),
.A2(n_432),
.B1(n_433),
.B2(n_434),
.Y(n_431)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_163),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_163),
.Y(n_414)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_163),
.Y(n_426)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_165),
.Y(n_169)
);

BUFx8_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g284 ( 
.A(n_166),
.Y(n_284)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_166),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_166),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_179),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_193),
.B2(n_194),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_185),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_186),
.B(n_358),
.Y(n_357)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_203),
.Y(n_263)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_208),
.A2(n_209),
.B1(n_236),
.B2(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_229),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_210),
.B(n_229),
.Y(n_260)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx4_ASAP7_75t_SL g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_224),
.Y(n_377)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_228),
.Y(n_373)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_232),
.Y(n_392)
);

INVx8_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_233),
.Y(n_381)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_236),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_243),
.C(n_251),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_237),
.B(n_251),
.Y(n_290)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

AOI32xp33_ASAP7_75t_L g457 ( 
.A1(n_241),
.A2(n_255),
.A3(n_453),
.B1(n_458),
.B2(n_460),
.Y(n_457)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_242),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_243),
.A2(n_244),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_257),
.B(n_272),
.C(n_285),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_272),
.B1(n_285),
.B2(n_286),
.Y(n_258)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_259),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_260),
.B(n_262),
.C(n_271),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_267),
.B1(n_270),
.B2(n_271),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_262),
.Y(n_270)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_267),
.Y(n_271)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_275),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_273),
.B(n_275),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_306),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_288),
.B(n_306),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_292),
.C(n_295),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_289),
.B(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_290),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_292),
.A2(n_293),
.B1(n_295),
.B2(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_295),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_298),
.C(n_305),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g472 ( 
.A(n_296),
.B(n_473),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_298),
.B(n_305),
.Y(n_473)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_299),
.Y(n_456)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx4_ASAP7_75t_SL g301 ( 
.A(n_302),
.Y(n_301)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NAND2xp33_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_362),
.Y(n_309)
);

A2O1A1Ixp33_ASAP7_75t_SL g482 ( 
.A1(n_310),
.A2(n_362),
.B(n_483),
.C(n_486),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_334),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_311),
.B(n_334),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_321),
.C(n_333),
.Y(n_311)
);

FAx1_ASAP7_75t_SL g364 ( 
.A(n_312),
.B(n_321),
.CI(n_333),
.CON(n_364),
.SN(n_364)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_313),
.B(n_315),
.C(n_320),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_320),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_316),
.Y(n_341)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_322),
.A2(n_323),
.B1(n_328),
.B2(n_332),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_323),
.B(n_328),
.Y(n_354)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_328),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_328),
.A2(n_332),
.B1(n_356),
.B2(n_357),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_328),
.A2(n_354),
.B(n_357),
.Y(n_491)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_335),
.B(n_338),
.C(n_352),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_338),
.B1(n_352),
.B2(n_353),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_348),
.B(n_351),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_340),
.B(n_349),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_342),
.Y(n_499)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

FAx1_ASAP7_75t_SL g490 ( 
.A(n_351),
.B(n_491),
.CI(n_492),
.CON(n_490),
.SN(n_490)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_351),
.B(n_491),
.C(n_492),
.Y(n_512)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_355),
.Y(n_353)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_359),
.Y(n_495)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_360),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_364),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_363),
.B(n_364),
.Y(n_486)
);

BUFx24_ASAP7_75t_SL g528 ( 
.A(n_364),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_366),
.A2(n_476),
.B(n_481),
.Y(n_365)
);

AO21x1_ASAP7_75t_SL g366 ( 
.A1(n_367),
.A2(n_465),
.B(n_475),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_368),
.A2(n_439),
.B(n_464),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_369),
.A2(n_402),
.B(n_438),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_382),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_370),
.B(n_382),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_371),
.B(n_375),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_371),
.A2(n_375),
.B1(n_376),
.B2(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_371),
.Y(n_436)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_378),
.Y(n_376)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_393),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_383),
.B(n_394),
.C(n_401),
.Y(n_440)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_384),
.Y(n_433)
);

INVx6_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx4_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_391),
.Y(n_388)
);

INVx4_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_394),
.A2(n_395),
.B1(n_400),
.B2(n_401),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_397),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_403),
.A2(n_430),
.B(n_437),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_404),
.A2(n_416),
.B(n_429),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_415),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_412),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_413),
.Y(n_434)
);

INVx8_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_417),
.B(n_428),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_417),
.B(n_428),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_418),
.A2(n_424),
.B(n_427),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_418),
.Y(n_432)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx5_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx5_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_426),
.A2(n_427),
.B(n_456),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_435),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_431),
.B(n_435),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_441),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_440),
.B(n_441),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_454),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_443),
.A2(n_444),
.B1(n_449),
.B2(n_450),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_444),
.B(n_449),
.C(n_454),
.Y(n_466)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVxp33_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_457),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_455),
.B(n_457),
.Y(n_471)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

NAND2xp33_ASAP7_75t_SL g460 ( 
.A(n_461),
.B(n_463),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_467),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_466),
.B(n_467),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_468),
.A2(n_469),
.B1(n_472),
.B2(n_474),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_SL g469 ( 
.A(n_470),
.B(n_471),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_470),
.B(n_471),
.C(n_474),
.Y(n_477)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_472),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_478),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_477),
.B(n_478),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_502),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_490),
.B(n_501),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_490),
.B(n_501),
.Y(n_514)
);

BUFx24_ASAP7_75t_SL g527 ( 
.A(n_490),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_493),
.A2(n_494),
.B1(n_496),
.B2(n_500),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_493),
.A2(n_494),
.B1(n_508),
.B2(n_509),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_493),
.B(n_504),
.C(n_508),
.Y(n_520)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_496),
.Y(n_500)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_502),
.A2(n_514),
.B(n_515),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_503),
.B(n_512),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_503),
.B(n_512),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_504),
.A2(n_505),
.B1(n_506),
.B2(n_507),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_520),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_517),
.B(n_520),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_519),
.Y(n_518)
);

INVx6_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx6_ASAP7_75t_L g525 ( 
.A(n_523),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_525),
.B(n_526),
.Y(n_524)
);


endmodule