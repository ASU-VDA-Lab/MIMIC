module fake_jpeg_10900_n_91 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_91);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_91;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_19),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_46),
.Y(n_52)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_43),
.Y(n_50)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_45),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_39),
.Y(n_53)
);

OR2x2_ASAP7_75t_SL g48 ( 
.A(n_42),
.B(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_48),
.B(n_51),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_47),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_4),
.Y(n_65)
);

AND2x4_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_0),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_3),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_38),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_17),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_35),
.B(n_33),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_59),
.A2(n_64),
.B(n_5),
.Y(n_78)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_52),
.A2(n_1),
.B(n_2),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_7),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_58),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_62),
.A2(n_56),
.B1(n_5),
.B2(n_8),
.Y(n_74)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_65),
.B(n_70),
.Y(n_73)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_69),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_4),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_75),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_59),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_79),
.C(n_64),
.Y(n_80)
);

OA21x2_ASAP7_75t_SL g84 ( 
.A1(n_80),
.A2(n_82),
.B(n_77),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_68),
.C(n_60),
.Y(n_82)
);

AOI221xp5_ASAP7_75t_L g83 ( 
.A1(n_81),
.A2(n_71),
.B1(n_79),
.B2(n_62),
.C(n_72),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_84),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_85),
.A2(n_76),
.B1(n_10),
.B2(n_13),
.Y(n_86)
);

AOI222xp33_ASAP7_75t_SL g87 ( 
.A1(n_86),
.A2(n_9),
.B1(n_14),
.B2(n_18),
.C1(n_20),
.C2(n_21),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_22),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_SL g90 ( 
.A1(n_89),
.A2(n_76),
.B(n_24),
.C(n_26),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_90),
.A2(n_23),
.B(n_29),
.Y(n_91)
);


endmodule