module fake_jpeg_24523_n_291 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_291);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_291;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx8_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_3),
.B(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_38),
.B(n_42),
.Y(n_68)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_39),
.B(n_41),
.Y(n_66)
);

NOR2xp67_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_0),
.Y(n_40)
);

NOR2x1_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_20),
.Y(n_56)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_0),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_51),
.Y(n_84)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_27),
.B1(n_17),
.B2(n_25),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_48),
.B1(n_53),
.B2(n_62),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_17),
.B1(n_27),
.B2(n_20),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_49),
.Y(n_80)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_50),
.A2(n_60),
.B1(n_63),
.B2(n_43),
.Y(n_71)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

AO22x1_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_20),
.B1(n_22),
.B2(n_24),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_31),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_65),
.Y(n_74)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_59),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_56),
.A2(n_26),
.B(n_30),
.C(n_32),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_19),
.Y(n_58)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_43),
.A2(n_17),
.B1(n_27),
.B2(n_33),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_17),
.B1(n_31),
.B2(n_33),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_19),
.Y(n_64)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_31),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_14),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_23),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_56),
.A2(n_43),
.B1(n_41),
.B2(n_39),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_69),
.A2(n_83),
.B1(n_28),
.B2(n_32),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g114 ( 
.A(n_70),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_71),
.A2(n_92),
.B(n_72),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVxp33_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_79),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_54),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_41),
.C(n_39),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_47),
.C(n_51),
.Y(n_108)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_82),
.B(n_89),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_48),
.A2(n_18),
.B1(n_33),
.B2(n_32),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_67),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_44),
.B(n_30),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_90),
.Y(n_95)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_49),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_41),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_91),
.Y(n_96)
);

AO22x2_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_37),
.B1(n_35),
.B2(n_39),
.Y(n_92)
);

OA21x2_ASAP7_75t_L g117 ( 
.A1(n_92),
.A2(n_63),
.B(n_45),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_93),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_97),
.A2(n_104),
.B1(n_119),
.B2(n_92),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_90),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_101),
.Y(n_123)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_103),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_68),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_107),
.Y(n_143)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_111),
.Y(n_137)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_108),
.B(n_121),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_L g109 ( 
.A1(n_84),
.A2(n_7),
.B(n_13),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_109),
.A2(n_28),
.B(n_29),
.Y(n_138)
);

NOR3xp33_ASAP7_75t_SL g111 ( 
.A(n_92),
.B(n_68),
.C(n_30),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_112),
.B(n_82),
.Y(n_125)
);

AO22x1_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_92),
.B1(n_61),
.B2(n_57),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_79),
.B(n_59),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_49),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_86),
.B(n_0),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_120),
.A2(n_29),
.B(n_21),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_81),
.B(n_37),
.C(n_35),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_95),
.A2(n_84),
.B(n_87),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_122),
.A2(n_124),
.B(n_125),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_95),
.A2(n_87),
.B(n_73),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_128),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_99),
.A2(n_76),
.B1(n_73),
.B2(n_69),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_127),
.A2(n_104),
.B1(n_99),
.B2(n_106),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_131),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_76),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_114),
.A2(n_70),
.B1(n_92),
.B2(n_50),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_132),
.A2(n_134),
.B1(n_142),
.B2(n_72),
.Y(n_157)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_135),
.Y(n_162)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_115),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_141),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_138),
.B(n_149),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_102),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_139),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_70),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_145),
.Y(n_153)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_144),
.B(n_23),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_77),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_146),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_77),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_148),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_97),
.B(n_120),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_118),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_121),
.C(n_108),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_160),
.C(n_172),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_157),
.A2(n_163),
.B1(n_164),
.B2(n_167),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_129),
.B(n_75),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_158),
.B(n_18),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_140),
.A2(n_117),
.B(n_112),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_159),
.A2(n_134),
.B(n_141),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_148),
.C(n_123),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_168),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_131),
.A2(n_114),
.B1(n_117),
.B2(n_116),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_123),
.B(n_97),
.Y(n_165)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_165),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_132),
.A2(n_114),
.B1(n_117),
.B2(n_96),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_129),
.Y(n_168)
);

OAI32xp33_ASAP7_75t_L g169 ( 
.A1(n_127),
.A2(n_96),
.A3(n_120),
.B1(n_103),
.B2(n_100),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_180),
.Y(n_181)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_170),
.B(n_179),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_124),
.B(n_110),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_122),
.B(n_110),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_175),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_89),
.C(n_80),
.Y(n_175)
);

NOR2xp67_ASAP7_75t_R g189 ( 
.A(n_177),
.B(n_138),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_134),
.A2(n_147),
.B1(n_145),
.B2(n_137),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_178),
.A2(n_57),
.B1(n_61),
.B2(n_52),
.Y(n_196)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_125),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_133),
.B(n_80),
.C(n_75),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_136),
.Y(n_182)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_182),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_162),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_183),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_139),
.Y(n_184)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_186),
.A2(n_166),
.B(n_174),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_159),
.A2(n_137),
.B1(n_72),
.B2(n_78),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_187),
.A2(n_196),
.B1(n_200),
.B2(n_164),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_144),
.Y(n_188)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_188),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_177),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_176),
.Y(n_190)
);

NOR3xp33_ASAP7_75t_L g191 ( 
.A(n_154),
.B(n_18),
.C(n_29),
.Y(n_191)
);

AOI322xp5_ASAP7_75t_L g216 ( 
.A1(n_191),
.A2(n_194),
.A3(n_26),
.B1(n_151),
.B2(n_165),
.C1(n_170),
.C2(n_166),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_199),
.Y(n_212)
);

NOR3xp33_ASAP7_75t_L g194 ( 
.A(n_154),
.B(n_21),
.C(n_28),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_153),
.B(n_128),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_153),
.A2(n_52),
.B1(n_135),
.B2(n_21),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_171),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_202),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_179),
.B(n_1),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_155),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_205),
.Y(n_228)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_175),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_207),
.B(n_189),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_156),
.C(n_160),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_218),
.C(n_227),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_209),
.A2(n_221),
.B1(n_224),
.B2(n_226),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_203),
.A2(n_176),
.B1(n_174),
.B2(n_168),
.Y(n_211)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_217),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_203),
.A2(n_169),
.B1(n_180),
.B2(n_167),
.Y(n_215)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_215),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_216),
.B(n_201),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_172),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_173),
.C(n_178),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_163),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_225),
.Y(n_234)
);

AOI322xp5_ASAP7_75t_L g220 ( 
.A1(n_181),
.A2(n_35),
.A3(n_128),
.B1(n_26),
.B2(n_24),
.C1(n_23),
.C2(n_22),
.Y(n_220)
);

AOI21xp33_ASAP7_75t_L g231 ( 
.A1(n_220),
.A2(n_204),
.B(n_183),
.Y(n_231)
);

OAI31xp33_ASAP7_75t_L g221 ( 
.A1(n_181),
.A2(n_24),
.A3(n_23),
.B(n_3),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_187),
.A2(n_24),
.B1(n_35),
.B2(n_3),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_35),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_190),
.A2(n_1),
.B(n_2),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_2),
.C(n_3),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_L g229 ( 
.A1(n_223),
.A2(n_199),
.B1(n_197),
.B2(n_182),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_229),
.A2(n_236),
.B1(n_239),
.B2(n_224),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_231),
.A2(n_212),
.B(n_214),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_184),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_238),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_200),
.Y(n_235)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_235),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_210),
.A2(n_206),
.B1(n_228),
.B2(n_198),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_228),
.A2(n_198),
.B1(n_196),
.B2(n_188),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_207),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_197),
.C(n_185),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_243),
.C(n_212),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_185),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_246),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_244),
.A2(n_221),
.B1(n_209),
.B2(n_225),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_247),
.A2(n_254),
.B1(n_257),
.B2(n_8),
.Y(n_267)
);

OAI21xp33_ASAP7_75t_L g248 ( 
.A1(n_241),
.A2(n_226),
.B(n_213),
.Y(n_248)
);

NOR5xp2_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_237),
.C(n_238),
.D(n_233),
.E(n_234),
.Y(n_258)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_256),
.C(n_230),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_227),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_253),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_217),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_236),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_4),
.C(n_5),
.Y(n_256)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

AND2x2_ASAP7_75t_SL g273 ( 
.A(n_258),
.B(n_266),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_260),
.C(n_264),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_234),
.C(n_232),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_248),
.A2(n_11),
.B(n_6),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_4),
.C(n_7),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_7),
.Y(n_266)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_267),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_262),
.B(n_255),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_271),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_254),
.Y(n_270)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_270),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_266),
.B(n_247),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_265),
.B(n_251),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_272),
.A2(n_275),
.B(n_16),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_252),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_272),
.A2(n_259),
.B1(n_260),
.B2(n_252),
.Y(n_276)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_276),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_269),
.A2(n_12),
.B(n_13),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_277),
.A2(n_278),
.B(n_281),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_16),
.C(n_12),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_280),
.A2(n_273),
.B(n_279),
.Y(n_284)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_284),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_281),
.A2(n_274),
.B(n_13),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_286),
.C(n_283),
.Y(n_287)
);

AOI21xp33_ASAP7_75t_SL g286 ( 
.A1(n_276),
.A2(n_12),
.B(n_16),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_289),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_282),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_288),
.Y(n_291)
);


endmodule