module fake_jpeg_15882_n_121 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_121);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx4f_ASAP7_75t_SL g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_21),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx6f_ASAP7_75t_SL g50 ( 
.A(n_12),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_18),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_0),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_55),
.B(n_58),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_46),
.B(n_0),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_61),
.Y(n_68)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_48),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_59),
.A2(n_53),
.B1(n_49),
.B2(n_48),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_63),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_55),
.A2(n_53),
.B1(n_49),
.B2(n_45),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_54),
.B1(n_43),
.B2(n_40),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_51),
.B1(n_47),
.B2(n_44),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_60),
.A2(n_41),
.B1(n_42),
.B2(n_19),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_69),
.A2(n_74),
.B1(n_1),
.B2(n_4),
.Y(n_75)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_42),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_73),
.B(n_56),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_61),
.A2(n_42),
.B1(n_2),
.B2(n_3),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_81),
.Y(n_95)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_70),
.A2(n_56),
.B1(n_4),
.B2(n_5),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_77),
.A2(n_83),
.B1(n_86),
.B2(n_71),
.Y(n_91)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_85),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_62),
.B(n_6),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_84),
.B(n_88),
.Y(n_90)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_72),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_87),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_7),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_91),
.A2(n_98),
.B1(n_8),
.B2(n_10),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_62),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_92),
.B(n_93),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_65),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_25),
.B1(n_35),
.B2(n_32),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_95),
.A2(n_77),
.B(n_86),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_103),
.Y(n_108)
);

AND2x6_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_24),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_102),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_78),
.C(n_26),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_104),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_98),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_100),
.C(n_90),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_110),
.C(n_105),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_10),
.Y(n_110)
);

BUFx24_ASAP7_75t_SL g111 ( 
.A(n_106),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_108),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_112),
.B(n_113),
.Y(n_114)
);

NAND4xp25_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_107),
.C(n_13),
.D(n_15),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_28),
.B1(n_17),
.B2(n_20),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_30),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_97),
.C(n_22),
.Y(n_118)
);

AOI322xp5_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_27),
.A3(n_29),
.B1(n_38),
.B2(n_97),
.C1(n_11),
.C2(n_89),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_89),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_11),
.Y(n_121)
);


endmodule