module fake_ariane_1167_n_35 (n_8, n_3, n_2, n_7, n_5, n_1, n_0, n_6, n_9, n_4, n_35);

input n_8;
input n_3;
input n_2;
input n_7;
input n_5;
input n_1;
input n_0;
input n_6;
input n_9;
input n_4;

output n_35;

wire n_24;
wire n_22;
wire n_13;
wire n_27;
wire n_20;
wire n_29;
wire n_17;
wire n_18;
wire n_32;
wire n_28;
wire n_11;
wire n_34;
wire n_26;
wire n_14;
wire n_33;
wire n_19;
wire n_30;
wire n_31;
wire n_16;
wire n_12;
wire n_15;
wire n_21;
wire n_23;
wire n_10;
wire n_25;

NOR2xp33_ASAP7_75t_R g10 ( 
.A(n_8),
.B(n_1),
.Y(n_10)
);

INVx2_ASAP7_75t_SL g11 ( 
.A(n_6),
.Y(n_11)
);

NAND3xp33_ASAP7_75t_L g12 ( 
.A(n_7),
.B(n_6),
.C(n_5),
.Y(n_12)
);

AO21x2_ASAP7_75t_L g13 ( 
.A1(n_2),
.A2(n_1),
.B(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_4),
.B(n_0),
.Y(n_15)
);

OR2x2_ASAP7_75t_L g16 ( 
.A(n_5),
.B(n_9),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_R g17 ( 
.A(n_0),
.B(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_2),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_3),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_18),
.B(n_15),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_22),
.Y(n_24)
);

AO31x2_ASAP7_75t_L g25 ( 
.A1(n_21),
.A2(n_18),
.A3(n_13),
.B(n_12),
.Y(n_25)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_21),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_26),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_24),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_19),
.Y(n_30)
);

AOI221xp5_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_20),
.B1(n_23),
.B2(n_17),
.C(n_13),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_30),
.B1(n_16),
.B2(n_28),
.Y(n_34)
);

AOI222xp33_ASAP7_75t_L g35 ( 
.A1(n_34),
.A2(n_25),
.B1(n_33),
.B2(n_32),
.C1(n_31),
.C2(n_12),
.Y(n_35)
);


endmodule