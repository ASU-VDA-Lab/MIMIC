module fake_jpeg_25560_n_315 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_315);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_315;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_31),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_33),
.Y(n_47)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_12),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_47),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_32),
.A2(n_19),
.B1(n_22),
.B2(n_21),
.Y(n_42)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_29),
.B1(n_21),
.B2(n_19),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_33),
.A2(n_19),
.B1(n_16),
.B2(n_23),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_44),
.A2(n_16),
.B1(n_19),
.B2(n_18),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_56),
.Y(n_72)
);

AO22x2_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_28),
.B1(n_33),
.B2(n_16),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_61),
.B1(n_66),
.B2(n_21),
.Y(n_67)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_47),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_28),
.Y(n_80)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_34),
.Y(n_57)
);

NAND3xp33_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_37),
.C(n_41),
.Y(n_75)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_64),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_45),
.Y(n_66)
);

OAI22x1_ASAP7_75t_L g101 ( 
.A1(n_67),
.A2(n_56),
.B1(n_40),
.B2(n_64),
.Y(n_101)
);

OR2x6_ASAP7_75t_SL g69 ( 
.A(n_49),
.B(n_41),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_69),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_56),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_75),
.A2(n_37),
.B1(n_16),
.B2(n_60),
.Y(n_104)
);

CKINVDCx12_ASAP7_75t_R g78 ( 
.A(n_49),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_86),
.B(n_87),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_49),
.B1(n_66),
.B2(n_53),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_91),
.B(n_92),
.Y(n_119)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

MAJx2_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_48),
.C(n_57),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_31),
.C(n_30),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_68),
.Y(n_94)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_95),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_96),
.A2(n_107),
.B(n_8),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_58),
.Y(n_97)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_58),
.Y(n_98)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_73),
.A2(n_42),
.B1(n_56),
.B2(n_66),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_99),
.A2(n_36),
.B1(n_83),
.B2(n_38),
.Y(n_134)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_103),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_101),
.A2(n_67),
.B1(n_76),
.B2(n_81),
.Y(n_110)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_71),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_67),
.A2(n_43),
.B1(n_36),
.B2(n_62),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_67),
.A2(n_82),
.B1(n_81),
.B2(n_83),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_88),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_108),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_110),
.A2(n_138),
.B1(n_136),
.B2(n_122),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_76),
.B1(n_54),
.B2(n_74),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_111),
.A2(n_115),
.B1(n_118),
.B2(n_128),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_87),
.A2(n_74),
.B1(n_50),
.B2(n_63),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_46),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_116),
.B(n_117),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_46),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_59),
.B1(n_55),
.B2(n_84),
.Y(n_118)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_122),
.B(n_132),
.Y(n_157)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_135),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_68),
.Y(n_125)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_125),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_102),
.A2(n_84),
.B1(n_43),
.B2(n_60),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_105),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_130),
.Y(n_149)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_71),
.C(n_39),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_94),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_127),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_134),
.A2(n_91),
.B1(n_100),
.B2(n_85),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_90),
.B(n_39),
.C(n_65),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_136),
.A2(n_17),
.B1(n_14),
.B2(n_23),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_90),
.B(n_12),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_12),
.Y(n_165)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_139),
.B(n_151),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_119),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_140),
.B(n_154),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_141),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_SL g142 ( 
.A1(n_113),
.A2(n_85),
.B(n_23),
.C(n_17),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_142),
.A2(n_158),
.B(n_160),
.Y(n_189)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_144),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_124),
.A2(n_36),
.B1(n_19),
.B2(n_38),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_150),
.A2(n_153),
.B1(n_155),
.B2(n_156),
.Y(n_176)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_110),
.A2(n_19),
.B1(n_38),
.B2(n_21),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_114),
.A2(n_21),
.B1(n_16),
.B2(n_51),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_114),
.A2(n_13),
.B1(n_18),
.B2(n_14),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_111),
.A2(n_7),
.B(n_10),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_138),
.A2(n_13),
.B1(n_18),
.B2(n_14),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_159),
.A2(n_169),
.B1(n_172),
.B2(n_17),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_129),
.A2(n_13),
.B1(n_18),
.B2(n_20),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_129),
.A2(n_13),
.B1(n_18),
.B2(n_20),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_134),
.A2(n_13),
.B1(n_15),
.B2(n_20),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_12),
.Y(n_164)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_165),
.B(n_27),
.Y(n_196)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_115),
.Y(n_167)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_167),
.Y(n_188)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_109),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_168),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_170),
.Y(n_200)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_109),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_171),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_121),
.A2(n_17),
.B1(n_23),
.B2(n_20),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_132),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_173),
.B(n_183),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_146),
.A2(n_123),
.B(n_121),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_174),
.A2(n_166),
.B(n_139),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_149),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_175),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_177),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_117),
.C(n_116),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_178),
.B(n_185),
.C(n_186),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_146),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_137),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_123),
.C(n_127),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_143),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_187),
.Y(n_215)
);

NAND2xp33_ASAP7_75t_SL g190 ( 
.A(n_142),
.B(n_40),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_190),
.B(n_155),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_126),
.C(n_31),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_192),
.C(n_193),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_147),
.B(n_126),
.C(n_30),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_147),
.B(n_27),
.C(n_25),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_198),
.Y(n_211)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_196),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_160),
.A2(n_20),
.B1(n_15),
.B2(n_25),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_197),
.A2(n_159),
.B1(n_156),
.B2(n_163),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_145),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_148),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_150),
.Y(n_212)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_202),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_181),
.Y(n_204)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_204),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_192),
.A2(n_154),
.B1(n_158),
.B2(n_141),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_207),
.A2(n_208),
.B1(n_225),
.B2(n_200),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_176),
.A2(n_171),
.B1(n_153),
.B2(n_162),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_209),
.B(n_10),
.Y(n_245)
);

INVx13_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_216),
.Y(n_231)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_212),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_213),
.A2(n_217),
.B1(n_218),
.B2(n_220),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_161),
.Y(n_214)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_214),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_182),
.B(n_12),
.Y(n_216)
);

NOR2xp67_ASAP7_75t_L g217 ( 
.A(n_174),
.B(n_142),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_179),
.A2(n_142),
.B1(n_20),
.B2(n_15),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_179),
.A2(n_20),
.B1(n_15),
.B2(n_24),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_182),
.B(n_12),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_223),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_11),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_189),
.A2(n_188),
.B(n_194),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_224),
.A2(n_184),
.B(n_194),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_176),
.A2(n_193),
.B1(n_189),
.B2(n_200),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_183),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_227),
.B(n_243),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_173),
.C(n_186),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_230),
.C(n_232),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_229),
.A2(n_214),
.B1(n_218),
.B2(n_220),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_226),
.B(n_178),
.C(n_191),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_185),
.C(n_196),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_180),
.Y(n_233)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_233),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_235),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_209),
.C(n_204),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_238),
.C(n_242),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_197),
.C(n_24),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_206),
.B(n_11),
.C(n_1),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_203),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_245),
.B(n_222),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_206),
.B(n_11),
.C(n_1),
.Y(n_246)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_246),
.Y(n_253)
);

XNOR2x1_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_224),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_251),
.Y(n_274)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_230),
.B(n_207),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_252),
.A2(n_255),
.B1(n_260),
.B2(n_205),
.Y(n_264)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_231),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_262),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_240),
.A2(n_211),
.B1(n_213),
.B2(n_225),
.Y(n_255)
);

FAx1_ASAP7_75t_SL g256 ( 
.A(n_245),
.B(n_217),
.CI(n_202),
.CON(n_256),
.SN(n_256)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_241),
.A2(n_215),
.B1(n_208),
.B2(n_205),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_259),
.A2(n_9),
.B1(n_8),
.B2(n_7),
.Y(n_270)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_237),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_235),
.Y(n_262)
);

OAI321xp33_ASAP7_75t_L g263 ( 
.A1(n_259),
.A2(n_239),
.A3(n_236),
.B1(n_234),
.B2(n_244),
.C(n_215),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_263),
.A2(n_269),
.B(n_9),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_264),
.B(n_266),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_250),
.A2(n_238),
.B1(n_210),
.B2(n_246),
.Y(n_266)
);

XNOR2x2_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_242),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_267),
.B(n_258),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_228),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_270),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_227),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_11),
.C(n_1),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_275),
.C(n_253),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_11),
.C(n_2),
.Y(n_275)
);

FAx1_ASAP7_75t_SL g276 ( 
.A(n_249),
.B(n_11),
.CI(n_9),
.CON(n_276),
.SN(n_276)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_9),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_280),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_247),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_278),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_281),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_267),
.A2(n_260),
.B1(n_256),
.B2(n_257),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_257),
.Y(n_281)
);

OAI321xp33_ASAP7_75t_L g292 ( 
.A1(n_282),
.A2(n_285),
.A3(n_7),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_292)
);

INVx11_ASAP7_75t_L g286 ( 
.A(n_276),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_275),
.Y(n_289)
);

NOR2xp67_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_8),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_287),
.A2(n_0),
.B(n_2),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_7),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_288),
.B(n_0),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_292),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_268),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_294),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_274),
.C(n_269),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_297),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_265),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_283),
.Y(n_303)
);

NAND3xp33_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_286),
.C(n_284),
.Y(n_300)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_300),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_303),
.B(n_304),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_290),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_296),
.C(n_291),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_302),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_299),
.B(n_300),
.Y(n_308)
);

OAI311xp33_ASAP7_75t_L g310 ( 
.A1(n_308),
.A2(n_309),
.A3(n_305),
.B1(n_3),
.C1(n_4),
.Y(n_310)
);

AOI21x1_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_0),
.B(n_3),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_0),
.C(n_3),
.Y(n_312)
);

MAJx2_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_3),
.C(n_4),
.Y(n_313)
);

AOI221xp5_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.C(n_243),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_4),
.C(n_6),
.Y(n_315)
);


endmodule