module fake_jpeg_25114_n_114 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_114);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_114;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

AOI21xp33_ASAP7_75t_L g31 ( 
.A1(n_23),
.A2(n_16),
.B(n_17),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_24),
.A2(n_10),
.B1(n_13),
.B2(n_12),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_19),
.A2(n_0),
.B(n_1),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_28),
.A2(n_31),
.B(n_32),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_18),
.A2(n_14),
.B1(n_10),
.B2(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_32),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_31),
.B(n_23),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_38),
.B(n_39),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_28),
.B(n_17),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_26),
.B(n_15),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_42),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_22),
.Y(n_42)
);

AO21x2_ASAP7_75t_SL g44 ( 
.A1(n_41),
.A2(n_27),
.B(n_30),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_46),
.B1(n_34),
.B2(n_30),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_30),
.B1(n_29),
.B2(n_18),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_42),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_51),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_49),
.Y(n_56)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_33),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_14),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_53),
.A2(n_55),
.B1(n_58),
.B2(n_62),
.Y(n_67)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_59),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_41),
.B1(n_29),
.B2(n_14),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_44),
.A2(n_49),
.B1(n_48),
.B2(n_47),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_21),
.Y(n_59)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_10),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_43),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_44),
.A2(n_33),
.B(n_25),
.Y(n_62)
);

OA21x2_ASAP7_75t_L g66 ( 
.A1(n_62),
.A2(n_53),
.B(n_54),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_44),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_68),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_56),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_64),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_24),
.B(n_20),
.C(n_19),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_29),
.B1(n_25),
.B2(n_13),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_57),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_72),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_52),
.C(n_50),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_22),
.C(n_21),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_43),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_74),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_52),
.C(n_43),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_82),
.C(n_11),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_16),
.B1(n_11),
.B2(n_20),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_11),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_81),
.A2(n_0),
.B(n_2),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_63),
.B(n_66),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_87),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_78),
.Y(n_84)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

MAJx2_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_66),
.C(n_24),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_2),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_89),
.A2(n_90),
.B1(n_3),
.B2(n_4),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_94),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_87),
.A2(n_79),
.B(n_81),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_77),
.C(n_82),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_96),
.C(n_3),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_97),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_92),
.B(n_86),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_99),
.B(n_5),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_91),
.B(n_8),
.Y(n_100)
);

AOI21x1_ASAP7_75t_L g106 ( 
.A1(n_100),
.A2(n_6),
.B(n_7),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_102),
.Y(n_105)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_103),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_104),
.B(n_106),
.Y(n_107)
);

NOR2xp67_ASAP7_75t_SL g108 ( 
.A(n_105),
.B(n_101),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_108),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_101),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_110),
.A2(n_109),
.B1(n_95),
.B2(n_8),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_111),
.Y(n_113)
);

BUFx24_ASAP7_75t_SL g114 ( 
.A(n_113),
.Y(n_114)
);


endmodule