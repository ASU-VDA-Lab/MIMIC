module real_jpeg_15311_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_292;
wire n_221;
wire n_249;
wire n_288;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_173;
wire n_40;
wire n_105;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_164;
wire n_48;
wire n_184;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_18;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_258;
wire n_205;
wire n_61;
wire n_110;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_150;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_244;
wire n_128;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_283;
wire n_85;
wire n_102;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;

INVx1_ASAP7_75t_L g90 ( 
.A(n_0),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_0),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_1),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_1),
.Y(n_176)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_1),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g229 ( 
.A(n_1),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_2),
.B(n_145),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_3),
.B(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_3),
.A2(n_14),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_3),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_3),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_3),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_3),
.B(n_195),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_3),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_3),
.B(n_236),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_4),
.B(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_4),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_4),
.B(n_173),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_4),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_4),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_4),
.B(n_226),
.Y(n_225)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_5),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_6),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_7),
.B(n_30),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_7),
.B(n_126),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_7),
.B(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_8),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_9),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_9),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_9),
.B(n_32),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_9),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_9),
.B(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_9),
.B(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_9),
.B(n_258),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_10),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_10),
.B(n_47),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_10),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_10),
.B(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_11),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_13),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_13),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_14),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_14),
.B(n_141),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_15),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_15),
.B(n_51),
.Y(n_50)
);

AND2x4_ASAP7_75t_SL g84 ( 
.A(n_15),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_15),
.B(n_101),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_15),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_15),
.B(n_138),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_15),
.B(n_145),
.Y(n_212)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_182),
.B1(n_292),
.B2(n_293),
.Y(n_17)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_18),
.Y(n_292)
);

NAND2xp33_ASAP7_75t_R g18 ( 
.A(n_19),
.B(n_179),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_130),
.Y(n_19)
);

NOR2xp67_ASAP7_75t_SL g181 ( 
.A(n_20),
.B(n_130),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_76),
.C(n_111),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_21),
.B(n_290),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_39),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_22),
.B(n_40),
.C(n_55),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_31),
.C(n_34),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_23),
.B(n_277),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

XNOR2x1_ASAP7_75t_SL g224 ( 
.A(n_24),
.B(n_28),
.Y(n_224)
);

INVxp67_ASAP7_75t_SL g234 ( 
.A(n_24),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_24),
.A2(n_234),
.B1(n_235),
.B2(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_27),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_31),
.A2(n_34),
.B1(n_35),
.B2(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_31),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_38),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_55),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_45),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_41),
.B(n_46),
.C(n_50),
.Y(n_170)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_49),
.B1(n_50),
.B2(n_54),
.Y(n_45)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_49),
.B(n_190),
.C(n_194),
.Y(n_217)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_50),
.B(n_189),
.Y(n_188)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_64),
.B(n_69),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_62),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_68),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_69),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_148)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_69),
.Y(n_151)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_77),
.B(n_111),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_92),
.C(n_103),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_78),
.B(n_283),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_83),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_84),
.C(n_87),
.Y(n_113)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_82),
.Y(n_161)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_82),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_86),
.B1(n_87),
.B2(n_91),
.Y(n_83)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_84),
.A2(n_91),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_84),
.B(n_240),
.C(n_244),
.Y(n_268)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_93),
.B(n_104),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.C(n_99),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_94),
.A2(n_99),
.B1(n_100),
.B2(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_94),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_95),
.B(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_99),
.A2(n_163),
.B1(n_167),
.B2(n_168),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_100),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_100),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_106),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_109),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_110),
.Y(n_261)
);

XNOR2x2_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_115),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_154),
.C(n_155),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_121),
.Y(n_115)
);

MAJx2_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_125),
.C(n_129),
.Y(n_150)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_120),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_125),
.B1(n_128),
.B2(n_129),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_122),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_125),
.Y(n_128)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_152),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_148),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_139),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_144),
.Y(n_139)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_143),
.Y(n_211)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_156),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_169),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_162),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_163),
.Y(n_168)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_175),
.B1(n_177),
.B2(n_178),
.Y(n_171)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_172),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_175),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_182),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_287),
.B(n_291),
.Y(n_183)
);

AOI21x1_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_271),
.B(n_286),
.Y(n_184)
);

OAI21x1_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_230),
.B(n_270),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_215),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_187),
.B(n_215),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_198),
.C(n_208),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_188),
.B(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_194),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_198),
.A2(n_199),
.B1(n_208),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_204),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_200),
.B(n_204),
.Y(n_241)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_207),
.Y(n_238)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_208),
.Y(n_267)
);

AO22x1_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_208)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_209),
.Y(n_213)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_212),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_213),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_214),
.B(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_221),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_217),
.B(n_221),
.C(n_285),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_218),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

MAJx2_ASAP7_75t_L g280 ( 
.A(n_222),
.B(n_224),
.C(n_225),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_229),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_264),
.B(n_269),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_247),
.B(n_263),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_239),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_239),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_235),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_256),
.B(n_262),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_254),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_254),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_268),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_268),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_284),
.Y(n_271)
);

NOR2x1_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_284),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_281),
.B2(n_282),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_279),
.B2(n_280),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_280),
.C(n_281),
.Y(n_288)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NOR2xp67_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_289),
.Y(n_291)
);


endmodule