module real_jpeg_32569_n_27 (n_17, n_8, n_0, n_21, n_2, n_188, n_196, n_191, n_10, n_186, n_9, n_12, n_24, n_189, n_187, n_6, n_190, n_194, n_192, n_23, n_11, n_14, n_25, n_195, n_7, n_22, n_18, n_3, n_193, n_5, n_4, n_1, n_26, n_20, n_19, n_16, n_15, n_13, n_27);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_188;
input n_196;
input n_191;
input n_10;
input n_186;
input n_9;
input n_12;
input n_24;
input n_189;
input n_187;
input n_6;
input n_190;
input n_194;
input n_192;
input n_23;
input n_11;
input n_14;
input n_25;
input n_195;
input n_7;
input n_22;
input n_18;
input n_3;
input n_193;
input n_5;
input n_4;
input n_1;
input n_26;
input n_20;
input n_19;
input n_16;
input n_15;
input n_13;

output n_27;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_174;
wire n_87;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_1),
.B(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_2),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_2),
.B(n_137),
.Y(n_155)
);

NOR2x1_ASAP7_75t_L g60 ( 
.A(n_3),
.B(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_3),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_4),
.Y(n_54)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_5),
.Y(n_133)
);

AOI322xp5_ASAP7_75t_L g156 ( 
.A1(n_5),
.A2(n_129),
.A3(n_131),
.B1(n_135),
.B2(n_157),
.C1(n_159),
.C2(n_196),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_6),
.B(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_8),
.B(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_9),
.Y(n_115)
);

AOI221xp5_ASAP7_75t_L g96 ( 
.A1(n_10),
.A2(n_20),
.B1(n_97),
.B2(n_101),
.C(n_103),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_10),
.B(n_97),
.C(n_101),
.Y(n_106)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_11),
.A2(n_38),
.B1(n_40),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_13),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_13),
.B(n_149),
.Y(n_158)
);

NOR2x1_ASAP7_75t_L g64 ( 
.A(n_14),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_14),
.B(n_65),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_15),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_15),
.B(n_142),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_16),
.B(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_16),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_17),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_17),
.B(n_77),
.Y(n_184)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_18),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_18),
.B(n_84),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_20),
.Y(n_105)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_21),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_22),
.B(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_22),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_23),
.B(n_85),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_26),
.B(n_72),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_35),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21x1_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_88),
.B(n_162),
.Y(n_36)
);

NAND4xp25_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_49),
.C(n_75),
.D(n_82),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_48),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR3xp33_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_60),
.C(n_62),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND3xp33_ASAP7_75t_L g172 ( 
.A(n_51),
.B(n_173),
.C(n_174),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_59),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_52),
.B(n_59),
.Y(n_177)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_100),
.Y(n_99)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_60),
.Y(n_171)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_61),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI21xp33_ASAP7_75t_L g164 ( 
.A1(n_63),
.A2(n_165),
.B(n_168),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_63),
.B(n_75),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_70),
.Y(n_63)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_64),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_69),
.Y(n_146)
);

INVxp67_ASAP7_75t_SL g170 ( 
.A(n_70),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_70),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_71),
.Y(n_181)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AOI21xp33_ASAP7_75t_L g178 ( 
.A1(n_75),
.A2(n_179),
.B(n_183),
.Y(n_178)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI221xp5_ASAP7_75t_L g163 ( 
.A1(n_76),
.A2(n_164),
.B1(n_175),
.B2(n_176),
.C(n_178),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_87),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI31xp33_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_121),
.A3(n_147),
.B(n_152),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_115),
.C(n_116),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_107),
.B(n_114),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_96),
.B1(n_105),
.B2(n_106),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_98),
.B(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_188),
.Y(n_101)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_113),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_113),
.Y(n_114)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_111),
.Y(n_120)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NOR3xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_134),
.C(n_141),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_122),
.A2(n_153),
.B(n_156),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_129),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NOR3xp33_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_141),
.C(n_158),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_125),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_133),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_192),
.Y(n_131)
);

OA21x2_ASAP7_75t_SL g153 ( 
.A1(n_134),
.A2(n_154),
.B(n_155),
.Y(n_153)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_140),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

NOR2x1_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_186),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_187),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_189),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_190),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_191),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_193),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_194),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_195),
.Y(n_150)
);


endmodule