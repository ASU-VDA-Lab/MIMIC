module real_aes_7255_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g115 ( .A(n_0), .Y(n_115) );
A2O1A1Ixp33_ASAP7_75t_L g233 ( .A1(n_1), .A2(n_151), .B(n_154), .C(n_234), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_2), .A2(n_180), .B(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g507 ( .A(n_3), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_4), .B(n_210), .Y(n_209) );
AOI21xp33_ASAP7_75t_L g490 ( .A1(n_5), .A2(n_180), .B(n_491), .Y(n_490) );
AND2x6_ASAP7_75t_L g151 ( .A(n_6), .B(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g247 ( .A(n_7), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_8), .B(n_43), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_9), .A2(n_179), .B(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_10), .B(n_163), .Y(n_236) );
INVx1_ASAP7_75t_L g495 ( .A(n_11), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_12), .B(n_204), .Y(n_530) );
OAI22xp5_ASAP7_75t_SL g449 ( .A1(n_13), .A2(n_450), .B1(n_451), .B2(n_457), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_13), .Y(n_457) );
INVx1_ASAP7_75t_L g143 ( .A(n_14), .Y(n_143) );
INVx1_ASAP7_75t_L g542 ( .A(n_15), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_16), .A2(n_81), .B1(n_455), .B2(n_456), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_16), .Y(n_455) );
A2O1A1Ixp33_ASAP7_75t_L g268 ( .A1(n_17), .A2(n_188), .B(n_269), .C(n_271), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_18), .B(n_210), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_19), .B(n_473), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_20), .B(n_180), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_21), .B(n_194), .Y(n_193) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_22), .A2(n_204), .B(n_255), .C(n_257), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_23), .B(n_210), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_24), .B(n_163), .Y(n_162) );
A2O1A1Ixp33_ASAP7_75t_L g540 ( .A1(n_25), .A2(n_190), .B(n_271), .C(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_26), .B(n_163), .Y(n_218) );
CKINVDCx16_ASAP7_75t_R g145 ( .A(n_27), .Y(n_145) );
INVx1_ASAP7_75t_L g217 ( .A(n_28), .Y(n_217) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_29), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g232 ( .A(n_30), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_31), .B(n_163), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g443 ( .A(n_32), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g186 ( .A(n_33), .Y(n_186) );
INVx1_ASAP7_75t_L g485 ( .A(n_34), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_35), .A2(n_452), .B1(n_453), .B2(n_454), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_35), .Y(n_452) );
INVx2_ASAP7_75t_L g149 ( .A(n_36), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g238 ( .A(n_37), .Y(n_238) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_38), .A2(n_204), .B(n_205), .C(n_207), .Y(n_203) );
INVxp67_ASAP7_75t_L g189 ( .A(n_39), .Y(n_189) );
CKINVDCx14_ASAP7_75t_R g202 ( .A(n_40), .Y(n_202) );
A2O1A1Ixp33_ASAP7_75t_L g215 ( .A1(n_41), .A2(n_154), .B(n_216), .C(n_220), .Y(n_215) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_42), .A2(n_151), .B(n_154), .C(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g484 ( .A(n_44), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_45), .A2(n_165), .B(n_245), .C(n_246), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_46), .B(n_163), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_47), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_48), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_49), .A2(n_105), .B1(n_117), .B2(n_752), .Y(n_104) );
INVx1_ASAP7_75t_L g253 ( .A(n_50), .Y(n_253) );
CKINVDCx16_ASAP7_75t_R g486 ( .A(n_51), .Y(n_486) );
AOI222xp33_ASAP7_75t_SL g447 ( .A1(n_52), .A2(n_448), .B1(n_449), .B2(n_458), .C1(n_745), .C2(n_748), .Y(n_447) );
OAI22xp5_ASAP7_75t_SL g434 ( .A1(n_53), .A2(n_62), .B1(n_435), .B2(n_436), .Y(n_434) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_53), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_54), .B(n_180), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_55), .A2(n_154), .B1(n_257), .B2(n_483), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_56), .Y(n_522) );
CKINVDCx16_ASAP7_75t_R g504 ( .A(n_57), .Y(n_504) );
CKINVDCx14_ASAP7_75t_R g243 ( .A(n_58), .Y(n_243) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_59), .A2(n_207), .B(n_245), .C(n_494), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g124 ( .A1(n_60), .A2(n_125), .B1(n_126), .B2(n_439), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_60), .Y(n_439) );
INVx1_ASAP7_75t_L g492 ( .A(n_61), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_62), .Y(n_436) );
INVx1_ASAP7_75t_L g152 ( .A(n_63), .Y(n_152) );
INVx1_ASAP7_75t_L g142 ( .A(n_64), .Y(n_142) );
INVx1_ASAP7_75t_SL g206 ( .A(n_65), .Y(n_206) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_66), .Y(n_122) );
OAI22xp5_ASAP7_75t_SL g433 ( .A1(n_67), .A2(n_434), .B1(n_437), .B2(n_438), .Y(n_433) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_67), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_68), .B(n_210), .Y(n_259) );
INVx1_ASAP7_75t_L g158 ( .A(n_69), .Y(n_158) );
A2O1A1Ixp33_ASAP7_75t_SL g472 ( .A1(n_70), .A2(n_207), .B(n_473), .C(n_474), .Y(n_472) );
INVxp67_ASAP7_75t_L g475 ( .A(n_71), .Y(n_475) );
INVx1_ASAP7_75t_L g110 ( .A(n_72), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_73), .A2(n_180), .B(n_242), .Y(n_241) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_74), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_75), .A2(n_180), .B(n_266), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_76), .Y(n_488) );
INVx1_ASAP7_75t_L g548 ( .A(n_77), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_78), .A2(n_179), .B(n_181), .Y(n_178) );
CKINVDCx16_ASAP7_75t_R g214 ( .A(n_79), .Y(n_214) );
INVx1_ASAP7_75t_L g267 ( .A(n_80), .Y(n_267) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_81), .Y(n_456) );
A2O1A1Ixp33_ASAP7_75t_L g549 ( .A1(n_82), .A2(n_151), .B(n_154), .C(n_550), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_83), .A2(n_180), .B(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g270 ( .A(n_84), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_85), .B(n_187), .Y(n_519) );
INVx2_ASAP7_75t_L g140 ( .A(n_86), .Y(n_140) );
INVx1_ASAP7_75t_L g235 ( .A(n_87), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_88), .B(n_473), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_89), .A2(n_151), .B(n_154), .C(n_506), .Y(n_505) );
OR2x2_ASAP7_75t_L g112 ( .A(n_90), .B(n_113), .Y(n_112) );
OR2x2_ASAP7_75t_L g459 ( .A(n_90), .B(n_114), .Y(n_459) );
INVx2_ASAP7_75t_L g744 ( .A(n_90), .Y(n_744) );
A2O1A1Ixp33_ASAP7_75t_L g153 ( .A1(n_91), .A2(n_154), .B(n_157), .C(n_167), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_92), .B(n_172), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_93), .Y(n_511) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_94), .A2(n_151), .B(n_154), .C(n_528), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_95), .Y(n_534) );
INVx1_ASAP7_75t_L g471 ( .A(n_96), .Y(n_471) );
CKINVDCx16_ASAP7_75t_R g539 ( .A(n_97), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_98), .B(n_187), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_99), .B(n_138), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_100), .B(n_138), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_101), .B(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g256 ( .A(n_102), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_103), .A2(n_180), .B(n_470), .Y(n_469) );
BUFx4f_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
CKINVDCx6p67_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g753 ( .A(n_107), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_111), .Y(n_107) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
INVx1_ASAP7_75t_SL g442 ( .A(n_112), .Y(n_442) );
BUFx2_ASAP7_75t_L g445 ( .A(n_112), .Y(n_445) );
NOR2x2_ASAP7_75t_L g747 ( .A(n_113), .B(n_744), .Y(n_747) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
OR2x2_ASAP7_75t_L g743 ( .A(n_114), .B(n_744), .Y(n_743) );
AND2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
OA21x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_123), .B(n_446), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_SL g751 ( .A(n_121), .Y(n_751) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OAI21xp5_ASAP7_75t_SL g123 ( .A1(n_124), .A2(n_440), .B(n_443), .Y(n_123) );
INVxp67_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
XOR2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_433), .Y(n_126) );
OAI22xp5_ASAP7_75t_SL g458 ( .A1(n_127), .A2(n_459), .B1(n_460), .B2(n_741), .Y(n_458) );
INVx2_ASAP7_75t_L g749 ( .A(n_127), .Y(n_749) );
OR2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_367), .Y(n_127) );
NAND5xp2_ASAP7_75t_L g128 ( .A(n_129), .B(n_296), .C(n_326), .D(n_347), .E(n_353), .Y(n_128) );
AOI221xp5_ASAP7_75t_SL g129 ( .A1(n_130), .A2(n_226), .B1(n_260), .B2(n_262), .C(n_273), .Y(n_129) );
INVxp67_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_132), .B(n_223), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g132 ( .A(n_133), .B(n_195), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
A2O1A1Ixp33_ASAP7_75t_SL g347 ( .A1(n_134), .A2(n_211), .B(n_348), .C(n_351), .Y(n_347) );
AND2x2_ASAP7_75t_L g417 ( .A(n_134), .B(n_212), .Y(n_417) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_173), .Y(n_134) );
AND2x2_ASAP7_75t_L g275 ( .A(n_135), .B(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g279 ( .A(n_135), .B(n_276), .Y(n_279) );
OR2x2_ASAP7_75t_L g305 ( .A(n_135), .B(n_212), .Y(n_305) );
AND2x2_ASAP7_75t_L g307 ( .A(n_135), .B(n_198), .Y(n_307) );
AND2x2_ASAP7_75t_L g325 ( .A(n_135), .B(n_197), .Y(n_325) );
INVx1_ASAP7_75t_L g358 ( .A(n_135), .Y(n_358) );
INVx2_ASAP7_75t_SL g135 ( .A(n_136), .Y(n_135) );
BUFx2_ASAP7_75t_L g225 ( .A(n_136), .Y(n_225) );
AND2x2_ASAP7_75t_L g261 ( .A(n_136), .B(n_198), .Y(n_261) );
AND2x2_ASAP7_75t_L g414 ( .A(n_136), .B(n_212), .Y(n_414) );
AO21x2_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_144), .B(n_169), .Y(n_136) );
INVx3_ASAP7_75t_L g210 ( .A(n_137), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_137), .B(n_222), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_137), .B(n_238), .Y(n_237) );
NOR2xp33_ASAP7_75t_SL g521 ( .A(n_137), .B(n_522), .Y(n_521) );
INVx4_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_138), .Y(n_199) );
OA21x2_ASAP7_75t_L g468 ( .A1(n_138), .A2(n_469), .B(n_476), .Y(n_468) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g176 ( .A(n_139), .Y(n_176) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x2_ASAP7_75t_SL g172 ( .A(n_140), .B(n_141), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
OAI21xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_146), .B(n_153), .Y(n_144) );
O2A1O1Ixp33_ASAP7_75t_L g213 ( .A1(n_146), .A2(n_172), .B(n_214), .C(n_215), .Y(n_213) );
OAI21xp5_ASAP7_75t_L g231 ( .A1(n_146), .A2(n_232), .B(n_233), .Y(n_231) );
OAI22xp33_ASAP7_75t_L g481 ( .A1(n_146), .A2(n_168), .B1(n_482), .B2(n_486), .Y(n_481) );
OAI21xp5_ASAP7_75t_L g503 ( .A1(n_146), .A2(n_504), .B(n_505), .Y(n_503) );
OAI21xp5_ASAP7_75t_L g547 ( .A1(n_146), .A2(n_548), .B(n_549), .Y(n_547) );
NAND2x1p5_ASAP7_75t_L g146 ( .A(n_147), .B(n_151), .Y(n_146) );
AND2x4_ASAP7_75t_L g180 ( .A(n_147), .B(n_151), .Y(n_180) );
AND2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_150), .Y(n_147) );
INVx1_ASAP7_75t_L g191 ( .A(n_148), .Y(n_191) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g155 ( .A(n_149), .Y(n_155) );
INVx1_ASAP7_75t_L g258 ( .A(n_149), .Y(n_258) );
INVx1_ASAP7_75t_L g156 ( .A(n_150), .Y(n_156) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_150), .Y(n_161) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_150), .Y(n_163) );
INVx3_ASAP7_75t_L g188 ( .A(n_150), .Y(n_188) );
INVx1_ASAP7_75t_L g473 ( .A(n_150), .Y(n_473) );
INVx4_ASAP7_75t_SL g168 ( .A(n_151), .Y(n_168) );
BUFx3_ASAP7_75t_L g220 ( .A(n_151), .Y(n_220) );
INVx5_ASAP7_75t_L g183 ( .A(n_154), .Y(n_183) );
AND2x6_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
BUFx3_ASAP7_75t_L g166 ( .A(n_155), .Y(n_166) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_155), .Y(n_208) );
O2A1O1Ixp33_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_159), .B(n_162), .C(n_164), .Y(n_157) );
O2A1O1Ixp5_ASAP7_75t_L g234 ( .A1(n_159), .A2(n_164), .B(n_235), .C(n_236), .Y(n_234) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
OAI22xp5_ASAP7_75t_SL g483 ( .A1(n_160), .A2(n_161), .B1(n_484), .B2(n_485), .Y(n_483) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx4_ASAP7_75t_L g190 ( .A(n_161), .Y(n_190) );
INVx4_ASAP7_75t_L g204 ( .A(n_163), .Y(n_204) );
INVx2_ASAP7_75t_L g245 ( .A(n_163), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_164), .A2(n_519), .B(n_520), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_164), .A2(n_551), .B(n_552), .Y(n_550) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g271 ( .A(n_166), .Y(n_271) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
O2A1O1Ixp33_ASAP7_75t_SL g181 ( .A1(n_168), .A2(n_182), .B(n_183), .C(n_184), .Y(n_181) );
O2A1O1Ixp33_ASAP7_75t_L g201 ( .A1(n_168), .A2(n_183), .B(n_202), .C(n_203), .Y(n_201) );
O2A1O1Ixp33_ASAP7_75t_SL g242 ( .A1(n_168), .A2(n_183), .B(n_243), .C(n_244), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_SL g252 ( .A1(n_168), .A2(n_183), .B(n_253), .C(n_254), .Y(n_252) );
O2A1O1Ixp33_ASAP7_75t_SL g266 ( .A1(n_168), .A2(n_183), .B(n_267), .C(n_268), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_L g470 ( .A1(n_168), .A2(n_183), .B(n_471), .C(n_472), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_168), .A2(n_183), .B(n_492), .C(n_493), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_L g538 ( .A1(n_168), .A2(n_183), .B(n_539), .C(n_540), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
INVx1_ASAP7_75t_L g194 ( .A(n_171), .Y(n_194) );
AO21x2_ASAP7_75t_L g525 ( .A1(n_171), .A2(n_526), .B(n_533), .Y(n_525) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g230 ( .A(n_172), .Y(n_230) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_172), .A2(n_241), .B(n_248), .Y(n_240) );
OA21x2_ASAP7_75t_L g536 ( .A1(n_172), .A2(n_537), .B(n_543), .Y(n_536) );
AND2x2_ASAP7_75t_L g295 ( .A(n_173), .B(n_196), .Y(n_295) );
OR2x2_ASAP7_75t_L g299 ( .A(n_173), .B(n_212), .Y(n_299) );
AND2x2_ASAP7_75t_L g324 ( .A(n_173), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_SL g371 ( .A(n_173), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_173), .B(n_333), .Y(n_419) );
AO21x2_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_177), .B(n_192), .Y(n_173) );
INVx1_ASAP7_75t_L g277 ( .A(n_174), .Y(n_277) );
AO21x2_ASAP7_75t_L g546 ( .A1(n_174), .A2(n_547), .B(n_553), .Y(n_546) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AOI21xp5_ASAP7_75t_SL g515 ( .A1(n_175), .A2(n_516), .B(n_517), .Y(n_515) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AO21x2_ASAP7_75t_L g480 ( .A1(n_176), .A2(n_481), .B(n_487), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_176), .B(n_488), .Y(n_487) );
AO21x2_ASAP7_75t_L g502 ( .A1(n_176), .A2(n_503), .B(n_510), .Y(n_502) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
OA21x2_ASAP7_75t_L g276 ( .A1(n_178), .A2(n_193), .B(n_277), .Y(n_276) );
BUFx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_185), .B(n_191), .Y(n_184) );
OAI22xp33_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B1(n_189), .B2(n_190), .Y(n_185) );
O2A1O1Ixp33_ASAP7_75t_L g216 ( .A1(n_187), .A2(n_217), .B(n_218), .C(n_219), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_L g506 ( .A1(n_187), .A2(n_507), .B(n_508), .C(n_509), .Y(n_506) );
INVx5_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_188), .B(n_247), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_188), .B(n_475), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_188), .B(n_495), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_190), .B(n_256), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_190), .B(n_270), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_190), .B(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g219 ( .A(n_191), .Y(n_219) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
OAI322xp33_ASAP7_75t_L g420 ( .A1(n_195), .A2(n_356), .A3(n_379), .B1(n_400), .B2(n_421), .C1(n_423), .C2(n_424), .Y(n_420) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_196), .B(n_276), .Y(n_423) );
AND2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_211), .Y(n_196) );
AND2x2_ASAP7_75t_L g224 ( .A(n_197), .B(n_225), .Y(n_224) );
AND2x4_ASAP7_75t_L g292 ( .A(n_197), .B(n_212), .Y(n_292) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g333 ( .A(n_198), .B(n_212), .Y(n_333) );
AND2x2_ASAP7_75t_L g377 ( .A(n_198), .B(n_211), .Y(n_377) );
OA21x2_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B(n_209), .Y(n_198) );
OA21x2_ASAP7_75t_L g250 ( .A1(n_199), .A2(n_251), .B(n_259), .Y(n_250) );
OA21x2_ASAP7_75t_L g264 ( .A1(n_199), .A2(n_265), .B(n_272), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_204), .B(n_206), .Y(n_205) );
INVx3_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
HB1xp67_ASAP7_75t_L g531 ( .A(n_208), .Y(n_531) );
OA21x2_ASAP7_75t_L g489 ( .A1(n_210), .A2(n_490), .B(n_496), .Y(n_489) );
AND2x2_ASAP7_75t_L g260 ( .A(n_211), .B(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g278 ( .A(n_211), .B(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_211), .B(n_307), .Y(n_431) );
INVx3_ASAP7_75t_SL g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g223 ( .A(n_212), .B(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_212), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g345 ( .A(n_212), .B(n_276), .Y(n_345) );
AND2x2_ASAP7_75t_L g372 ( .A(n_212), .B(n_307), .Y(n_372) );
OR2x2_ASAP7_75t_L g428 ( .A(n_212), .B(n_279), .Y(n_428) );
OR2x6_ASAP7_75t_L g212 ( .A(n_213), .B(n_221), .Y(n_212) );
INVx1_ASAP7_75t_SL g314 ( .A(n_223), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_224), .B(n_345), .Y(n_346) );
AND2x2_ASAP7_75t_L g380 ( .A(n_224), .B(n_370), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_224), .B(n_303), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_224), .B(n_425), .Y(n_424) );
OAI31xp33_ASAP7_75t_L g398 ( .A1(n_226), .A2(n_260), .A3(n_399), .B(n_401), .Y(n_398) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_239), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g365 ( .A(n_227), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g381 ( .A(n_227), .B(n_316), .Y(n_381) );
OR2x2_ASAP7_75t_L g388 ( .A(n_227), .B(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g400 ( .A(n_227), .B(n_289), .Y(n_400) );
CKINVDCx16_ASAP7_75t_R g227 ( .A(n_228), .Y(n_227) );
OR2x2_ASAP7_75t_L g334 ( .A(n_228), .B(n_335), .Y(n_334) );
BUFx3_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g262 ( .A(n_229), .B(n_263), .Y(n_262) );
INVx4_ASAP7_75t_L g283 ( .A(n_229), .Y(n_283) );
AND2x2_ASAP7_75t_L g320 ( .A(n_229), .B(n_264), .Y(n_320) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_237), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_230), .B(n_511), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_230), .B(n_534), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_230), .B(n_439), .Y(n_553) );
AND2x2_ASAP7_75t_L g319 ( .A(n_239), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_SL g389 ( .A(n_239), .Y(n_389) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_249), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_240), .B(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g289 ( .A(n_240), .B(n_250), .Y(n_289) );
INVx2_ASAP7_75t_L g309 ( .A(n_240), .Y(n_309) );
AND2x2_ASAP7_75t_L g323 ( .A(n_240), .B(n_250), .Y(n_323) );
AND2x2_ASAP7_75t_L g330 ( .A(n_240), .B(n_286), .Y(n_330) );
BUFx3_ASAP7_75t_L g340 ( .A(n_240), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_240), .B(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g285 ( .A(n_249), .Y(n_285) );
AND2x2_ASAP7_75t_L g293 ( .A(n_249), .B(n_283), .Y(n_293) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g263 ( .A(n_250), .B(n_264), .Y(n_263) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_250), .Y(n_317) );
INVx2_ASAP7_75t_L g509 ( .A(n_257), .Y(n_509) );
INVx3_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx2_ASAP7_75t_SL g300 ( .A(n_261), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_261), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_261), .B(n_370), .Y(n_391) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_262), .B(n_340), .Y(n_393) );
INVx1_ASAP7_75t_SL g427 ( .A(n_262), .Y(n_427) );
INVx1_ASAP7_75t_SL g335 ( .A(n_263), .Y(n_335) );
INVx1_ASAP7_75t_SL g286 ( .A(n_264), .Y(n_286) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_264), .Y(n_297) );
OR2x2_ASAP7_75t_L g308 ( .A(n_264), .B(n_283), .Y(n_308) );
AND2x2_ASAP7_75t_L g322 ( .A(n_264), .B(n_283), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_264), .B(n_312), .Y(n_374) );
A2O1A1Ixp33_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_278), .B(n_280), .C(n_291), .Y(n_273) );
AOI31xp33_ASAP7_75t_L g390 ( .A1(n_274), .A2(n_391), .A3(n_392), .B(n_393), .Y(n_390) );
AND2x2_ASAP7_75t_L g363 ( .A(n_275), .B(n_292), .Y(n_363) );
BUFx3_ASAP7_75t_L g303 ( .A(n_276), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_276), .B(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g339 ( .A(n_276), .B(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_276), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_SL g294 ( .A(n_279), .Y(n_294) );
OAI222xp33_ASAP7_75t_L g403 ( .A1(n_279), .A2(n_404), .B1(n_407), .B2(n_408), .C1(n_409), .C2(n_410), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_281), .B(n_287), .Y(n_280) );
INVx1_ASAP7_75t_L g409 ( .A(n_281), .Y(n_409) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_283), .B(n_286), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_283), .B(n_309), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_283), .B(n_284), .Y(n_379) );
INVx1_ASAP7_75t_L g430 ( .A(n_283), .Y(n_430) );
NAND2xp5_ASAP7_75t_SL g360 ( .A(n_284), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g432 ( .A(n_284), .Y(n_432) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVx2_ASAP7_75t_L g312 ( .A(n_285), .Y(n_312) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_286), .Y(n_355) );
AOI32xp33_ASAP7_75t_L g291 ( .A1(n_287), .A2(n_292), .A3(n_293), .B1(n_294), .B2(n_295), .Y(n_291) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_289), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g366 ( .A(n_289), .Y(n_366) );
OR2x2_ASAP7_75t_L g407 ( .A(n_289), .B(n_308), .Y(n_407) );
INVx1_ASAP7_75t_L g343 ( .A(n_290), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_292), .B(n_303), .Y(n_328) );
INVx3_ASAP7_75t_L g337 ( .A(n_292), .Y(n_337) );
AOI322xp5_ASAP7_75t_L g353 ( .A1(n_292), .A2(n_337), .A3(n_354), .B1(n_356), .B2(n_359), .C1(n_363), .C2(n_364), .Y(n_353) );
AND2x2_ASAP7_75t_L g329 ( .A(n_293), .B(n_330), .Y(n_329) );
INVxp67_ASAP7_75t_L g406 ( .A(n_293), .Y(n_406) );
A2O1A1O1Ixp25_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_298), .B(n_301), .C(n_309), .D(n_310), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_297), .B(n_340), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
OAI221xp5_ASAP7_75t_L g310 ( .A1(n_299), .A2(n_311), .B1(n_314), .B2(n_315), .C(n_318), .Y(n_310) );
INVx1_ASAP7_75t_SL g425 ( .A(n_299), .Y(n_425) );
AOI21xp33_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_306), .B(n_308), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
NAND2xp5_ASAP7_75t_SL g413 ( .A(n_303), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OAI221xp5_ASAP7_75t_SL g395 ( .A1(n_305), .A2(n_389), .B1(n_396), .B2(n_397), .C(n_398), .Y(n_395) );
OAI222xp33_ASAP7_75t_L g426 ( .A1(n_306), .A2(n_427), .B1(n_428), .B2(n_429), .C1(n_431), .C2(n_432), .Y(n_426) );
AND2x2_ASAP7_75t_L g384 ( .A(n_307), .B(n_370), .Y(n_384) );
AOI21xp5_ASAP7_75t_L g396 ( .A1(n_307), .A2(n_322), .B(n_369), .Y(n_396) );
INVx1_ASAP7_75t_L g410 ( .A(n_307), .Y(n_410) );
INVx2_ASAP7_75t_SL g313 ( .A(n_308), .Y(n_313) );
AND2x2_ASAP7_75t_L g316 ( .A(n_309), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx1_ASAP7_75t_SL g350 ( .A(n_312), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_312), .B(n_322), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_313), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_313), .B(n_323), .Y(n_352) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OAI21xp5_ASAP7_75t_SL g318 ( .A1(n_319), .A2(n_321), .B(n_324), .Y(n_318) );
INVx1_ASAP7_75t_SL g336 ( .A(n_320), .Y(n_336) );
AND2x2_ASAP7_75t_L g383 ( .A(n_320), .B(n_366), .Y(n_383) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
AND2x2_ASAP7_75t_L g422 ( .A(n_322), .B(n_340), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_323), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_SL g408 ( .A(n_324), .Y(n_408) );
AOI221xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_329), .B1(n_331), .B2(n_338), .C(n_341), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OAI22xp5_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_334), .B1(n_336), .B2(n_337), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OAI22xp33_ASAP7_75t_L g341 ( .A1(n_335), .A2(n_342), .B1(n_344), .B2(n_346), .Y(n_341) );
OR2x2_ASAP7_75t_L g412 ( .A(n_336), .B(n_340), .Y(n_412) );
OR2x2_ASAP7_75t_L g415 ( .A(n_336), .B(n_350), .Y(n_415) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OAI221xp5_ASAP7_75t_L g411 ( .A1(n_357), .A2(n_412), .B1(n_413), .B2(n_415), .C(n_416), .Y(n_411) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVxp67_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND3xp33_ASAP7_75t_SL g367 ( .A(n_368), .B(n_382), .C(n_394), .Y(n_367) );
AOI222xp33_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_373), .B1(n_375), .B2(n_378), .C1(n_380), .C2(n_381), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_372), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_370), .B(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g392 ( .A(n_372), .Y(n_392) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVxp67_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AOI221xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_384), .B1(n_385), .B2(n_387), .C(n_390), .Y(n_382) );
INVx1_ASAP7_75t_L g397 ( .A(n_383), .Y(n_397) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
OAI21xp33_ASAP7_75t_L g416 ( .A1(n_387), .A2(n_417), .B(n_418), .Y(n_416) );
INVx1_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
NOR5xp2_ASAP7_75t_L g394 ( .A(n_395), .B(n_403), .C(n_411), .D(n_420), .E(n_426), .Y(n_394) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
OR2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
INVxp67_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_434), .Y(n_438) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
NAND3xp33_ASAP7_75t_L g446 ( .A(n_443), .B(n_447), .C(n_750), .Y(n_446) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OAI22xp5_ASAP7_75t_SL g748 ( .A1(n_459), .A2(n_461), .B1(n_741), .B2(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_SL g461 ( .A(n_462), .B(n_678), .Y(n_461) );
NOR4xp25_ASAP7_75t_L g462 ( .A(n_463), .B(n_608), .C(n_639), .D(n_658), .Y(n_462) );
NAND4xp25_ASAP7_75t_L g463 ( .A(n_464), .B(n_566), .C(n_581), .D(n_599), .Y(n_463) );
AOI222xp33_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_512), .B1(n_544), .B2(n_554), .C1(n_559), .C2(n_561), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_497), .Y(n_465) );
INVx1_ASAP7_75t_L g622 ( .A(n_466), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_477), .Y(n_466) );
AND2x2_ASAP7_75t_L g498 ( .A(n_467), .B(n_489), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_467), .B(n_501), .Y(n_651) );
INVx3_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
OR2x2_ASAP7_75t_L g558 ( .A(n_468), .B(n_479), .Y(n_558) );
AND2x2_ASAP7_75t_L g567 ( .A(n_468), .B(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g593 ( .A(n_468), .Y(n_593) );
AND2x2_ASAP7_75t_L g614 ( .A(n_468), .B(n_479), .Y(n_614) );
BUFx2_ASAP7_75t_L g637 ( .A(n_468), .Y(n_637) );
AND2x2_ASAP7_75t_L g661 ( .A(n_468), .B(n_480), .Y(n_661) );
AND2x2_ASAP7_75t_L g725 ( .A(n_468), .B(n_489), .Y(n_725) );
AND2x2_ASAP7_75t_L g626 ( .A(n_477), .B(n_557), .Y(n_626) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_478), .B(n_651), .Y(n_650) );
OR2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_489), .Y(n_478) );
OR2x2_ASAP7_75t_L g586 ( .A(n_479), .B(n_502), .Y(n_586) );
AND2x2_ASAP7_75t_L g598 ( .A(n_479), .B(n_557), .Y(n_598) );
BUFx2_ASAP7_75t_L g730 ( .A(n_479), .Y(n_730) );
INVx3_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
OR2x2_ASAP7_75t_L g500 ( .A(n_480), .B(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g580 ( .A(n_480), .B(n_502), .Y(n_580) );
AND2x2_ASAP7_75t_L g633 ( .A(n_480), .B(n_489), .Y(n_633) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_480), .Y(n_669) );
AND2x2_ASAP7_75t_L g556 ( .A(n_489), .B(n_557), .Y(n_556) );
INVx1_ASAP7_75t_SL g568 ( .A(n_489), .Y(n_568) );
INVx2_ASAP7_75t_L g579 ( .A(n_489), .Y(n_579) );
BUFx2_ASAP7_75t_L g603 ( .A(n_489), .Y(n_603) );
AND2x2_ASAP7_75t_SL g660 ( .A(n_489), .B(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
AOI332xp33_ASAP7_75t_L g581 ( .A1(n_498), .A2(n_582), .A3(n_586), .B1(n_587), .B2(n_591), .B3(n_594), .C1(n_595), .C2(n_597), .Y(n_581) );
NAND2x1_ASAP7_75t_L g666 ( .A(n_498), .B(n_557), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_498), .B(n_571), .Y(n_717) );
A2O1A1Ixp33_ASAP7_75t_SL g599 ( .A1(n_499), .A2(n_600), .B(n_603), .C(n_604), .Y(n_599) );
AND2x2_ASAP7_75t_L g738 ( .A(n_499), .B(n_579), .Y(n_738) );
INVx3_ASAP7_75t_SL g499 ( .A(n_500), .Y(n_499) );
OR2x2_ASAP7_75t_L g635 ( .A(n_500), .B(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g640 ( .A(n_500), .B(n_637), .Y(n_640) );
INVx1_ASAP7_75t_L g571 ( .A(n_501), .Y(n_571) );
AND2x2_ASAP7_75t_L g674 ( .A(n_501), .B(n_633), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_501), .B(n_614), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_501), .B(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_501), .B(n_592), .Y(n_700) );
INVx3_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx3_ASAP7_75t_L g557 ( .A(n_502), .Y(n_557) );
OAI31xp33_ASAP7_75t_L g739 ( .A1(n_512), .A2(n_660), .A3(n_667), .B(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_523), .Y(n_512) );
AND2x2_ASAP7_75t_L g544 ( .A(n_513), .B(n_545), .Y(n_544) );
NAND2x1_ASAP7_75t_SL g562 ( .A(n_513), .B(n_563), .Y(n_562) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_513), .Y(n_649) );
AND2x2_ASAP7_75t_L g654 ( .A(n_513), .B(n_565), .Y(n_654) );
INVx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g566 ( .A1(n_514), .A2(n_567), .B(n_569), .C(n_572), .Y(n_566) );
OR2x2_ASAP7_75t_L g583 ( .A(n_514), .B(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g596 ( .A(n_514), .Y(n_596) );
AND2x2_ASAP7_75t_L g602 ( .A(n_514), .B(n_546), .Y(n_602) );
INVx2_ASAP7_75t_L g620 ( .A(n_514), .Y(n_620) );
AND2x2_ASAP7_75t_L g631 ( .A(n_514), .B(n_585), .Y(n_631) );
AND2x2_ASAP7_75t_L g663 ( .A(n_514), .B(n_621), .Y(n_663) );
AND2x2_ASAP7_75t_L g667 ( .A(n_514), .B(n_590), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_514), .B(n_523), .Y(n_672) );
AND2x2_ASAP7_75t_L g706 ( .A(n_514), .B(n_707), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_514), .B(n_609), .Y(n_740) );
OR2x6_ASAP7_75t_L g514 ( .A(n_515), .B(n_521), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_523), .B(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g648 ( .A(n_523), .Y(n_648) );
AND2x2_ASAP7_75t_L g710 ( .A(n_523), .B(n_631), .Y(n_710) );
AND2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_535), .Y(n_523) );
OR2x2_ASAP7_75t_L g564 ( .A(n_524), .B(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g574 ( .A(n_524), .B(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_524), .B(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g682 ( .A(n_524), .Y(n_682) );
AND2x2_ASAP7_75t_L g699 ( .A(n_524), .B(n_546), .Y(n_699) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g590 ( .A(n_525), .B(n_535), .Y(n_590) );
AND2x2_ASAP7_75t_L g619 ( .A(n_525), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g630 ( .A(n_525), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_525), .B(n_585), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_532), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_530), .B(n_531), .Y(n_528) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g545 ( .A(n_536), .B(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g565 ( .A(n_536), .Y(n_565) );
AND2x2_ASAP7_75t_L g621 ( .A(n_536), .B(n_585), .Y(n_621) );
INVx1_ASAP7_75t_L g723 ( .A(n_544), .Y(n_723) );
INVx1_ASAP7_75t_L g727 ( .A(n_545), .Y(n_727) );
INVx2_ASAP7_75t_L g585 ( .A(n_546), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_555), .B(n_558), .Y(n_554) );
INVx1_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_556), .B(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_556), .B(n_661), .Y(n_719) );
OR2x2_ASAP7_75t_L g560 ( .A(n_557), .B(n_558), .Y(n_560) );
INVx1_ASAP7_75t_SL g612 ( .A(n_557), .Y(n_612) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AOI221xp5_ASAP7_75t_L g615 ( .A1(n_563), .A2(n_616), .B1(n_618), .B2(n_622), .C(n_623), .Y(n_615) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
OR2x2_ASAP7_75t_L g643 ( .A(n_564), .B(n_607), .Y(n_643) );
INVx2_ASAP7_75t_L g575 ( .A(n_565), .Y(n_575) );
INVx1_ASAP7_75t_L g601 ( .A(n_565), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_565), .B(n_585), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_565), .B(n_588), .Y(n_695) );
INVx1_ASAP7_75t_L g703 ( .A(n_565), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_567), .B(n_571), .Y(n_617) );
AND2x4_ASAP7_75t_L g592 ( .A(n_568), .B(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g705 ( .A(n_571), .B(n_661), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_576), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_574), .B(n_606), .Y(n_605) );
INVxp67_ASAP7_75t_L g713 ( .A(n_575), .Y(n_713) );
INVxp67_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_580), .Y(n_577) );
INVx1_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g613 ( .A(n_579), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g685 ( .A(n_579), .B(n_661), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_579), .B(n_598), .Y(n_691) );
AOI322xp5_ASAP7_75t_L g645 ( .A1(n_580), .A2(n_614), .A3(n_621), .B1(n_646), .B2(n_649), .C1(n_650), .C2(n_652), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_580), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g711 ( .A(n_583), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g657 ( .A(n_584), .Y(n_657) );
INVx2_ASAP7_75t_L g588 ( .A(n_585), .Y(n_588) );
INVx1_ASAP7_75t_L g647 ( .A(n_585), .Y(n_647) );
CKINVDCx16_ASAP7_75t_R g594 ( .A(n_586), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
AND2x2_ASAP7_75t_L g683 ( .A(n_588), .B(n_596), .Y(n_683) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g595 ( .A(n_590), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g638 ( .A(n_590), .B(n_631), .Y(n_638) );
AND2x2_ASAP7_75t_L g642 ( .A(n_590), .B(n_602), .Y(n_642) );
OAI21xp33_ASAP7_75t_SL g652 ( .A1(n_591), .A2(n_653), .B(n_655), .Y(n_652) );
OAI22xp33_ASAP7_75t_L g722 ( .A1(n_591), .A2(n_723), .B1(n_724), .B2(n_726), .Y(n_722) );
INVx3_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g597 ( .A(n_592), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_592), .B(n_612), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_594), .B(n_732), .Y(n_731) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx1_ASAP7_75t_L g734 ( .A(n_601), .Y(n_734) );
INVx4_ASAP7_75t_L g607 ( .A(n_602), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_602), .B(n_629), .Y(n_677) );
INVx1_ASAP7_75t_SL g689 ( .A(n_603), .Y(n_689) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NOR2xp67_ASAP7_75t_L g702 ( .A(n_607), .B(n_703), .Y(n_702) );
OAI211xp5_ASAP7_75t_SL g608 ( .A1(n_609), .A2(n_610), .B(n_615), .C(n_632), .Y(n_608) );
OAI221xp5_ASAP7_75t_SL g728 ( .A1(n_610), .A2(n_648), .B1(n_727), .B2(n_729), .C(n_731), .Y(n_728) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_612), .B(n_725), .Y(n_724) );
OAI31xp33_ASAP7_75t_L g704 ( .A1(n_613), .A2(n_690), .A3(n_705), .B(n_706), .Y(n_704) );
INVx1_ASAP7_75t_L g644 ( .A(n_614), .Y(n_644) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
INVx1_ASAP7_75t_L g694 ( .A(n_619), .Y(n_694) );
AND2x2_ASAP7_75t_L g707 ( .A(n_621), .B(n_630), .Y(n_707) );
AOI21xp33_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_625), .B(n_627), .Y(n_623) );
INVx1_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
INVxp67_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_631), .B(n_734), .Y(n_733) );
OAI21xp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_634), .B(n_638), .Y(n_632) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OAI221xp5_ASAP7_75t_SL g639 ( .A1(n_640), .A2(n_641), .B1(n_643), .B2(n_644), .C(n_645), .Y(n_639) );
A2O1A1Ixp33_ASAP7_75t_L g708 ( .A1(n_640), .A2(n_709), .B(n_711), .C(n_714), .Y(n_708) );
CKINVDCx16_ASAP7_75t_R g641 ( .A(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g692 ( .A(n_643), .B(n_693), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
INVx1_ASAP7_75t_L g670 ( .A(n_651), .Y(n_670) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g656 ( .A(n_654), .B(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g698 ( .A(n_654), .B(n_699), .Y(n_698) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OAI211xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_662), .B(n_664), .C(n_673), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OAI221xp5_ASAP7_75t_L g735 ( .A1(n_662), .A2(n_672), .B1(n_736), .B2(n_737), .C(n_739), .Y(n_735) );
INVx1_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_667), .B1(n_668), .B2(n_671), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OAI21xp5_ASAP7_75t_SL g673 ( .A1(n_674), .A2(n_675), .B(n_676), .Y(n_673) );
INVx1_ASAP7_75t_SL g736 ( .A(n_675), .Y(n_736) );
INVxp67_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NOR4xp25_ASAP7_75t_L g678 ( .A(n_679), .B(n_708), .C(n_728), .D(n_735), .Y(n_678) );
OAI211xp5_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_684), .B(n_686), .C(n_704), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_683), .Y(n_680) );
INVxp67_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
O2A1O1Ixp33_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_690), .B(n_692), .C(n_696), .Y(n_686) );
INVx1_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_SL g715 ( .A(n_693), .Y(n_715) );
OR2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
OR2x2_ASAP7_75t_L g726 ( .A(n_694), .B(n_727), .Y(n_726) );
OAI21xp33_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_700), .B(n_701), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AOI221xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_716), .B1(n_718), .B2(n_720), .C(n_722), .Y(n_714) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVxp67_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_725), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
endmodule