module fake_jpeg_2618_n_191 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_191);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_191;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_27),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_49),
.Y(n_51)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

CKINVDCx6p67_ASAP7_75t_R g57 ( 
.A(n_46),
.Y(n_57)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_23),
.Y(n_62)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_27),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_50),
.A2(n_28),
.B1(n_20),
.B2(n_26),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_17),
.B1(n_30),
.B2(n_23),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_52),
.A2(n_68),
.B1(n_21),
.B2(n_6),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_30),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_60),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_32),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_58),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_32),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_17),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_1),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_19),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_35),
.B(n_19),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_7),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_46),
.A2(n_28),
.B1(n_20),
.B2(n_18),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_70),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_25),
.Y(n_71)
);

CKINVDCx5p33_ASAP7_75t_R g81 ( 
.A(n_71),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_41),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_72),
.Y(n_84)
);

O2A1O1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_47),
.A2(n_29),
.B(n_26),
.C(n_21),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_76),
.A2(n_26),
.B(n_25),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_78),
.A2(n_87),
.B(n_88),
.Y(n_113)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_55),
.A2(n_29),
.B1(n_21),
.B2(n_5),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_SL g110 ( 
.A1(n_82),
.A2(n_85),
.B(n_57),
.C(n_76),
.Y(n_110)
);

INVx3_ASAP7_75t_SL g83 ( 
.A(n_63),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_60),
.A2(n_21),
.B1(n_3),
.B2(n_6),
.Y(n_85)
);

NOR2x1_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_21),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_98),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_66),
.C(n_77),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_94),
.Y(n_120)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_1),
.C(n_6),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_99),
.Y(n_106)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_7),
.C(n_8),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_8),
.Y(n_99)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_100),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_11),
.Y(n_109)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_103),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_118),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_111),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_96),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_81),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_54),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_124),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_12),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_122),
.B(n_123),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_13),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_78),
.A2(n_65),
.B(n_53),
.C(n_73),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_108),
.A2(n_86),
.B1(n_84),
.B2(n_90),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_133),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_121),
.A2(n_85),
.B1(n_92),
.B2(n_82),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_129),
.A2(n_130),
.B1(n_106),
.B2(n_110),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_113),
.A2(n_88),
.B1(n_99),
.B2(n_61),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_120),
.A2(n_88),
.B1(n_75),
.B2(n_61),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_135),
.Y(n_146)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_81),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_136),
.B(n_137),
.Y(n_145)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_98),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_138),
.B(n_139),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_94),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_93),
.C(n_97),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_140),
.B(n_120),
.Y(n_142)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_141),
.B(n_116),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_149),
.Y(n_162)
);

NOR2xp67_ASAP7_75t_SL g144 ( 
.A(n_135),
.B(n_110),
.Y(n_144)
);

INVx13_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_114),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_125),
.A2(n_106),
.B1(n_110),
.B2(n_124),
.Y(n_148)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

OAI32xp33_ASAP7_75t_L g149 ( 
.A1(n_128),
.A2(n_131),
.A3(n_140),
.B1(n_110),
.B2(n_129),
.Y(n_149)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_151),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_136),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_152),
.B(n_112),
.Y(n_156)
);

OAI32xp33_ASAP7_75t_L g154 ( 
.A1(n_128),
.A2(n_114),
.A3(n_102),
.B1(n_105),
.B2(n_107),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_154),
.A2(n_103),
.B1(n_100),
.B2(n_53),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_107),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_141),
.C(n_127),
.Y(n_159)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_146),
.A2(n_131),
.B1(n_130),
.B2(n_133),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_163),
.B1(n_166),
.B2(n_83),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_145),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_79),
.C(n_117),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_165),
.C(n_155),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_105),
.C(n_89),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_158),
.A2(n_149),
.B(n_154),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_167),
.A2(n_173),
.B(n_163),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_169),
.C(n_171),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_153),
.C(n_146),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_165),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_174),
.Y(n_179)
);

AOI322xp5_ASAP7_75t_L g173 ( 
.A1(n_161),
.A2(n_153),
.A3(n_143),
.B1(n_126),
.B2(n_134),
.C1(n_59),
.C2(n_73),
.Y(n_173)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_170),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_177),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_160),
.Y(n_177)
);

NAND4xp25_ASAP7_75t_L g178 ( 
.A(n_173),
.B(n_160),
.C(n_161),
.D(n_164),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_159),
.Y(n_184)
);

AO21x1_ASAP7_75t_L g183 ( 
.A1(n_180),
.A2(n_179),
.B(n_157),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_162),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_182),
.B(n_176),
.Y(n_185)
);

AO21x1_ASAP7_75t_L g187 ( 
.A1(n_183),
.A2(n_65),
.B(n_59),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_184),
.A2(n_175),
.B(n_13),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_185),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_186),
.A2(n_187),
.B(n_181),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_183),
.C(n_73),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_188),
.Y(n_191)
);


endmodule