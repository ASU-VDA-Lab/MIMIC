module fake_jpeg_19973_n_165 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_165);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_8),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_32),
.Y(n_43)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_8),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_41),
.Y(n_48)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_34),
.B(n_19),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_46),
.B(n_55),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_30),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_60),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_24),
.B1(n_15),
.B2(n_27),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_50),
.A2(n_57),
.B1(n_1),
.B2(n_3),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_15),
.B(n_27),
.C(n_30),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_51),
.A2(n_21),
.B1(n_23),
.B2(n_4),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_16),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_53),
.A2(n_3),
.B(n_6),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_41),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_32),
.A2(n_19),
.B1(n_29),
.B2(n_26),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_23),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_29),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_64),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_40),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_65),
.A2(n_69),
.B1(n_85),
.B2(n_52),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_46),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_66),
.B(n_74),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_43),
.A2(n_17),
.B(n_18),
.C(n_20),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_70),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_40),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_43),
.A2(n_17),
.B(n_18),
.C(n_20),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_51),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_84),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_53),
.A2(n_39),
.B(n_2),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_73),
.A2(n_11),
.B(n_12),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_26),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_75),
.A2(n_82),
.B1(n_55),
.B2(n_47),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_14),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_76),
.B(n_79),
.Y(n_91)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_1),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_14),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_83),
.Y(n_102)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_3),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_88),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_61),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_90),
.A2(n_104),
.B1(n_77),
.B2(n_80),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_61),
.C(n_52),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_105),
.C(n_109),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_95),
.A2(n_73),
.B(n_65),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_L g96 ( 
.A1(n_72),
.A2(n_6),
.B(n_7),
.Y(n_96)
);

NOR3xp33_ASAP7_75t_SL g121 ( 
.A(n_96),
.B(n_63),
.C(n_108),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_78),
.B(n_9),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_91),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_71),
.A2(n_54),
.B1(n_62),
.B2(n_47),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_54),
.C(n_62),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_87),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_106),
.A2(n_69),
.B1(n_67),
.B2(n_70),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_108),
.A2(n_81),
.B1(n_83),
.B2(n_63),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_85),
.B(n_86),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_88),
.Y(n_111)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

HAxp5_ASAP7_75t_SL g132 ( 
.A(n_112),
.B(n_121),
.CON(n_132),
.SN(n_132)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_93),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_123),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_100),
.A2(n_75),
.B1(n_69),
.B2(n_84),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_115),
.A2(n_117),
.B1(n_99),
.B2(n_103),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_81),
.Y(n_116)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_124),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_97),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_95),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_125),
.A2(n_92),
.B1(n_113),
.B2(n_106),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_102),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_114),
.A2(n_90),
.B1(n_104),
.B2(n_92),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_134),
.A2(n_117),
.B1(n_131),
.B2(n_126),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_118),
.Y(n_140)
);

AO21x1_ASAP7_75t_L g137 ( 
.A1(n_127),
.A2(n_112),
.B(n_123),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_138),
.Y(n_146)
);

AOI321xp33_ASAP7_75t_L g138 ( 
.A1(n_131),
.A2(n_121),
.A3(n_124),
.B1(n_118),
.B2(n_109),
.C(n_119),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_127),
.A2(n_132),
.B(n_135),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_140),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_129),
.A2(n_120),
.B(n_110),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_145),
.Y(n_148)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_143),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_122),
.B(n_103),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_144),
.A2(n_137),
.B(n_133),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_102),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_144),
.A2(n_130),
.B1(n_128),
.B2(n_134),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_151),
.B(n_136),
.Y(n_155)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_150),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_154),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_143),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_156),
.Y(n_160)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_151),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_148),
.C(n_149),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_158),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_160),
.A2(n_146),
.B(n_147),
.C(n_155),
.Y(n_162)
);

NOR3xp33_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_152),
.C(n_148),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_147),
.C(n_159),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_164),
.Y(n_165)
);


endmodule