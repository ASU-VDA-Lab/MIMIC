module real_jpeg_5625_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_233;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_11;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_188;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_1),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_53)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_1),
.B(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_1),
.A2(n_75),
.B1(n_76),
.B2(n_79),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_1),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_1),
.A2(n_75),
.B1(n_121),
.B2(n_123),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_1),
.B(n_49),
.C(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_1),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_1),
.Y(n_144)
);

O2A1O1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_1),
.A2(n_179),
.B(n_182),
.C(n_185),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_1),
.B(n_176),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_1),
.B(n_118),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_1),
.B(n_102),
.C(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_1),
.B(n_220),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_2),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_2),
.Y(n_86)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_2),
.Y(n_114)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_4),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_4),
.Y(n_176)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_5),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_5),
.Y(n_181)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_7),
.A2(n_19),
.B1(n_25),
.B2(n_26),
.Y(n_18)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_7),
.A2(n_25),
.B1(n_69),
.B2(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_7),
.A2(n_25),
.B1(n_92),
.B2(n_96),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_7),
.A2(n_25),
.B1(n_142),
.B2(n_158),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g143 ( 
.A(n_8),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_8),
.Y(n_145)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_8),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_8),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_8),
.Y(n_160)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_8),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_9),
.Y(n_102)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_9),
.Y(n_104)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_9),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_189),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_188),
.Y(n_11)
);

INVxp67_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_137),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_14),
.B(n_137),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_89),
.C(n_127),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_15),
.A2(n_16),
.B1(n_233),
.B2(n_235),
.Y(n_232)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_58),
.B1(n_59),
.B2(n_88),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_17),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_29),
.B1(n_41),
.B2(n_53),
.Y(n_17)
);

OA22x2_ASAP7_75t_L g165 ( 
.A1(n_18),
.A2(n_29),
.B1(n_41),
.B2(n_53),
.Y(n_165)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2x1_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_41),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_35),
.B1(n_38),
.B2(n_40),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_36),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_41),
.Y(n_220)
);

AOI22x1_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_46),
.B1(n_49),
.B2(n_51),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_45),
.Y(n_126)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_47),
.Y(n_132)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_62)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_54),
.Y(n_184)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp33_ASAP7_75t_L g182 ( 
.A1(n_56),
.A2(n_180),
.B(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_67),
.B2(n_87),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_60),
.B(n_87),
.C(n_88),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_62),
.B(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_62),
.Y(n_161)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_66),
.Y(n_156)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_67),
.B(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_74),
.B1(n_80),
.B2(n_83),
.Y(n_67)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_68),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_68),
.A2(n_74),
.B1(n_83),
.B2(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_73),
.Y(n_68)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_69),
.Y(n_198)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_74),
.B(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_78),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_81),
.B(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_86),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_87),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_87),
.B(n_204),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_89),
.A2(n_219),
.B1(n_221),
.B2(n_222),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_89),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_89),
.B(n_175),
.C(n_219),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_89),
.A2(n_127),
.B1(n_221),
.B2(n_234),
.Y(n_233)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_97),
.B1(n_117),
.B2(n_119),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_91),
.B(n_118),
.Y(n_208)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_95),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_95),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_97),
.B(n_117),
.Y(n_167)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_98),
.B(n_120),
.Y(n_207)
);

NOR2x1_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_107),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_103),
.B2(n_105),
.Y(n_99)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_110),
.B1(n_111),
.B2(n_115),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_120),
.B(n_167),
.Y(n_166)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx5_ASAP7_75t_SL g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_127),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_133),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_128),
.A2(n_129),
.B1(n_133),
.B2(n_134),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_169),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_162),
.B2(n_163),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_140),
.Y(n_139)
);

OA22x2_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_146),
.B1(n_157),
.B2(n_161),
.Y(n_140)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_150),
.B1(n_153),
.B2(n_155),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_168),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_164),
.A2(n_165),
.B1(n_205),
.B2(n_206),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_164),
.B(n_205),
.C(n_228),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_166),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_177),
.B2(n_178),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_174),
.A2(n_175),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_175),
.B(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_201),
.Y(n_202)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

AOI21x1_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_231),
.B(n_237),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_225),
.B(n_230),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_215),
.B(n_224),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_203),
.B(n_214),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_200),
.B(n_202),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_199),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_209),
.B2(n_213),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_213),
.Y(n_223)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

AND2x2_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_209),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_223),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_223),
.Y(n_224)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_219),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_226),
.B(n_227),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_236),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_236),
.Y(n_237)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_233),
.Y(n_235)
);


endmodule