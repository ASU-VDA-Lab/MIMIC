module real_aes_6647_n_350 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_350);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_350;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_800;
wire n_778;
wire n_618;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_357;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_364;
wire n_555;
wire n_766;
wire n_852;
wire n_974;
wire n_919;
wire n_857;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_491;
wire n_1034;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_353;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_537;
wire n_884;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_856;
wire n_594;
wire n_983;
wire n_767;
wire n_889;
wire n_696;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_453;
wire n_374;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1046;
wire n_677;
wire n_958;
wire n_1021;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_961;
wire n_870;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_356;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_994;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_875;
wire n_467;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_746;
wire n_656;
wire n_755;
wire n_532;
wire n_1025;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_725;
wire n_960;
wire n_671;
wire n_973;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1017;
wire n_1013;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_867;
wire n_722;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1037;
wire n_1031;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_985;
wire n_777;
wire n_488;
wire n_501;
wire n_1041;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_713;
wire n_756;
wire n_598;
wire n_735;
wire n_728;
wire n_997;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1000;
wire n_1028;
wire n_1003;
wire n_366;
wire n_727;
wire n_1014;
wire n_649;
wire n_358;
wire n_385;
wire n_397;
wire n_663;
wire n_749;
wire n_588;
wire n_914;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_354;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_978;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_762;
wire n_575;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_836;
wire n_793;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_911;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1024;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx20_ASAP7_75t_R g897 ( .A(n_0), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_1), .A2(n_153), .B1(n_440), .B2(n_444), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_2), .A2(n_157), .B1(n_538), .B2(n_579), .Y(n_933) );
INVx1_ASAP7_75t_L g967 ( .A(n_3), .Y(n_967) );
AOI22xp33_ASAP7_75t_SL g844 ( .A1(n_4), .A2(n_322), .B1(n_400), .B2(n_473), .Y(n_844) );
AOI22xp33_ASAP7_75t_SL g1012 ( .A1(n_5), .A2(n_124), .B1(n_439), .B2(n_444), .Y(n_1012) );
CKINVDCx20_ASAP7_75t_R g1034 ( .A(n_6), .Y(n_1034) );
AOI222xp33_ASAP7_75t_L g804 ( .A1(n_7), .A2(n_178), .B1(n_276), .B2(n_470), .C1(n_487), .C2(n_546), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_8), .A2(n_89), .B1(n_566), .B2(n_649), .Y(n_648) );
AO22x2_ASAP7_75t_L g387 ( .A1(n_9), .A2(n_207), .B1(n_378), .B2(n_383), .Y(n_387) );
INVx1_ASAP7_75t_L g998 ( .A(n_9), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_10), .A2(n_141), .B1(n_499), .B2(n_500), .Y(n_498) );
AOI222xp33_ASAP7_75t_L g1016 ( .A1(n_11), .A2(n_299), .B1(n_309), .B2(n_488), .C1(n_608), .C2(n_678), .Y(n_1016) );
CKINVDCx20_ASAP7_75t_R g981 ( .A(n_12), .Y(n_981) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_13), .A2(n_42), .B1(n_535), .B2(n_980), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_14), .A2(n_119), .B1(n_530), .B2(n_872), .Y(n_902) );
AOI22xp33_ASAP7_75t_SL g689 ( .A1(n_15), .A2(n_112), .B1(n_572), .B2(n_690), .Y(n_689) );
AOI22xp33_ASAP7_75t_SL g677 ( .A1(n_16), .A2(n_265), .B1(n_488), .B2(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g962 ( .A(n_17), .Y(n_962) );
AOI22xp5_ASAP7_75t_SL g813 ( .A1(n_18), .A2(n_181), .B1(n_538), .B2(n_814), .Y(n_813) );
AOI22xp33_ASAP7_75t_SL g686 ( .A1(n_19), .A2(n_242), .B1(n_656), .B2(n_687), .Y(n_686) );
AOI22xp33_ASAP7_75t_SL g654 ( .A1(n_20), .A2(n_195), .B1(n_655), .B2(n_656), .Y(n_654) );
AOI22xp33_ASAP7_75t_SL g968 ( .A1(n_21), .A2(n_182), .B1(n_490), .B2(n_545), .Y(n_968) );
AOI221xp5_ASAP7_75t_L g785 ( .A1(n_22), .A2(n_102), .B1(n_399), .B2(n_476), .C(n_786), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g1015 ( .A1(n_23), .A2(n_145), .B1(n_570), .B2(n_741), .Y(n_1015) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_24), .A2(n_293), .B1(n_533), .B2(n_535), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_25), .A2(n_104), .B1(n_697), .B2(n_956), .Y(n_955) );
AOI22xp33_ASAP7_75t_SL g651 ( .A1(n_26), .A2(n_128), .B1(n_502), .B2(n_652), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_27), .A2(n_232), .B1(n_444), .B2(n_602), .Y(n_601) );
AO22x2_ASAP7_75t_L g385 ( .A1(n_28), .A2(n_111), .B1(n_378), .B2(n_379), .Y(n_385) );
AOI22xp33_ASAP7_75t_SL g841 ( .A1(n_29), .A2(n_251), .B1(n_482), .B2(n_500), .Y(n_841) );
AOI222xp33_ASAP7_75t_L g513 ( .A1(n_30), .A2(n_179), .B1(n_275), .B2(n_443), .C1(n_490), .C2(n_514), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_31), .A2(n_287), .B1(n_511), .B2(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_32), .B(n_647), .Y(n_646) );
CKINVDCx20_ASAP7_75t_R g898 ( .A(n_33), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_34), .A2(n_61), .B1(n_482), .B2(n_528), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_35), .A2(n_241), .B1(n_570), .B2(n_571), .Y(n_569) );
CKINVDCx20_ASAP7_75t_R g943 ( .A(n_36), .Y(n_943) );
AOI221xp5_ASAP7_75t_L g797 ( .A1(n_37), .A2(n_192), .B1(n_798), .B2(n_799), .C(n_800), .Y(n_797) );
AOI22xp33_ASAP7_75t_SL g684 ( .A1(n_38), .A2(n_113), .B1(n_476), .B2(n_685), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_39), .A2(n_164), .B1(n_528), .B2(n_659), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g895 ( .A(n_40), .B(n_641), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_41), .A2(n_85), .B1(n_482), .B2(n_484), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_43), .A2(n_132), .B1(n_697), .B2(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g868 ( .A(n_44), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_45), .A2(n_73), .B1(n_538), .B2(n_655), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_46), .A2(n_95), .B1(n_511), .B2(n_524), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g978 ( .A1(n_47), .A2(n_213), .B1(n_482), .B2(n_875), .Y(n_978) );
AOI222xp33_ASAP7_75t_L g447 ( .A1(n_48), .A2(n_165), .B1(n_318), .B2(n_448), .C1(n_449), .C2(n_453), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_49), .A2(n_84), .B1(n_537), .B2(n_1008), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_50), .A2(n_286), .B1(n_616), .B2(n_875), .Y(n_959) );
INVx1_ASAP7_75t_L g795 ( .A(n_51), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_52), .A2(n_173), .B1(n_602), .B2(n_649), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_53), .A2(n_69), .B1(n_507), .B2(n_541), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_54), .A2(n_338), .B1(n_537), .B2(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g846 ( .A(n_55), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g1011 ( .A(n_56), .B(n_507), .Y(n_1011) );
AOI22xp33_ASAP7_75t_SL g658 ( .A1(n_57), .A2(n_348), .B1(n_399), .B2(n_659), .Y(n_658) );
AOI22xp33_ASAP7_75t_SL g845 ( .A1(n_58), .A2(n_211), .B1(n_484), .B2(n_511), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_59), .A2(n_313), .B1(n_409), .B2(n_416), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_60), .A2(n_305), .B1(n_624), .B2(n_625), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_62), .A2(n_344), .B1(n_443), .B2(n_602), .Y(n_863) );
CKINVDCx20_ASAP7_75t_R g951 ( .A(n_63), .Y(n_951) );
CKINVDCx20_ASAP7_75t_R g1037 ( .A(n_64), .Y(n_1037) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_65), .A2(n_189), .B1(n_535), .B2(n_624), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_66), .A2(n_106), .B1(n_487), .B2(n_526), .Y(n_1041) );
AOI22xp33_ASAP7_75t_SL g842 ( .A1(n_67), .A2(n_238), .B1(n_476), .B2(n_503), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_68), .A2(n_260), .B1(n_444), .B2(n_543), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g919 ( .A(n_70), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_71), .A2(n_187), .B1(n_655), .B2(n_656), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_72), .A2(n_234), .B1(n_482), .B2(n_741), .Y(n_740) );
AOI221xp5_ASAP7_75t_L g791 ( .A1(n_74), .A2(n_98), .B1(n_528), .B2(n_616), .C(n_792), .Y(n_791) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_75), .Y(n_388) );
AO22x2_ASAP7_75t_L g382 ( .A1(n_76), .A2(n_240), .B1(n_378), .B2(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g995 ( .A(n_76), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_77), .A2(n_81), .B1(n_530), .B2(n_582), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_78), .A2(n_94), .B1(n_528), .B2(n_530), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_79), .A2(n_137), .B1(n_565), .B2(n_566), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_80), .A2(n_219), .B1(n_476), .B2(n_523), .Y(n_772) );
AOI211xp5_ASAP7_75t_L g350 ( .A1(n_82), .A2(n_351), .B(n_360), .C(n_1000), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_83), .A2(n_202), .B1(n_558), .B2(n_566), .Y(n_822) );
AOI22xp33_ASAP7_75t_SL g838 ( .A1(n_86), .A2(n_254), .B1(n_440), .B2(n_545), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_87), .A2(n_174), .B1(n_644), .B2(n_702), .Y(n_701) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_88), .Y(n_723) );
AOI22xp5_ASAP7_75t_L g366 ( .A1(n_90), .A2(n_367), .B1(n_457), .B2(n_458), .Y(n_366) );
CKINVDCx16_ASAP7_75t_R g457 ( .A(n_90), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_91), .Y(n_756) );
AOI222xp33_ASAP7_75t_L g486 ( .A1(n_92), .A2(n_107), .B1(n_167), .B2(n_487), .C1(n_488), .C2(n_491), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_93), .A2(n_341), .B1(n_439), .B2(n_470), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_96), .A2(n_592), .B1(n_628), .B2(n_629), .Y(n_591) );
CKINVDCx20_ASAP7_75t_R g628 ( .A(n_96), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_97), .A2(n_244), .B1(n_511), .B2(n_524), .Y(n_769) );
CKINVDCx20_ASAP7_75t_R g1038 ( .A(n_99), .Y(n_1038) );
CKINVDCx20_ASAP7_75t_R g1032 ( .A(n_100), .Y(n_1032) );
INVx1_ASAP7_75t_L g801 ( .A(n_101), .Y(n_801) );
XOR2x2_ASAP7_75t_L g549 ( .A(n_103), .B(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g825 ( .A(n_105), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_108), .A2(n_259), .B1(n_404), .B2(n_685), .Y(n_1014) );
CKINVDCx20_ASAP7_75t_R g833 ( .A(n_109), .Y(n_833) );
AOI22xp5_ASAP7_75t_L g812 ( .A1(n_110), .A2(n_249), .B1(n_374), .B2(n_473), .Y(n_812) );
INVx1_ASAP7_75t_L g999 ( .A(n_111), .Y(n_999) );
AOI22xp5_ASAP7_75t_L g817 ( .A1(n_114), .A2(n_279), .B1(n_399), .B2(n_818), .Y(n_817) );
CKINVDCx20_ASAP7_75t_R g888 ( .A(n_115), .Y(n_888) );
XOR2x2_ASAP7_75t_L g671 ( .A(n_116), .B(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_117), .B(n_563), .Y(n_562) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_118), .Y(n_432) );
AO22x1_ASAP7_75t_L g518 ( .A1(n_120), .A2(n_519), .B1(n_520), .B2(n_547), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_120), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_121), .A2(n_139), .B1(n_421), .B2(n_424), .Y(n_957) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_122), .B(n_561), .Y(n_560) );
CKINVDCx20_ASAP7_75t_R g766 ( .A(n_123), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_125), .A2(n_311), .B1(n_455), .B2(n_566), .Y(n_1035) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_126), .A2(n_321), .B1(n_400), .B2(n_413), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g597 ( .A(n_127), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g783 ( .A1(n_129), .A2(n_784), .B1(n_805), .B2(n_806), .Y(n_783) );
INVx1_ASAP7_75t_L g805 ( .A(n_129), .Y(n_805) );
OAI22xp5_ASAP7_75t_SL g883 ( .A1(n_130), .A2(n_884), .B1(n_885), .B2(n_907), .Y(n_883) );
CKINVDCx20_ASAP7_75t_R g907 ( .A(n_130), .Y(n_907) );
INVx1_ASAP7_75t_L g793 ( .A(n_131), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_133), .A2(n_319), .B1(n_583), .B2(n_687), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_134), .A2(n_151), .B1(n_624), .B2(n_932), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_135), .A2(n_210), .B1(n_625), .B2(n_692), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_136), .A2(n_149), .B1(n_537), .B2(n_538), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_138), .A2(n_331), .B1(n_416), .B2(n_574), .Y(n_573) );
CKINVDCx20_ASAP7_75t_R g894 ( .A(n_140), .Y(n_894) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_142), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_143), .A2(n_194), .B1(n_439), .B2(n_443), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_144), .A2(n_280), .B1(n_530), .B2(n_956), .Y(n_1006) );
AND2x6_ASAP7_75t_L g355 ( .A(n_146), .B(n_356), .Y(n_355) );
HB1xp67_ASAP7_75t_L g992 ( .A(n_146), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_147), .A2(n_264), .B1(n_579), .B2(n_583), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_148), .A2(n_306), .B1(n_470), .B2(n_490), .Y(n_949) );
AOI22xp33_ASAP7_75t_SL g637 ( .A1(n_150), .A2(n_245), .B1(n_638), .B2(n_641), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_152), .A2(n_177), .B1(n_500), .B2(n_980), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_154), .A2(n_253), .B1(n_449), .B2(n_741), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_155), .A2(n_297), .B1(n_579), .B2(n_621), .Y(n_738) );
AOI222xp33_ASAP7_75t_L g876 ( .A1(n_156), .A2(n_224), .B1(n_239), .B2(n_448), .C1(n_470), .C2(n_641), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_158), .A2(n_285), .B1(n_697), .B2(n_698), .Y(n_696) );
AOI22xp33_ASAP7_75t_SL g661 ( .A1(n_159), .A2(n_316), .B1(n_372), .B2(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g877 ( .A(n_160), .Y(n_877) );
AOI22xp33_ASAP7_75t_SL g976 ( .A1(n_161), .A2(n_333), .B1(n_421), .B2(n_503), .Y(n_976) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_162), .A2(n_290), .B1(n_662), .B2(n_698), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_163), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_166), .A2(n_229), .B1(n_578), .B2(n_579), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_168), .A2(n_324), .B1(n_404), .B2(n_961), .Y(n_960) );
AO22x2_ASAP7_75t_L g377 ( .A1(n_169), .A2(n_230), .B1(n_378), .B2(n_379), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g996 ( .A(n_169), .B(n_997), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_170), .A2(n_200), .B1(n_582), .B2(n_583), .Y(n_581) );
CKINVDCx20_ASAP7_75t_R g1010 ( .A(n_171), .Y(n_1010) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_172), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_175), .A2(n_340), .B1(n_578), .B2(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g636 ( .A(n_176), .Y(n_636) );
CKINVDCx20_ASAP7_75t_R g676 ( .A(n_180), .Y(n_676) );
AOI222xp33_ASAP7_75t_L g544 ( .A1(n_183), .A2(n_304), .B1(n_315), .B2(n_487), .C1(n_545), .C2(n_546), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_184), .B(n_454), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_185), .A2(n_233), .B1(n_526), .B2(n_530), .Y(n_705) );
CKINVDCx20_ASAP7_75t_R g890 ( .A(n_186), .Y(n_890) );
XOR2x2_ASAP7_75t_L g460 ( .A(n_188), .B(n_461), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_190), .A2(n_282), .B1(n_464), .B2(n_644), .Y(n_821) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_191), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_193), .Y(n_437) );
INVx1_ASAP7_75t_L g870 ( .A(n_196), .Y(n_870) );
CKINVDCx20_ASAP7_75t_R g619 ( .A(n_197), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_198), .A2(n_278), .B1(n_464), .B2(n_467), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_199), .B(n_464), .Y(n_836) );
CKINVDCx20_ASAP7_75t_R g370 ( .A(n_201), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_203), .A2(n_248), .B1(n_400), .B2(n_421), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_204), .B(n_644), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_205), .A2(n_272), .B1(n_476), .B2(n_478), .Y(n_475) );
AOI22xp33_ASAP7_75t_SL g834 ( .A1(n_206), .A2(n_228), .B1(n_454), .B2(n_649), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_208), .A2(n_263), .B1(n_502), .B2(n_503), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_209), .A2(n_273), .B1(n_491), .B2(n_602), .Y(n_682) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_212), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_214), .A2(n_339), .B1(n_424), .B2(n_473), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g397 ( .A(n_215), .Y(n_397) );
CKINVDCx20_ASAP7_75t_R g914 ( .A(n_216), .Y(n_914) );
INVx1_ASAP7_75t_L g866 ( .A(n_217), .Y(n_866) );
INVx1_ASAP7_75t_L g1024 ( .A(n_218), .Y(n_1024) );
OA22x2_ASAP7_75t_L g1027 ( .A1(n_218), .A2(n_1024), .B1(n_1028), .B2(n_1046), .Y(n_1027) );
INVx1_ASAP7_75t_L g803 ( .A(n_220), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_221), .A2(n_308), .B1(n_439), .B2(n_470), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_222), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_223), .A2(n_243), .B1(n_421), .B2(n_424), .Y(n_420) );
AOI222xp33_ASAP7_75t_L g708 ( .A1(n_225), .A2(n_323), .B1(n_334), .B2(n_448), .C1(n_545), .C2(n_546), .Y(n_708) );
INVx2_ASAP7_75t_L g359 ( .A(n_226), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_227), .A2(n_261), .B1(n_454), .B2(n_556), .Y(n_555) );
CKINVDCx20_ASAP7_75t_R g606 ( .A(n_231), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_235), .A2(n_277), .B1(n_449), .B2(n_490), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_236), .A2(n_337), .B1(n_523), .B2(n_524), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_237), .Y(n_758) );
INVx1_ASAP7_75t_L g952 ( .A(n_246), .Y(n_952) );
CKINVDCx20_ASAP7_75t_R g892 ( .A(n_247), .Y(n_892) );
CKINVDCx20_ASAP7_75t_R g610 ( .A(n_250), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g751 ( .A1(n_252), .A2(n_752), .B1(n_774), .B2(n_775), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_252), .Y(n_774) );
AOI22xp33_ASAP7_75t_SL g691 ( .A1(n_255), .A2(n_347), .B1(n_499), .B2(n_692), .Y(n_691) );
XOR2x2_ASAP7_75t_L g632 ( .A(n_256), .B(n_633), .Y(n_632) );
CKINVDCx20_ASAP7_75t_R g1031 ( .A(n_257), .Y(n_1031) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_258), .Y(n_721) );
INVx1_ASAP7_75t_L g378 ( .A(n_262), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_262), .Y(n_380) );
CKINVDCx20_ASAP7_75t_R g617 ( .A(n_266), .Y(n_617) );
CKINVDCx20_ASAP7_75t_R g600 ( .A(n_267), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_268), .B(n_507), .Y(n_681) );
CKINVDCx20_ASAP7_75t_R g915 ( .A(n_269), .Y(n_915) );
INVx1_ASAP7_75t_L g790 ( .A(n_270), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_271), .B(n_467), .Y(n_970) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_274), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g922 ( .A(n_281), .Y(n_922) );
CKINVDCx20_ASAP7_75t_R g402 ( .A(n_283), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g971 ( .A(n_284), .B(n_798), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_288), .A2(n_346), .B1(n_468), .B2(n_507), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_289), .A2(n_325), .B1(n_743), .B2(n_745), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_291), .Y(n_737) );
INVx1_ASAP7_75t_L g358 ( .A(n_292), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_294), .B(n_762), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g918 ( .A(n_295), .Y(n_918) );
INVx1_ASAP7_75t_L g356 ( .A(n_296), .Y(n_356) );
INVx1_ASAP7_75t_L g827 ( .A(n_298), .Y(n_827) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_300), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_301), .A2(n_307), .B1(n_473), .B2(n_511), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g947 ( .A(n_302), .Y(n_947) );
INVx1_ASAP7_75t_L g873 ( .A(n_303), .Y(n_873) );
XOR2xp5_ASAP7_75t_L g1001 ( .A(n_310), .B(n_1002), .Y(n_1001) );
CKINVDCx20_ASAP7_75t_R g924 ( .A(n_312), .Y(n_924) );
INVx1_ASAP7_75t_L g787 ( .A(n_314), .Y(n_787) );
CKINVDCx20_ASAP7_75t_R g612 ( .A(n_317), .Y(n_612) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_320), .Y(n_764) );
INVx1_ASAP7_75t_L g859 ( .A(n_326), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_327), .B(n_467), .Y(n_837) );
AOI22xp33_ASAP7_75t_SL g975 ( .A1(n_328), .A2(n_343), .B1(n_526), .B2(n_961), .Y(n_975) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_329), .B(n_644), .Y(n_680) );
XOR2x2_ASAP7_75t_L g693 ( .A(n_330), .B(n_694), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_332), .A2(n_710), .B1(n_746), .B2(n_747), .Y(n_709) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_332), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_335), .B(n_862), .Y(n_861) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_336), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_342), .Y(n_717) );
AOI22xp5_ASAP7_75t_L g910 ( .A1(n_345), .A2(n_911), .B1(n_934), .B2(n_935), .Y(n_910) );
INVx1_ASAP7_75t_L g934 ( .A(n_345), .Y(n_934) );
CKINVDCx20_ASAP7_75t_R g945 ( .A(n_349), .Y(n_945) );
CKINVDCx20_ASAP7_75t_R g351 ( .A(n_352), .Y(n_351) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_353), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x4_ASAP7_75t_L g354 ( .A(n_355), .B(n_357), .Y(n_354) );
HB1xp67_ASAP7_75t_L g991 ( .A(n_356), .Y(n_991) );
OAI21xp5_ASAP7_75t_L g1022 ( .A1(n_357), .A2(n_990), .B(n_1023), .Y(n_1022) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
AOI221xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_779), .B1(n_985), .B2(n_986), .C(n_987), .Y(n_360) );
INVx1_ASAP7_75t_L g985 ( .A(n_361), .Y(n_985) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_363), .B1(n_587), .B2(n_778), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_365), .B1(n_494), .B2(n_586), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_459), .B1(n_492), .B2(n_493), .Y(n_365) );
INVx1_ASAP7_75t_L g492 ( .A(n_366), .Y(n_492) );
INVx2_ASAP7_75t_SL g458 ( .A(n_367), .Y(n_458) );
AND4x1_ASAP7_75t_L g367 ( .A(n_368), .B(n_407), .C(n_427), .D(n_447), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_369), .B(n_396), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_371), .B1(n_388), .B2(n_389), .Y(n_369) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g578 ( .A(n_373), .Y(n_578) );
INVx2_ASAP7_75t_L g625 ( .A(n_373), .Y(n_625) );
INVx3_ASAP7_75t_L g875 ( .A(n_373), .Y(n_875) );
INVx6_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
BUFx3_ASAP7_75t_L g484 ( .A(n_374), .Y(n_484) );
BUFx3_ASAP7_75t_L g499 ( .A(n_374), .Y(n_499) );
BUFx3_ASAP7_75t_L g741 ( .A(n_374), .Y(n_741) );
AND2x4_ASAP7_75t_L g374 ( .A(n_375), .B(n_384), .Y(n_374) );
AND2x2_ASAP7_75t_L g401 ( .A(n_375), .B(n_394), .Y(n_401) );
AND2x6_ASAP7_75t_L g413 ( .A(n_375), .B(n_414), .Y(n_413) );
AND2x6_ASAP7_75t_L g448 ( .A(n_375), .B(n_446), .Y(n_448) );
AND2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_381), .Y(n_375) );
AND2x2_ASAP7_75t_L g406 ( .A(n_376), .B(n_382), .Y(n_406) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g392 ( .A(n_377), .B(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_377), .B(n_382), .Y(n_419) );
AND2x2_ASAP7_75t_L g442 ( .A(n_377), .B(n_387), .Y(n_442) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g383 ( .A(n_380), .Y(n_383) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g393 ( .A(n_382), .Y(n_393) );
INVx1_ASAP7_75t_L g452 ( .A(n_382), .Y(n_452) );
AND2x2_ASAP7_75t_L g423 ( .A(n_384), .B(n_392), .Y(n_423) );
NAND2x1p5_ASAP7_75t_L g436 ( .A(n_384), .B(n_406), .Y(n_436) );
AND2x6_ASAP7_75t_L g468 ( .A(n_384), .B(n_406), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g789 ( .A(n_384), .B(n_392), .Y(n_789) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
INVx2_ASAP7_75t_L g395 ( .A(n_385), .Y(n_395) );
OR2x2_ASAP7_75t_L g415 ( .A(n_385), .B(n_386), .Y(n_415) );
INVx1_ASAP7_75t_L g426 ( .A(n_385), .Y(n_426) );
AND2x2_ASAP7_75t_L g446 ( .A(n_385), .B(n_387), .Y(n_446) );
AND2x2_ASAP7_75t_L g394 ( .A(n_386), .B(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g865 ( .A1(n_389), .A2(n_866), .B1(n_867), .B2(n_868), .Y(n_865) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g794 ( .A(n_390), .Y(n_794) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_392), .B(n_394), .Y(n_391) );
AND2x2_ASAP7_75t_L g474 ( .A(n_392), .B(n_394), .Y(n_474) );
INVx1_ASAP7_75t_L g445 ( .A(n_393), .Y(n_445) );
AND2x4_ASAP7_75t_L g405 ( .A(n_394), .B(n_406), .Y(n_405) );
AND2x4_ASAP7_75t_L g417 ( .A(n_394), .B(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g451 ( .A(n_395), .B(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g504 ( .A(n_395), .Y(n_504) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_398), .B1(n_402), .B2(n_403), .Y(n_396) );
INVx1_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
BUFx3_ASAP7_75t_L g523 ( .A(n_400), .Y(n_523) );
BUFx3_ASAP7_75t_L g624 ( .A(n_400), .Y(n_624) );
BUFx6f_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g575 ( .A(n_401), .Y(n_575) );
BUFx2_ASAP7_75t_SL g685 ( .A(n_401), .Y(n_685) );
BUFx2_ASAP7_75t_SL g697 ( .A(n_401), .Y(n_697) );
INVxp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx3_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g477 ( .A(n_405), .Y(n_477) );
BUFx6f_ASAP7_75t_L g502 ( .A(n_405), .Y(n_502) );
BUFx3_ASAP7_75t_L g535 ( .A(n_405), .Y(n_535) );
BUFx3_ASAP7_75t_L g582 ( .A(n_405), .Y(n_582) );
INVx1_ASAP7_75t_L g431 ( .A(n_406), .Y(n_431) );
AND2x4_ASAP7_75t_L g466 ( .A(n_406), .B(n_414), .Y(n_466) );
AND2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_420), .Y(n_407) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx5_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_412), .Y(n_534) );
INVx2_ASAP7_75t_SL g570 ( .A(n_412), .Y(n_570) );
INVx4_ASAP7_75t_L g616 ( .A(n_412), .Y(n_616) );
INVx1_ASAP7_75t_L g707 ( .A(n_412), .Y(n_707) );
INVx2_ASAP7_75t_L g818 ( .A(n_412), .Y(n_818) );
INVx11_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx11_ASAP7_75t_L g483 ( .A(n_413), .Y(n_483) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g430 ( .A(n_415), .B(n_431), .Y(n_430) );
BUFx3_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g479 ( .A(n_417), .Y(n_479) );
BUFx3_ASAP7_75t_L g511 ( .A(n_417), .Y(n_511) );
BUFx3_ASAP7_75t_L g530 ( .A(n_417), .Y(n_530) );
BUFx2_ASAP7_75t_SL g662 ( .A(n_417), .Y(n_662) );
BUFx2_ASAP7_75t_SL g690 ( .A(n_417), .Y(n_690) );
BUFx3_ASAP7_75t_L g745 ( .A(n_417), .Y(n_745) );
BUFx2_ASAP7_75t_L g961 ( .A(n_417), .Y(n_961) );
AND2x2_ASAP7_75t_L g503 ( .A(n_418), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
OR2x6_ASAP7_75t_L g425 ( .A(n_419), .B(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx5_ASAP7_75t_L g500 ( .A(n_422), .Y(n_500) );
INVx3_ASAP7_75t_L g537 ( .A(n_422), .Y(n_537) );
BUFx3_ASAP7_75t_L g580 ( .A(n_422), .Y(n_580) );
INVx4_ASAP7_75t_L g815 ( .A(n_422), .Y(n_815) );
INVx8_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx2_ASAP7_75t_L g538 ( .A(n_424), .Y(n_538) );
BUFx2_ASAP7_75t_L g583 ( .A(n_424), .Y(n_583) );
BUFx2_ASAP7_75t_L g656 ( .A(n_424), .Y(n_656) );
BUFx2_ASAP7_75t_L g1008 ( .A(n_424), .Y(n_1008) );
INVx6_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_SL g621 ( .A(n_425), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g786 ( .A1(n_425), .A2(n_787), .B1(n_788), .B2(n_790), .Y(n_786) );
OAI22xp5_ASAP7_75t_L g1036 ( .A1(n_425), .A2(n_730), .B1(n_1037), .B2(n_1038), .Y(n_1036) );
INVx1_ASAP7_75t_L g441 ( .A(n_426), .Y(n_441) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OAI221xp5_ASAP7_75t_SL g428 ( .A1(n_429), .A2(n_432), .B1(n_433), .B2(n_437), .C(n_438), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_429), .A2(n_433), .B1(n_713), .B2(n_714), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g913 ( .A1(n_429), .A2(n_914), .B1(n_915), .B2(n_916), .Y(n_913) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g596 ( .A(n_430), .Y(n_596) );
BUFx3_ASAP7_75t_L g944 ( .A(n_430), .Y(n_944) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_433), .A2(n_595), .B1(n_755), .B2(n_756), .Y(n_754) );
OAI22xp5_ASAP7_75t_L g887 ( .A1(n_433), .A2(n_888), .B1(n_889), .B2(n_890), .Y(n_887) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx3_ASAP7_75t_L g860 ( .A(n_435), .Y(n_860) );
BUFx3_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g599 ( .A(n_436), .Y(n_599) );
BUFx3_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx2_ASAP7_75t_L g543 ( .A(n_440), .Y(n_543) );
BUFx2_ASAP7_75t_L g566 ( .A(n_440), .Y(n_566) );
INVx1_ASAP7_75t_L g603 ( .A(n_440), .Y(n_603) );
AND2x4_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
AND2x4_ASAP7_75t_L g450 ( .A(n_442), .B(n_451), .Y(n_450) );
AND2x4_ASAP7_75t_L g455 ( .A(n_442), .B(n_456), .Y(n_455) );
NAND2x1p5_ASAP7_75t_L g726 ( .A(n_442), .B(n_504), .Y(n_726) );
BUFx3_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
BUFx2_ASAP7_75t_SL g491 ( .A(n_444), .Y(n_491) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_444), .Y(n_558) );
BUFx2_ASAP7_75t_SL g649 ( .A(n_444), .Y(n_649) );
AND2x4_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
INVx1_ASAP7_75t_L g732 ( .A(n_445), .Y(n_732) );
INVx1_ASAP7_75t_L g731 ( .A(n_446), .Y(n_731) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_448), .Y(n_487) );
BUFx3_ASAP7_75t_L g514 ( .A(n_448), .Y(n_514) );
INVx2_ASAP7_75t_SL g553 ( .A(n_448), .Y(n_553) );
INVx4_ASAP7_75t_L g609 ( .A(n_448), .Y(n_609) );
INVx2_ASAP7_75t_L g832 ( .A(n_448), .Y(n_832) );
BUFx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_450), .Y(n_470) );
BUFx4f_ASAP7_75t_SL g545 ( .A(n_450), .Y(n_545) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_450), .Y(n_565) );
BUFx6f_ASAP7_75t_L g640 ( .A(n_450), .Y(n_640) );
INVx1_ASAP7_75t_L g456 ( .A(n_452), .Y(n_456) );
BUFx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g720 ( .A(n_454), .Y(n_720) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx12f_ASAP7_75t_L g490 ( .A(n_455), .Y(n_490) );
BUFx6f_ASAP7_75t_L g641 ( .A(n_455), .Y(n_641) );
INVxp67_ASAP7_75t_L g493 ( .A(n_459), .Y(n_493) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
XOR2x2_ASAP7_75t_L g548 ( .A(n_460), .B(n_549), .Y(n_548) );
NAND4xp75_ASAP7_75t_L g461 ( .A(n_462), .B(n_471), .C(n_480), .D(n_486), .Y(n_461) );
AND2x2_ASAP7_75t_SL g462 ( .A(n_463), .B(n_469), .Y(n_462) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx5_ASAP7_75t_L g507 ( .A(n_465), .Y(n_507) );
INVx2_ASAP7_75t_L g647 ( .A(n_465), .Y(n_647) );
INVx2_ASAP7_75t_L g798 ( .A(n_465), .Y(n_798) );
INVx4_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
BUFx4f_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
BUFx2_ASAP7_75t_L g541 ( .A(n_468), .Y(n_541) );
BUFx2_ASAP7_75t_L g563 ( .A(n_468), .Y(n_563) );
INVx1_ASAP7_75t_SL g645 ( .A(n_468), .Y(n_645) );
BUFx6f_ASAP7_75t_L g678 ( .A(n_470), .Y(n_678) );
AND2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_475), .Y(n_471) );
INVx1_ASAP7_75t_L g660 ( .A(n_473), .Y(n_660) );
BUFx3_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx3_ASAP7_75t_L g526 ( .A(n_474), .Y(n_526) );
BUFx3_ASAP7_75t_L g572 ( .A(n_474), .Y(n_572) );
BUFx3_ASAP7_75t_L g956 ( .A(n_474), .Y(n_956) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_485), .Y(n_480) );
INVx4_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_SL g692 ( .A(n_483), .Y(n_692) );
INVx3_ASAP7_75t_L g872 ( .A(n_483), .Y(n_872) );
OAI21xp33_ASAP7_75t_SL g1033 ( .A1(n_483), .A2(n_1034), .B(n_1035), .Y(n_1033) );
INVx2_ASAP7_75t_SL g675 ( .A(n_487), .Y(n_675) );
INVx2_ASAP7_75t_L g718 ( .A(n_487), .Y(n_718) );
INVx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx4f_ASAP7_75t_SL g546 ( .A(n_490), .Y(n_546) );
INVx1_ASAP7_75t_L g586 ( .A(n_494), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_516), .B1(n_584), .B2(n_585), .Y(n_494) );
INVx2_ASAP7_75t_SL g584 ( .A(n_495), .Y(n_584) );
XOR2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_515), .Y(n_495) );
NAND4xp75_ASAP7_75t_L g496 ( .A(n_497), .B(n_505), .C(n_509), .D(n_513), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_501), .Y(n_497) );
INVx3_ASAP7_75t_L g529 ( .A(n_499), .Y(n_529) );
BUFx2_ASAP7_75t_L g655 ( .A(n_500), .Y(n_655) );
BUFx6f_ASAP7_75t_L g687 ( .A(n_500), .Y(n_687) );
INVx4_ASAP7_75t_L g618 ( .A(n_502), .Y(n_618) );
AND2x2_ASAP7_75t_SL g505 ( .A(n_506), .B(n_508), .Y(n_505) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_507), .Y(n_561) );
BUFx6f_ASAP7_75t_L g702 ( .A(n_507), .Y(n_702) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_512), .Y(n_509) );
INVx3_ASAP7_75t_L g948 ( .A(n_514), .Y(n_948) );
INVx2_ASAP7_75t_L g585 ( .A(n_516), .Y(n_585) );
XNOR2x1_ASAP7_75t_L g516 ( .A(n_517), .B(n_548), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_SL g519 ( .A(n_520), .Y(n_519) );
NAND4xp75_ASAP7_75t_SL g520 ( .A(n_521), .B(n_531), .C(n_539), .D(n_544), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_527), .Y(n_521) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx2_ASAP7_75t_L g627 ( .A(n_526), .Y(n_627) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVxp67_ASAP7_75t_L g867 ( .A(n_530), .Y(n_867) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_536), .Y(n_531) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_SL g539 ( .A(n_540), .B(n_542), .Y(n_539) );
INVx1_ASAP7_75t_L g716 ( .A(n_545), .Y(n_716) );
INVx1_ASAP7_75t_L g759 ( .A(n_545), .Y(n_759) );
INVx1_ASAP7_75t_L g611 ( .A(n_546), .Y(n_611) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_551), .B(n_567), .Y(n_550) );
NOR2xp33_ASAP7_75t_SL g551 ( .A(n_552), .B(n_559), .Y(n_551) );
OAI21xp5_ASAP7_75t_SL g552 ( .A1(n_553), .A2(n_554), .B(n_555), .Y(n_552) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
NAND3xp33_ASAP7_75t_L g559 ( .A(n_560), .B(n_562), .C(n_564), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g605 ( .A(n_565), .Y(n_605) );
NOR2x1_ASAP7_75t_L g567 ( .A(n_568), .B(n_576), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_573), .Y(n_568) );
INVx1_ASAP7_75t_L g653 ( .A(n_570), .Y(n_653) );
BUFx4f_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g744 ( .A(n_572), .Y(n_744) );
INVx3_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx3_ASAP7_75t_L g980 ( .A(n_575), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_581), .Y(n_576) );
INVx3_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
HB1xp67_ASAP7_75t_L g932 ( .A(n_582), .Y(n_932) );
INVx1_ASAP7_75t_L g778 ( .A(n_587), .Y(n_778) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_589), .B1(n_665), .B2(n_666), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OAI22xp5_ASAP7_75t_SL g589 ( .A1(n_590), .A2(n_630), .B1(n_663), .B2(n_664), .Y(n_589) );
INVx1_ASAP7_75t_L g663 ( .A(n_590), .Y(n_663) );
INVx1_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g629 ( .A(n_592), .Y(n_629) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_613), .Y(n_592) );
NOR2xp33_ASAP7_75t_SL g593 ( .A(n_594), .B(n_604), .Y(n_593) );
OAI221xp5_ASAP7_75t_SL g594 ( .A1(n_595), .A2(n_597), .B1(n_598), .B2(n_600), .C(n_601), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_SL g889 ( .A(n_596), .Y(n_889) );
OAI22xp5_ASAP7_75t_L g942 ( .A1(n_598), .A2(n_943), .B1(n_944), .B2(n_945), .Y(n_942) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_SL g916 ( .A(n_599), .Y(n_916) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OAI222xp33_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_606), .B1(n_607), .B2(n_610), .C1(n_611), .C2(n_612), .Y(n_604) );
OAI21xp5_ASAP7_75t_SL g635 ( .A1(n_607), .A2(n_636), .B(n_637), .Y(n_635) );
OAI221xp5_ASAP7_75t_SL g891 ( .A1(n_607), .A2(n_892), .B1(n_893), .B2(n_894), .C(n_895), .Y(n_891) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx4_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
BUFx2_ASAP7_75t_L g824 ( .A(n_609), .Y(n_824) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_614), .B(n_622), .Y(n_613) );
OAI221xp5_ASAP7_75t_SL g614 ( .A1(n_615), .A2(n_617), .B1(n_618), .B2(n_619), .C(n_620), .Y(n_614) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
INVx4_ASAP7_75t_L g698 ( .A(n_618), .Y(n_698) );
OAI221xp5_ASAP7_75t_SL g734 ( .A1(n_618), .A2(n_735), .B1(n_736), .B2(n_737), .C(n_738), .Y(n_734) );
INVx3_ASAP7_75t_L g856 ( .A(n_618), .Y(n_856) );
NAND2xp33_ASAP7_75t_SL g622 ( .A(n_623), .B(n_626), .Y(n_622) );
INVx1_ASAP7_75t_L g664 ( .A(n_630), .Y(n_664) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND3x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_650), .C(n_657), .Y(n_633) );
NOR2x1_ASAP7_75t_SL g634 ( .A(n_635), .B(n_642), .Y(n_634) );
INVx3_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx4_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
BUFx4f_ASAP7_75t_L g762 ( .A(n_641), .Y(n_762) );
NAND3xp33_ASAP7_75t_L g642 ( .A(n_643), .B(n_646), .C(n_648), .Y(n_642) );
INVx1_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_SL g799 ( .A(n_645), .Y(n_799) );
AND2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_654), .Y(n_650) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_661), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_668), .B1(n_749), .B2(n_750), .Y(n_666) );
INVx1_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_670), .B1(n_709), .B2(n_748), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
XNOR2xp5_ASAP7_75t_L g670 ( .A(n_671), .B(n_693), .Y(n_670) );
NAND3xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_683), .C(n_688), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_674), .B(n_679), .Y(n_673) );
OAI21xp5_ASAP7_75t_SL g674 ( .A1(n_675), .A2(n_676), .B(n_677), .Y(n_674) );
OAI221xp5_ASAP7_75t_L g757 ( .A1(n_675), .A2(n_758), .B1(n_759), .B2(n_760), .C(n_761), .Y(n_757) );
INVx2_ASAP7_75t_SL g893 ( .A(n_678), .Y(n_893) );
NAND3xp33_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .C(n_682), .Y(n_679) );
AND2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_686), .Y(n_683) );
AND2x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_691), .Y(n_688) );
INVx1_ASAP7_75t_SL g796 ( .A(n_690), .Y(n_796) );
OA22x2_ASAP7_75t_L g750 ( .A1(n_693), .A2(n_751), .B1(n_776), .B2(n_777), .Y(n_750) );
INVx1_ASAP7_75t_L g777 ( .A(n_693), .Y(n_777) );
NAND4xp75_ASAP7_75t_L g694 ( .A(n_695), .B(n_700), .C(n_704), .D(n_708), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_699), .Y(n_695) );
INVx1_ASAP7_75t_L g735 ( .A(n_697), .Y(n_735) );
AND2x2_ASAP7_75t_SL g700 ( .A(n_701), .B(n_703), .Y(n_700) );
AND2x2_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .Y(n_704) );
INVx1_ASAP7_75t_L g748 ( .A(n_709), .Y(n_748) );
INVx1_ASAP7_75t_L g747 ( .A(n_710), .Y(n_747) );
AND2x2_ASAP7_75t_L g710 ( .A(n_711), .B(n_733), .Y(n_710) );
NOR3xp33_ASAP7_75t_L g711 ( .A(n_712), .B(n_715), .C(n_722), .Y(n_711) );
OAI222xp33_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_717), .B1(n_718), .B2(n_719), .C1(n_720), .C2(n_721), .Y(n_715) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_724), .B1(n_727), .B2(n_728), .Y(n_722) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx3_ASAP7_75t_SL g923 ( .A(n_725), .Y(n_923) );
INVx4_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_726), .Y(n_765) );
BUFx3_ASAP7_75t_L g802 ( .A(n_726), .Y(n_802) );
OAI22xp5_ASAP7_75t_L g763 ( .A1(n_728), .A2(n_764), .B1(n_765), .B2(n_766), .Y(n_763) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g899 ( .A(n_729), .Y(n_899) );
CKINVDCx16_ASAP7_75t_R g729 ( .A(n_730), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g800 ( .A1(n_730), .A2(n_801), .B1(n_802), .B2(n_803), .Y(n_800) );
BUFx2_ASAP7_75t_L g925 ( .A(n_730), .Y(n_925) );
OAI22xp5_ASAP7_75t_L g950 ( .A1(n_730), .A2(n_802), .B1(n_951), .B2(n_952), .Y(n_950) );
OR2x6_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_734), .B(n_739), .Y(n_733) );
NAND2xp5_ASAP7_75t_SL g739 ( .A(n_740), .B(n_742), .Y(n_739) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx3_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g776 ( .A(n_751), .Y(n_776) );
INVx2_ASAP7_75t_L g775 ( .A(n_752), .Y(n_775) );
AND2x2_ASAP7_75t_L g752 ( .A(n_753), .B(n_767), .Y(n_752) );
NOR3xp33_ASAP7_75t_L g753 ( .A(n_754), .B(n_757), .C(n_763), .Y(n_753) );
OAI221xp5_ASAP7_75t_SL g917 ( .A1(n_759), .A2(n_824), .B1(n_918), .B2(n_919), .C(n_920), .Y(n_917) );
NOR2xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_771), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_769), .B(n_770), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_772), .B(n_773), .Y(n_771) );
INVx1_ASAP7_75t_L g986 ( .A(n_779), .Y(n_986) );
AOI22xp5_ASAP7_75t_SL g779 ( .A1(n_780), .A2(n_878), .B1(n_879), .B2(n_984), .Y(n_779) );
INVx1_ASAP7_75t_L g984 ( .A(n_780), .Y(n_984) );
OAI22xp5_ASAP7_75t_SL g780 ( .A1(n_781), .A2(n_782), .B1(n_850), .B2(n_851), .Y(n_780) );
INVx2_ASAP7_75t_SL g781 ( .A(n_782), .Y(n_781) );
OA22x2_ASAP7_75t_L g782 ( .A1(n_783), .A2(n_807), .B1(n_808), .B2(n_849), .Y(n_782) );
INVx1_ASAP7_75t_L g849 ( .A(n_783), .Y(n_849) );
INVx1_ASAP7_75t_L g806 ( .A(n_784), .Y(n_806) );
AND4x1_ASAP7_75t_L g784 ( .A(n_785), .B(n_791), .C(n_797), .D(n_804), .Y(n_784) );
BUFx2_ASAP7_75t_R g788 ( .A(n_789), .Y(n_788) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_794), .B1(n_795), .B2(n_796), .Y(n_792) );
BUFx2_ASAP7_75t_L g862 ( .A(n_798), .Y(n_862) );
OAI22xp5_ASAP7_75t_L g896 ( .A1(n_802), .A2(n_897), .B1(n_898), .B2(n_899), .Y(n_896) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
AOI22xp5_ASAP7_75t_L g808 ( .A1(n_809), .A2(n_828), .B1(n_847), .B2(n_848), .Y(n_808) );
INVx2_ASAP7_75t_SL g847 ( .A(n_809), .Y(n_847) );
XOR2x2_ASAP7_75t_L g809 ( .A(n_810), .B(n_827), .Y(n_809) );
NOR4xp75_ASAP7_75t_L g810 ( .A(n_811), .B(n_816), .C(n_820), .D(n_823), .Y(n_810) );
NAND2xp5_ASAP7_75t_SL g811 ( .A(n_812), .B(n_813), .Y(n_811) );
BUFx6f_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
NAND2x1_ASAP7_75t_L g816 ( .A(n_817), .B(n_819), .Y(n_816) );
NAND2xp5_ASAP7_75t_SL g820 ( .A(n_821), .B(n_822), .Y(n_820) );
OAI21xp5_ASAP7_75t_SL g823 ( .A1(n_824), .A2(n_825), .B(n_826), .Y(n_823) );
INVx1_ASAP7_75t_L g848 ( .A(n_828), .Y(n_848) );
XOR2x2_ASAP7_75t_L g828 ( .A(n_829), .B(n_846), .Y(n_828) );
NAND2x1_ASAP7_75t_L g829 ( .A(n_830), .B(n_839), .Y(n_829) );
NOR2xp33_ASAP7_75t_L g830 ( .A(n_831), .B(n_835), .Y(n_830) );
OAI21xp5_ASAP7_75t_SL g831 ( .A1(n_832), .A2(n_833), .B(n_834), .Y(n_831) );
NAND3xp33_ASAP7_75t_L g835 ( .A(n_836), .B(n_837), .C(n_838), .Y(n_835) );
NOR2x1_ASAP7_75t_L g839 ( .A(n_840), .B(n_843), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_841), .B(n_842), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_844), .B(n_845), .Y(n_843) );
INVx1_ASAP7_75t_SL g850 ( .A(n_851), .Y(n_850) );
INVx2_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
XOR2x2_ASAP7_75t_L g852 ( .A(n_853), .B(n_877), .Y(n_852) );
NAND4xp75_ASAP7_75t_L g853 ( .A(n_854), .B(n_858), .C(n_864), .D(n_876), .Y(n_853) );
AND2x2_ASAP7_75t_L g854 ( .A(n_855), .B(n_857), .Y(n_854) );
OA211x2_ASAP7_75t_L g858 ( .A1(n_859), .A2(n_860), .B(n_861), .C(n_863), .Y(n_858) );
OA211x2_ASAP7_75t_L g1009 ( .A1(n_860), .A2(n_1010), .B(n_1011), .C(n_1012), .Y(n_1009) );
NOR2xp33_ASAP7_75t_L g864 ( .A(n_865), .B(n_869), .Y(n_864) );
OAI22xp5_ASAP7_75t_L g869 ( .A1(n_870), .A2(n_871), .B1(n_873), .B2(n_874), .Y(n_869) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx1_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
AOI22xp5_ASAP7_75t_L g880 ( .A1(n_881), .A2(n_882), .B1(n_908), .B2(n_983), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
BUFx2_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx1_ASAP7_75t_SL g884 ( .A(n_885), .Y(n_884) );
AND2x2_ASAP7_75t_L g885 ( .A(n_886), .B(n_900), .Y(n_885) );
NOR3xp33_ASAP7_75t_L g886 ( .A(n_887), .B(n_891), .C(n_896), .Y(n_886) );
NOR2xp33_ASAP7_75t_L g900 ( .A(n_901), .B(n_904), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_902), .B(n_903), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_905), .B(n_906), .Y(n_904) );
INVx1_ASAP7_75t_L g983 ( .A(n_908), .Y(n_983) );
AOI22xp5_ASAP7_75t_L g908 ( .A1(n_909), .A2(n_910), .B1(n_936), .B2(n_937), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
INVx2_ASAP7_75t_L g935 ( .A(n_911), .Y(n_935) );
AND2x2_ASAP7_75t_SL g911 ( .A(n_912), .B(n_926), .Y(n_911) );
NOR3xp33_ASAP7_75t_L g912 ( .A(n_913), .B(n_917), .C(n_921), .Y(n_912) );
OAI22xp5_ASAP7_75t_L g1030 ( .A1(n_916), .A2(n_944), .B1(n_1031), .B2(n_1032), .Y(n_1030) );
OAI22xp5_ASAP7_75t_L g921 ( .A1(n_922), .A2(n_923), .B1(n_924), .B2(n_925), .Y(n_921) );
NOR2xp33_ASAP7_75t_L g926 ( .A(n_927), .B(n_930), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_928), .B(n_929), .Y(n_927) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_931), .B(n_933), .Y(n_930) );
INVx1_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
AO22x1_ASAP7_75t_L g937 ( .A1(n_938), .A2(n_939), .B1(n_963), .B2(n_982), .Y(n_937) );
INVx2_ASAP7_75t_SL g938 ( .A(n_939), .Y(n_938) );
XOR2x2_ASAP7_75t_L g939 ( .A(n_940), .B(n_962), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_941), .B(n_953), .Y(n_940) );
NOR3xp33_ASAP7_75t_L g941 ( .A(n_942), .B(n_946), .C(n_950), .Y(n_941) );
OAI21xp33_ASAP7_75t_L g946 ( .A1(n_947), .A2(n_948), .B(n_949), .Y(n_946) );
OAI21xp5_ASAP7_75t_SL g966 ( .A1(n_948), .A2(n_967), .B(n_968), .Y(n_966) );
NOR2xp33_ASAP7_75t_L g953 ( .A(n_954), .B(n_958), .Y(n_953) );
NAND2xp5_ASAP7_75t_L g954 ( .A(n_955), .B(n_957), .Y(n_954) );
NAND2xp5_ASAP7_75t_L g958 ( .A(n_959), .B(n_960), .Y(n_958) );
INVx3_ASAP7_75t_SL g982 ( .A(n_963), .Y(n_982) );
XOR2x2_ASAP7_75t_L g963 ( .A(n_964), .B(n_981), .Y(n_963) );
NAND2xp5_ASAP7_75t_SL g964 ( .A(n_965), .B(n_973), .Y(n_964) );
NOR2xp33_ASAP7_75t_L g965 ( .A(n_966), .B(n_969), .Y(n_965) );
NAND3xp33_ASAP7_75t_L g969 ( .A(n_970), .B(n_971), .C(n_972), .Y(n_969) );
NOR2xp33_ASAP7_75t_L g973 ( .A(n_974), .B(n_977), .Y(n_973) );
NAND2xp5_ASAP7_75t_L g974 ( .A(n_975), .B(n_976), .Y(n_974) );
NAND2xp5_ASAP7_75t_L g977 ( .A(n_978), .B(n_979), .Y(n_977) );
INVx1_ASAP7_75t_SL g987 ( .A(n_988), .Y(n_987) );
NOR2x1_ASAP7_75t_L g988 ( .A(n_989), .B(n_993), .Y(n_988) );
OR2x2_ASAP7_75t_SL g1049 ( .A(n_989), .B(n_994), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g989 ( .A(n_990), .B(n_992), .Y(n_989) );
CKINVDCx20_ASAP7_75t_R g1018 ( .A(n_990), .Y(n_1018) );
INVx1_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
NAND2xp5_ASAP7_75t_L g1023 ( .A(n_991), .B(n_1020), .Y(n_1023) );
CKINVDCx16_ASAP7_75t_R g1020 ( .A(n_992), .Y(n_1020) );
CKINVDCx20_ASAP7_75t_R g993 ( .A(n_994), .Y(n_993) );
NAND2xp5_ASAP7_75t_L g994 ( .A(n_995), .B(n_996), .Y(n_994) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_998), .B(n_999), .Y(n_997) );
OAI322xp33_ASAP7_75t_L g1000 ( .A1(n_1001), .A2(n_1017), .A3(n_1019), .B1(n_1021), .B2(n_1024), .C1(n_1025), .C2(n_1047), .Y(n_1000) );
CKINVDCx20_ASAP7_75t_R g1002 ( .A(n_1003), .Y(n_1002) );
HB1xp67_ASAP7_75t_L g1003 ( .A(n_1004), .Y(n_1003) );
NAND4xp75_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1009), .C(n_1013), .D(n_1016), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_1006), .B(n_1007), .Y(n_1005) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1015), .Y(n_1013) );
HB1xp67_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
INVx1_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
CKINVDCx16_ASAP7_75t_R g1021 ( .A(n_1022), .Y(n_1021) );
INVx1_ASAP7_75t_L g1025 ( .A(n_1026), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
INVx2_ASAP7_75t_L g1046 ( .A(n_1028), .Y(n_1046) );
NAND2xp5_ASAP7_75t_L g1028 ( .A(n_1029), .B(n_1039), .Y(n_1028) );
NOR3xp33_ASAP7_75t_L g1029 ( .A(n_1030), .B(n_1033), .C(n_1036), .Y(n_1029) );
NOR2xp33_ASAP7_75t_L g1039 ( .A(n_1040), .B(n_1043), .Y(n_1039) );
NAND2xp5_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1042), .Y(n_1040) );
NAND2xp5_ASAP7_75t_L g1043 ( .A(n_1044), .B(n_1045), .Y(n_1043) );
CKINVDCx20_ASAP7_75t_R g1047 ( .A(n_1048), .Y(n_1047) );
CKINVDCx20_ASAP7_75t_R g1048 ( .A(n_1049), .Y(n_1048) );
endmodule