module fake_jpeg_26326_n_288 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_288);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_288;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_13),
.B(n_6),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_31),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_13),
.B(n_6),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_35),
.Y(n_40)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_12),
.Y(n_33)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_21),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_29),
.B(n_19),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_46),
.B(n_21),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_47),
.B(n_51),
.Y(n_66)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_27),
.B1(n_15),
.B2(n_28),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_62),
.B(n_33),
.Y(n_74)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_53),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_44),
.B(n_27),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_14),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_56),
.Y(n_81)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_14),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_60),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_22),
.B1(n_16),
.B2(n_19),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_61),
.A2(n_64),
.B1(n_38),
.B2(n_39),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_35),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_63),
.B(n_65),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_38),
.A2(n_22),
.B1(n_16),
.B2(n_19),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_72),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_70),
.A2(n_65),
.B1(n_45),
.B2(n_28),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_55),
.Y(n_71)
);

BUFx2_ASAP7_75t_SL g103 ( 
.A(n_71),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_74),
.A2(n_82),
.B(n_62),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_50),
.A2(n_39),
.B1(n_43),
.B2(n_45),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_75),
.A2(n_57),
.B1(n_43),
.B2(n_45),
.Y(n_89)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_77),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_63),
.B(n_35),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_84),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_49),
.Y(n_82)
);

NOR2x1_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_32),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_34),
.C(n_30),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_34),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_84),
.A2(n_55),
.B1(n_43),
.B2(n_57),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_86),
.A2(n_98),
.B1(n_102),
.B2(n_104),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_88),
.A2(n_82),
.B(n_79),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_90),
.B1(n_96),
.B2(n_104),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_68),
.A2(n_48),
.B1(n_59),
.B2(n_42),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_60),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_93),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_56),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_53),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_99),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_47),
.B1(n_58),
.B2(n_35),
.Y(n_96)
);

INVxp67_ASAP7_75t_SL g97 ( 
.A(n_71),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_102),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_82),
.A2(n_58),
.B1(n_34),
.B2(n_30),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_80),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_100),
.Y(n_109)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_41),
.B1(n_30),
.B2(n_26),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_85),
.C(n_74),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_106),
.C(n_120),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_85),
.C(n_81),
.Y(n_106)
);

NAND2x1_ASAP7_75t_SL g107 ( 
.A(n_98),
.B(n_84),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_107),
.A2(n_125),
.B(n_94),
.Y(n_131)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_108),
.B(n_115),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_113),
.A2(n_73),
.B(n_97),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_70),
.B1(n_75),
.B2(n_82),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_100),
.B1(n_77),
.B2(n_101),
.Y(n_134)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_118),
.Y(n_146)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_78),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_83),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_78),
.C(n_66),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_93),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_121),
.Y(n_130)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_73),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_95),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_123),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_87),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_127),
.Y(n_148)
);

NOR3xp33_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_83),
.C(n_66),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_122),
.A2(n_89),
.B1(n_87),
.B2(n_86),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_128),
.A2(n_137),
.B1(n_151),
.B2(n_108),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_114),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_131),
.A2(n_138),
.B(n_111),
.Y(n_158)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_135),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_113),
.A2(n_101),
.B(n_100),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_134),
.A2(n_152),
.B1(n_20),
.B2(n_26),
.Y(n_178)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_115),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_112),
.A2(n_100),
.B1(n_101),
.B2(n_77),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_106),
.A2(n_105),
.B(n_107),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_141),
.Y(n_170)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_121),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_143),
.Y(n_167)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_144),
.B(n_147),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_123),
.Y(n_147)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_110),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_154),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_125),
.A2(n_67),
.B1(n_69),
.B2(n_80),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_111),
.A2(n_67),
.B1(n_69),
.B2(n_71),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_52),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_153),
.B(n_67),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_107),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_119),
.C(n_120),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_176),
.C(n_179),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_156),
.B(n_174),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_158),
.B(n_160),
.Y(n_192)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_161),
.B(n_162),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_148),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_52),
.Y(n_163)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_163),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_164),
.A2(n_166),
.B1(n_171),
.B2(n_172),
.Y(n_185)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_165),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_128),
.A2(n_109),
.B1(n_118),
.B2(n_116),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_151),
.A2(n_69),
.B1(n_71),
.B2(n_73),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_154),
.A2(n_141),
.B1(n_144),
.B2(n_131),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_180),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_32),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_26),
.Y(n_175)
);

MAJx2_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_137),
.C(n_18),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_129),
.B(n_136),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_178),
.A2(n_164),
.B1(n_175),
.B2(n_176),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_25),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_168),
.A2(n_133),
.B(n_145),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_184),
.A2(n_9),
.B(n_11),
.Y(n_210)
);

INVx13_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_187),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_132),
.C(n_140),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_24),
.C(n_23),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_139),
.Y(n_189)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_189),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_168),
.A2(n_147),
.B1(n_130),
.B2(n_143),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_191),
.A2(n_202),
.B1(n_203),
.B2(n_156),
.Y(n_205)
);

OAI221xp5_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_139),
.B1(n_172),
.B2(n_157),
.C(n_155),
.Y(n_193)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

NOR3xp33_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_145),
.C(n_134),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_196),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_179),
.B(n_135),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_152),
.Y(n_198)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_166),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_201),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_18),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_20),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_171),
.Y(n_202)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_192),
.B(n_25),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_208),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_199),
.A2(n_20),
.B1(n_17),
.B2(n_24),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_209),
.A2(n_190),
.B1(n_186),
.B2(n_187),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_211),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_25),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_192),
.B(n_18),
.Y(n_213)
);

MAJx2_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_191),
.C(n_181),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_219),
.C(n_18),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_20),
.C(n_23),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_200),
.C(n_184),
.Y(n_225)
);

FAx1_ASAP7_75t_SL g217 ( 
.A(n_198),
.B(n_183),
.CI(n_182),
.CON(n_217),
.SN(n_217)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_221),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_185),
.A2(n_24),
.B1(n_23),
.B2(n_17),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_218),
.A2(n_201),
.B1(n_24),
.B2(n_23),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_183),
.B(n_18),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_194),
.A2(n_7),
.B(n_10),
.Y(n_221)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_223),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_227),
.C(n_229),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_226),
.A2(n_234),
.B1(n_4),
.B2(n_8),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_197),
.C(n_203),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_185),
.C(n_181),
.Y(n_229)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_230),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_215),
.A2(n_17),
.B1(n_18),
.B2(n_6),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_232),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_17),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_233),
.A2(n_237),
.B(n_0),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_204),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_0),
.C(n_1),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_4),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_224),
.Y(n_238)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_238),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_228),
.A2(n_222),
.B1(n_220),
.B2(n_218),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_239),
.A2(n_240),
.B1(n_244),
.B2(n_246),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_229),
.A2(n_217),
.B1(n_209),
.B2(n_207),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_234),
.A2(n_217),
.B(n_208),
.Y(n_243)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_243),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_225),
.A2(n_213),
.B1(n_211),
.B2(n_219),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_227),
.A2(n_4),
.B1(n_8),
.B2(n_7),
.Y(n_246)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_248),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_5),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_226),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_235),
.Y(n_251)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_251),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_259),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_244),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_258),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_235),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_247),
.B(n_231),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_0),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_231),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_4),
.Y(n_268)
);

INVxp33_ASAP7_75t_L g262 ( 
.A(n_251),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_270),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_242),
.C(n_238),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_266),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_245),
.C(n_250),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_248),
.C(n_5),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_269),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_268),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_5),
.C(n_8),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_261),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_273),
.B(n_10),
.Y(n_280)
);

AOI21x1_ASAP7_75t_L g276 ( 
.A1(n_263),
.A2(n_3),
.B(n_7),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_276),
.A2(n_3),
.B(n_7),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_275),
.A2(n_271),
.B(n_268),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_278),
.A2(n_272),
.B(n_277),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_279),
.A2(n_280),
.B(n_274),
.Y(n_281)
);

AOI21x1_ASAP7_75t_L g283 ( 
.A1(n_281),
.A2(n_282),
.B(n_10),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_10),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_284),
.A2(n_0),
.B(n_1),
.Y(n_285)
);

AOI321xp33_ASAP7_75t_L g286 ( 
.A1(n_285),
.A2(n_1),
.A3(n_2),
.B1(n_167),
.B2(n_274),
.C(n_215),
.Y(n_286)
);

BUFx24_ASAP7_75t_SL g287 ( 
.A(n_286),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_1),
.Y(n_288)
);


endmodule