module fake_jpeg_31560_n_127 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_127);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_127;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_37),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_1),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_18),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_27),
.Y(n_53)
);

INVx11_ASAP7_75t_SL g54 ( 
.A(n_19),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_0),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_57),
.Y(n_72)
);

BUFx4f_ASAP7_75t_SL g56 ( 
.A(n_44),
.Y(n_56)
);

INVx5_ASAP7_75t_SL g64 ( 
.A(n_56),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_0),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_1),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_61),
.Y(n_65)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_62),
.A2(n_56),
.B1(n_53),
.B2(n_52),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_57),
.A2(n_51),
.B1(n_49),
.B2(n_54),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_63),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_46),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_69),
.B(n_4),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_47),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_45),
.B1(n_43),
.B2(n_42),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_41),
.B1(n_48),
.B2(n_22),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_55),
.B(n_2),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_3),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_76),
.B(n_79),
.Y(n_98)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_11),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_5),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_5),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_88),
.Y(n_91)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

BUFx2_ASAP7_75t_SL g92 ( 
.A(n_84),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_67),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_6),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_6),
.Y(n_88)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_96),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_86),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_95),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_7),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_81),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_99),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_81),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_100),
.A2(n_16),
.B1(n_20),
.B2(n_21),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_91),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_SL g104 ( 
.A1(n_81),
.A2(n_12),
.B(n_14),
.C(n_15),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_104),
.A2(n_31),
.B(n_32),
.Y(n_114)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_108),
.Y(n_118)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_114),
.B1(n_92),
.B2(n_103),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_23),
.C(n_24),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_111),
.A2(n_112),
.B1(n_115),
.B2(n_104),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_101),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_117),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_119),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_120),
.B(n_110),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_110),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_98),
.C(n_118),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

A2O1A1O1Ixp25_ASAP7_75t_L g126 ( 
.A1(n_125),
.A2(n_121),
.B(n_118),
.C(n_113),
.D(n_104),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_126),
.B(n_113),
.Y(n_127)
);


endmodule