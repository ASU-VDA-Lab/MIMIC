module fake_jpeg_22970_n_258 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_258);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_258;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_33),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_34),
.B(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_38),
.Y(n_45)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_42),
.B(n_29),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_25),
.B1(n_28),
.B2(n_27),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_61)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_16),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_52),
.Y(n_57)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_53),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_25),
.B1(n_28),
.B2(n_27),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_36),
.B1(n_35),
.B2(n_40),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_25),
.B1(n_17),
.B2(n_32),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_50),
.A2(n_22),
.B(n_20),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_51),
.B(n_54),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_22),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_55),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_65),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_34),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_69),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_61),
.B(n_71),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_36),
.B1(n_35),
.B2(n_40),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_62),
.A2(n_79),
.B1(n_83),
.B2(n_33),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_31),
.Y(n_63)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

FAx1_ASAP7_75t_SL g64 ( 
.A(n_47),
.B(n_27),
.CI(n_32),
.CON(n_64),
.SN(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_64),
.A2(n_22),
.B(n_20),
.C(n_33),
.Y(n_91)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_75),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_17),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_85),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_55),
.A2(n_18),
.B1(n_21),
.B2(n_30),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_68),
.A2(n_74),
.B1(n_81),
.B2(n_89),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_42),
.B(n_36),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_33),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_33),
.Y(n_100)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_51),
.B(n_23),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_73),
.B(n_82),
.Y(n_116)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_45),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_78),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_41),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_SL g79 ( 
.A1(n_43),
.A2(n_33),
.B(n_16),
.C(n_18),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_23),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_84),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_55),
.A2(n_21),
.B1(n_31),
.B2(n_26),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_50),
.B(n_26),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_55),
.A2(n_33),
.B1(n_29),
.B2(n_24),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_0),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

BUFx4f_ASAP7_75t_SL g94 ( 
.A(n_86),
.Y(n_94)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_88),
.Y(n_114)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_97),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_91),
.B(n_82),
.Y(n_117)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_111),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_102),
.A2(n_107),
.B1(n_109),
.B2(n_79),
.Y(n_131)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_106),
.Y(n_135)
);

MAJx2_ASAP7_75t_L g104 ( 
.A(n_57),
.B(n_33),
.C(n_2),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_84),
.C(n_58),
.Y(n_143)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_66),
.A2(n_33),
.B1(n_1),
.B2(n_4),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_87),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_109)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

INVxp33_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_57),
.B(n_1),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_57),
.B(n_4),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_85),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_117),
.A2(n_118),
.B(n_5),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_111),
.A2(n_92),
.B(n_115),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_123),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_94),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_122),
.B(n_124),
.Y(n_154)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_70),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_125),
.A2(n_127),
.B(n_129),
.Y(n_146)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_134),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_91),
.A2(n_89),
.B(n_77),
.Y(n_127)
);

AOI322xp5_ASAP7_75t_L g128 ( 
.A1(n_99),
.A2(n_67),
.A3(n_64),
.B1(n_62),
.B2(n_72),
.C1(n_69),
.C2(n_78),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_116),
.C(n_104),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_94),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_131),
.A2(n_132),
.B1(n_139),
.B2(n_110),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_103),
.A2(n_79),
.B1(n_71),
.B2(n_64),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_94),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_133),
.A2(n_140),
.B(n_142),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_92),
.B(n_72),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_67),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_137),
.Y(n_167)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_96),
.A2(n_74),
.B1(n_88),
.B2(n_60),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_99),
.B(n_85),
.Y(n_141)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_141),
.Y(n_149)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_124),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_162),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_131),
.A2(n_105),
.B1(n_96),
.B2(n_102),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_145),
.A2(n_148),
.B1(n_153),
.B2(n_156),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_105),
.C(n_101),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_161),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_127),
.A2(n_101),
.B1(n_116),
.B2(n_65),
.Y(n_148)
);

INVxp33_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_138),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_135),
.A2(n_117),
.B(n_140),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_152),
.A2(n_160),
.B(n_166),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_130),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_155),
.B(n_158),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_142),
.A2(n_65),
.B1(n_106),
.B2(n_83),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_139),
.A2(n_83),
.B1(n_97),
.B2(n_113),
.Y(n_157)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_157),
.Y(n_182)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_141),
.A2(n_83),
.B(n_73),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_143),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_98),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_165),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_118),
.B(n_98),
.C(n_112),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_132),
.A2(n_90),
.B1(n_112),
.B2(n_8),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_168),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_134),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_169)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_133),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_176),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_163),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_125),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_178),
.Y(n_205)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_163),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_151),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_180),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_125),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_181),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_152),
.A2(n_128),
.B(n_123),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_184),
.A2(n_188),
.B(n_149),
.Y(n_201)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

BUFx24_ASAP7_75t_SL g204 ( 
.A(n_185),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_148),
.B(n_125),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_154),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_189),
.A2(n_167),
.B1(n_160),
.B2(n_168),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g190 ( 
.A(n_146),
.Y(n_190)
);

AOI21xp33_ASAP7_75t_L g196 ( 
.A1(n_190),
.A2(n_167),
.B(n_158),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_178),
.A2(n_145),
.B1(n_157),
.B2(n_156),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_193),
.A2(n_196),
.B1(n_174),
.B2(n_182),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_161),
.C(n_146),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_199),
.C(n_203),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_207),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_164),
.C(n_165),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_162),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_201),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_144),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_206),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_149),
.C(n_147),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_166),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_129),
.C(n_122),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_193),
.A2(n_174),
.B1(n_186),
.B2(n_190),
.Y(n_208)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_208),
.Y(n_232)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_209),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_192),
.A2(n_182),
.B1(n_187),
.B2(n_186),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_214),
.A2(n_219),
.B1(n_207),
.B2(n_188),
.Y(n_229)
);

NOR3xp33_ASAP7_75t_SL g215 ( 
.A(n_201),
.B(n_184),
.C(n_183),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_215),
.B(n_217),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_194),
.B(n_137),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_216),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_191),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_120),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_220),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_198),
.A2(n_181),
.B1(n_187),
.B2(n_188),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_175),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_183),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_195),
.Y(n_224)
);

XNOR2x1_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_221),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_222),
.A2(n_211),
.B1(n_169),
.B2(n_119),
.Y(n_239)
);

MAJx2_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_206),
.C(n_202),
.Y(n_223)
);

AOI321xp33_ASAP7_75t_L g240 ( 
.A1(n_223),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_211),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_229),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_203),
.C(n_200),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_231),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_119),
.C(n_126),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_224),
.Y(n_242)
);

INVxp33_ASAP7_75t_L g234 ( 
.A(n_225),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_234),
.A2(n_236),
.B(n_239),
.Y(n_243)
);

OAI321xp33_ASAP7_75t_L g236 ( 
.A1(n_226),
.A2(n_215),
.A3(n_209),
.B1(n_214),
.B2(n_219),
.C(n_228),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_212),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_238),
.B(n_231),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_240),
.A2(n_232),
.B(n_222),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_234),
.B(n_227),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_241),
.B(n_242),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_245),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_237),
.B(n_230),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_246),
.B(n_6),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_243),
.A2(n_235),
.B1(n_223),
.B2(n_233),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_248),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_251)
);

A2O1A1Ixp33_ASAP7_75t_L g252 ( 
.A1(n_249),
.A2(n_11),
.B(n_12),
.C(n_14),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_251),
.A2(n_253),
.B(n_250),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_252),
.A2(n_248),
.B1(n_12),
.B2(n_14),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_247),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_254),
.B(n_255),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_11),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_257),
.B(n_14),
.Y(n_258)
);


endmodule