module fake_ibex_1907_n_21 (n_3, n_1, n_5, n_4, n_2, n_0, n_6, n_21);

input n_3;
input n_1;
input n_5;
input n_4;
input n_2;
input n_0;
input n_6;

output n_21;



endmodule