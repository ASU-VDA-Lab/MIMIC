module real_jpeg_11995_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_195;
wire n_61;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_202;
wire n_128;
wire n_179;
wire n_167;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_4),
.A2(n_43),
.B1(n_45),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_4),
.A2(n_29),
.B1(n_36),
.B2(n_53),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_4),
.A2(n_53),
.B1(n_59),
.B2(n_63),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_5),
.A2(n_65),
.B1(n_66),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_5),
.A2(n_59),
.B1(n_63),
.B2(n_71),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_5),
.A2(n_43),
.B1(n_45),
.B2(n_71),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_5),
.A2(n_29),
.B1(n_36),
.B2(n_71),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_6),
.A2(n_65),
.B1(n_66),
.B2(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_6),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_6),
.A2(n_59),
.B1(n_63),
.B2(n_110),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_6),
.A2(n_43),
.B1(n_45),
.B2(n_110),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_6),
.A2(n_29),
.B1(n_36),
.B2(n_110),
.Y(n_214)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_8),
.A2(n_65),
.B1(n_66),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_8),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_8),
.A2(n_59),
.B1(n_63),
.B2(n_69),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_8),
.A2(n_43),
.B1(n_45),
.B2(n_69),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_8),
.A2(n_29),
.B1(n_36),
.B2(n_69),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_9),
.A2(n_29),
.B1(n_36),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_9),
.A2(n_38),
.B1(n_43),
.B2(n_45),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_10),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_10),
.A2(n_42),
.B1(n_59),
.B2(n_63),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_10),
.A2(n_29),
.B1(n_36),
.B2(n_42),
.Y(n_158)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_11),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_12),
.A2(n_29),
.B1(n_36),
.B2(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_12),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_13),
.A2(n_59),
.B1(n_63),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_13),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_13),
.A2(n_65),
.B1(n_66),
.B2(n_80),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_13),
.A2(n_43),
.B1(n_45),
.B2(n_80),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_13),
.A2(n_29),
.B1(n_36),
.B2(n_80),
.Y(n_181)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_15),
.Y(n_101)
);

AOI21xp33_ASAP7_75t_L g140 ( 
.A1(n_15),
.A2(n_65),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_15),
.B(n_113),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_L g192 ( 
.A1(n_15),
.A2(n_43),
.B1(n_45),
.B2(n_101),
.Y(n_192)
);

O2A1O1Ixp33_ASAP7_75t_L g194 ( 
.A1(n_15),
.A2(n_45),
.B(n_49),
.C(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_15),
.B(n_106),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_15),
.B(n_32),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_15),
.B(n_87),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_15),
.A2(n_63),
.B(n_74),
.C(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_16),
.A2(n_29),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_16),
.A2(n_35),
.B1(n_43),
.B2(n_45),
.Y(n_86)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_134),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_132),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_114),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_21),
.B(n_114),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_82),
.C(n_93),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_22),
.A2(n_23),
.B1(n_82),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_54),
.B2(n_55),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_24),
.B(n_56),
.C(n_72),
.Y(n_115)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_39),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_26),
.B(n_39),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_31),
.B1(n_33),
.B2(n_37),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_27),
.A2(n_31),
.B1(n_206),
.B2(n_208),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_28),
.A2(n_32),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_28),
.A2(n_32),
.B1(n_34),
.B2(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_28),
.A2(n_32),
.B(n_90),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_28),
.A2(n_32),
.B1(n_97),
.B2(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_28),
.A2(n_32),
.B1(n_158),
.B2(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_28),
.A2(n_32),
.B1(n_181),
.B2(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_28),
.A2(n_32),
.B1(n_101),
.B2(n_214),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_28),
.A2(n_32),
.B1(n_207),
.B2(n_214),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_29),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_29),
.A2(n_36),
.B1(n_49),
.B2(n_50),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_29),
.B(n_216),
.Y(n_215)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

OAI21xp33_ASAP7_75t_L g195 ( 
.A1(n_36),
.A2(n_50),
.B(n_101),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_46),
.B1(n_51),
.B2(n_52),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_41),
.A2(n_47),
.B1(n_87),
.B2(n_146),
.Y(n_145)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_45),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_43),
.A2(n_45),
.B1(n_76),
.B2(n_77),
.Y(n_78)
);

OAI32xp33_ASAP7_75t_L g177 ( 
.A1(n_43),
.A2(n_63),
.A3(n_76),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_45),
.B(n_77),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_46),
.A2(n_51),
.B1(n_173),
.B2(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_47),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_47),
.A2(n_86),
.B1(n_87),
.B2(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_47),
.A2(n_87),
.B1(n_146),
.B2(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_47),
.A2(n_87),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_47),
.A2(n_87),
.B1(n_193),
.B2(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_72),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_68),
.B2(n_70),
.Y(n_56)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_57),
.A2(n_58),
.B1(n_70),
.B2(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_57),
.A2(n_58),
.B1(n_109),
.B2(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_64),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_58),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_59),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_59),
.A2(n_63),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

OAI32xp33_ASAP7_75t_L g98 ( 
.A1(n_59),
.A2(n_62),
.A3(n_65),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_59),
.B(n_101),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_61),
.A2(n_62),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_63),
.Y(n_99)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_66),
.B(n_101),
.Y(n_100)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_78),
.B1(n_79),
.B2(n_81),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_73),
.A2(n_78),
.B1(n_81),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_73),
.A2(n_78),
.B1(n_104),
.B2(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_74),
.A2(n_103),
.B1(n_105),
.B2(n_106),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_74),
.A2(n_106),
.B1(n_153),
.B2(n_155),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_78),
.A2(n_154),
.B(n_228),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_82),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_88),
.B2(n_92),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_92),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_93),
.B(n_246),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_102),
.C(n_107),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_94),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_98),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_95),
.A2(n_96),
.B1(n_98),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_98),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_102),
.B(n_107),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_123),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_120),
.B2(n_122),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_130),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_165),
.B(n_243),
.C(n_248),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_159),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_136),
.B(n_159),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_149),
.C(n_151),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_137),
.A2(n_138),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_142),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_143),
.C(n_148),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_145),
.B1(n_147),
.B2(n_148),
.Y(n_142)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_143),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_145),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_149),
.B(n_151),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_156),
.C(n_157),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_152),
.B(n_170),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_157),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_161),
.B(n_162),
.C(n_163),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_242),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_185),
.B(n_241),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_182),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_168),
.B(n_182),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_171),
.C(n_174),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_169),
.B(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_171),
.A2(n_174),
.B1(n_175),
.B2(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_171),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_180),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_176),
.A2(n_177),
.B1(n_180),
.B2(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_178),
.Y(n_229)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_180),
.Y(n_233)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_183),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_235),
.B(n_240),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_223),
.B(n_234),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_203),
.B(n_222),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_196),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_189),
.B(n_196),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_194),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_190),
.A2(n_191),
.B1(n_194),
.B2(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_201),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_199),
.C(n_201),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_200),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_202),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_211),
.B(n_221),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_209),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_205),
.B(n_209),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_217),
.B(n_220),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_218),
.B(n_219),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_224),
.B(n_225),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_232),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_230),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_230),
.C(n_232),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_236),
.B(n_237),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_245),
.Y(n_248)
);


endmodule