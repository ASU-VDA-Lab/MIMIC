module fake_netlist_1_7666_n_664 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_664);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_664;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_472;
wire n_212;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g80 ( .A(n_10), .Y(n_80) );
CKINVDCx16_ASAP7_75t_R g81 ( .A(n_13), .Y(n_81) );
INVxp33_ASAP7_75t_SL g82 ( .A(n_74), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_11), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_49), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_79), .Y(n_85) );
INVxp33_ASAP7_75t_L g86 ( .A(n_38), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_20), .Y(n_87) );
INVxp67_ASAP7_75t_SL g88 ( .A(n_46), .Y(n_88) );
INVxp67_ASAP7_75t_SL g89 ( .A(n_36), .Y(n_89) );
INVxp33_ASAP7_75t_SL g90 ( .A(n_1), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_64), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_4), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_65), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_2), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_9), .Y(n_95) );
INVxp33_ASAP7_75t_SL g96 ( .A(n_12), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_18), .Y(n_97) );
INVx1_ASAP7_75t_SL g98 ( .A(n_51), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_55), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_17), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_30), .Y(n_101) );
HB1xp67_ASAP7_75t_L g102 ( .A(n_62), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_4), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_15), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_16), .Y(n_105) );
INVxp67_ASAP7_75t_SL g106 ( .A(n_20), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_63), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_14), .Y(n_108) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_47), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_54), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_23), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_67), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_45), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_37), .Y(n_114) );
CKINVDCx14_ASAP7_75t_R g115 ( .A(n_33), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_53), .Y(n_116) );
CKINVDCx14_ASAP7_75t_R g117 ( .A(n_77), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_11), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_12), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_29), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_8), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_58), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_19), .Y(n_123) );
INVxp33_ASAP7_75t_SL g124 ( .A(n_3), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_18), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_7), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_35), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_24), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_15), .Y(n_129) );
BUFx2_ASAP7_75t_L g130 ( .A(n_103), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_102), .B(n_0), .Y(n_131) );
INVx3_ASAP7_75t_L g132 ( .A(n_80), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_80), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_115), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_83), .Y(n_135) );
INVxp67_ASAP7_75t_L g136 ( .A(n_129), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_83), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_117), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_87), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_87), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_85), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_92), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_81), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_103), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_92), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_94), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_93), .Y(n_147) );
OAI21x1_ASAP7_75t_L g148 ( .A1(n_85), .A2(n_39), .B(n_76), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g149 ( .A(n_123), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_109), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_84), .Y(n_151) );
NOR2xp33_ASAP7_75t_R g152 ( .A(n_93), .B(n_34), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_127), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_94), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_95), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_127), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_109), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_84), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_122), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_109), .Y(n_160) );
BUFx3_ASAP7_75t_L g161 ( .A(n_91), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_128), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_82), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_119), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_109), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_95), .Y(n_166) );
AND2x6_ASAP7_75t_L g167 ( .A(n_91), .B(n_32), .Y(n_167) );
BUFx2_ASAP7_75t_L g168 ( .A(n_97), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g169 ( .A(n_97), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_126), .Y(n_170) );
HB1xp67_ASAP7_75t_L g171 ( .A(n_100), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_109), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_90), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_126), .Y(n_174) );
OR2x2_ASAP7_75t_SL g175 ( .A(n_171), .B(n_100), .Y(n_175) );
INVx4_ASAP7_75t_L g176 ( .A(n_167), .Y(n_176) );
OAI22xp5_ASAP7_75t_SL g177 ( .A1(n_149), .A2(n_124), .B1(n_96), .B2(n_106), .Y(n_177) );
BUFx3_ASAP7_75t_L g178 ( .A(n_167), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_141), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_141), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_168), .B(n_86), .Y(n_181) );
AND2x4_ASAP7_75t_L g182 ( .A(n_168), .B(n_125), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_150), .Y(n_183) );
OAI221xp5_ASAP7_75t_L g184 ( .A1(n_136), .A2(n_125), .B1(n_121), .B2(n_118), .C(n_105), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_134), .B(n_112), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_151), .Y(n_186) );
BUFx2_ASAP7_75t_L g187 ( .A(n_130), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_151), .Y(n_188) );
AND2x4_ASAP7_75t_L g189 ( .A(n_161), .B(n_121), .Y(n_189) );
NAND2x1p5_ASAP7_75t_L g190 ( .A(n_161), .B(n_120), .Y(n_190) );
AND2x6_ASAP7_75t_L g191 ( .A(n_158), .B(n_120), .Y(n_191) );
INVx4_ASAP7_75t_L g192 ( .A(n_167), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_158), .Y(n_193) );
BUFx3_ASAP7_75t_L g194 ( .A(n_167), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_134), .B(n_107), .Y(n_195) );
AND2x4_ASAP7_75t_L g196 ( .A(n_132), .B(n_118), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_147), .B(n_110), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_147), .B(n_113), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_135), .Y(n_199) );
OR2x6_ASAP7_75t_L g200 ( .A(n_148), .B(n_105), .Y(n_200) );
BUFx3_ASAP7_75t_L g201 ( .A(n_167), .Y(n_201) );
INVx4_ASAP7_75t_L g202 ( .A(n_167), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_150), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_137), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_139), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_148), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_140), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_153), .B(n_101), .Y(n_208) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_150), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_142), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_145), .Y(n_211) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_150), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_146), .Y(n_213) );
AO22x2_ASAP7_75t_L g214 ( .A1(n_154), .A2(n_116), .B1(n_114), .B2(n_99), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_155), .B(n_104), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_150), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_170), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_157), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_153), .B(n_111), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_157), .Y(n_220) );
NAND2x1p5_ASAP7_75t_L g221 ( .A(n_174), .B(n_116), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_132), .Y(n_222) );
AND2x2_ASAP7_75t_L g223 ( .A(n_156), .B(n_108), .Y(n_223) );
NOR2xp33_ASAP7_75t_SL g224 ( .A(n_156), .B(n_98), .Y(n_224) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_157), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_132), .B(n_114), .Y(n_226) );
AOI22xp5_ASAP7_75t_L g227 ( .A1(n_144), .A2(n_89), .B1(n_88), .B2(n_99), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_138), .B(n_0), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_138), .B(n_163), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_133), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_157), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_133), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_163), .B(n_40), .Y(n_233) );
INVx1_ASAP7_75t_SL g234 ( .A(n_144), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_164), .Y(n_235) );
OAI221xp5_ASAP7_75t_L g236 ( .A1(n_131), .A2(n_1), .B1(n_2), .B2(n_3), .C(n_5), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_133), .B(n_5), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_157), .Y(n_238) );
OAI22xp33_ASAP7_75t_SL g239 ( .A1(n_173), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_167), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_160), .Y(n_241) );
INVx3_ASAP7_75t_SL g242 ( .A(n_234), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_181), .B(n_173), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_176), .B(n_152), .Y(n_244) );
CKINVDCx20_ASAP7_75t_R g245 ( .A(n_235), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_237), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_206), .Y(n_247) );
NOR2xp33_ASAP7_75t_R g248 ( .A(n_235), .B(n_143), .Y(n_248) );
AND2x4_ASAP7_75t_L g249 ( .A(n_182), .B(n_143), .Y(n_249) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_187), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_181), .B(n_169), .Y(n_251) );
AOI22xp5_ASAP7_75t_L g252 ( .A1(n_182), .A2(n_166), .B1(n_162), .B2(n_159), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_237), .Y(n_253) );
NOR3xp33_ASAP7_75t_SL g254 ( .A(n_177), .B(n_159), .C(n_162), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_206), .Y(n_255) );
CKINVDCx20_ASAP7_75t_R g256 ( .A(n_187), .Y(n_256) );
INVxp67_ASAP7_75t_SL g257 ( .A(n_190), .Y(n_257) );
NOR2xp33_ASAP7_75t_R g258 ( .A(n_224), .B(n_6), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_182), .B(n_9), .Y(n_259) );
BUFx2_ASAP7_75t_L g260 ( .A(n_190), .Y(n_260) );
BUFx2_ASAP7_75t_L g261 ( .A(n_190), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_189), .B(n_172), .Y(n_262) );
NOR3xp33_ASAP7_75t_SL g263 ( .A(n_236), .B(n_10), .C(n_13), .Y(n_263) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_178), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_176), .B(n_165), .Y(n_265) );
BUFx2_ASAP7_75t_L g266 ( .A(n_221), .Y(n_266) );
BUFx2_ASAP7_75t_L g267 ( .A(n_221), .Y(n_267) );
CKINVDCx8_ASAP7_75t_R g268 ( .A(n_191), .Y(n_268) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_221), .Y(n_269) );
INVx1_ASAP7_75t_SL g270 ( .A(n_223), .Y(n_270) );
BUFx10_ASAP7_75t_L g271 ( .A(n_233), .Y(n_271) );
INVx4_ASAP7_75t_L g272 ( .A(n_189), .Y(n_272) );
NOR3xp33_ASAP7_75t_SL g273 ( .A(n_184), .B(n_14), .C(n_16), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_200), .Y(n_274) );
INVxp67_ASAP7_75t_SL g275 ( .A(n_207), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_200), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_200), .Y(n_277) );
BUFx2_ASAP7_75t_L g278 ( .A(n_214), .Y(n_278) );
AND2x4_ASAP7_75t_L g279 ( .A(n_223), .B(n_215), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_200), .Y(n_280) );
OR2x2_ASAP7_75t_L g281 ( .A(n_175), .B(n_17), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_186), .Y(n_282) );
INVx3_ASAP7_75t_L g283 ( .A(n_179), .Y(n_283) );
NOR2xp33_ASAP7_75t_R g284 ( .A(n_178), .B(n_19), .Y(n_284) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_194), .Y(n_285) );
NAND2xp33_ASAP7_75t_R g286 ( .A(n_240), .B(n_21), .Y(n_286) );
BUFx3_ASAP7_75t_L g287 ( .A(n_194), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_189), .B(n_172), .Y(n_288) );
AND2x6_ASAP7_75t_SL g289 ( .A(n_197), .B(n_21), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_215), .B(n_22), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_186), .Y(n_291) );
BUFx3_ASAP7_75t_L g292 ( .A(n_201), .Y(n_292) );
AND2x4_ASAP7_75t_L g293 ( .A(n_185), .B(n_22), .Y(n_293) );
BUFx2_ASAP7_75t_SL g294 ( .A(n_176), .Y(n_294) );
BUFx4f_ASAP7_75t_L g295 ( .A(n_191), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_207), .B(n_172), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_210), .B(n_199), .Y(n_297) );
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_192), .B(n_165), .Y(n_298) );
NOR2x2_ASAP7_75t_L g299 ( .A(n_175), .B(n_25), .Y(n_299) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_214), .Y(n_300) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_201), .Y(n_301) );
AND2x4_ASAP7_75t_L g302 ( .A(n_196), .B(n_172), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_188), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_188), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_193), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_210), .B(n_172), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_192), .B(n_160), .Y(n_307) );
AND2x4_ASAP7_75t_L g308 ( .A(n_195), .B(n_26), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_193), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_204), .B(n_165), .Y(n_310) );
OR2x2_ASAP7_75t_L g311 ( .A(n_227), .B(n_165), .Y(n_311) );
INVx1_ASAP7_75t_SL g312 ( .A(n_214), .Y(n_312) );
AOI22xp5_ASAP7_75t_L g313 ( .A1(n_259), .A2(n_198), .B1(n_208), .B2(n_219), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_275), .Y(n_314) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_250), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_247), .A2(n_202), .B(n_192), .Y(n_316) );
OR2x2_ASAP7_75t_L g317 ( .A(n_242), .B(n_229), .Y(n_317) );
BUFx2_ASAP7_75t_L g318 ( .A(n_256), .Y(n_318) );
INVx3_ASAP7_75t_SL g319 ( .A(n_242), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_302), .Y(n_320) );
INVx3_ASAP7_75t_SL g321 ( .A(n_256), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_297), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_246), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_253), .Y(n_324) );
INVx2_ASAP7_75t_SL g325 ( .A(n_269), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_279), .B(n_213), .Y(n_326) );
INVxp67_ASAP7_75t_L g327 ( .A(n_250), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_279), .B(n_211), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_266), .B(n_217), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_290), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_267), .B(n_205), .Y(n_331) );
AND2x4_ASAP7_75t_L g332 ( .A(n_269), .B(n_226), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_248), .Y(n_333) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_287), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_247), .Y(n_335) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_287), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_270), .B(n_272), .Y(n_337) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_292), .Y(n_338) );
AOI21xp5_ASAP7_75t_L g339 ( .A1(n_255), .A2(n_202), .B(n_214), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_282), .Y(n_340) );
INVx3_ASAP7_75t_L g341 ( .A(n_302), .Y(n_341) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_292), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_272), .B(n_226), .Y(n_343) );
INVxp67_ASAP7_75t_SL g344 ( .A(n_257), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_255), .Y(n_345) );
AND2x4_ASAP7_75t_L g346 ( .A(n_259), .B(n_226), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_296), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_290), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_248), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_260), .B(n_196), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_311), .Y(n_351) );
AND2x4_ASAP7_75t_L g352 ( .A(n_261), .B(n_196), .Y(n_352) );
OR2x6_ASAP7_75t_L g353 ( .A(n_278), .B(n_202), .Y(n_353) );
AOI21xp5_ASAP7_75t_SL g354 ( .A1(n_274), .A2(n_239), .B(n_180), .Y(n_354) );
CKINVDCx6p67_ASAP7_75t_R g355 ( .A(n_249), .Y(n_355) );
BUFx2_ASAP7_75t_L g356 ( .A(n_300), .Y(n_356) );
AOI21xp5_ASAP7_75t_L g357 ( .A1(n_265), .A2(n_180), .B(n_222), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_300), .A2(n_191), .B1(n_228), .B2(n_232), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_291), .Y(n_359) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_249), .Y(n_360) );
INVx3_ASAP7_75t_L g361 ( .A(n_302), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_243), .B(n_191), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_251), .B(n_230), .Y(n_363) );
INVx2_ASAP7_75t_SL g364 ( .A(n_284), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_312), .A2(n_191), .B1(n_179), .B2(n_230), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_293), .A2(n_191), .B1(n_179), .B2(n_222), .Y(n_366) );
INVx3_ASAP7_75t_L g367 ( .A(n_264), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_315), .A2(n_293), .B1(n_281), .B2(n_308), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_335), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_340), .Y(n_370) );
INVxp67_ASAP7_75t_SL g371 ( .A(n_325), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_356), .A2(n_308), .B1(n_252), .B2(n_258), .Y(n_372) );
AO31x2_ASAP7_75t_L g373 ( .A1(n_339), .A2(n_276), .A3(n_277), .B(n_280), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_322), .B(n_303), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_321), .B(n_304), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_340), .B(n_305), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_359), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_314), .B(n_309), .Y(n_378) );
INVx2_ASAP7_75t_SL g379 ( .A(n_325), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_335), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_345), .Y(n_381) );
AND2x4_ASAP7_75t_L g382 ( .A(n_332), .B(n_274), .Y(n_382) );
INVx4_ASAP7_75t_L g383 ( .A(n_353), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_346), .B(n_263), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_345), .Y(n_385) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_319), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_332), .B(n_273), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_356), .A2(n_258), .B1(n_283), .B2(n_277), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_360), .A2(n_283), .B1(n_280), .B2(n_276), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_347), .Y(n_390) );
NAND2x1p5_ASAP7_75t_L g391 ( .A(n_332), .B(n_264), .Y(n_391) );
AO21x2_ASAP7_75t_L g392 ( .A1(n_354), .A2(n_284), .B(n_306), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_323), .B(n_254), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_355), .B(n_245), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_327), .A2(n_271), .B1(n_245), .B2(n_295), .Y(n_395) );
INVx2_ASAP7_75t_SL g396 ( .A(n_346), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_324), .Y(n_397) );
AOI211xp5_ASAP7_75t_L g398 ( .A1(n_354), .A2(n_299), .B(n_289), .C(n_262), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_346), .A2(n_271), .B1(n_295), .B2(n_294), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_355), .A2(n_244), .B1(n_288), .B2(n_301), .Y(n_400) );
AOI22xp5_ASAP7_75t_L g401 ( .A1(n_363), .A2(n_286), .B1(n_244), .B2(n_299), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_390), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_384), .B(n_321), .Y(n_403) );
OAI22xp33_ASAP7_75t_L g404 ( .A1(n_401), .A2(n_319), .B1(n_318), .B2(n_313), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_390), .B(n_352), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_374), .A2(n_351), .B1(n_366), .B2(n_348), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_374), .A2(n_330), .B1(n_344), .B2(n_353), .Y(n_407) );
AOI222xp33_ASAP7_75t_L g408 ( .A1(n_384), .A2(n_318), .B1(n_326), .B2(n_328), .C1(n_329), .C2(n_331), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_368), .B(n_352), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_390), .B(n_352), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_370), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_370), .B(n_347), .Y(n_412) );
AO31x2_ASAP7_75t_L g413 ( .A1(n_369), .A2(n_357), .A3(n_310), .B(n_362), .Y(n_413) );
INVx3_ASAP7_75t_L g414 ( .A(n_383), .Y(n_414) );
OAI211xp5_ASAP7_75t_L g415 ( .A1(n_398), .A2(n_349), .B(n_333), .C(n_317), .Y(n_415) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_393), .A2(n_349), .B1(n_333), .B2(n_337), .C(n_350), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_380), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g418 ( .A1(n_376), .A2(n_316), .B(n_307), .Y(n_418) );
OA21x2_ASAP7_75t_L g419 ( .A1(n_380), .A2(n_365), .B(n_358), .Y(n_419) );
BUFx2_ASAP7_75t_L g420 ( .A(n_383), .Y(n_420) );
OAI211xp5_ASAP7_75t_L g421 ( .A1(n_398), .A2(n_317), .B(n_343), .C(n_361), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_386), .Y(n_422) );
NOR2x1_ASAP7_75t_SL g423 ( .A(n_383), .B(n_353), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_387), .A2(n_364), .B1(n_341), .B2(n_361), .Y(n_424) );
INVx3_ASAP7_75t_L g425 ( .A(n_383), .Y(n_425) );
BUFx12f_ASAP7_75t_L g426 ( .A(n_375), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_381), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_381), .Y(n_428) );
A2O1A1Ixp33_ASAP7_75t_L g429 ( .A1(n_401), .A2(n_364), .B(n_361), .C(n_320), .Y(n_429) );
AOI21xp5_ASAP7_75t_L g430 ( .A1(n_376), .A2(n_265), .B(n_298), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_412), .B(n_385), .Y(n_431) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_426), .Y(n_432) );
AOI21xp33_ASAP7_75t_L g433 ( .A1(n_408), .A2(n_392), .B(n_372), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_407), .A2(n_388), .B1(n_371), .B2(n_379), .Y(n_434) );
INVx3_ASAP7_75t_L g435 ( .A(n_414), .Y(n_435) );
AND2x4_ASAP7_75t_L g436 ( .A(n_414), .B(n_385), .Y(n_436) );
NAND3xp33_ASAP7_75t_L g437 ( .A(n_408), .B(n_286), .C(n_400), .Y(n_437) );
OAI21xp33_ASAP7_75t_L g438 ( .A1(n_429), .A2(n_393), .B(n_379), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_407), .A2(n_353), .B1(n_375), .B2(n_395), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_411), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_402), .Y(n_441) );
OAI221xp5_ASAP7_75t_L g442 ( .A1(n_416), .A2(n_394), .B1(n_396), .B2(n_397), .C(n_389), .Y(n_442) );
INVx4_ASAP7_75t_L g443 ( .A(n_414), .Y(n_443) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_426), .Y(n_444) );
AOI33xp33_ASAP7_75t_L g445 ( .A1(n_404), .A2(n_397), .A3(n_377), .B1(n_396), .B2(n_399), .B3(n_382), .Y(n_445) );
INVxp67_ASAP7_75t_SL g446 ( .A(n_402), .Y(n_446) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_426), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_417), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_406), .A2(n_392), .B(n_369), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g450 ( .A1(n_409), .A2(n_378), .B1(n_369), .B2(n_377), .Y(n_450) );
INVx4_ASAP7_75t_L g451 ( .A(n_414), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_406), .A2(n_392), .B(n_378), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_417), .Y(n_453) );
INVx1_ASAP7_75t_SL g454 ( .A(n_422), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_412), .B(n_382), .Y(n_455) );
AOI22xp33_ASAP7_75t_SL g456 ( .A1(n_423), .A2(n_392), .B1(n_382), .B2(n_391), .Y(n_456) );
BUFx4f_ASAP7_75t_L g457 ( .A(n_420), .Y(n_457) );
AOI221xp5_ASAP7_75t_L g458 ( .A1(n_403), .A2(n_320), .B1(n_341), .B2(n_382), .C(n_391), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_427), .Y(n_459) );
OR2x6_ASAP7_75t_L g460 ( .A(n_420), .B(n_391), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_427), .Y(n_461) );
AOI221xp5_ASAP7_75t_L g462 ( .A1(n_421), .A2(n_320), .B1(n_341), .B2(n_160), .C(n_165), .Y(n_462) );
OAI221xp5_ASAP7_75t_L g463 ( .A1(n_424), .A2(n_268), .B1(n_298), .B2(n_307), .C(n_367), .Y(n_463) );
CKINVDCx5p33_ASAP7_75t_R g464 ( .A(n_405), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_428), .B(n_373), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_405), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_446), .B(n_428), .Y(n_467) );
AND2x4_ASAP7_75t_L g468 ( .A(n_465), .B(n_425), .Y(n_468) );
BUFx2_ASAP7_75t_L g469 ( .A(n_457), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_465), .B(n_425), .Y(n_470) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_454), .Y(n_471) );
INVx2_ASAP7_75t_SL g472 ( .A(n_457), .Y(n_472) );
INVx1_ASAP7_75t_SL g473 ( .A(n_432), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_441), .B(n_410), .Y(n_474) );
AOI33xp33_ASAP7_75t_L g475 ( .A1(n_440), .A2(n_410), .A3(n_415), .B1(n_238), .B2(n_231), .B3(n_183), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_437), .A2(n_425), .B1(n_419), .B2(n_423), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_441), .Y(n_477) );
NAND2x1_ASAP7_75t_L g478 ( .A(n_443), .B(n_425), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_448), .B(n_373), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_448), .B(n_373), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_453), .B(n_373), .Y(n_481) );
OAI211xp5_ASAP7_75t_L g482 ( .A1(n_433), .A2(n_430), .B(n_418), .C(n_419), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_444), .B(n_419), .Y(n_483) );
INVx3_ASAP7_75t_L g484 ( .A(n_443), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_440), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_461), .Y(n_486) );
NAND3xp33_ASAP7_75t_L g487 ( .A(n_445), .B(n_160), .C(n_419), .Y(n_487) );
OAI221xp5_ASAP7_75t_L g488 ( .A1(n_442), .A2(n_367), .B1(n_160), .B2(n_334), .C(n_342), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_453), .Y(n_489) );
AOI221xp5_ASAP7_75t_L g490 ( .A1(n_439), .A2(n_437), .B1(n_450), .B2(n_438), .C(n_461), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_431), .B(n_373), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_464), .A2(n_336), .B1(n_342), .B2(n_338), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_431), .B(n_373), .Y(n_493) );
INVx1_ASAP7_75t_SL g494 ( .A(n_447), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_459), .B(n_413), .Y(n_495) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_457), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_459), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_435), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_466), .B(n_413), .Y(n_499) );
AND2x4_ASAP7_75t_L g500 ( .A(n_443), .B(n_413), .Y(n_500) );
BUFx2_ASAP7_75t_L g501 ( .A(n_451), .Y(n_501) );
INVxp67_ASAP7_75t_SL g502 ( .A(n_436), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_436), .B(n_413), .Y(n_503) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_449), .A2(n_413), .B(n_231), .Y(n_504) );
NAND4xp25_ASAP7_75t_L g505 ( .A(n_458), .B(n_218), .C(n_241), .D(n_238), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_435), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_436), .B(n_464), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_455), .B(n_413), .Y(n_508) );
INVx4_ASAP7_75t_L g509 ( .A(n_451), .Y(n_509) );
INVxp67_ASAP7_75t_SL g510 ( .A(n_452), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_451), .B(n_367), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_435), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_460), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_456), .B(n_27), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_460), .B(n_28), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_438), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_483), .A2(n_434), .B1(n_462), .B2(n_460), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_473), .B(n_460), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_471), .B(n_463), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_503), .B(n_31), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_470), .B(n_41), .Y(n_521) );
AND2x4_ASAP7_75t_L g522 ( .A(n_500), .B(n_42), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_470), .B(n_43), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_474), .B(n_342), .Y(n_524) );
NAND2xp33_ASAP7_75t_SL g525 ( .A(n_469), .B(n_342), .Y(n_525) );
BUFx4f_ASAP7_75t_L g526 ( .A(n_469), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_474), .B(n_342), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_503), .B(n_44), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_491), .B(n_48), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_477), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_491), .B(n_50), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_508), .B(n_52), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_485), .B(n_338), .Y(n_533) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_501), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_499), .B(n_56), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_468), .A2(n_338), .B1(n_336), .B2(n_334), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_486), .Y(n_537) );
NOR2xp33_ASAP7_75t_R g538 ( .A(n_472), .B(n_57), .Y(n_538) );
INVx1_ASAP7_75t_SL g539 ( .A(n_494), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_477), .Y(n_540) );
AND2x2_ASAP7_75t_SL g541 ( .A(n_509), .B(n_338), .Y(n_541) );
BUFx2_ASAP7_75t_L g542 ( .A(n_501), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_493), .B(n_59), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_468), .A2(n_336), .B1(n_334), .B2(n_209), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_490), .A2(n_334), .B1(n_336), .B2(n_203), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_477), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_467), .B(n_60), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_507), .B(n_336), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_493), .B(n_61), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_496), .B(n_66), .Y(n_550) );
OAI21xp33_ASAP7_75t_SL g551 ( .A1(n_509), .A2(n_68), .B(n_69), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_472), .B(n_513), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_495), .B(n_70), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_495), .B(n_71), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_468), .B(n_72), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_467), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_479), .B(n_73), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_497), .B(n_75), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_468), .B(n_500), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_497), .Y(n_560) );
AOI31xp33_ASAP7_75t_L g561 ( .A1(n_515), .A2(n_78), .A3(n_183), .B(n_203), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_489), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_502), .B(n_241), .Y(n_563) );
NOR4xp25_ASAP7_75t_SL g564 ( .A(n_488), .B(n_516), .C(n_510), .D(n_506), .Y(n_564) );
AO22x1_ASAP7_75t_L g565 ( .A1(n_509), .A2(n_220), .B1(n_218), .B2(n_216), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_480), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_500), .B(n_216), .Y(n_567) );
OAI22xp33_ASAP7_75t_SL g568 ( .A1(n_526), .A2(n_509), .B1(n_478), .B2(n_484), .Y(n_568) );
AOI321xp33_ASAP7_75t_L g569 ( .A1(n_519), .A2(n_476), .A3(n_514), .B1(n_500), .B2(n_515), .C(n_482), .Y(n_569) );
NOR2xp33_ASAP7_75t_R g570 ( .A(n_526), .B(n_484), .Y(n_570) );
NAND2xp33_ASAP7_75t_SL g571 ( .A(n_538), .B(n_478), .Y(n_571) );
INVxp67_ASAP7_75t_SL g572 ( .A(n_534), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_556), .B(n_481), .Y(n_573) );
NOR2x1_ASAP7_75t_L g574 ( .A(n_539), .B(n_484), .Y(n_574) );
NAND2x1p5_ASAP7_75t_L g575 ( .A(n_526), .B(n_484), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_566), .B(n_481), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_517), .A2(n_487), .B1(n_514), .B2(n_513), .Y(n_577) );
AOI322xp5_ASAP7_75t_L g578 ( .A1(n_551), .A2(n_492), .A3(n_498), .B1(n_511), .B2(n_512), .C1(n_487), .C2(n_475), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_537), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_542), .B(n_480), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_560), .B(n_512), .Y(n_581) );
OAI21xp33_ASAP7_75t_SL g582 ( .A1(n_541), .A2(n_492), .B(n_511), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_562), .Y(n_583) );
AOI22xp33_ASAP7_75t_SL g584 ( .A1(n_538), .A2(n_528), .B1(n_520), .B2(n_531), .Y(n_584) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_530), .Y(n_585) );
AOI221xp5_ASAP7_75t_L g586 ( .A1(n_518), .A2(n_505), .B1(n_504), .B2(n_225), .C(n_209), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_552), .B(n_505), .Y(n_587) );
NOR3xp33_ASAP7_75t_L g588 ( .A(n_561), .B(n_504), .C(n_212), .Y(n_588) );
OAI21xp5_ASAP7_75t_SL g589 ( .A1(n_522), .A2(n_209), .B(n_212), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_540), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_528), .A2(n_209), .B1(n_212), .B2(n_225), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_529), .B(n_225), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_531), .B(n_285), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_540), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_546), .Y(n_595) );
AOI21xp5_ASAP7_75t_L g596 ( .A1(n_525), .A2(n_285), .B(n_301), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_546), .Y(n_597) );
NAND3xp33_ASAP7_75t_SL g598 ( .A(n_564), .B(n_301), .C(n_547), .Y(n_598) );
INVxp67_ASAP7_75t_L g599 ( .A(n_543), .Y(n_599) );
AND2x4_ASAP7_75t_SL g600 ( .A(n_559), .B(n_522), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_535), .B(n_548), .Y(n_601) );
AOI33xp33_ASAP7_75t_L g602 ( .A1(n_549), .A2(n_554), .A3(n_553), .B1(n_555), .B2(n_522), .B3(n_567), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_580), .B(n_572), .Y(n_603) );
NAND2xp33_ASAP7_75t_SL g604 ( .A(n_570), .B(n_535), .Y(n_604) );
NAND2xp5_ASAP7_75t_SL g605 ( .A(n_568), .B(n_557), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_587), .B(n_532), .Y(n_606) );
OAI22xp33_ASAP7_75t_L g607 ( .A1(n_599), .A2(n_521), .B1(n_523), .B2(n_557), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_576), .B(n_524), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_600), .B(n_554), .Y(n_609) );
XNOR2xp5_ASAP7_75t_L g610 ( .A(n_584), .B(n_521), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_599), .B(n_523), .Y(n_611) );
INVx1_ASAP7_75t_SL g612 ( .A(n_571), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_602), .B(n_527), .Y(n_613) );
AOI21xp33_ASAP7_75t_L g614 ( .A1(n_582), .A2(n_550), .B(n_558), .Y(n_614) );
NOR2x1_ASAP7_75t_L g615 ( .A(n_589), .B(n_574), .Y(n_615) );
XNOR2x1_ASAP7_75t_L g616 ( .A(n_575), .B(n_565), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_579), .Y(n_617) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_588), .B(n_545), .Y(n_618) );
INVx4_ASAP7_75t_L g619 ( .A(n_575), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_585), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_583), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_584), .A2(n_536), .B1(n_544), .B2(n_533), .Y(n_622) );
O2A1O1Ixp33_ASAP7_75t_SL g623 ( .A1(n_569), .A2(n_563), .B(n_578), .C(n_598), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g624 ( .A1(n_588), .A2(n_598), .B(n_586), .Y(n_624) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_585), .Y(n_625) );
XNOR2xp5_ASAP7_75t_L g626 ( .A(n_577), .B(n_573), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_581), .Y(n_627) );
BUFx2_ASAP7_75t_L g628 ( .A(n_625), .Y(n_628) );
AND2x4_ASAP7_75t_SL g629 ( .A(n_619), .B(n_601), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g630 ( .A(n_612), .B(n_596), .Y(n_630) );
NOR3xp33_ASAP7_75t_SL g631 ( .A(n_624), .B(n_592), .C(n_593), .Y(n_631) );
OAI31xp33_ASAP7_75t_SL g632 ( .A1(n_610), .A2(n_590), .A3(n_594), .B(n_595), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_626), .B(n_597), .Y(n_633) );
NOR3xp33_ASAP7_75t_L g634 ( .A(n_623), .B(n_591), .C(n_618), .Y(n_634) );
AOI221xp5_ASAP7_75t_L g635 ( .A1(n_606), .A2(n_613), .B1(n_627), .B2(n_611), .C(n_617), .Y(n_635) );
A2O1A1Ixp33_ASAP7_75t_L g636 ( .A1(n_604), .A2(n_615), .B(n_605), .C(n_606), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_621), .B(n_608), .Y(n_637) );
NAND2x1_ASAP7_75t_L g638 ( .A(n_609), .B(n_620), .Y(n_638) );
OAI21xp33_ASAP7_75t_L g639 ( .A1(n_605), .A2(n_603), .B(n_618), .Y(n_639) );
NOR3xp33_ASAP7_75t_L g640 ( .A(n_614), .B(n_622), .C(n_604), .Y(n_640) );
AOI21xp33_ASAP7_75t_L g641 ( .A1(n_639), .A2(n_616), .B(n_611), .Y(n_641) );
NOR2x1_ASAP7_75t_L g642 ( .A(n_636), .B(n_607), .Y(n_642) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_628), .Y(n_643) );
INVx2_ASAP7_75t_SL g644 ( .A(n_629), .Y(n_644) );
OAI21xp5_ASAP7_75t_SL g645 ( .A1(n_636), .A2(n_632), .B(n_634), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g646 ( .A1(n_640), .A2(n_635), .B1(n_633), .B2(n_637), .C(n_631), .Y(n_646) );
AND2x4_ASAP7_75t_L g647 ( .A(n_629), .B(n_638), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g648 ( .A1(n_640), .A2(n_639), .B1(n_635), .B2(n_634), .C(n_636), .Y(n_648) );
OAI21xp33_ASAP7_75t_SL g649 ( .A1(n_632), .A2(n_630), .B(n_605), .Y(n_649) );
NAND4xp25_ASAP7_75t_SL g650 ( .A(n_636), .B(n_640), .C(n_634), .D(n_584), .Y(n_650) );
NAND3xp33_ASAP7_75t_SL g651 ( .A(n_636), .B(n_634), .C(n_640), .Y(n_651) );
INVx1_ASAP7_75t_SL g652 ( .A(n_644), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_643), .Y(n_653) );
CKINVDCx5p33_ASAP7_75t_R g654 ( .A(n_644), .Y(n_654) );
CKINVDCx5p33_ASAP7_75t_R g655 ( .A(n_651), .Y(n_655) );
INVx1_ASAP7_75t_SL g656 ( .A(n_647), .Y(n_656) );
NOR4xp25_ASAP7_75t_L g657 ( .A(n_652), .B(n_650), .C(n_645), .D(n_648), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_653), .Y(n_658) );
AOI22xp33_ASAP7_75t_SL g659 ( .A1(n_657), .A2(n_655), .B1(n_652), .B2(n_656), .Y(n_659) );
OR2x2_ASAP7_75t_L g660 ( .A(n_658), .B(n_654), .Y(n_660) );
INVxp67_ASAP7_75t_SL g661 ( .A(n_660), .Y(n_661) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_659), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_662), .A2(n_661), .B1(n_642), .B2(n_649), .Y(n_663) );
AOI21xp5_ASAP7_75t_L g664 ( .A1(n_663), .A2(n_646), .B(n_641), .Y(n_664) );
endmodule