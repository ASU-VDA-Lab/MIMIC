module real_aes_8594_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_505;
wire n_434;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_712;
wire n_183;
wire n_312;
wire n_266;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_719;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g109 ( .A(n_0), .Y(n_109) );
A2O1A1Ixp33_ASAP7_75t_L g451 ( .A1(n_1), .A2(n_140), .B(n_152), .C(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g259 ( .A(n_2), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_3), .A2(n_167), .B(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_4), .B(n_163), .Y(n_496) );
AOI21xp33_ASAP7_75t_L g166 ( .A1(n_5), .A2(n_167), .B(n_168), .Y(n_166) );
AND2x6_ASAP7_75t_L g140 ( .A(n_6), .B(n_141), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_7), .A2(n_235), .B(n_236), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g110 ( .A(n_8), .B(n_40), .Y(n_110) );
INVx1_ASAP7_75t_L g467 ( .A(n_9), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_10), .B(n_173), .Y(n_455) );
INVx1_ASAP7_75t_L g175 ( .A(n_11), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_12), .B(n_227), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_13), .A2(n_100), .B1(n_111), .B2(n_723), .Y(n_99) );
INVx1_ASAP7_75t_L g137 ( .A(n_14), .Y(n_137) );
INVx1_ASAP7_75t_L g241 ( .A(n_15), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g475 ( .A1(n_16), .A2(n_176), .B(n_242), .C(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_17), .B(n_163), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_18), .B(n_186), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_19), .B(n_167), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_20), .B(n_509), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_L g483 ( .A1(n_21), .A2(n_143), .B(n_227), .C(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_22), .B(n_163), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_23), .B(n_173), .Y(n_530) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_24), .A2(n_239), .B(n_240), .C(n_242), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_25), .B(n_173), .Y(n_517) );
CKINVDCx16_ASAP7_75t_R g526 ( .A(n_26), .Y(n_526) );
INVx1_ASAP7_75t_L g516 ( .A(n_27), .Y(n_516) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_28), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_29), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_30), .B(n_173), .Y(n_260) );
INVx1_ASAP7_75t_L g505 ( .A(n_31), .Y(n_505) );
INVx1_ASAP7_75t_L g151 ( .A(n_32), .Y(n_151) );
INVx2_ASAP7_75t_L g145 ( .A(n_33), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_34), .Y(n_457) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_35), .A2(n_177), .B(n_227), .C(n_494), .Y(n_493) );
INVxp67_ASAP7_75t_L g506 ( .A(n_36), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_37), .A2(n_140), .B(n_152), .C(n_197), .Y(n_196) );
CKINVDCx14_ASAP7_75t_R g492 ( .A(n_38), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g514 ( .A1(n_39), .A2(n_152), .B(n_515), .C(n_519), .Y(n_514) );
INVx1_ASAP7_75t_L g149 ( .A(n_41), .Y(n_149) );
A2O1A1Ixp33_ASAP7_75t_L g465 ( .A1(n_42), .A2(n_172), .B(n_202), .C(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_43), .B(n_173), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_44), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_45), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_46), .Y(n_121) );
INVx1_ASAP7_75t_L g482 ( .A(n_47), .Y(n_482) );
CKINVDCx16_ASAP7_75t_R g155 ( .A(n_48), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_49), .B(n_167), .Y(n_229) );
AOI222xp33_ASAP7_75t_SL g122 ( .A1(n_50), .A2(n_59), .B1(n_123), .B2(n_709), .C1(n_710), .C2(n_714), .Y(n_122) );
AOI22xp5_ASAP7_75t_L g142 ( .A1(n_51), .A2(n_143), .B1(n_146), .B2(n_152), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g206 ( .A(n_52), .Y(n_206) );
CKINVDCx16_ASAP7_75t_R g256 ( .A(n_53), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_L g171 ( .A1(n_54), .A2(n_172), .B(n_174), .C(n_177), .Y(n_171) );
CKINVDCx14_ASAP7_75t_R g464 ( .A(n_55), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_56), .Y(n_216) );
INVx1_ASAP7_75t_L g169 ( .A(n_57), .Y(n_169) );
INVx1_ASAP7_75t_L g141 ( .A(n_58), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_59), .Y(n_709) );
INVx1_ASAP7_75t_L g136 ( .A(n_60), .Y(n_136) );
INVx1_ASAP7_75t_SL g495 ( .A(n_61), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_62), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_63), .B(n_163), .Y(n_486) );
OAI22xp5_ASAP7_75t_SL g719 ( .A1(n_64), .A2(n_441), .B1(n_711), .B2(n_720), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_64), .Y(n_720) );
INVx1_ASAP7_75t_L g529 ( .A(n_65), .Y(n_529) );
A2O1A1Ixp33_ASAP7_75t_SL g185 ( .A1(n_66), .A2(n_177), .B(n_186), .C(n_187), .Y(n_185) );
INVxp67_ASAP7_75t_L g188 ( .A(n_67), .Y(n_188) );
INVx1_ASAP7_75t_L g104 ( .A(n_68), .Y(n_104) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_69), .A2(n_167), .B(n_463), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_70), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_71), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_72), .A2(n_167), .B(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g209 ( .A(n_73), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_74), .A2(n_235), .B(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g474 ( .A(n_75), .Y(n_474) );
CKINVDCx16_ASAP7_75t_R g513 ( .A(n_76), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g210 ( .A1(n_77), .A2(n_140), .B(n_152), .C(n_211), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_78), .A2(n_167), .B(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g477 ( .A(n_79), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_80), .B(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g134 ( .A(n_81), .Y(n_134) );
INVx1_ASAP7_75t_L g453 ( .A(n_82), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_83), .B(n_186), .Y(n_200) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_84), .A2(n_140), .B(n_152), .C(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g106 ( .A(n_85), .B(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g440 ( .A(n_85), .Y(n_440) );
OR2x2_ASAP7_75t_L g708 ( .A(n_85), .B(n_108), .Y(n_708) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_86), .A2(n_152), .B(n_528), .C(n_531), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_87), .B(n_180), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g263 ( .A(n_88), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_89), .A2(n_140), .B(n_152), .C(n_224), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g231 ( .A(n_90), .Y(n_231) );
INVx1_ASAP7_75t_L g184 ( .A(n_91), .Y(n_184) );
CKINVDCx16_ASAP7_75t_R g237 ( .A(n_92), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_93), .B(n_199), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_94), .B(n_165), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_95), .B(n_165), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_96), .B(n_104), .Y(n_103) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_97), .A2(n_167), .B(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g485 ( .A(n_98), .Y(n_485) );
INVx2_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g724 ( .A(n_101), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g101 ( .A(n_102), .B(n_105), .Y(n_101) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_SL g120 ( .A(n_106), .Y(n_120) );
INVx1_ASAP7_75t_SL g722 ( .A(n_106), .Y(n_722) );
NOR2x2_ASAP7_75t_L g716 ( .A(n_107), .B(n_440), .Y(n_716) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
OR2x2_ASAP7_75t_L g439 ( .A(n_108), .B(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AOI22xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_122), .B1(n_717), .B2(n_718), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_114), .B(n_118), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_SL g717 ( .A(n_115), .Y(n_717) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g718 ( .A1(n_118), .A2(n_719), .B(n_721), .Y(n_718) );
NOR2xp33_ASAP7_75t_SL g118 ( .A(n_119), .B(n_121), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_124), .A2(n_437), .B1(n_441), .B2(n_708), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OAI22xp5_ASAP7_75t_SL g710 ( .A1(n_125), .A2(n_437), .B1(n_711), .B2(n_712), .Y(n_710) );
AND3x1_ASAP7_75t_L g125 ( .A(n_126), .B(n_362), .C(n_411), .Y(n_125) );
NOR3xp33_ASAP7_75t_SL g126 ( .A(n_127), .B(n_269), .C(n_307), .Y(n_126) );
OAI222xp33_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_190), .B1(n_244), .B2(n_250), .C1(n_264), .C2(n_267), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_161), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_129), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_129), .B(n_312), .Y(n_403) );
BUFx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OR2x2_ASAP7_75t_L g280 ( .A(n_130), .B(n_181), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_130), .B(n_162), .Y(n_288) );
AND2x2_ASAP7_75t_L g323 ( .A(n_130), .B(n_300), .Y(n_323) );
OR2x2_ASAP7_75t_L g347 ( .A(n_130), .B(n_162), .Y(n_347) );
OR2x2_ASAP7_75t_L g355 ( .A(n_130), .B(n_254), .Y(n_355) );
AND2x2_ASAP7_75t_L g358 ( .A(n_130), .B(n_181), .Y(n_358) );
INVx3_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OR2x2_ASAP7_75t_L g252 ( .A(n_131), .B(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g266 ( .A(n_131), .B(n_181), .Y(n_266) );
AND2x2_ASAP7_75t_L g316 ( .A(n_131), .B(n_254), .Y(n_316) );
AND2x2_ASAP7_75t_L g329 ( .A(n_131), .B(n_162), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_131), .B(n_415), .Y(n_436) );
AO21x2_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_138), .B(n_159), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_132), .B(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g204 ( .A(n_132), .Y(n_204) );
AO21x2_ASAP7_75t_L g254 ( .A1(n_132), .A2(n_255), .B(n_262), .Y(n_254) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_133), .Y(n_165) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
AND2x2_ASAP7_75t_SL g180 ( .A(n_134), .B(n_135), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
OAI22xp33_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_142), .B1(n_155), .B2(n_156), .Y(n_138) );
O2A1O1Ixp33_ASAP7_75t_L g168 ( .A1(n_139), .A2(n_169), .B(n_170), .C(n_171), .Y(n_168) );
O2A1O1Ixp33_ASAP7_75t_L g183 ( .A1(n_139), .A2(n_170), .B(n_184), .C(n_185), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_L g236 ( .A1(n_139), .A2(n_170), .B(n_237), .C(n_238), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_SL g463 ( .A1(n_139), .A2(n_170), .B(n_464), .C(n_465), .Y(n_463) );
O2A1O1Ixp33_ASAP7_75t_SL g473 ( .A1(n_139), .A2(n_170), .B(n_474), .C(n_475), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_SL g481 ( .A1(n_139), .A2(n_170), .B(n_482), .C(n_483), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_139), .A2(n_170), .B(n_492), .C(n_493), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_SL g501 ( .A1(n_139), .A2(n_170), .B(n_502), .C(n_503), .Y(n_501) );
INVx1_ASAP7_75t_L g531 ( .A(n_139), .Y(n_531) );
INVx4_ASAP7_75t_SL g139 ( .A(n_140), .Y(n_139) );
NAND2x1p5_ASAP7_75t_L g156 ( .A(n_140), .B(n_157), .Y(n_156) );
AND2x4_ASAP7_75t_L g167 ( .A(n_140), .B(n_157), .Y(n_167) );
BUFx3_ASAP7_75t_L g519 ( .A(n_140), .Y(n_519) );
INVx2_ASAP7_75t_L g261 ( .A(n_143), .Y(n_261) );
INVx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g153 ( .A(n_145), .Y(n_153) );
INVx1_ASAP7_75t_L g158 ( .A(n_145), .Y(n_158) );
OAI22xp5_ASAP7_75t_SL g146 ( .A1(n_147), .A2(n_149), .B1(n_150), .B2(n_151), .Y(n_146) );
INVx2_ASAP7_75t_L g150 ( .A(n_147), .Y(n_150) );
INVx4_ASAP7_75t_L g239 ( .A(n_147), .Y(n_239) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g154 ( .A(n_148), .Y(n_154) );
AND2x2_ASAP7_75t_L g157 ( .A(n_148), .B(n_158), .Y(n_157) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_148), .Y(n_173) );
INVx3_ASAP7_75t_L g176 ( .A(n_148), .Y(n_176) );
INVx1_ASAP7_75t_L g186 ( .A(n_148), .Y(n_186) );
INVx2_ASAP7_75t_L g454 ( .A(n_150), .Y(n_454) );
INVx5_ASAP7_75t_L g170 ( .A(n_152), .Y(n_170) );
AND2x6_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_153), .Y(n_178) );
BUFx3_ASAP7_75t_L g203 ( .A(n_153), .Y(n_203) );
OAI21xp5_ASAP7_75t_L g208 ( .A1(n_156), .A2(n_209), .B(n_210), .Y(n_208) );
OAI21xp5_ASAP7_75t_L g255 ( .A1(n_156), .A2(n_256), .B(n_257), .Y(n_255) );
OAI21xp5_ASAP7_75t_L g449 ( .A1(n_156), .A2(n_450), .B(n_451), .Y(n_449) );
O2A1O1Ixp33_ASAP7_75t_L g512 ( .A1(n_156), .A2(n_180), .B(n_513), .C(n_514), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g525 ( .A1(n_156), .A2(n_526), .B(n_527), .Y(n_525) );
INVx1_ASAP7_75t_L g507 ( .A(n_158), .Y(n_507) );
O2A1O1Ixp33_ASAP7_75t_L g354 ( .A1(n_161), .A2(n_355), .B(n_356), .C(n_359), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_161), .B(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_161), .B(n_299), .Y(n_421) );
AND2x2_ASAP7_75t_L g161 ( .A(n_162), .B(n_181), .Y(n_161) );
AND2x2_ASAP7_75t_SL g265 ( .A(n_162), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g279 ( .A(n_162), .Y(n_279) );
AND2x2_ASAP7_75t_L g306 ( .A(n_162), .B(n_300), .Y(n_306) );
INVx1_ASAP7_75t_SL g314 ( .A(n_162), .Y(n_314) );
AND2x2_ASAP7_75t_L g337 ( .A(n_162), .B(n_338), .Y(n_337) );
BUFx2_ASAP7_75t_L g415 ( .A(n_162), .Y(n_415) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_166), .B(n_179), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NOR2xp33_ASAP7_75t_SL g205 ( .A(n_164), .B(n_206), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_164), .B(n_457), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_164), .B(n_521), .Y(n_520) );
AO21x2_ASAP7_75t_L g524 ( .A1(n_164), .A2(n_525), .B(n_532), .Y(n_524) );
INVx4_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
OA21x2_ASAP7_75t_L g181 ( .A1(n_165), .A2(n_182), .B(n_189), .Y(n_181) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_165), .Y(n_471) );
BUFx2_ASAP7_75t_L g235 ( .A(n_167), .Y(n_235) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx4_ASAP7_75t_L g227 ( .A(n_173), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_175), .B(n_176), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_176), .B(n_188), .Y(n_187) );
INVx5_ASAP7_75t_L g199 ( .A(n_176), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_176), .B(n_467), .Y(n_466) );
INVx3_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_178), .Y(n_228) );
INVx1_ASAP7_75t_L g217 ( .A(n_180), .Y(n_217) );
INVx2_ASAP7_75t_L g221 ( .A(n_180), .Y(n_221) );
OA21x2_ASAP7_75t_L g233 ( .A1(n_180), .A2(n_234), .B(n_243), .Y(n_233) );
OA21x2_ASAP7_75t_L g461 ( .A1(n_180), .A2(n_462), .B(n_468), .Y(n_461) );
BUFx2_ASAP7_75t_L g251 ( .A(n_181), .Y(n_251) );
INVx1_ASAP7_75t_L g313 ( .A(n_181), .Y(n_313) );
INVx3_ASAP7_75t_L g338 ( .A(n_181), .Y(n_338) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_190), .B(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_218), .Y(n_190) );
INVx1_ASAP7_75t_L g334 ( .A(n_191), .Y(n_334) );
OAI32xp33_ASAP7_75t_L g340 ( .A1(n_191), .A2(n_279), .A3(n_341), .B1(n_342), .B2(n_343), .Y(n_340) );
OAI22xp5_ASAP7_75t_L g344 ( .A1(n_191), .A2(n_345), .B1(n_348), .B2(n_353), .Y(n_344) );
INVx4_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_L g282 ( .A(n_192), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g360 ( .A(n_192), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g430 ( .A(n_192), .B(n_376), .Y(n_430) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_207), .Y(n_192) );
AND2x2_ASAP7_75t_L g245 ( .A(n_193), .B(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g275 ( .A(n_193), .Y(n_275) );
INVx1_ASAP7_75t_L g294 ( .A(n_193), .Y(n_294) );
OR2x2_ASAP7_75t_L g302 ( .A(n_193), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g309 ( .A(n_193), .B(n_283), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_193), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g330 ( .A(n_193), .B(n_248), .Y(n_330) );
INVx3_ASAP7_75t_L g352 ( .A(n_193), .Y(n_352) );
AND2x2_ASAP7_75t_L g377 ( .A(n_193), .B(n_249), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_193), .B(n_342), .Y(n_425) );
OR2x6_ASAP7_75t_L g193 ( .A(n_194), .B(n_205), .Y(n_193) );
AOI21xp5_ASAP7_75t_SL g194 ( .A1(n_195), .A2(n_196), .B(n_204), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_200), .B(n_201), .Y(n_197) );
O2A1O1Ixp33_ASAP7_75t_L g258 ( .A1(n_199), .A2(n_259), .B(n_260), .C(n_261), .Y(n_258) );
OAI22xp33_ASAP7_75t_L g504 ( .A1(n_199), .A2(n_239), .B1(n_505), .B2(n_506), .Y(n_504) );
O2A1O1Ixp33_ASAP7_75t_L g515 ( .A1(n_199), .A2(n_516), .B(n_517), .C(n_518), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_201), .A2(n_212), .B(n_213), .Y(n_211) );
O2A1O1Ixp5_ASAP7_75t_L g452 ( .A1(n_201), .A2(n_453), .B(n_454), .C(n_455), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_L g528 ( .A1(n_201), .A2(n_454), .B(n_529), .C(n_530), .Y(n_528) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g242 ( .A(n_203), .Y(n_242) );
INVx1_ASAP7_75t_L g214 ( .A(n_204), .Y(n_214) );
INVx2_ASAP7_75t_L g249 ( .A(n_207), .Y(n_249) );
AND2x2_ASAP7_75t_L g381 ( .A(n_207), .B(n_219), .Y(n_381) );
AO21x2_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_214), .B(n_215), .Y(n_207) );
INVx1_ASAP7_75t_L g499 ( .A(n_214), .Y(n_499) );
AO21x2_ASAP7_75t_L g551 ( .A1(n_214), .A2(n_552), .B(n_553), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_216), .B(n_217), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_217), .B(n_231), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_217), .B(n_263), .Y(n_262) );
AO21x2_ASAP7_75t_L g448 ( .A1(n_217), .A2(n_449), .B(n_456), .Y(n_448) );
INVx2_ASAP7_75t_L g423 ( .A(n_218), .Y(n_423) );
OR2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_232), .Y(n_218) );
INVx1_ASAP7_75t_L g268 ( .A(n_219), .Y(n_268) );
AND2x2_ASAP7_75t_L g295 ( .A(n_219), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_219), .B(n_249), .Y(n_303) );
AND2x2_ASAP7_75t_L g361 ( .A(n_219), .B(n_284), .Y(n_361) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g247 ( .A(n_220), .Y(n_247) );
AND2x2_ASAP7_75t_L g274 ( .A(n_220), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g283 ( .A(n_220), .B(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_220), .B(n_249), .Y(n_349) );
AO21x2_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_230), .Y(n_220) );
INVx1_ASAP7_75t_L g509 ( .A(n_221), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_221), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_223), .B(n_229), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_228), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_227), .B(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_232), .B(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g296 ( .A(n_232), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_232), .B(n_249), .Y(n_342) );
AND2x2_ASAP7_75t_L g351 ( .A(n_232), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g376 ( .A(n_232), .Y(n_376) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g248 ( .A(n_233), .B(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g284 ( .A(n_233), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_239), .B(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_239), .B(n_477), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_239), .B(n_485), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_244), .A2(n_254), .B1(n_413), .B2(n_416), .Y(n_412) );
INVx1_ASAP7_75t_SL g244 ( .A(n_245), .Y(n_244) );
OAI21xp5_ASAP7_75t_SL g435 ( .A1(n_246), .A2(n_357), .B(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_247), .B(n_352), .Y(n_369) );
INVx1_ASAP7_75t_L g394 ( .A(n_247), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_248), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g321 ( .A(n_248), .B(n_274), .Y(n_321) );
INVx2_ASAP7_75t_L g277 ( .A(n_249), .Y(n_277) );
INVx1_ASAP7_75t_L g327 ( .A(n_249), .Y(n_327) );
OAI221xp5_ASAP7_75t_L g418 ( .A1(n_250), .A2(n_402), .B1(n_419), .B2(n_422), .C(n_424), .Y(n_418) );
OR2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
INVx1_ASAP7_75t_L g289 ( .A(n_251), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_251), .B(n_300), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_252), .B(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g343 ( .A(n_252), .B(n_289), .Y(n_343) );
INVx3_ASAP7_75t_SL g384 ( .A(n_252), .Y(n_384) );
AND2x2_ASAP7_75t_L g328 ( .A(n_253), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g357 ( .A(n_253), .B(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_253), .B(n_266), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_253), .B(n_312), .Y(n_398) );
INVx3_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx3_ASAP7_75t_L g300 ( .A(n_254), .Y(n_300) );
OAI322xp33_ASAP7_75t_L g395 ( .A1(n_254), .A2(n_326), .A3(n_348), .B1(n_396), .B2(n_398), .C1(n_399), .C2(n_400), .Y(n_395) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AOI21xp33_ASAP7_75t_L g419 ( .A1(n_265), .A2(n_268), .B(n_420), .Y(n_419) );
NOR2xp33_ASAP7_75t_SL g345 ( .A(n_266), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g367 ( .A(n_266), .B(n_279), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_266), .B(n_306), .Y(n_382) );
INVxp67_ASAP7_75t_L g333 ( .A(n_268), .Y(n_333) );
AOI211xp5_ASAP7_75t_L g339 ( .A1(n_268), .A2(n_340), .B(n_344), .C(n_354), .Y(n_339) );
OAI221xp5_ASAP7_75t_SL g269 ( .A1(n_270), .A2(n_278), .B1(n_281), .B2(n_285), .C(n_290), .Y(n_269) );
INVxp67_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_276), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g293 ( .A(n_277), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g410 ( .A(n_277), .Y(n_410) );
OAI221xp5_ASAP7_75t_L g426 ( .A1(n_278), .A2(n_427), .B1(n_432), .B2(n_433), .C(n_435), .Y(n_426) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_279), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_SL g326 ( .A(n_279), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_279), .B(n_357), .Y(n_364) );
AND2x2_ASAP7_75t_L g406 ( .A(n_279), .B(n_384), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g304 ( .A(n_280), .B(n_305), .Y(n_304) );
OAI22xp33_ASAP7_75t_L g401 ( .A1(n_280), .A2(n_292), .B1(n_402), .B2(n_403), .Y(n_401) );
OR2x2_ASAP7_75t_L g432 ( .A(n_280), .B(n_300), .Y(n_432) );
CKINVDCx16_ASAP7_75t_R g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g409 ( .A(n_283), .Y(n_409) );
AND2x2_ASAP7_75t_L g434 ( .A(n_283), .B(n_377), .Y(n_434) );
INVxp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NOR2xp33_ASAP7_75t_SL g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g298 ( .A(n_288), .B(n_299), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_297), .B1(n_301), .B2(n_304), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
INVx1_ASAP7_75t_L g365 ( .A(n_293), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_293), .B(n_333), .Y(n_400) );
AOI322xp5_ASAP7_75t_L g324 ( .A1(n_295), .A2(n_325), .A3(n_327), .B1(n_328), .B2(n_330), .C1(n_331), .C2(n_335), .Y(n_324) );
INVxp67_ASAP7_75t_L g318 ( .A(n_296), .Y(n_318) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OAI22xp5_ASAP7_75t_L g319 ( .A1(n_298), .A2(n_303), .B1(n_320), .B2(n_322), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_299), .B(n_312), .Y(n_399) );
INVx1_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_300), .B(n_338), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_300), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g396 ( .A(n_302), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
NAND3xp33_ASAP7_75t_SL g307 ( .A(n_308), .B(n_324), .C(n_339), .Y(n_307) );
AOI221xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_310), .B1(n_315), .B2(n_317), .C(n_319), .Y(n_308) );
AND2x2_ASAP7_75t_L g315 ( .A(n_311), .B(n_316), .Y(n_315) );
INVx3_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
AND2x4_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
AND2x2_ASAP7_75t_L g325 ( .A(n_316), .B(n_326), .Y(n_325) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_318), .Y(n_397) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_323), .B(n_337), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_326), .B(n_384), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_327), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_SL g402 ( .A(n_330), .Y(n_402) );
AND2x2_ASAP7_75t_L g417 ( .A(n_330), .B(n_394), .Y(n_417) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AOI211xp5_ASAP7_75t_L g411 ( .A1(n_341), .A2(n_412), .B(n_418), .C(n_426), .Y(n_411) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g380 ( .A(n_351), .B(n_381), .Y(n_380) );
NAND2x1_ASAP7_75t_SL g422 ( .A(n_352), .B(n_423), .Y(n_422) );
CKINVDCx16_ASAP7_75t_R g392 ( .A(n_355), .Y(n_392) );
INVx1_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g387 ( .A(n_361), .Y(n_387) );
AND2x2_ASAP7_75t_L g391 ( .A(n_361), .B(n_377), .Y(n_391) );
NOR5xp2_ASAP7_75t_L g362 ( .A(n_363), .B(n_378), .C(n_395), .D(n_401), .E(n_404), .Y(n_362) );
OAI221xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_365), .B1(n_366), .B2(n_368), .C(n_370), .Y(n_363) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_367), .B(n_425), .Y(n_424) );
INVxp67_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_373), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_375), .B(n_377), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g393 ( .A(n_377), .B(n_394), .Y(n_393) );
OAI221xp5_ASAP7_75t_SL g378 ( .A1(n_379), .A2(n_382), .B1(n_383), .B2(n_385), .C(n_388), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_391), .B1(n_392), .B2(n_393), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g431 ( .A(n_391), .Y(n_431) );
AOI211xp5_ASAP7_75t_SL g404 ( .A1(n_405), .A2(n_407), .B(n_409), .C(n_410), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVxp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_431), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
CKINVDCx14_ASAP7_75t_R g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g711 ( .A(n_441), .Y(n_711) );
OR2x2_ASAP7_75t_SL g441 ( .A(n_442), .B(n_663), .Y(n_441) );
NAND5xp2_ASAP7_75t_L g442 ( .A(n_443), .B(n_575), .C(n_613), .D(n_634), .E(n_651), .Y(n_442) );
NOR3xp33_ASAP7_75t_L g443 ( .A(n_444), .B(n_547), .C(n_568), .Y(n_443) );
OAI221xp5_ASAP7_75t_SL g444 ( .A1(n_445), .A2(n_487), .B1(n_510), .B2(n_534), .C(n_538), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_458), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_447), .B(n_536), .Y(n_555) );
OR2x2_ASAP7_75t_L g582 ( .A(n_447), .B(n_470), .Y(n_582) );
AND2x2_ASAP7_75t_L g596 ( .A(n_447), .B(n_470), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_447), .B(n_461), .Y(n_610) );
AND2x2_ASAP7_75t_L g648 ( .A(n_447), .B(n_612), .Y(n_648) );
AND2x2_ASAP7_75t_L g677 ( .A(n_447), .B(n_587), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_447), .B(n_559), .Y(n_694) );
INVx4_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g574 ( .A(n_448), .B(n_469), .Y(n_574) );
BUFx3_ASAP7_75t_L g599 ( .A(n_448), .Y(n_599) );
AND2x2_ASAP7_75t_L g628 ( .A(n_448), .B(n_470), .Y(n_628) );
AND3x2_ASAP7_75t_L g641 ( .A(n_448), .B(n_642), .C(n_643), .Y(n_641) );
INVx1_ASAP7_75t_L g564 ( .A(n_458), .Y(n_564) );
AND2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_469), .Y(n_458) );
AOI32xp33_ASAP7_75t_L g619 ( .A1(n_459), .A2(n_571), .A3(n_620), .B1(n_623), .B2(n_624), .Y(n_619) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g546 ( .A(n_460), .B(n_469), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g617 ( .A(n_460), .B(n_574), .Y(n_617) );
AND2x2_ASAP7_75t_L g624 ( .A(n_460), .B(n_596), .Y(n_624) );
OR2x2_ASAP7_75t_L g630 ( .A(n_460), .B(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_460), .B(n_585), .Y(n_655) );
OR2x2_ASAP7_75t_L g673 ( .A(n_460), .B(n_498), .Y(n_673) );
BUFx3_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g537 ( .A(n_461), .B(n_479), .Y(n_537) );
INVx2_ASAP7_75t_L g559 ( .A(n_461), .Y(n_559) );
OR2x2_ASAP7_75t_L g581 ( .A(n_461), .B(n_479), .Y(n_581) );
AND2x2_ASAP7_75t_L g586 ( .A(n_461), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_461), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g642 ( .A(n_461), .B(n_536), .Y(n_642) );
INVx1_ASAP7_75t_SL g693 ( .A(n_469), .Y(n_693) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_479), .Y(n_469) );
INVx1_ASAP7_75t_SL g536 ( .A(n_470), .Y(n_536) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_470), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_470), .B(n_622), .Y(n_621) );
NAND3xp33_ASAP7_75t_L g688 ( .A(n_470), .B(n_559), .C(n_677), .Y(n_688) );
OA21x2_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B(n_478), .Y(n_470) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_471), .A2(n_480), .B(n_486), .Y(n_479) );
OA21x2_ASAP7_75t_L g489 ( .A1(n_471), .A2(n_490), .B(n_496), .Y(n_489) );
INVx2_ASAP7_75t_L g587 ( .A(n_479), .Y(n_587) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_479), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_488), .B(n_497), .Y(n_487) );
INVx1_ASAP7_75t_L g623 ( .A(n_488), .Y(n_623) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g541 ( .A(n_489), .B(n_523), .Y(n_541) );
INVx2_ASAP7_75t_L g558 ( .A(n_489), .Y(n_558) );
AND2x2_ASAP7_75t_L g563 ( .A(n_489), .B(n_524), .Y(n_563) );
AND2x2_ASAP7_75t_L g578 ( .A(n_489), .B(n_511), .Y(n_578) );
AND2x2_ASAP7_75t_L g590 ( .A(n_489), .B(n_562), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_497), .B(n_606), .Y(n_605) );
NAND2x1p5_ASAP7_75t_L g662 ( .A(n_497), .B(n_563), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_497), .B(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_497), .B(n_557), .Y(n_685) );
BUFx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
OR2x2_ASAP7_75t_L g522 ( .A(n_498), .B(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_498), .B(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g567 ( .A(n_498), .B(n_511), .Y(n_567) );
AND2x2_ASAP7_75t_L g593 ( .A(n_498), .B(n_523), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_498), .B(n_633), .Y(n_632) );
OA21x2_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_500), .B(n_508), .Y(n_498) );
INVx1_ASAP7_75t_L g552 ( .A(n_500), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_504), .B(n_507), .Y(n_503) );
INVx2_ASAP7_75t_L g518 ( .A(n_507), .Y(n_518) );
INVx1_ASAP7_75t_L g553 ( .A(n_508), .Y(n_553) );
OR2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_522), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_511), .B(n_544), .Y(n_543) );
AND2x4_ASAP7_75t_L g557 ( .A(n_511), .B(n_558), .Y(n_557) );
INVx3_ASAP7_75t_SL g562 ( .A(n_511), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_511), .B(n_549), .Y(n_615) );
OR2x2_ASAP7_75t_L g625 ( .A(n_511), .B(n_551), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_511), .B(n_593), .Y(n_653) );
OR2x2_ASAP7_75t_L g683 ( .A(n_511), .B(n_523), .Y(n_683) );
AND2x2_ASAP7_75t_L g687 ( .A(n_511), .B(n_524), .Y(n_687) );
NAND2xp5_ASAP7_75t_SL g700 ( .A(n_511), .B(n_563), .Y(n_700) );
AND2x2_ASAP7_75t_L g707 ( .A(n_511), .B(n_589), .Y(n_707) );
OR2x6_ASAP7_75t_L g511 ( .A(n_512), .B(n_520), .Y(n_511) );
INVx1_ASAP7_75t_SL g650 ( .A(n_522), .Y(n_650) );
AND2x2_ASAP7_75t_L g589 ( .A(n_523), .B(n_551), .Y(n_589) );
AND2x2_ASAP7_75t_L g603 ( .A(n_523), .B(n_558), .Y(n_603) );
AND2x2_ASAP7_75t_L g606 ( .A(n_523), .B(n_562), .Y(n_606) );
INVx1_ASAP7_75t_L g633 ( .A(n_523), .Y(n_633) );
INVx2_ASAP7_75t_SL g523 ( .A(n_524), .Y(n_523) );
BUFx2_ASAP7_75t_L g545 ( .A(n_524), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_537), .Y(n_534) );
A2O1A1Ixp33_ASAP7_75t_L g704 ( .A1(n_535), .A2(n_581), .B(n_705), .C(n_706), .Y(n_704) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g611 ( .A(n_536), .B(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_537), .B(n_554), .Y(n_569) );
AND2x2_ASAP7_75t_L g595 ( .A(n_537), .B(n_596), .Y(n_595) );
OAI21xp5_ASAP7_75t_SL g538 ( .A1(n_539), .A2(n_542), .B(n_546), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_540), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g566 ( .A(n_541), .B(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_541), .B(n_562), .Y(n_607) );
AND2x2_ASAP7_75t_L g698 ( .A(n_541), .B(n_549), .Y(n_698) );
INVxp67_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g571 ( .A(n_545), .B(n_558), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_545), .B(n_556), .Y(n_572) );
OAI322xp33_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_555), .A3(n_556), .B1(n_559), .B2(n_560), .C1(n_564), .C2(n_565), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_554), .Y(n_548) );
AND2x2_ASAP7_75t_L g659 ( .A(n_549), .B(n_571), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_549), .B(n_623), .Y(n_705) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g602 ( .A(n_551), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OR2x2_ASAP7_75t_L g668 ( .A(n_555), .B(n_581), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_556), .B(n_650), .Y(n_649) );
INVx3_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_557), .B(n_589), .Y(n_646) );
AND2x2_ASAP7_75t_L g592 ( .A(n_558), .B(n_562), .Y(n_592) );
AND2x2_ASAP7_75t_L g600 ( .A(n_559), .B(n_601), .Y(n_600) );
A2O1A1Ixp33_ASAP7_75t_L g697 ( .A1(n_559), .A2(n_638), .B(n_698), .C(n_699), .Y(n_697) );
AOI21xp33_ASAP7_75t_L g670 ( .A1(n_560), .A2(n_573), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_562), .B(n_589), .Y(n_629) );
AND2x2_ASAP7_75t_L g635 ( .A(n_562), .B(n_603), .Y(n_635) );
AND2x2_ASAP7_75t_L g669 ( .A(n_562), .B(n_571), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_563), .B(n_578), .Y(n_577) );
INVx2_ASAP7_75t_SL g679 ( .A(n_563), .Y(n_679) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_567), .A2(n_595), .B1(n_597), .B2(n_602), .Y(n_594) );
OAI22xp5_ASAP7_75t_SL g568 ( .A1(n_569), .A2(n_570), .B1(n_572), .B2(n_573), .Y(n_568) );
OAI22xp33_ASAP7_75t_L g604 ( .A1(n_569), .A2(n_605), .B1(n_607), .B2(n_608), .Y(n_604) );
INVxp67_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
AOI221xp5_ASAP7_75t_L g675 ( .A1(n_574), .A2(n_676), .B1(n_678), .B2(n_680), .C(n_684), .Y(n_675) );
AOI211xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_579), .B(n_583), .C(n_604), .Y(n_575) );
INVxp67_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
OR2x2_ASAP7_75t_L g645 ( .A(n_581), .B(n_598), .Y(n_645) );
INVx1_ASAP7_75t_L g696 ( .A(n_581), .Y(n_696) );
OAI221xp5_ASAP7_75t_L g583 ( .A1(n_582), .A2(n_584), .B1(n_588), .B2(n_591), .C(n_594), .Y(n_583) );
INVx2_ASAP7_75t_SL g638 ( .A(n_582), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
INVx1_ASAP7_75t_L g703 ( .A(n_585), .Y(n_703) );
AND2x2_ASAP7_75t_L g627 ( .A(n_586), .B(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g612 ( .A(n_587), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
INVx1_ASAP7_75t_L g674 ( .A(n_590), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_598), .B(n_700), .Y(n_699) );
CKINVDCx16_ASAP7_75t_R g598 ( .A(n_599), .Y(n_598) );
INVxp67_ASAP7_75t_L g643 ( .A(n_601), .Y(n_643) );
O2A1O1Ixp33_ASAP7_75t_L g613 ( .A1(n_602), .A2(n_614), .B(n_616), .C(n_618), .Y(n_613) );
INVx1_ASAP7_75t_L g691 ( .A(n_605), .Y(n_691) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_609), .B(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx2_ASAP7_75t_L g622 ( .A(n_612), .Y(n_622) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OAI222xp33_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_625), .B1(n_626), .B2(n_629), .C1(n_630), .C2(n_632), .Y(n_618) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_SL g658 ( .A(n_622), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_625), .B(n_679), .Y(n_678) );
NAND2xp33_ASAP7_75t_SL g656 ( .A(n_626), .B(n_657), .Y(n_656) );
INVx1_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_SL g631 ( .A(n_628), .Y(n_631) );
AND2x2_ASAP7_75t_L g695 ( .A(n_628), .B(n_696), .Y(n_695) );
OR2x2_ASAP7_75t_L g661 ( .A(n_631), .B(n_658), .Y(n_661) );
INVx1_ASAP7_75t_L g690 ( .A(n_632), .Y(n_690) );
AOI211xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_636), .B(n_639), .C(n_644), .Y(n_634) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_638), .B(n_658), .Y(n_657) );
INVx2_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
AOI322xp5_ASAP7_75t_L g689 ( .A1(n_641), .A2(n_669), .A3(n_674), .B1(n_690), .B2(n_691), .C1(n_692), .C2(n_695), .Y(n_689) );
AND2x2_ASAP7_75t_L g676 ( .A(n_642), .B(n_677), .Y(n_676) );
OAI22xp33_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_646), .B1(n_647), .B2(n_649), .Y(n_644) );
INVxp33_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_654), .B1(n_656), .B2(n_659), .C(n_660), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
NAND5xp2_ASAP7_75t_L g663 ( .A(n_664), .B(n_675), .C(n_689), .D(n_697), .E(n_701), .Y(n_663) );
AOI21xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_669), .B(n_670), .Y(n_664) );
INVxp67_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVxp33_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
A2O1A1Ixp33_ASAP7_75t_L g701 ( .A1(n_677), .A2(n_702), .B(n_703), .C(n_704), .Y(n_701) );
AOI31xp33_ASAP7_75t_L g684 ( .A1(n_679), .A2(n_685), .A3(n_686), .B(n_688), .Y(n_684) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
INVx1_ASAP7_75t_L g702 ( .A(n_700), .Y(n_702) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g713 ( .A(n_708), .Y(n_713) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
endmodule