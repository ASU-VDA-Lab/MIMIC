module fake_netlist_6_885_n_4524 (n_52, n_1, n_91, n_326, n_256, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_396, n_350, n_78, n_84, n_392, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_421, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_141, n_383, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_413, n_377, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_397, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_414, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_9, n_107, n_6, n_417, n_14, n_89, n_374, n_366, n_407, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_395, n_323, n_393, n_411, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_406, n_102, n_204, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_422, n_135, n_165, n_351, n_259, n_177, n_391, n_364, n_295, n_385, n_388, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_4524);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_350;
input n_78;
input n_84;
input n_392;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_421;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_141;
input n_383;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_397;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_9;
input n_107;
input n_6;
input n_417;
input n_14;
input n_89;
input n_374;
input n_366;
input n_407;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_102;
input n_204;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_422;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_391;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_4524;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_3660;
wire n_3813;
wire n_801;
wire n_4452;
wire n_3766;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_3254;
wire n_3684;
wire n_1199;
wire n_1674;
wire n_3392;
wire n_741;
wire n_1027;
wire n_1351;
wire n_3266;
wire n_3574;
wire n_625;
wire n_1189;
wire n_3152;
wire n_4154;
wire n_3579;
wire n_1212;
wire n_4251;
wire n_726;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_4177;
wire n_3773;
wire n_700;
wire n_3783;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_3849;
wire n_4127;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_4504;
wire n_3844;
wire n_4395;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_3301;
wire n_4388;
wire n_4099;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_3741;
wire n_4517;
wire n_4168;
wire n_783;
wire n_4372;
wire n_2451;
wire n_1738;
wire n_4490;
wire n_2243;
wire n_798;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_3088;
wire n_3443;
wire n_1923;
wire n_3257;
wire n_509;
wire n_1342;
wire n_1348;
wire n_1209;
wire n_2260;
wire n_1387;
wire n_3222;
wire n_1708;
wire n_677;
wire n_805;
wire n_1151;
wire n_2977;
wire n_3952;
wire n_1739;
wire n_2051;
wire n_4370;
wire n_2317;
wire n_1380;
wire n_3911;
wire n_2359;
wire n_442;
wire n_2847;
wire n_480;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_4285;
wire n_3465;
wire n_1975;
wire n_1009;
wire n_1930;
wire n_1743;
wire n_2405;
wire n_3706;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_4092;
wire n_1724;
wire n_1032;
wire n_3708;
wire n_2336;
wire n_1247;
wire n_3668;
wire n_4078;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_3801;
wire n_4249;
wire n_1264;
wire n_1192;
wire n_471;
wire n_3564;
wire n_1844;
wire n_424;
wire n_3619;
wire n_4359;
wire n_4087;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_4302;
wire n_2291;
wire n_830;
wire n_2299;
wire n_3340;
wire n_4179;
wire n_873;
wire n_1371;
wire n_1285;
wire n_461;
wire n_2886;
wire n_2974;
wire n_3946;
wire n_1985;
wire n_4213;
wire n_2989;
wire n_447;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_4474;
wire n_852;
wire n_2509;
wire n_4065;
wire n_4026;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_3626;
wire n_3757;
wire n_3904;
wire n_4178;
wire n_1393;
wire n_1867;
wire n_1517;
wire n_2926;
wire n_1704;
wire n_2247;
wire n_544;
wire n_1711;
wire n_1078;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_4273;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_4446;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_4029;
wire n_836;
wire n_3345;
wire n_2074;
wire n_4417;
wire n_2447;
wire n_522;
wire n_2919;
wire n_4501;
wire n_3678;
wire n_3440;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_4010;
wire n_3879;
wire n_2286;
wire n_1649;
wire n_2094;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_4308;
wire n_616;
wire n_658;
wire n_1874;
wire n_4347;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_2739;
wire n_3023;
wire n_822;
wire n_3232;
wire n_693;
wire n_1313;
wire n_2791;
wire n_3607;
wire n_3750;
wire n_3251;
wire n_1056;
wire n_4325;
wire n_3316;
wire n_3877;
wire n_2212;
wire n_3929;
wire n_758;
wire n_516;
wire n_3494;
wire n_3063;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3048;
wire n_4311;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_1798;
wire n_943;
wire n_4060;
wire n_1550;
wire n_2703;
wire n_491;
wire n_3998;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_772;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_666;
wire n_4187;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2090;
wire n_2058;
wire n_2603;
wire n_2660;
wire n_3028;
wire n_538;
wire n_3829;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_4164;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_3737;
wire n_3624;
wire n_3077;
wire n_3979;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3655;
wire n_3452;
wire n_494;
wire n_539;
wire n_493;
wire n_3107;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_4117;
wire n_454;
wire n_3948;
wire n_1421;
wire n_2836;
wire n_3664;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_4327;
wire n_1961;
wire n_3047;
wire n_4414;
wire n_1280;
wire n_3765;
wire n_713;
wire n_2655;
wire n_4125;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_4221;
wire n_1467;
wire n_3297;
wire n_4250;
wire n_976;
wire n_3760;
wire n_3067;
wire n_2155;
wire n_3906;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_4262;
wire n_4392;
wire n_1894;
wire n_2996;
wire n_1231;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_3803;
wire n_2085;
wire n_3963;
wire n_3368;
wire n_917;
wire n_574;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_3792;
wire n_907;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_2591;
wire n_3507;
wire n_4334;
wire n_659;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_4253;
wire n_913;
wire n_4110;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_4071;
wire n_4255;
wire n_4403;
wire n_3506;
wire n_4268;
wire n_3568;
wire n_3269;
wire n_4047;
wire n_3531;
wire n_1230;
wire n_3413;
wire n_3850;
wire n_473;
wire n_1193;
wire n_1967;
wire n_3999;
wire n_1054;
wire n_3928;
wire n_559;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_3791;
wire n_4139;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_3943;
wire n_4320;
wire n_4305;
wire n_564;
wire n_2397;
wire n_3931;
wire n_3884;
wire n_4349;
wire n_451;
wire n_824;
wire n_686;
wire n_4102;
wire n_4297;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_3603;
wire n_3871;
wire n_2907;
wire n_577;
wire n_3438;
wire n_2735;
wire n_4141;
wire n_1843;
wire n_619;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_2778;
wire n_4227;
wire n_2850;
wire n_572;
wire n_4314;
wire n_1909;
wire n_2080;
wire n_813;
wire n_1481;
wire n_3822;
wire n_4163;
wire n_1441;
wire n_606;
wire n_818;
wire n_3373;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_2961;
wire n_3910;
wire n_1699;
wire n_3812;
wire n_916;
wire n_3934;
wire n_2093;
wire n_4033;
wire n_4415;
wire n_4296;
wire n_4009;
wire n_2633;
wire n_483;
wire n_3883;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_608;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_630;
wire n_2059;
wire n_4507;
wire n_2198;
wire n_3319;
wire n_541;
wire n_512;
wire n_2669;
wire n_2925;
wire n_3728;
wire n_4094;
wire n_4499;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_433;
wire n_3748;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_792;
wire n_2522;
wire n_476;
wire n_3949;
wire n_4364;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_4354;
wire n_2616;
wire n_3912;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_3923;
wire n_2529;
wire n_3900;
wire n_4393;
wire n_1162;
wire n_860;
wire n_1530;
wire n_3798;
wire n_788;
wire n_939;
wire n_3488;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_3732;
wire n_982;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_2832;
wire n_4226;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_932;
wire n_2831;
wire n_2998;
wire n_4318;
wire n_4366;
wire n_3446;
wire n_4158;
wire n_4377;
wire n_3317;
wire n_3857;
wire n_3978;
wire n_1876;
wire n_4107;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_4074;
wire n_3716;
wire n_1873;
wire n_4294;
wire n_905;
wire n_3630;
wire n_3518;
wire n_4445;
wire n_3824;
wire n_3859;
wire n_1866;
wire n_4013;
wire n_1680;
wire n_2692;
wire n_993;
wire n_3842;
wire n_689;
wire n_3248;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_3714;
wire n_3514;
wire n_2228;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_547;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_558;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_4032;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_634;
wire n_2355;
wire n_3927;
wire n_4147;
wire n_4477;
wire n_966;
wire n_3888;
wire n_4511;
wire n_2908;
wire n_3168;
wire n_764;
wire n_4468;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_4130;
wire n_4337;
wire n_4161;
wire n_2895;
wire n_2009;
wire n_4172;
wire n_692;
wire n_3403;
wire n_733;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_3882;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_487;
wire n_3092;
wire n_3055;
wire n_3492;
wire n_3895;
wire n_3966;
wire n_4369;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_4454;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_1014;
wire n_3734;
wire n_4331;
wire n_3686;
wire n_4520;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_4118;
wire n_4502;
wire n_882;
wire n_4503;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_1354;
wire n_2821;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_2459;
wire n_3746;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_4375;
wire n_715;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_3935;
wire n_1265;
wire n_4277;
wire n_2711;
wire n_3490;
wire n_4291;
wire n_4199;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1912;
wire n_1563;
wire n_2434;
wire n_4319;
wire n_3369;
wire n_3419;
wire n_4441;
wire n_1982;
wire n_3872;
wire n_2878;
wire n_618;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_3772;
wire n_3875;
wire n_4478;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3581;
wire n_3794;
wire n_674;
wire n_3247;
wire n_871;
wire n_3069;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_2641;
wire n_612;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_1165;
wire n_3933;
wire n_702;
wire n_2008;
wire n_2749;
wire n_3298;
wire n_2192;
wire n_3281;
wire n_2254;
wire n_2345;
wire n_3346;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_4467;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_3691;
wire n_4427;
wire n_780;
wire n_3861;
wire n_675;
wire n_2624;
wire n_4066;
wire n_903;
wire n_4386;
wire n_4485;
wire n_4146;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_4340;
wire n_3891;
wire n_2193;
wire n_3961;
wire n_2676;
wire n_1655;
wire n_3940;
wire n_4072;
wire n_4220;
wire n_4523;
wire n_835;
wire n_1214;
wire n_1801;
wire n_690;
wire n_850;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_928;
wire n_1654;
wire n_816;
wire n_4371;
wire n_1157;
wire n_3453;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3428;
wire n_3153;
wire n_3410;
wire n_1188;
wire n_3689;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_3768;
wire n_2206;
wire n_604;
wire n_4004;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_4043;
wire n_825;
wire n_728;
wire n_4353;
wire n_2916;
wire n_3415;
wire n_1063;
wire n_4292;
wire n_1588;
wire n_3785;
wire n_3942;
wire n_3997;
wire n_2963;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_4381;
wire n_1124;
wire n_1624;
wire n_3873;
wire n_3983;
wire n_515;
wire n_2096;
wire n_2980;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_598;
wire n_3434;
wire n_4510;
wire n_696;
wire n_1515;
wire n_4473;
wire n_961;
wire n_4356;
wire n_3510;
wire n_437;
wire n_1317;
wire n_1082;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_593;
wire n_4169;
wire n_514;
wire n_4055;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_3271;
wire n_950;
wire n_4248;
wire n_2812;
wire n_4518;
wire n_484;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_4361;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_3827;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_3889;
wire n_2687;
wire n_3237;
wire n_949;
wire n_1630;
wire n_678;
wire n_2887;
wire n_3809;
wire n_3500;
wire n_3834;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_3707;
wire n_2075;
wire n_4045;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_4367;
wire n_2763;
wire n_2762;
wire n_4070;
wire n_1987;
wire n_3545;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_3578;
wire n_3885;
wire n_881;
wire n_2271;
wire n_1008;
wire n_3192;
wire n_760;
wire n_3993;
wire n_1546;
wire n_2583;
wire n_590;
wire n_4394;
wire n_4116;
wire n_2606;
wire n_4031;
wire n_2279;
wire n_462;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_3805;
wire n_2431;
wire n_3073;
wire n_4018;
wire n_2987;
wire n_694;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_3696;
wire n_3780;
wire n_4082;
wire n_1634;
wire n_2078;
wire n_3252;
wire n_2932;
wire n_595;
wire n_1767;
wire n_627;
wire n_1779;
wire n_524;
wire n_1465;
wire n_3253;
wire n_3337;
wire n_3450;
wire n_3209;
wire n_4002;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_4329;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_449;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_2893;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2954;
wire n_3477;
wire n_4289;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_3763;
wire n_4288;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_495;
wire n_815;
wire n_3953;
wire n_1100;
wire n_585;
wire n_1487;
wire n_4435;
wire n_2691;
wire n_3421;
wire n_840;
wire n_2913;
wire n_3614;
wire n_874;
wire n_4471;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_2230;
wire n_2705;
wire n_673;
wire n_1969;
wire n_4019;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_898;
wire n_4385;
wire n_1952;
wire n_865;
wire n_3616;
wire n_4228;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_4044;
wire n_3436;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_3366;
wire n_3442;
wire n_2631;
wire n_4191;
wire n_1364;
wire n_4322;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_3937;
wire n_2870;
wire n_615;
wire n_1249;
wire n_2706;
wire n_3838;
wire n_4287;
wire n_1293;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_3941;
wire n_963;
wire n_639;
wire n_2767;
wire n_794;
wire n_3793;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_3789;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_3385;
wire n_4350;
wire n_3747;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_872;
wire n_1714;
wire n_1139;
wire n_3922;
wire n_3179;
wire n_718;
wire n_1018;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_4330;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_2537;
wire n_2897;
wire n_3970;
wire n_4389;
wire n_4483;
wire n_4345;
wire n_2554;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_1513;
wire n_2747;
wire n_3924;
wire n_3171;
wire n_791;
wire n_1913;
wire n_4216;
wire n_3608;
wire n_510;
wire n_837;
wire n_4315;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_4156;
wire n_3491;
wire n_4240;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_704;
wire n_2148;
wire n_4284;
wire n_4162;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_536;
wire n_3158;
wire n_1788;
wire n_3426;
wire n_1999;
wire n_2731;
wire n_622;
wire n_2643;
wire n_2590;
wire n_3150;
wire n_3018;
wire n_3353;
wire n_3782;
wire n_3975;
wire n_1469;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_4011;
wire n_1835;
wire n_3470;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_581;
wire n_2650;
wire n_2138;
wire n_4098;
wire n_4021;
wire n_4476;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_3700;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_4058;
wire n_4103;
wire n_3104;
wire n_631;
wire n_720;
wire n_3435;
wire n_842;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_3348;
wire n_4022;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_3611;
wire n_4310;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_4481;
wire n_1246;
wire n_3799;
wire n_1878;
wire n_2574;
wire n_4475;
wire n_899;
wire n_2012;
wire n_738;
wire n_3497;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_499;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_705;
wire n_3580;
wire n_3775;
wire n_3537;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_4443;
wire n_3887;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_3704;
wire n_2362;
wire n_425;
wire n_684;
wire n_2539;
wire n_2698;
wire n_2667;
wire n_4123;
wire n_1431;
wire n_4096;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_3835;
wire n_4286;
wire n_1809;
wire n_3119;
wire n_4280;
wire n_2958;
wire n_1577;
wire n_2948;
wire n_3735;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_4379;
wire n_3731;
wire n_1822;
wire n_486;
wire n_947;
wire n_2936;
wire n_3224;
wire n_1117;
wire n_2489;
wire n_1448;
wire n_1087;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_648;
wire n_657;
wire n_1049;
wire n_3223;
wire n_3996;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_3770;
wire n_2605;
wire n_4097;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_4218;
wire n_4440;
wire n_4402;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_3557;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_3880;
wire n_1849;
wire n_2848;
wire n_919;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_478;
wire n_4100;
wire n_2231;
wire n_3609;
wire n_929;
wire n_3832;
wire n_2520;
wire n_1228;
wire n_4264;
wire n_4484;
wire n_2857;
wire n_446;
wire n_3693;
wire n_4497;
wire n_3788;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_4459;
wire n_1299;
wire n_2896;
wire n_526;
wire n_3837;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_3674;
wire n_2494;
wire n_2959;
wire n_4079;
wire n_2501;
wire n_3203;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_2368;
wire n_4464;
wire n_458;
wire n_1070;
wire n_2403;
wire n_3342;
wire n_2837;
wire n_4175;
wire n_998;
wire n_717;
wire n_3200;
wire n_1665;
wire n_4306;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_4224;
wire n_3390;
wire n_3656;
wire n_4339;
wire n_1178;
wire n_2338;
wire n_1424;
wire n_2127;
wire n_3324;
wire n_3593;
wire n_3341;
wire n_3867;
wire n_4455;
wire n_4453;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_3559;
wire n_4514;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_4005;
wire n_1507;
wire n_2482;
wire n_3810;
wire n_552;
wire n_3546;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3661;
wire n_3006;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_912;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_3201;
wire n_3633;
wire n_3447;
wire n_4487;
wire n_3971;
wire n_1142;
wire n_2849;
wire n_716;
wire n_1475;
wire n_1774;
wire n_1048;
wire n_1398;
wire n_1201;
wire n_884;
wire n_2354;
wire n_2682;
wire n_623;
wire n_3032;
wire n_3103;
wire n_3638;
wire n_2589;
wire n_1395;
wire n_2199;
wire n_2110;
wire n_2661;
wire n_731;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_3393;
wire n_527;
wire n_811;
wire n_474;
wire n_1207;
wire n_2442;
wire n_683;
wire n_3627;
wire n_1791;
wire n_1368;
wire n_3451;
wire n_3480;
wire n_1418;
wire n_958;
wire n_1250;
wire n_3331;
wire n_1137;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_880;
wire n_3087;
wire n_3072;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_4222;
wire n_2545;
wire n_3540;
wire n_3577;
wire n_4401;
wire n_889;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_4368;
wire n_1478;
wire n_589;
wire n_3606;
wire n_1310;
wire n_3142;
wire n_3598;
wire n_819;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_3591;
wire n_767;
wire n_3641;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_2218;
wire n_1837;
wire n_2788;
wire n_477;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_954;
wire n_4419;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_4120;
wire n_1382;
wire n_1534;
wire n_3892;
wire n_1564;
wire n_1736;
wire n_4069;
wire n_2748;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2860;
wire n_2292;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_505;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_537;
wire n_2511;
wire n_3964;
wire n_1993;
wire n_2281;
wire n_4167;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_596;
wire n_3944;
wire n_3909;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2784;
wire n_2301;
wire n_2209;
wire n_3582;
wire n_3605;
wire n_3287;
wire n_4223;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_4431;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_4387;
wire n_2618;
wire n_2357;
wire n_2025;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_970;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_3481;
wire n_2237;
wire n_3026;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_4299;
wire n_444;
wire n_3033;
wire n_3724;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_3571;
wire n_1223;
wire n_3913;
wire n_4276;
wire n_4362;
wire n_511;
wire n_2990;
wire n_3847;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_4430;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_4348;
wire n_520;
wire n_1093;
wire n_4428;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3364;
wire n_3226;
wire n_3323;
wire n_4020;
wire n_4176;
wire n_4489;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_775;
wire n_4404;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_3407;
wire n_518;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_3856;
wire n_453;
wire n_4236;
wire n_3425;
wire n_2384;
wire n_3894;
wire n_4204;
wire n_4261;
wire n_1745;
wire n_914;
wire n_759;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_426;
wire n_4496;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_4063;
wire n_1625;
wire n_3986;
wire n_4237;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_4513;
wire n_1453;
wire n_2146;
wire n_4006;
wire n_2226;
wire n_2131;
wire n_488;
wire n_2502;
wire n_2801;
wire n_3646;
wire n_497;
wire n_2920;
wire n_4015;
wire n_773;
wire n_3547;
wire n_1901;
wire n_3869;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_3188;
wire n_3742;
wire n_4410;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_2889;
wire n_3243;
wire n_3683;
wire n_4034;
wire n_1617;
wire n_4056;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_3816;
wire n_3960;
wire n_1470;
wire n_2550;
wire n_463;
wire n_3093;
wire n_3175;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_3736;
wire n_848;
wire n_2732;
wire n_2928;
wire n_4206;
wire n_4448;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_3862;
wire n_4267;
wire n_1580;
wire n_2227;
wire n_4247;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_4180;
wire n_3284;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_3205;
wire n_983;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_427;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1733;
wire n_2315;
wire n_1077;
wire n_1419;
wire n_2863;
wire n_3299;
wire n_3663;
wire n_4132;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_3360;
wire n_4438;
wire n_2135;
wire n_3956;
wire n_3367;
wire n_1645;
wire n_1832;
wire n_4001;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_858;
wire n_2049;
wire n_4149;
wire n_1331;
wire n_613;
wire n_736;
wire n_2627;
wire n_4355;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_3234;
wire n_4422;
wire n_3917;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_2993;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_3016;
wire n_3566;
wire n_3688;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_4003;
wire n_1129;
wire n_3870;
wire n_4030;
wire n_4126;
wire n_554;
wire n_602;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_2181;
wire n_1594;
wire n_3845;
wire n_1869;
wire n_664;
wire n_2911;
wire n_3625;
wire n_3751;
wire n_3804;
wire n_1764;
wire n_4207;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_4113;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_4470;
wire n_587;
wire n_3466;
wire n_3554;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_3901;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_1635;
wire n_2942;
wire n_4014;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_4067;
wire n_4252;
wire n_4357;
wire n_607;
wire n_1551;
wire n_4028;
wire n_4054;
wire n_4509;
wire n_2448;
wire n_2875;
wire n_1103;
wire n_3907;
wire n_2555;
wire n_4048;
wire n_4444;
wire n_3338;
wire n_4217;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_1203;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_820;
wire n_2327;
wire n_951;
wire n_4374;
wire n_2201;
wire n_725;
wire n_952;
wire n_3919;
wire n_999;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_2984;
wire n_575;
wire n_994;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_4024;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_3194;
wire n_3276;
wire n_1934;
wire n_3250;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_4214;
wire n_1728;
wire n_3973;
wire n_557;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_4338;
wire n_617;
wire n_3886;
wire n_845;
wire n_807;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_485;
wire n_1549;
wire n_4420;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_3637;
wire n_3120;
wire n_1468;
wire n_3991;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_3797;
wire n_3926;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_4405;
wire n_610;
wire n_4304;
wire n_4234;
wire n_4413;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_4488;
wire n_4101;
wire n_3548;
wire n_3767;
wire n_1024;
wire n_3864;
wire n_4036;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_3974;
wire n_2052;
wire n_1847;
wire n_3634;
wire n_2302;
wire n_517;
wire n_4211;
wire n_4182;
wire n_1667;
wire n_667;
wire n_1206;
wire n_3230;
wire n_4016;
wire n_621;
wire n_1037;
wire n_1397;
wire n_3268;
wire n_3236;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_3592;
wire n_468;
wire n_2755;
wire n_3141;
wire n_923;
wire n_504;
wire n_1409;
wire n_4230;
wire n_1841;
wire n_3839;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_3967;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_4328;
wire n_3195;
wire n_466;
wire n_2526;
wire n_3041;
wire n_4274;
wire n_2423;
wire n_1057;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_603;
wire n_991;
wire n_2785;
wire n_1657;
wire n_4270;
wire n_4189;
wire n_4151;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_3817;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_2439;
wire n_710;
wire n_1818;
wire n_1108;
wire n_3730;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_4124;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_3399;
wire n_4397;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_785;
wire n_4155;
wire n_2740;
wire n_746;
wire n_4238;
wire n_609;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2401;
wire n_2337;
wire n_3042;
wire n_1356;
wire n_1589;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_4472;
wire n_1216;
wire n_1943;
wire n_3228;
wire n_1320;
wire n_2716;
wire n_3249;
wire n_3081;
wire n_3657;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3672;
wire n_3010;
wire n_2499;
wire n_4152;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_3382;
wire n_4406;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_4380;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_4398;
wire n_2498;
wire n_4219;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3238;
wire n_2235;
wire n_3529;
wire n_4193;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_3828;
wire n_2232;
wire n_1715;
wire n_3536;
wire n_4109;
wire n_4192;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_3424;
wire n_3957;
wire n_4038;
wire n_2790;
wire n_4131;
wire n_2037;
wire n_2808;
wire n_3710;
wire n_4159;
wire n_4195;
wire n_3784;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_3594;
wire n_809;
wire n_1043;
wire n_3819;
wire n_4090;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_4165;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_3628;
wire n_4144;
wire n_1870;
wire n_2964;
wire n_4174;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3475;
wire n_662;
wire n_3501;
wire n_4442;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_3905;
wire n_4434;
wire n_450;
wire n_3262;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_4008;
wire n_2244;
wire n_4290;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_937;
wire n_2257;
wire n_3692;
wire n_4515;
wire n_1682;
wire n_2017;
wire n_4516;
wire n_4258;
wire n_1695;
wire n_1828;
wire n_2699;
wire n_2272;
wire n_2046;
wire n_2200;
wire n_3029;
wire n_650;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_3826;
wire n_1406;
wire n_456;
wire n_3790;
wire n_3878;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_4323;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_3134;
wire n_3647;
wire n_1569;
wire n_3681;
wire n_936;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_3821;
wire n_1288;
wire n_4300;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_3676;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_4017;
wire n_4260;
wire n_3320;
wire n_2541;
wire n_654;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_1974;
wire n_3988;
wire n_4122;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_482;
wire n_934;
wire n_1637;
wire n_2635;
wire n_3439;
wire n_3307;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_3588;
wire n_4135;
wire n_2871;
wire n_4209;
wire n_4279;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_3858;
wire n_4183;
wire n_1489;
wire n_4321;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_4128;
wire n_543;
wire n_2229;
wire n_1964;
wire n_4133;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_4145;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_4271;
wire n_1946;
wire n_1355;
wire n_4181;
wire n_1225;
wire n_3184;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_4040;
wire n_804;
wire n_4461;
wire n_1846;
wire n_464;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_4111;
wire n_533;
wire n_2390;
wire n_4007;
wire n_806;
wire n_3712;
wire n_879;
wire n_959;
wire n_2310;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_4239;
wire n_2734;
wire n_548;
wire n_1782;
wire n_2383;
wire n_4184;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_4037;
wire n_523;
wire n_1319;
wire n_707;
wire n_2986;
wire n_1900;
wire n_3930;
wire n_3246;
wire n_799;
wire n_1548;
wire n_3381;
wire n_3044;
wire n_3562;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_3915;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_787;
wire n_2172;
wire n_3528;
wire n_3489;
wire n_4343;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_4215;
wire n_1282;
wire n_2561;
wire n_550;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2962;
wire n_2727;
wire n_2154;
wire n_652;
wire n_3377;
wire n_2939;
wire n_560;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_2533;
wire n_3157;
wire n_3530;
wire n_4185;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_3752;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_4378;
wire n_4407;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_3457;
wire n_1229;
wire n_2759;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_3893;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_3762;
wire n_3932;
wire n_3469;
wire n_3958;
wire n_2266;
wire n_2960;
wire n_3005;
wire n_3985;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_1029;
wire n_4196;
wire n_3779;
wire n_1447;
wire n_4519;
wire n_2388;
wire n_3984;
wire n_2056;
wire n_790;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_4358;
wire n_1706;
wire n_4242;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_4232;
wire n_4190;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_4052;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_3375;
wire n_3899;
wire n_4084;
wire n_3558;
wire n_4469;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3713;
wire n_431;
wire n_3379;
wire n_4326;
wire n_3156;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_502;
wire n_2668;
wire n_672;
wire n_4424;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_3939;
wire n_1941;
wire n_1375;
wire n_3613;
wire n_3483;
wire n_3972;
wire n_4153;
wire n_2128;
wire n_655;
wire n_706;
wire n_1650;
wire n_1045;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_2398;
wire n_1725;
wire n_1928;
wire n_1559;
wire n_3743;
wire n_3855;
wire n_1872;
wire n_3091;
wire n_4317;
wire n_834;
wire n_4493;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_4269;
wire n_743;
wire n_766;
wire n_3124;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_4088;
wire n_1949;
wire n_3398;
wire n_3761;
wire n_3759;
wire n_545;
wire n_3524;
wire n_2671;
wire n_489;
wire n_2761;
wire n_2885;
wire n_2793;
wire n_2715;
wire n_2923;
wire n_1804;
wire n_2888;
wire n_3711;
wire n_3776;
wire n_4235;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_4301;
wire n_3511;
wire n_2054;
wire n_4143;
wire n_4170;
wire n_729;
wire n_876;
wire n_774;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_2062;
wire n_660;
wire n_2041;
wire n_2975;
wire n_438;
wire n_1477;
wire n_4421;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_4498;
wire n_2070;
wire n_2588;
wire n_479;
wire n_3814;
wire n_1607;
wire n_3781;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_3831;
wire n_869;
wire n_1154;
wire n_4492;
wire n_3308;
wire n_1113;
wire n_1600;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_3843;
wire n_2366;
wire n_646;
wire n_528;
wire n_1098;
wire n_3694;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_4423;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_3602;
wire n_897;
wire n_846;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_841;
wire n_1476;
wire n_3621;
wire n_2516;
wire n_3391;
wire n_4376;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_3777;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_3458;
wire n_4203;
wire n_3515;
wire n_1150;
wire n_4505;
wire n_3808;
wire n_3190;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_4365;
wire n_1826;
wire n_566;
wire n_1882;
wire n_1023;
wire n_2951;
wire n_1118;
wire n_1076;
wire n_4512;
wire n_2949;
wire n_3726;
wire n_1807;
wire n_1007;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_591;
wire n_3758;
wire n_1879;
wire n_853;
wire n_440;
wire n_695;
wire n_3806;
wire n_4081;
wire n_1542;
wire n_2587;
wire n_3199;
wire n_2931;
wire n_875;
wire n_680;
wire n_4462;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_3866;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_671;
wire n_3565;
wire n_1953;
wire n_4450;
wire n_933;
wire n_740;
wire n_703;
wire n_3343;
wire n_3303;
wire n_978;
wire n_4157;
wire n_2752;
wire n_4173;
wire n_3135;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_4229;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_3990;
wire n_751;
wire n_749;
wire n_3865;
wire n_1824;
wire n_3954;
wire n_1628;
wire n_4073;
wire n_1324;
wire n_3890;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_969;
wire n_988;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_3658;
wire n_1516;
wire n_1536;
wire n_3846;
wire n_2186;
wire n_2163;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3951;
wire n_3034;
wire n_823;
wire n_4408;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_4439;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_955;
wire n_739;
wire n_3874;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2969;
wire n_2395;
wire n_935;
wire n_3027;
wire n_781;
wire n_789;
wire n_1554;
wire n_3231;
wire n_4083;
wire n_4494;
wire n_1130;
wire n_3083;
wire n_4212;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_4295;
wire n_1120;
wire n_832;
wire n_1583;
wire n_4480;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_4225;
wire n_4171;
wire n_2048;
wire n_3652;
wire n_3830;
wire n_3679;
wire n_2005;
wire n_747;
wire n_3541;
wire n_2565;
wire n_4023;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_721;
wire n_1461;
wire n_742;
wire n_3432;
wire n_535;
wire n_691;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_3583;
wire n_3860;
wire n_1408;
wire n_3851;
wire n_3567;
wire n_1196;
wire n_4282;
wire n_1598;
wire n_3493;
wire n_4344;
wire n_2935;
wire n_4046;
wire n_3807;
wire n_863;
wire n_3015;
wire n_2175;
wire n_601;
wire n_2182;
wire n_3774;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_918;
wire n_748;
wire n_506;
wire n_1785;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1114;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3701;
wire n_3154;
wire n_4027;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_3473;
wire n_895;
wire n_866;
wire n_1227;
wire n_2485;
wire n_2450;
wire n_3739;
wire n_2284;
wire n_3898;
wire n_4432;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_452;
wire n_4352;
wire n_744;
wire n_971;
wire n_4391;
wire n_4416;
wire n_2702;
wire n_3241;
wire n_946;
wire n_2906;
wire n_761;
wire n_1303;
wire n_2769;
wire n_4342;
wire n_4465;
wire n_3622;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_3778;
wire n_4095;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_4495;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_611;
wire n_1219;
wire n_3551;
wire n_4436;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3897;
wire n_3721;
wire n_1689;
wire n_2180;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_3573;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_4106;
wire n_795;
wire n_1501;
wire n_3604;
wire n_1221;
wire n_3334;
wire n_4373;
wire n_1245;
wire n_838;
wire n_3215;
wire n_3969;
wire n_3336;
wire n_647;
wire n_4160;
wire n_4231;
wire n_844;
wire n_448;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_3853;
wire n_2117;
wire n_2234;
wire n_4256;
wire n_2779;
wire n_2685;
wire n_3823;
wire n_1083;
wire n_445;
wire n_3553;
wire n_1561;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_3811;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_653;
wire n_2430;
wire n_3486;
wire n_1414;
wire n_3584;
wire n_4086;
wire n_752;
wire n_908;
wire n_2721;
wire n_2649;
wire n_944;
wire n_4335;
wire n_3556;
wire n_2034;
wire n_576;
wire n_1028;
wire n_3836;
wire n_2106;
wire n_472;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_563;
wire n_4068;
wire n_2032;
wire n_4409;
wire n_2744;
wire n_4309;
wire n_4363;
wire n_1011;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_4521;
wire n_2444;
wire n_2437;
wire n_1215;
wire n_839;
wire n_2743;
wire n_3962;
wire n_708;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_668;
wire n_4166;
wire n_626;
wire n_990;
wire n_1821;
wire n_779;
wire n_1537;
wire n_1500;
wire n_2205;
wire n_3699;
wire n_4243;
wire n_3204;
wire n_1104;
wire n_854;
wire n_1058;
wire n_3378;
wire n_4025;
wire n_2312;
wire n_498;
wire n_3404;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_3362;
wire n_3745;
wire n_4059;
wire n_1509;
wire n_4188;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_4121;
wire n_1109;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3256;
wire n_1276;
wire n_3802;
wire n_3868;
wire n_3176;
wire n_3309;
wire n_3671;
wire n_4142;
wire n_2015;
wire n_2118;
wire n_4313;
wire n_2111;
wire n_2466;
wire n_3982;
wire n_4266;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2505;
wire n_2188;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_3796;
wire n_2999;
wire n_4115;
wire n_3840;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_3643;
wire n_3697;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_3461;
wire n_3408;
wire n_1582;
wire n_492;
wire n_3680;
wire n_4265;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_2408;
wire n_4246;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_3690;
wire n_1184;
wire n_3645;
wire n_2483;
wire n_2950;
wire n_719;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_3771;
wire n_1525;
wire n_4383;
wire n_4491;
wire n_3098;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_455;
wire n_2666;
wire n_4105;
wire n_1851;
wire n_1585;
wire n_1799;
wire n_1090;
wire n_2564;
wire n_2147;
wire n_592;
wire n_4244;
wire n_4486;
wire n_1816;
wire n_4064;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_4049;
wire n_829;
wire n_1362;
wire n_1156;
wire n_4259;
wire n_3123;
wire n_984;
wire n_2600;
wire n_3380;
wire n_1829;
wire n_503;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_868;
wire n_3038;
wire n_570;
wire n_859;
wire n_2033;
wire n_3086;
wire n_735;
wire n_4104;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_3285;
wire n_519;
wire n_4208;
wire n_2523;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_3769;
wire n_1482;
wire n_3361;
wire n_981;
wire n_3596;
wire n_714;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_4089;
wire n_4346;
wire n_4351;
wire n_1144;
wire n_2071;
wire n_3669;
wire n_3863;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_985;
wire n_4316;
wire n_2723;
wire n_2440;
wire n_2233;
wire n_481;
wire n_3521;
wire n_3233;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_3496;
wire n_4437;
wire n_1301;
wire n_2805;
wire n_802;
wire n_561;
wire n_3310;
wire n_980;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_4390;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_3764;
wire n_2047;
wire n_4061;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_436;
wire n_4075;
wire n_3344;
wire n_2334;
wire n_3902;
wire n_4062;
wire n_3881;
wire n_3295;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_4396;
wire n_4508;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_3989;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_4233;
wire n_4451;
wire n_1606;
wire n_4332;
wire n_810;
wire n_4108;
wire n_1133;
wire n_4460;
wire n_635;
wire n_1194;
wire n_3374;
wire n_4429;
wire n_4506;
wire n_3786;
wire n_3841;
wire n_2742;
wire n_2640;
wire n_3695;
wire n_4254;
wire n_1051;
wire n_3976;
wire n_4051;
wire n_1552;
wire n_2918;
wire n_583;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_3992;
wire n_2367;
wire n_4307;
wire n_3876;
wire n_2867;
wire n_3198;
wire n_1039;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_4303;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_754;
wire n_4293;
wire n_941;
wire n_3552;
wire n_975;
wire n_3206;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_553;
wire n_849;
wire n_2662;
wire n_3116;
wire n_3147;
wire n_3383;
wire n_3709;
wire n_753;
wire n_3925;
wire n_4091;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_4186;
wire n_467;
wire n_3187;
wire n_2540;
wire n_4412;
wire n_973;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_3330;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_2879;
wire n_861;
wire n_3717;
wire n_857;
wire n_967;
wire n_4522;
wire n_4148;
wire n_571;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_4341;
wire n_1884;
wire n_2040;
wire n_679;
wire n_4057;
wire n_2968;
wire n_4336;
wire n_4201;
wire n_633;
wire n_1170;
wire n_1629;
wire n_2221;
wire n_665;
wire n_588;
wire n_4263;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_3555;
wire n_1010;
wire n_3444;
wire n_4210;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_4447;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_3955;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_2280;
wire n_1557;
wire n_1833;
wire n_3945;
wire n_730;
wire n_1311;
wire n_3903;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_3854;
wire n_2308;
wire n_4205;
wire n_2162;
wire n_3908;
wire n_2333;
wire n_1868;
wire n_2079;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1089;
wire n_4278;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_3795;
wire n_2512;
wire n_3950;
wire n_3433;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_4463;
wire n_1417;
wire n_1242;
wire n_2185;
wire n_2086;
wire n_2927;
wire n_3673;
wire n_1836;
wire n_3833;
wire n_4281;
wire n_3896;
wire n_2774;
wire n_3815;
wire n_3039;
wire n_681;
wire n_1226;
wire n_3740;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3274;
wire n_3333;
wire n_3186;
wire n_640;
wire n_1322;
wire n_4129;
wire n_4457;
wire n_965;
wire n_1899;
wire n_1428;
wire n_4093;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_3965;
wire n_2632;
wire n_2579;
wire n_722;
wire n_4500;
wire n_862;
wire n_2105;
wire n_3079;
wire n_4360;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_540;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_4039;
wire n_3387;
wire n_2027;
wire n_457;
wire n_3070;
wire n_3800;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_3431;
wire n_4197;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_629;
wire n_1621;
wire n_4275;
wire n_4482;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_4283;
wire n_900;
wire n_3504;
wire n_4194;
wire n_1449;
wire n_4426;
wire n_531;
wire n_827;
wire n_2912;
wire n_4272;
wire n_2659;
wire n_2930;
wire n_4425;
wire n_1025;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_4449;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_1742;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_L g423 ( 
.A(n_26),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_391),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_44),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_122),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_52),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_352),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_178),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_26),
.Y(n_430)
);

BUFx10_ASAP7_75t_L g431 ( 
.A(n_155),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_255),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_398),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_299),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_70),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_72),
.Y(n_436)
);

BUFx5_ASAP7_75t_L g437 ( 
.A(n_42),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_316),
.Y(n_438)
);

CKINVDCx14_ASAP7_75t_R g439 ( 
.A(n_329),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_253),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_102),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_60),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_266),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_146),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_406),
.Y(n_445)
);

CKINVDCx14_ASAP7_75t_R g446 ( 
.A(n_293),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_142),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_371),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_146),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_222),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_104),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_229),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_181),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_415),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_5),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_411),
.Y(n_456)
);

BUFx10_ASAP7_75t_L g457 ( 
.A(n_159),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_418),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_127),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_364),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_251),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_283),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_65),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_389),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g465 ( 
.A(n_359),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_35),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_126),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_30),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_281),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_66),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_388),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_349),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_176),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_209),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_416),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_137),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_133),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_35),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_422),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_308),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_404),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_130),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_387),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_381),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_63),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_210),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_161),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_386),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_86),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_242),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_323),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_152),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_394),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_333),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_338),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_225),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_51),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_403),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_6),
.Y(n_499)
);

BUFx10_ASAP7_75t_L g500 ( 
.A(n_79),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_245),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_72),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_132),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_119),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_300),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_337),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_358),
.Y(n_507)
);

CKINVDCx14_ASAP7_75t_R g508 ( 
.A(n_208),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_95),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_248),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_66),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_219),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_92),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_365),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_288),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_59),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_262),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_280),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_113),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_102),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_80),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_396),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_0),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_363),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_113),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_150),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_111),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_408),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_327),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_152),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_263),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_226),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_45),
.Y(n_533)
);

BUFx10_ASAP7_75t_L g534 ( 
.A(n_186),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_38),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_413),
.Y(n_536)
);

INVxp67_ASAP7_75t_SL g537 ( 
.A(n_315),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_111),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_11),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_23),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_325),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_50),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_64),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_244),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_218),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_230),
.Y(n_546)
);

INVxp67_ASAP7_75t_L g547 ( 
.A(n_56),
.Y(n_547)
);

BUFx10_ASAP7_75t_L g548 ( 
.A(n_298),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_252),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_233),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_241),
.Y(n_551)
);

INVx1_ASAP7_75t_SL g552 ( 
.A(n_273),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_228),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_223),
.Y(n_554)
);

CKINVDCx16_ASAP7_75t_R g555 ( 
.A(n_48),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_154),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_374),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_390),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_4),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_112),
.Y(n_560)
);

CKINVDCx16_ASAP7_75t_R g561 ( 
.A(n_144),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_297),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_49),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_107),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_243),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_62),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_328),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_242),
.Y(n_568)
);

BUFx10_ASAP7_75t_L g569 ( 
.A(n_399),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_138),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_402),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_216),
.Y(n_572)
);

BUFx5_ASAP7_75t_L g573 ( 
.A(n_392),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_194),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_265),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_96),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_175),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_264),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_401),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_285),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_166),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_64),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_6),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_320),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_410),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_29),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_148),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_257),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_228),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_290),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_307),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_421),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_419),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_256),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_180),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_90),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_310),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_400),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_140),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_123),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_177),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_164),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_133),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_131),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_60),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_261),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_195),
.Y(n_607)
);

BUFx8_ASAP7_75t_SL g608 ( 
.A(n_149),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_79),
.Y(n_609)
);

INVx1_ASAP7_75t_SL g610 ( 
.A(n_238),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_409),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_369),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_169),
.Y(n_613)
);

INVxp67_ASAP7_75t_L g614 ( 
.A(n_373),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_318),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_197),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_147),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_417),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_69),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_380),
.Y(n_620)
);

CKINVDCx14_ASAP7_75t_R g621 ( 
.A(n_216),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_183),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_302),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_185),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_204),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_225),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_291),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_237),
.Y(n_628)
);

CKINVDCx14_ASAP7_75t_R g629 ( 
.A(n_181),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_247),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_36),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_195),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_38),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_122),
.Y(n_634)
);

BUFx10_ASAP7_75t_L g635 ( 
.A(n_348),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_345),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_11),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_43),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_88),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_19),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_97),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_126),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_30),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_49),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_86),
.Y(n_645)
);

BUFx10_ASAP7_75t_L g646 ( 
.A(n_110),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_18),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_172),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_362),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_149),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_186),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_202),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_260),
.Y(n_653)
);

BUFx2_ASAP7_75t_L g654 ( 
.A(n_153),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_74),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_407),
.Y(n_656)
);

INVx1_ASAP7_75t_SL g657 ( 
.A(n_129),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_27),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_397),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_305),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_210),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_91),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_277),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_10),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_227),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_167),
.Y(n_666)
);

CKINVDCx16_ASAP7_75t_R g667 ( 
.A(n_100),
.Y(n_667)
);

BUFx5_ASAP7_75t_L g668 ( 
.A(n_393),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_71),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_97),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_267),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_229),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_206),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_148),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_125),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_227),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_420),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_412),
.Y(n_678)
);

INVx1_ASAP7_75t_SL g679 ( 
.A(n_304),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_58),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_89),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_378),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_384),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_90),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_153),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_209),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_169),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_326),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_372),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_23),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_63),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_274),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_166),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_405),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_211),
.Y(n_695)
);

INVx1_ASAP7_75t_SL g696 ( 
.A(n_347),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_351),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_15),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_176),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_109),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_77),
.Y(n_701)
);

CKINVDCx20_ASAP7_75t_R g702 ( 
.A(n_232),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_118),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_368),
.Y(n_704)
);

CKINVDCx20_ASAP7_75t_R g705 ( 
.A(n_103),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_178),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_142),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_312),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_87),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_331),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_382),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_68),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_217),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_47),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_350),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_89),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_78),
.Y(n_717)
);

BUFx5_ASAP7_75t_L g718 ( 
.A(n_161),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_56),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_160),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_139),
.Y(n_721)
);

CKINVDCx14_ASAP7_75t_R g722 ( 
.A(n_27),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_118),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_105),
.Y(n_724)
);

BUFx10_ASAP7_75t_L g725 ( 
.A(n_140),
.Y(n_725)
);

CKINVDCx20_ASAP7_75t_R g726 ( 
.A(n_383),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_1),
.Y(n_727)
);

INVx1_ASAP7_75t_SL g728 ( 
.A(n_194),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_53),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_226),
.Y(n_730)
);

CKINVDCx20_ASAP7_75t_R g731 ( 
.A(n_375),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_385),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_7),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_240),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_289),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_341),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_239),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_414),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_158),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_16),
.Y(n_740)
);

CKINVDCx14_ASAP7_75t_R g741 ( 
.A(n_366),
.Y(n_741)
);

INVx1_ASAP7_75t_SL g742 ( 
.A(n_135),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_189),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_395),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_353),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_98),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_25),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_32),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_339),
.Y(n_749)
);

INVxp67_ASAP7_75t_SL g750 ( 
.A(n_379),
.Y(n_750)
);

CKINVDCx20_ASAP7_75t_R g751 ( 
.A(n_336),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_206),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_145),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_437),
.Y(n_754)
);

CKINVDCx16_ASAP7_75t_R g755 ( 
.A(n_555),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_437),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_437),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_437),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_437),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_584),
.Y(n_760)
);

INVxp67_ASAP7_75t_L g761 ( 
.A(n_477),
.Y(n_761)
);

INVx1_ASAP7_75t_SL g762 ( 
.A(n_589),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_437),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_437),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_608),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_508),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_437),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_718),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_718),
.Y(n_769)
);

INVxp67_ASAP7_75t_L g770 ( 
.A(n_654),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_718),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_621),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_718),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_718),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_718),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_718),
.Y(n_776)
);

CKINVDCx16_ASAP7_75t_R g777 ( 
.A(n_561),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_718),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_629),
.Y(n_779)
);

BUFx3_ASAP7_75t_L g780 ( 
.A(n_584),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_604),
.Y(n_781)
);

BUFx3_ASAP7_75t_L g782 ( 
.A(n_594),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_604),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_722),
.Y(n_784)
);

INVxp67_ASAP7_75t_SL g785 ( 
.A(n_544),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_636),
.B(n_0),
.Y(n_786)
);

BUFx8_ASAP7_75t_SL g787 ( 
.A(n_426),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_604),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_560),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_667),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_560),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_485),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_492),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_492),
.Y(n_794)
);

INVx3_ASAP7_75t_L g795 ( 
.A(n_492),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_492),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_487),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_492),
.Y(n_798)
);

BUFx2_ASAP7_75t_L g799 ( 
.A(n_425),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_516),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_436),
.B(n_1),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_489),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_516),
.Y(n_803)
);

INVxp67_ASAP7_75t_SL g804 ( 
.A(n_710),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_490),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_499),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_512),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_516),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_520),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_521),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_516),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_516),
.Y(n_812)
);

INVxp67_ASAP7_75t_L g813 ( 
.A(n_502),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_525),
.Y(n_814)
);

INVx4_ASAP7_75t_R g815 ( 
.A(n_594),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_472),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_523),
.Y(n_817)
);

OR2x2_ASAP7_75t_L g818 ( 
.A(n_441),
.B(n_2),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_472),
.Y(n_819)
);

CKINVDCx16_ASAP7_75t_R g820 ( 
.A(n_439),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_525),
.Y(n_821)
);

INVx1_ASAP7_75t_SL g822 ( 
.A(n_435),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_525),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_527),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_525),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_530),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_533),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_535),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_525),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_581),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_538),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_540),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_581),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_581),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_581),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_472),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_581),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_628),
.Y(n_838)
);

CKINVDCx20_ASAP7_75t_R g839 ( 
.A(n_428),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_628),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_543),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_546),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_550),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_553),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_628),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_628),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_554),
.Y(n_847)
);

BUFx2_ASAP7_75t_L g848 ( 
.A(n_425),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_556),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_628),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_642),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_563),
.Y(n_852)
);

INVxp67_ASAP7_75t_SL g853 ( 
.A(n_614),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_570),
.Y(n_854)
);

CKINVDCx14_ASAP7_75t_R g855 ( 
.A(n_446),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_642),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_472),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_642),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_572),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_548),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_642),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_574),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_642),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_423),
.Y(n_864)
);

CKINVDCx16_ASAP7_75t_R g865 ( 
.A(n_741),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_509),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_472),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_577),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_423),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_511),
.Y(n_870)
);

CKINVDCx20_ASAP7_75t_R g871 ( 
.A(n_434),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_444),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_573),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_447),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_586),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_451),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_459),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_468),
.Y(n_878)
);

INVx1_ASAP7_75t_SL g879 ( 
.A(n_476),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_486),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_573),
.Y(n_881)
);

BUFx2_ASAP7_75t_L g882 ( 
.A(n_427),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_497),
.Y(n_883)
);

CKINVDCx20_ASAP7_75t_R g884 ( 
.A(n_529),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_595),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_532),
.Y(n_886)
);

INVx4_ASAP7_75t_R g887 ( 
.A(n_450),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_596),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_600),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_539),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_573),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_545),
.Y(n_892)
);

INVxp67_ASAP7_75t_SL g893 ( 
.A(n_440),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_551),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_564),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_576),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_582),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_548),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_603),
.Y(n_899)
);

CKINVDCx14_ASAP7_75t_R g900 ( 
.A(n_431),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_605),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_602),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_609),
.Y(n_903)
);

HB1xp67_ASAP7_75t_L g904 ( 
.A(n_427),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_607),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_431),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_616),
.Y(n_907)
);

INVxp67_ASAP7_75t_SL g908 ( 
.A(n_458),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_626),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_613),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_632),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_637),
.Y(n_912)
);

INVxp67_ASAP7_75t_L g913 ( 
.A(n_431),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_640),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_645),
.Y(n_915)
);

CKINVDCx20_ASAP7_75t_R g916 ( 
.A(n_659),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_647),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_650),
.Y(n_918)
);

BUFx3_ASAP7_75t_L g919 ( 
.A(n_548),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_573),
.Y(n_920)
);

NOR2xp67_ASAP7_75t_L g921 ( 
.A(n_547),
.B(n_2),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_573),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_655),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_617),
.Y(n_924)
);

BUFx2_ASAP7_75t_L g925 ( 
.A(n_429),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_675),
.Y(n_926)
);

CKINVDCx16_ASAP7_75t_R g927 ( 
.A(n_457),
.Y(n_927)
);

INVxp33_ASAP7_75t_L g928 ( 
.A(n_676),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_573),
.Y(n_929)
);

INVxp67_ASAP7_75t_SL g930 ( 
.A(n_460),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_622),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_624),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_573),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_680),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_685),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_569),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_625),
.Y(n_937)
);

CKINVDCx20_ASAP7_75t_R g938 ( 
.A(n_726),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_686),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_633),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_634),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_638),
.Y(n_942)
);

INVxp67_ASAP7_75t_L g943 ( 
.A(n_457),
.Y(n_943)
);

INVxp67_ASAP7_75t_L g944 ( 
.A(n_457),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_691),
.Y(n_945)
);

CKINVDCx20_ASAP7_75t_R g946 ( 
.A(n_731),
.Y(n_946)
);

CKINVDCx20_ASAP7_75t_R g947 ( 
.A(n_732),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_700),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_701),
.Y(n_949)
);

CKINVDCx20_ASAP7_75t_R g950 ( 
.A(n_751),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_643),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_706),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_644),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_709),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_648),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_712),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_716),
.Y(n_957)
);

CKINVDCx20_ASAP7_75t_R g958 ( 
.A(n_481),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_720),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_734),
.Y(n_960)
);

BUFx3_ASAP7_75t_L g961 ( 
.A(n_569),
.Y(n_961)
);

CKINVDCx20_ASAP7_75t_R g962 ( 
.A(n_484),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_740),
.Y(n_963)
);

CKINVDCx14_ASAP7_75t_R g964 ( 
.A(n_500),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_743),
.Y(n_965)
);

BUFx3_ASAP7_75t_L g966 ( 
.A(n_569),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_746),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_747),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_462),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_469),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_573),
.Y(n_971)
);

CKINVDCx20_ASAP7_75t_R g972 ( 
.A(n_488),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_471),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_687),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_483),
.Y(n_975)
);

CKINVDCx20_ASAP7_75t_R g976 ( 
.A(n_491),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_668),
.Y(n_977)
);

INVxp67_ASAP7_75t_L g978 ( 
.A(n_500),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_494),
.Y(n_979)
);

CKINVDCx16_ASAP7_75t_R g980 ( 
.A(n_500),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_690),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_498),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_510),
.Y(n_983)
);

INVxp33_ASAP7_75t_L g984 ( 
.A(n_511),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_522),
.Y(n_985)
);

INVxp67_ASAP7_75t_SL g986 ( 
.A(n_528),
.Y(n_986)
);

CKINVDCx20_ASAP7_75t_R g987 ( 
.A(n_493),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_693),
.Y(n_988)
);

INVxp67_ASAP7_75t_L g989 ( 
.A(n_534),
.Y(n_989)
);

BUFx10_ASAP7_75t_L g990 ( 
.A(n_450),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_698),
.Y(n_991)
);

INVxp67_ASAP7_75t_L g992 ( 
.A(n_534),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_541),
.Y(n_993)
);

CKINVDCx16_ASAP7_75t_R g994 ( 
.A(n_534),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_699),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_549),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_703),
.Y(n_997)
);

INVx2_ASAP7_75t_SL g998 ( 
.A(n_646),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_707),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_714),
.Y(n_1000)
);

INVxp67_ASAP7_75t_SL g1001 ( 
.A(n_557),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_565),
.Y(n_1002)
);

BUFx2_ASAP7_75t_L g1003 ( 
.A(n_429),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_717),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_719),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_571),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_578),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_579),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_588),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_668),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_590),
.Y(n_1011)
);

INVxp67_ASAP7_75t_SL g1012 ( 
.A(n_592),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_593),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_495),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_653),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_682),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_721),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_723),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_724),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_430),
.Y(n_1020)
);

CKINVDCx20_ASAP7_75t_R g1021 ( 
.A(n_501),
.Y(n_1021)
);

INVxp67_ASAP7_75t_L g1022 ( 
.A(n_646),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_668),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_519),
.Y(n_1024)
);

CKINVDCx16_ASAP7_75t_R g1025 ( 
.A(n_646),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_688),
.Y(n_1026)
);

NOR2xp67_ASAP7_75t_L g1027 ( 
.A(n_496),
.B(n_3),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_689),
.Y(n_1028)
);

INVx1_ASAP7_75t_SL g1029 ( 
.A(n_482),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_711),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_745),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_727),
.Y(n_1032)
);

CKINVDCx20_ASAP7_75t_R g1033 ( 
.A(n_506),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_505),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_729),
.Y(n_1035)
);

INVxp33_ASAP7_75t_SL g1036 ( 
.A(n_430),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_505),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_697),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_697),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_730),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_733),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_704),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_442),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_704),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_737),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_668),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_708),
.Y(n_1047)
);

CKINVDCx20_ASAP7_75t_R g1048 ( 
.A(n_507),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_708),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_442),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_519),
.Y(n_1051)
);

CKINVDCx20_ASAP7_75t_R g1052 ( 
.A(n_514),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_526),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_526),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_635),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_449),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_449),
.Y(n_1057)
);

BUFx2_ASAP7_75t_SL g1058 ( 
.A(n_496),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_568),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_568),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_452),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_587),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_668),
.Y(n_1063)
);

INVx1_ASAP7_75t_SL g1064 ( 
.A(n_503),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_452),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_515),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_587),
.Y(n_1067)
);

INVxp67_ASAP7_75t_SL g1068 ( 
.A(n_537),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_601),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_601),
.Y(n_1070)
);

CKINVDCx20_ASAP7_75t_R g1071 ( 
.A(n_517),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_695),
.Y(n_1072)
);

CKINVDCx20_ASAP7_75t_R g1073 ( 
.A(n_518),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_453),
.Y(n_1074)
);

CKINVDCx20_ASAP7_75t_R g1075 ( 
.A(n_524),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_695),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_713),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_713),
.Y(n_1078)
);

CKINVDCx14_ASAP7_75t_R g1079 ( 
.A(n_725),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_753),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_453),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_753),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_725),
.Y(n_1083)
);

CKINVDCx16_ASAP7_75t_R g1084 ( 
.A(n_725),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_566),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_566),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_669),
.Y(n_1087)
);

INVxp67_ASAP7_75t_SL g1088 ( 
.A(n_750),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_669),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_455),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_475),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_475),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_475),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_475),
.Y(n_1094)
);

CKINVDCx20_ASAP7_75t_R g1095 ( 
.A(n_531),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_455),
.Y(n_1096)
);

BUFx3_ASAP7_75t_L g1097 ( 
.A(n_635),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_475),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_562),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_463),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_562),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_668),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_668),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_562),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_562),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_463),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_466),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_466),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_562),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_467),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_424),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_424),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_635),
.Y(n_1113)
);

NOR2xp67_ASAP7_75t_L g1114 ( 
.A(n_467),
.B(n_3),
.Y(n_1114)
);

INVx1_ASAP7_75t_SL g1115 ( 
.A(n_504),
.Y(n_1115)
);

INVxp33_ASAP7_75t_SL g1116 ( 
.A(n_470),
.Y(n_1116)
);

INVxp67_ASAP7_75t_L g1117 ( 
.A(n_752),
.Y(n_1117)
);

CKINVDCx20_ASAP7_75t_R g1118 ( 
.A(n_839),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_793),
.Y(n_1119)
);

INVxp67_ASAP7_75t_SL g1120 ( 
.A(n_1113),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_794),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_796),
.Y(n_1122)
);

INVxp67_ASAP7_75t_SL g1123 ( 
.A(n_1113),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_760),
.Y(n_1124)
);

INVxp67_ASAP7_75t_SL g1125 ( 
.A(n_1113),
.Y(n_1125)
);

CKINVDCx16_ASAP7_75t_R g1126 ( 
.A(n_755),
.Y(n_1126)
);

INVxp33_ASAP7_75t_SL g1127 ( 
.A(n_766),
.Y(n_1127)
);

CKINVDCx20_ASAP7_75t_R g1128 ( 
.A(n_871),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_798),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_1113),
.B(n_465),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_958),
.Y(n_1131)
);

OR2x2_ASAP7_75t_L g1132 ( 
.A(n_762),
.B(n_513),
.Y(n_1132)
);

INVxp67_ASAP7_75t_SL g1133 ( 
.A(n_1113),
.Y(n_1133)
);

CKINVDCx20_ASAP7_75t_R g1134 ( 
.A(n_884),
.Y(n_1134)
);

INVxp67_ASAP7_75t_SL g1135 ( 
.A(n_1111),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_962),
.Y(n_1136)
);

BUFx3_ASAP7_75t_L g1137 ( 
.A(n_760),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_972),
.Y(n_1138)
);

CKINVDCx20_ASAP7_75t_R g1139 ( 
.A(n_916),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_1112),
.B(n_552),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_766),
.B(n_679),
.Y(n_1141)
);

INVxp67_ASAP7_75t_SL g1142 ( 
.A(n_780),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_976),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_800),
.Y(n_1144)
);

CKINVDCx16_ASAP7_75t_R g1145 ( 
.A(n_777),
.Y(n_1145)
);

INVxp67_ASAP7_75t_L g1146 ( 
.A(n_904),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_803),
.Y(n_1147)
);

HB1xp67_ASAP7_75t_L g1148 ( 
.A(n_790),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_808),
.Y(n_1149)
);

HB1xp67_ASAP7_75t_L g1150 ( 
.A(n_790),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_811),
.Y(n_1151)
);

HB1xp67_ASAP7_75t_L g1152 ( 
.A(n_792),
.Y(n_1152)
);

INVxp67_ASAP7_75t_L g1153 ( 
.A(n_799),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_812),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_987),
.Y(n_1155)
);

CKINVDCx20_ASAP7_75t_R g1156 ( 
.A(n_938),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_1014),
.Y(n_1157)
);

BUFx6f_ASAP7_75t_SL g1158 ( 
.A(n_860),
.Y(n_1158)
);

INVxp33_ASAP7_75t_SL g1159 ( 
.A(n_772),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_772),
.B(n_696),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_814),
.Y(n_1161)
);

CKINVDCx20_ASAP7_75t_R g1162 ( 
.A(n_946),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_1021),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_821),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_1033),
.Y(n_1165)
);

NAND2xp33_ASAP7_75t_R g1166 ( 
.A(n_792),
.B(n_432),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_823),
.Y(n_1167)
);

HB1xp67_ASAP7_75t_L g1168 ( 
.A(n_797),
.Y(n_1168)
);

CKINVDCx20_ASAP7_75t_R g1169 ( 
.A(n_947),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_794),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_825),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_829),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_795),
.Y(n_1173)
);

OR2x2_ASAP7_75t_L g1174 ( 
.A(n_906),
.B(n_610),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_797),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_779),
.B(n_432),
.Y(n_1176)
);

CKINVDCx20_ASAP7_75t_R g1177 ( 
.A(n_950),
.Y(n_1177)
);

CKINVDCx20_ASAP7_75t_R g1178 ( 
.A(n_787),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_830),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_795),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_833),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_1048),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_1052),
.Y(n_1183)
);

CKINVDCx20_ASAP7_75t_R g1184 ( 
.A(n_1066),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_1071),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_833),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_1073),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_834),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_834),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_835),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_835),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_837),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1068),
.B(n_536),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_837),
.Y(n_1194)
);

CKINVDCx20_ASAP7_75t_R g1195 ( 
.A(n_1075),
.Y(n_1195)
);

INVxp67_ASAP7_75t_L g1196 ( 
.A(n_799),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_838),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_838),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_840),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_840),
.Y(n_1200)
);

HB1xp67_ASAP7_75t_L g1201 ( 
.A(n_802),
.Y(n_1201)
);

INVxp67_ASAP7_75t_L g1202 ( 
.A(n_848),
.Y(n_1202)
);

CKINVDCx20_ASAP7_75t_R g1203 ( 
.A(n_1095),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_765),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_765),
.Y(n_1205)
);

OR2x2_ASAP7_75t_L g1206 ( 
.A(n_906),
.B(n_657),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_845),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_845),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_846),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_846),
.Y(n_1210)
);

CKINVDCx20_ASAP7_75t_R g1211 ( 
.A(n_900),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_850),
.Y(n_1212)
);

INVxp67_ASAP7_75t_L g1213 ( 
.A(n_848),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_802),
.Y(n_1214)
);

CKINVDCx20_ASAP7_75t_R g1215 ( 
.A(n_964),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_850),
.Y(n_1216)
);

CKINVDCx20_ASAP7_75t_R g1217 ( 
.A(n_1079),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_816),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_851),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_851),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_805),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_856),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_856),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_858),
.Y(n_1224)
);

INVxp67_ASAP7_75t_SL g1225 ( 
.A(n_780),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_805),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_858),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_806),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_861),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_861),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_795),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_863),
.Y(n_1232)
);

CKINVDCx20_ASAP7_75t_R g1233 ( 
.A(n_927),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_806),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_855),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_863),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_779),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_781),
.Y(n_1238)
);

CKINVDCx20_ASAP7_75t_R g1239 ( 
.A(n_980),
.Y(n_1239)
);

NOR2xp67_ASAP7_75t_L g1240 ( 
.A(n_1117),
.B(n_433),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_807),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_807),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_809),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_783),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_788),
.Y(n_1245)
);

CKINVDCx20_ASAP7_75t_R g1246 ( 
.A(n_994),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_809),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_969),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_970),
.Y(n_1249)
);

CKINVDCx16_ASAP7_75t_R g1250 ( 
.A(n_1025),
.Y(n_1250)
);

CKINVDCx20_ASAP7_75t_R g1251 ( 
.A(n_1084),
.Y(n_1251)
);

CKINVDCx16_ASAP7_75t_R g1252 ( 
.A(n_820),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_810),
.Y(n_1253)
);

CKINVDCx20_ASAP7_75t_R g1254 ( 
.A(n_822),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_810),
.Y(n_1255)
);

CKINVDCx20_ASAP7_75t_R g1256 ( 
.A(n_879),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_973),
.Y(n_1257)
);

INVxp67_ASAP7_75t_SL g1258 ( 
.A(n_782),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_817),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_768),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_782),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_975),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_817),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_979),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_982),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_824),
.Y(n_1266)
);

INVxp33_ASAP7_75t_SL g1267 ( 
.A(n_784),
.Y(n_1267)
);

CKINVDCx20_ASAP7_75t_R g1268 ( 
.A(n_1029),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_824),
.Y(n_1269)
);

INVxp67_ASAP7_75t_L g1270 ( 
.A(n_882),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_983),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_768),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_SL g1273 ( 
.A(n_860),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_784),
.B(n_433),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_985),
.Y(n_1275)
);

CKINVDCx20_ASAP7_75t_R g1276 ( 
.A(n_1064),
.Y(n_1276)
);

CKINVDCx20_ASAP7_75t_R g1277 ( 
.A(n_1115),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_826),
.Y(n_1278)
);

CKINVDCx20_ASAP7_75t_R g1279 ( 
.A(n_826),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_993),
.Y(n_1280)
);

NOR2xp67_ASAP7_75t_L g1281 ( 
.A(n_827),
.B(n_438),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_996),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_827),
.Y(n_1283)
);

HB1xp67_ASAP7_75t_L g1284 ( 
.A(n_828),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_828),
.Y(n_1285)
);

HB1xp67_ASAP7_75t_L g1286 ( 
.A(n_831),
.Y(n_1286)
);

CKINVDCx20_ASAP7_75t_R g1287 ( 
.A(n_831),
.Y(n_1287)
);

BUFx2_ASAP7_75t_L g1288 ( 
.A(n_832),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1002),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1006),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1007),
.Y(n_1291)
);

CKINVDCx20_ASAP7_75t_R g1292 ( 
.A(n_832),
.Y(n_1292)
);

CKINVDCx20_ASAP7_75t_R g1293 ( 
.A(n_841),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1008),
.Y(n_1294)
);

NOR2xp67_ASAP7_75t_L g1295 ( 
.A(n_841),
.B(n_438),
.Y(n_1295)
);

CKINVDCx20_ASAP7_75t_R g1296 ( 
.A(n_842),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1088),
.B(n_443),
.Y(n_1297)
);

CKINVDCx16_ASAP7_75t_R g1298 ( 
.A(n_865),
.Y(n_1298)
);

CKINVDCx16_ASAP7_75t_R g1299 ( 
.A(n_898),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1009),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_842),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1011),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_843),
.Y(n_1303)
);

CKINVDCx20_ASAP7_75t_R g1304 ( 
.A(n_843),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1013),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1015),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1016),
.Y(n_1307)
);

INVxp67_ASAP7_75t_SL g1308 ( 
.A(n_786),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_844),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1026),
.Y(n_1310)
);

NOR2xp67_ASAP7_75t_L g1311 ( 
.A(n_844),
.B(n_443),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_785),
.B(n_445),
.Y(n_1312)
);

XNOR2xp5_ASAP7_75t_L g1313 ( 
.A(n_866),
.B(n_542),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1028),
.Y(n_1314)
);

INVxp67_ASAP7_75t_SL g1315 ( 
.A(n_893),
.Y(n_1315)
);

INVxp67_ASAP7_75t_SL g1316 ( 
.A(n_908),
.Y(n_1316)
);

CKINVDCx20_ASAP7_75t_R g1317 ( 
.A(n_847),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_847),
.Y(n_1318)
);

INVxp67_ASAP7_75t_SL g1319 ( 
.A(n_930),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1030),
.Y(n_1320)
);

INVxp67_ASAP7_75t_SL g1321 ( 
.A(n_986),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1031),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_872),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_874),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_849),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_876),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_877),
.Y(n_1327)
);

INVxp67_ASAP7_75t_L g1328 ( 
.A(n_882),
.Y(n_1328)
);

HB1xp67_ASAP7_75t_L g1329 ( 
.A(n_849),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_878),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_852),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_852),
.Y(n_1332)
);

BUFx3_ASAP7_75t_L g1333 ( 
.A(n_789),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_880),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_883),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_854),
.Y(n_1336)
);

INVx1_ASAP7_75t_SL g1337 ( 
.A(n_898),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_854),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_886),
.Y(n_1339)
);

CKINVDCx20_ASAP7_75t_R g1340 ( 
.A(n_859),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_859),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_862),
.Y(n_1342)
);

CKINVDCx16_ASAP7_75t_R g1343 ( 
.A(n_919),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_890),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_862),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_892),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_868),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_894),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_895),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_868),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_896),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_897),
.Y(n_1352)
);

CKINVDCx20_ASAP7_75t_R g1353 ( 
.A(n_875),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_899),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_901),
.Y(n_1355)
);

BUFx2_ASAP7_75t_SL g1356 ( 
.A(n_919),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_875),
.Y(n_1357)
);

NOR2xp67_ASAP7_75t_L g1358 ( 
.A(n_885),
.B(n_445),
.Y(n_1358)
);

INVxp67_ASAP7_75t_L g1359 ( 
.A(n_925),
.Y(n_1359)
);

CKINVDCx16_ASAP7_75t_R g1360 ( 
.A(n_936),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_903),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_907),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_909),
.Y(n_1363)
);

INVxp33_ASAP7_75t_SL g1364 ( 
.A(n_885),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_888),
.Y(n_1365)
);

CKINVDCx16_ASAP7_75t_R g1366 ( 
.A(n_936),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_911),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_888),
.Y(n_1368)
);

CKINVDCx20_ASAP7_75t_R g1369 ( 
.A(n_889),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_889),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_912),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_914),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_915),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_917),
.Y(n_1374)
);

CKINVDCx20_ASAP7_75t_R g1375 ( 
.A(n_902),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_804),
.B(n_448),
.Y(n_1376)
);

NOR2xp67_ASAP7_75t_L g1377 ( 
.A(n_902),
.B(n_448),
.Y(n_1377)
);

NOR2xp67_ASAP7_75t_L g1378 ( 
.A(n_905),
.B(n_454),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_918),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_923),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_926),
.Y(n_1381)
);

INVx1_ASAP7_75t_SL g1382 ( 
.A(n_961),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_934),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_905),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_910),
.Y(n_1385)
);

CKINVDCx14_ASAP7_75t_R g1386 ( 
.A(n_961),
.Y(n_1386)
);

CKINVDCx20_ASAP7_75t_R g1387 ( 
.A(n_910),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_791),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_935),
.Y(n_1389)
);

BUFx3_ASAP7_75t_L g1390 ( 
.A(n_1085),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_939),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_924),
.Y(n_1392)
);

INVxp67_ASAP7_75t_SL g1393 ( 
.A(n_1001),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_924),
.Y(n_1394)
);

CKINVDCx20_ASAP7_75t_R g1395 ( 
.A(n_931),
.Y(n_1395)
);

CKINVDCx20_ASAP7_75t_R g1396 ( 
.A(n_931),
.Y(n_1396)
);

INVxp67_ASAP7_75t_SL g1397 ( 
.A(n_1012),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_945),
.Y(n_1398)
);

CKINVDCx20_ASAP7_75t_R g1399 ( 
.A(n_932),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_932),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_937),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_937),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_853),
.B(n_454),
.Y(n_1403)
);

NOR2xp33_ASAP7_75t_R g1404 ( 
.A(n_940),
.B(n_558),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_940),
.Y(n_1405)
);

CKINVDCx16_ASAP7_75t_R g1406 ( 
.A(n_966),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_948),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_941),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_949),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_952),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_954),
.Y(n_1411)
);

CKINVDCx20_ASAP7_75t_R g1412 ( 
.A(n_941),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_956),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_957),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_959),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_754),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_960),
.Y(n_1417)
);

INVxp33_ASAP7_75t_SL g1418 ( 
.A(n_942),
.Y(n_1418)
);

CKINVDCx20_ASAP7_75t_R g1419 ( 
.A(n_942),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_951),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_951),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_963),
.Y(n_1422)
);

CKINVDCx20_ASAP7_75t_R g1423 ( 
.A(n_953),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1121),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1323),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_SL g1426 ( 
.A1(n_1313),
.A2(n_599),
.B1(n_619),
.B2(n_559),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1121),
.Y(n_1427)
);

INVx3_ASAP7_75t_L g1428 ( 
.A(n_1218),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1120),
.B(n_756),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1324),
.Y(n_1430)
);

BUFx6f_ASAP7_75t_L g1431 ( 
.A(n_1218),
.Y(n_1431)
);

BUFx2_ASAP7_75t_L g1432 ( 
.A(n_1254),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1124),
.B(n_965),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_1193),
.B(n_1036),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_SL g1435 ( 
.A1(n_1254),
.A2(n_639),
.B1(n_641),
.B2(n_631),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1170),
.Y(n_1436)
);

BUFx3_ASAP7_75t_L g1437 ( 
.A(n_1124),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1123),
.B(n_1125),
.Y(n_1438)
);

AOI22xp5_ASAP7_75t_SL g1439 ( 
.A1(n_1279),
.A2(n_705),
.B1(n_702),
.B2(n_1036),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1133),
.B(n_757),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_L g1441 ( 
.A(n_1337),
.B(n_1382),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1326),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_SL g1443 ( 
.A(n_1130),
.B(n_953),
.Y(n_1443)
);

AOI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1308),
.A2(n_974),
.B1(n_981),
.B2(n_955),
.Y(n_1444)
);

INVx6_ASAP7_75t_L g1445 ( 
.A(n_1218),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1170),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1260),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1238),
.B(n_1058),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1327),
.Y(n_1449)
);

INVx3_ASAP7_75t_L g1450 ( 
.A(n_1218),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_1218),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1260),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1272),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1330),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1272),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_SL g1456 ( 
.A(n_1140),
.B(n_955),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1334),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1244),
.B(n_1058),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1335),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1256),
.Y(n_1460)
);

INVx5_ASAP7_75t_L g1461 ( 
.A(n_1416),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1135),
.B(n_758),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_SL g1463 ( 
.A(n_1281),
.B(n_974),
.Y(n_1463)
);

BUFx6f_ASAP7_75t_L g1464 ( 
.A(n_1416),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1339),
.Y(n_1465)
);

BUFx6f_ASAP7_75t_L g1466 ( 
.A(n_1333),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1245),
.B(n_1034),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_1131),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1344),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1315),
.B(n_759),
.Y(n_1470)
);

BUFx6f_ASAP7_75t_L g1471 ( 
.A(n_1173),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1346),
.Y(n_1472)
);

INVx6_ASAP7_75t_L g1473 ( 
.A(n_1137),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1142),
.B(n_1037),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1348),
.Y(n_1475)
);

AND2x6_ASAP7_75t_L g1476 ( 
.A(n_1297),
.B(n_873),
.Y(n_1476)
);

INVx3_ASAP7_75t_L g1477 ( 
.A(n_1173),
.Y(n_1477)
);

INVx4_ASAP7_75t_L g1478 ( 
.A(n_1180),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1349),
.Y(n_1479)
);

INVxp67_ASAP7_75t_L g1480 ( 
.A(n_1132),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1180),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1351),
.Y(n_1482)
);

AOI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1166),
.A2(n_988),
.B1(n_991),
.B2(n_981),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1352),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1231),
.Y(n_1485)
);

AND2x6_ASAP7_75t_L g1486 ( 
.A(n_1248),
.B(n_873),
.Y(n_1486)
);

AND2x4_ASAP7_75t_L g1487 ( 
.A(n_1137),
.B(n_967),
.Y(n_1487)
);

AND2x6_ASAP7_75t_L g1488 ( 
.A(n_1249),
.B(n_881),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1231),
.Y(n_1489)
);

BUFx2_ASAP7_75t_L g1490 ( 
.A(n_1256),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1354),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1181),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_1136),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1186),
.Y(n_1494)
);

BUFx6f_ASAP7_75t_L g1495 ( 
.A(n_1188),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1355),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1316),
.A2(n_1056),
.B1(n_1057),
.B2(n_1050),
.Y(n_1497)
);

INVx3_ASAP7_75t_L g1498 ( 
.A(n_1189),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_1138),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1361),
.Y(n_1500)
);

INVx3_ASAP7_75t_L g1501 ( 
.A(n_1190),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1362),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1363),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_SL g1504 ( 
.A(n_1295),
.B(n_988),
.Y(n_1504)
);

INVxp67_ASAP7_75t_L g1505 ( 
.A(n_1174),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_SL g1506 ( 
.A1(n_1268),
.A2(n_1116),
.B1(n_473),
.B2(n_474),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1225),
.B(n_1038),
.Y(n_1507)
);

NOR2x1_ASAP7_75t_L g1508 ( 
.A(n_1356),
.B(n_966),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1258),
.B(n_1039),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1367),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1371),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1191),
.Y(n_1512)
);

BUFx6f_ASAP7_75t_L g1513 ( 
.A(n_1333),
.Y(n_1513)
);

INVx2_ASAP7_75t_SL g1514 ( 
.A(n_1261),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1388),
.B(n_1042),
.Y(n_1515)
);

AND2x6_ASAP7_75t_L g1516 ( 
.A(n_1257),
.B(n_881),
.Y(n_1516)
);

BUFx6f_ASAP7_75t_L g1517 ( 
.A(n_1388),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1372),
.Y(n_1518)
);

AND2x4_ASAP7_75t_L g1519 ( 
.A(n_1261),
.B(n_968),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1373),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1319),
.B(n_1321),
.Y(n_1521)
);

AOI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1141),
.A2(n_995),
.B1(n_997),
.B2(n_991),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1374),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1379),
.Y(n_1524)
);

OAI21x1_ASAP7_75t_L g1525 ( 
.A1(n_1192),
.A2(n_764),
.B(n_763),
.Y(n_1525)
);

OA21x2_ASAP7_75t_L g1526 ( 
.A1(n_1194),
.A2(n_769),
.B(n_767),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1197),
.Y(n_1527)
);

BUFx2_ASAP7_75t_L g1528 ( 
.A(n_1268),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1198),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1393),
.B(n_771),
.Y(n_1530)
);

NOR2xp33_ASAP7_75t_SL g1531 ( 
.A(n_1211),
.B(n_1116),
.Y(n_1531)
);

BUFx6f_ASAP7_75t_L g1532 ( 
.A(n_1262),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1380),
.Y(n_1533)
);

OAI22x1_ASAP7_75t_L g1534 ( 
.A1(n_1153),
.A2(n_770),
.B1(n_761),
.B2(n_913),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1381),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_L g1536 ( 
.A(n_1397),
.B(n_1160),
.Y(n_1536)
);

OAI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1196),
.A2(n_1202),
.B1(n_1270),
.B2(n_1213),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1199),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1383),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1264),
.B(n_864),
.Y(n_1540)
);

BUFx6f_ASAP7_75t_L g1541 ( 
.A(n_1265),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1328),
.A2(n_1050),
.B1(n_1057),
.B2(n_1056),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_R g1543 ( 
.A(n_1155),
.B(n_995),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1200),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1389),
.Y(n_1545)
);

AND2x4_ASAP7_75t_L g1546 ( 
.A(n_1271),
.B(n_864),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_SL g1547 ( 
.A1(n_1276),
.A2(n_473),
.B1(n_474),
.B2(n_470),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1391),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1403),
.B(n_773),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1207),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1398),
.Y(n_1551)
);

INVx3_ASAP7_75t_L g1552 ( 
.A(n_1208),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1275),
.B(n_869),
.Y(n_1553)
);

BUFx6f_ASAP7_75t_L g1554 ( 
.A(n_1209),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1312),
.B(n_774),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1407),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_L g1557 ( 
.A(n_1210),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1409),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1212),
.Y(n_1559)
);

BUFx6f_ASAP7_75t_L g1560 ( 
.A(n_1216),
.Y(n_1560)
);

BUFx6f_ASAP7_75t_L g1561 ( 
.A(n_1219),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1359),
.A2(n_1061),
.B1(n_1074),
.B2(n_1065),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1220),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1280),
.B(n_1044),
.Y(n_1564)
);

INVx6_ASAP7_75t_L g1565 ( 
.A(n_1390),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1222),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1410),
.Y(n_1567)
);

INVx3_ASAP7_75t_L g1568 ( 
.A(n_1223),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1224),
.Y(n_1569)
);

AND2x4_ASAP7_75t_L g1570 ( 
.A(n_1282),
.B(n_869),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1411),
.Y(n_1571)
);

AOI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1146),
.A2(n_997),
.B1(n_1000),
.B2(n_999),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1289),
.B(n_870),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1206),
.B(n_925),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1290),
.B(n_1047),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1413),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1291),
.B(n_870),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1414),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1294),
.B(n_1024),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1376),
.B(n_775),
.Y(n_1580)
);

NAND2xp33_ASAP7_75t_L g1581 ( 
.A(n_1300),
.B(n_668),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1415),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1227),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1417),
.Y(n_1584)
);

INVx3_ASAP7_75t_L g1585 ( 
.A(n_1229),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1230),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1422),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1302),
.B(n_1049),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1232),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1240),
.B(n_776),
.Y(n_1590)
);

INVx2_ASAP7_75t_SL g1591 ( 
.A(n_1148),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1236),
.B(n_778),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1305),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1119),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1306),
.Y(n_1595)
);

INVx3_ASAP7_75t_L g1596 ( 
.A(n_1122),
.Y(n_1596)
);

BUFx6f_ASAP7_75t_L g1597 ( 
.A(n_1129),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1144),
.Y(n_1598)
);

BUFx6f_ASAP7_75t_L g1599 ( 
.A(n_1147),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1149),
.B(n_1099),
.Y(n_1600)
);

BUFx3_ASAP7_75t_L g1601 ( 
.A(n_1390),
.Y(n_1601)
);

NOR2x1_ASAP7_75t_L g1602 ( 
.A(n_1311),
.B(n_1358),
.Y(n_1602)
);

BUFx6f_ASAP7_75t_L g1603 ( 
.A(n_1151),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1276),
.Y(n_1604)
);

BUFx6f_ASAP7_75t_L g1605 ( 
.A(n_1154),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1307),
.B(n_1310),
.Y(n_1606)
);

INVxp67_ASAP7_75t_L g1607 ( 
.A(n_1176),
.Y(n_1607)
);

CKINVDCx20_ASAP7_75t_R g1608 ( 
.A(n_1277),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1314),
.B(n_1320),
.Y(n_1609)
);

BUFx6f_ASAP7_75t_L g1610 ( 
.A(n_1161),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1322),
.Y(n_1611)
);

CKINVDCx20_ASAP7_75t_R g1612 ( 
.A(n_1277),
.Y(n_1612)
);

BUFx6f_ASAP7_75t_L g1613 ( 
.A(n_1164),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1167),
.Y(n_1614)
);

BUFx6f_ASAP7_75t_L g1615 ( 
.A(n_1171),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1172),
.B(n_1101),
.Y(n_1616)
);

AOI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1377),
.A2(n_999),
.B1(n_1004),
.B2(n_1000),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1274),
.B(n_1004),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1179),
.Y(n_1619)
);

BUFx6f_ASAP7_75t_L g1620 ( 
.A(n_1288),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1386),
.B(n_984),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_1143),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1364),
.B(n_1005),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1158),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1378),
.B(n_1104),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1404),
.B(n_1105),
.Y(n_1626)
);

AND2x6_ASAP7_75t_L g1627 ( 
.A(n_1158),
.B(n_891),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1158),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1299),
.B(n_1024),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1343),
.B(n_1109),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1360),
.B(n_1005),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1152),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1273),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1168),
.B(n_1051),
.Y(n_1634)
);

BUFx3_ASAP7_75t_L g1635 ( 
.A(n_1214),
.Y(n_1635)
);

INVx3_ASAP7_75t_L g1636 ( 
.A(n_1273),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1175),
.Y(n_1637)
);

BUFx6f_ASAP7_75t_L g1638 ( 
.A(n_1221),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1273),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1201),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1242),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_1163),
.Y(n_1642)
);

INVx6_ASAP7_75t_L g1643 ( 
.A(n_1366),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1243),
.Y(n_1644)
);

BUFx6f_ASAP7_75t_L g1645 ( 
.A(n_1226),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1284),
.Y(n_1646)
);

AND2x2_ASAP7_75t_SL g1647 ( 
.A(n_1286),
.B(n_801),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1406),
.B(n_1053),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1329),
.B(n_1054),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1228),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1252),
.B(n_1059),
.Y(n_1651)
);

OA21x2_ASAP7_75t_L g1652 ( 
.A1(n_1345),
.A2(n_1092),
.B(n_1091),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1150),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1126),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1234),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1241),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1235),
.B(n_1060),
.Y(n_1657)
);

INVx4_ASAP7_75t_L g1658 ( 
.A(n_1235),
.Y(n_1658)
);

OA21x2_ASAP7_75t_L g1659 ( 
.A1(n_1345),
.A2(n_1092),
.B(n_1091),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1145),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1247),
.Y(n_1661)
);

BUFx2_ASAP7_75t_L g1662 ( 
.A(n_1279),
.Y(n_1662)
);

AND2x4_ASAP7_75t_L g1663 ( 
.A(n_1253),
.B(n_1062),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1255),
.Y(n_1664)
);

BUFx6f_ASAP7_75t_L g1665 ( 
.A(n_1259),
.Y(n_1665)
);

INVx6_ASAP7_75t_L g1666 ( 
.A(n_1298),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1263),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1266),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1269),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1364),
.B(n_1017),
.Y(n_1670)
);

OA21x2_ASAP7_75t_L g1671 ( 
.A1(n_1347),
.A2(n_1094),
.B(n_1093),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1418),
.B(n_1017),
.Y(n_1672)
);

BUFx2_ASAP7_75t_L g1673 ( 
.A(n_1287),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1278),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1283),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1285),
.Y(n_1676)
);

BUFx3_ASAP7_75t_L g1677 ( 
.A(n_1301),
.Y(n_1677)
);

AND2x4_ASAP7_75t_L g1678 ( 
.A(n_1303),
.B(n_1067),
.Y(n_1678)
);

INVx3_ASAP7_75t_L g1679 ( 
.A(n_1309),
.Y(n_1679)
);

BUFx6f_ASAP7_75t_L g1680 ( 
.A(n_1318),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1325),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1331),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1332),
.B(n_1069),
.Y(n_1683)
);

BUFx2_ASAP7_75t_L g1684 ( 
.A(n_1287),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1418),
.B(n_1018),
.Y(n_1685)
);

BUFx6f_ASAP7_75t_L g1686 ( 
.A(n_1336),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1338),
.Y(n_1687)
);

BUFx3_ASAP7_75t_L g1688 ( 
.A(n_1341),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1342),
.Y(n_1689)
);

OAI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1127),
.A2(n_1061),
.B1(n_1074),
.B2(n_1065),
.Y(n_1690)
);

INVx2_ASAP7_75t_SL g1691 ( 
.A(n_1421),
.Y(n_1691)
);

OAI21x1_ASAP7_75t_L g1692 ( 
.A1(n_1127),
.A2(n_920),
.B(n_891),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1347),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1350),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1350),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1357),
.B(n_1070),
.Y(n_1696)
);

INVx3_ASAP7_75t_L g1697 ( 
.A(n_1357),
.Y(n_1697)
);

AND2x6_ASAP7_75t_L g1698 ( 
.A(n_1159),
.B(n_920),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1368),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1368),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1370),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1370),
.Y(n_1702)
);

AOI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1159),
.A2(n_1018),
.B1(n_1032),
.B2(n_1019),
.Y(n_1703)
);

INVxp67_ASAP7_75t_L g1704 ( 
.A(n_1384),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1384),
.B(n_1019),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1385),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1385),
.Y(n_1707)
);

INVx3_ASAP7_75t_L g1708 ( 
.A(n_1392),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1392),
.Y(n_1709)
);

AND2x4_ASAP7_75t_L g1710 ( 
.A(n_1394),
.B(n_1072),
.Y(n_1710)
);

AOI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1267),
.A2(n_1032),
.B1(n_1040),
.B2(n_1035),
.Y(n_1711)
);

HB1xp67_ASAP7_75t_L g1712 ( 
.A(n_1394),
.Y(n_1712)
);

CKINVDCx5p33_ASAP7_75t_R g1713 ( 
.A(n_1468),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_1468),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1447),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1467),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1447),
.Y(n_1717)
);

INVx1_ASAP7_75t_SL g1718 ( 
.A(n_1608),
.Y(n_1718)
);

CKINVDCx20_ASAP7_75t_R g1719 ( 
.A(n_1493),
.Y(n_1719)
);

CKINVDCx5p33_ASAP7_75t_R g1720 ( 
.A(n_1493),
.Y(n_1720)
);

CKINVDCx20_ASAP7_75t_R g1721 ( 
.A(n_1499),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1452),
.Y(n_1722)
);

CKINVDCx5p33_ASAP7_75t_R g1723 ( 
.A(n_1499),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_R g1724 ( 
.A(n_1622),
.B(n_1155),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1467),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_R g1726 ( 
.A(n_1622),
.B(n_1157),
.Y(n_1726)
);

INVx3_ASAP7_75t_L g1727 ( 
.A(n_1692),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_1642),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_SL g1729 ( 
.A(n_1441),
.B(n_1400),
.Y(n_1729)
);

NOR2xp33_ASAP7_75t_SL g1730 ( 
.A(n_1658),
.B(n_1400),
.Y(n_1730)
);

CKINVDCx5p33_ASAP7_75t_R g1731 ( 
.A(n_1642),
.Y(n_1731)
);

CKINVDCx20_ASAP7_75t_R g1732 ( 
.A(n_1608),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1452),
.Y(n_1733)
);

CKINVDCx5p33_ASAP7_75t_R g1734 ( 
.A(n_1543),
.Y(n_1734)
);

INVx3_ASAP7_75t_L g1735 ( 
.A(n_1692),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_1612),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1607),
.B(n_1401),
.Y(n_1737)
);

CKINVDCx5p33_ASAP7_75t_R g1738 ( 
.A(n_1612),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1540),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_1666),
.Y(n_1740)
);

NOR2xp67_ASAP7_75t_L g1741 ( 
.A(n_1658),
.B(n_1704),
.Y(n_1741)
);

BUFx6f_ASAP7_75t_SL g1742 ( 
.A(n_1658),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_1666),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_SL g1744 ( 
.A(n_1536),
.B(n_1401),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_1666),
.Y(n_1745)
);

CKINVDCx16_ASAP7_75t_R g1746 ( 
.A(n_1654),
.Y(n_1746)
);

CKINVDCx5p33_ASAP7_75t_R g1747 ( 
.A(n_1666),
.Y(n_1747)
);

CKINVDCx5p33_ASAP7_75t_R g1748 ( 
.A(n_1643),
.Y(n_1748)
);

CKINVDCx5p33_ASAP7_75t_R g1749 ( 
.A(n_1643),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_1643),
.Y(n_1750)
);

CKINVDCx20_ASAP7_75t_R g1751 ( 
.A(n_1660),
.Y(n_1751)
);

INVxp67_ASAP7_75t_L g1752 ( 
.A(n_1621),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_1643),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1540),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1540),
.Y(n_1755)
);

CKINVDCx20_ASAP7_75t_R g1756 ( 
.A(n_1635),
.Y(n_1756)
);

CKINVDCx20_ASAP7_75t_R g1757 ( 
.A(n_1635),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1546),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_1680),
.Y(n_1759)
);

CKINVDCx5p33_ASAP7_75t_R g1760 ( 
.A(n_1680),
.Y(n_1760)
);

CKINVDCx5p33_ASAP7_75t_R g1761 ( 
.A(n_1680),
.Y(n_1761)
);

CKINVDCx5p33_ASAP7_75t_R g1762 ( 
.A(n_1680),
.Y(n_1762)
);

CKINVDCx20_ASAP7_75t_R g1763 ( 
.A(n_1677),
.Y(n_1763)
);

HB1xp67_ASAP7_75t_L g1764 ( 
.A(n_1629),
.Y(n_1764)
);

XNOR2xp5_ASAP7_75t_L g1765 ( 
.A(n_1439),
.B(n_1118),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1546),
.Y(n_1766)
);

CKINVDCx5p33_ASAP7_75t_R g1767 ( 
.A(n_1638),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_1638),
.Y(n_1768)
);

CKINVDCx5p33_ASAP7_75t_R g1769 ( 
.A(n_1638),
.Y(n_1769)
);

BUFx2_ASAP7_75t_L g1770 ( 
.A(n_1432),
.Y(n_1770)
);

INVx3_ASAP7_75t_L g1771 ( 
.A(n_1478),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_R g1772 ( 
.A(n_1636),
.B(n_1157),
.Y(n_1772)
);

INVx1_ASAP7_75t_SL g1773 ( 
.A(n_1621),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1546),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_R g1775 ( 
.A(n_1636),
.B(n_1165),
.Y(n_1775)
);

INVx3_ASAP7_75t_L g1776 ( 
.A(n_1478),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1553),
.Y(n_1777)
);

CKINVDCx5p33_ASAP7_75t_R g1778 ( 
.A(n_1677),
.Y(n_1778)
);

CKINVDCx5p33_ASAP7_75t_R g1779 ( 
.A(n_1688),
.Y(n_1779)
);

CKINVDCx5p33_ASAP7_75t_R g1780 ( 
.A(n_1638),
.Y(n_1780)
);

BUFx2_ASAP7_75t_L g1781 ( 
.A(n_1432),
.Y(n_1781)
);

CKINVDCx5p33_ASAP7_75t_R g1782 ( 
.A(n_1688),
.Y(n_1782)
);

CKINVDCx20_ASAP7_75t_R g1783 ( 
.A(n_1490),
.Y(n_1783)
);

CKINVDCx20_ASAP7_75t_R g1784 ( 
.A(n_1490),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_1638),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_R g1786 ( 
.A(n_1636),
.B(n_1165),
.Y(n_1786)
);

CKINVDCx5p33_ASAP7_75t_R g1787 ( 
.A(n_1645),
.Y(n_1787)
);

CKINVDCx5p33_ASAP7_75t_R g1788 ( 
.A(n_1645),
.Y(n_1788)
);

NAND2x1p5_ASAP7_75t_L g1789 ( 
.A(n_1652),
.B(n_816),
.Y(n_1789)
);

CKINVDCx5p33_ASAP7_75t_R g1790 ( 
.A(n_1645),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1553),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1553),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1549),
.B(n_1035),
.Y(n_1793)
);

CKINVDCx5p33_ASAP7_75t_R g1794 ( 
.A(n_1645),
.Y(n_1794)
);

CKINVDCx5p33_ASAP7_75t_R g1795 ( 
.A(n_1645),
.Y(n_1795)
);

NOR2xp67_ASAP7_75t_L g1796 ( 
.A(n_1480),
.B(n_1204),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_1665),
.Y(n_1797)
);

HB1xp67_ASAP7_75t_L g1798 ( 
.A(n_1629),
.Y(n_1798)
);

CKINVDCx5p33_ASAP7_75t_R g1799 ( 
.A(n_1665),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1453),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_1665),
.Y(n_1801)
);

CKINVDCx5p33_ASAP7_75t_R g1802 ( 
.A(n_1665),
.Y(n_1802)
);

CKINVDCx6p67_ASAP7_75t_R g1803 ( 
.A(n_1665),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1570),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1570),
.Y(n_1805)
);

CKINVDCx5p33_ASAP7_75t_R g1806 ( 
.A(n_1686),
.Y(n_1806)
);

CKINVDCx5p33_ASAP7_75t_R g1807 ( 
.A(n_1686),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1570),
.Y(n_1808)
);

CKINVDCx5p33_ASAP7_75t_R g1809 ( 
.A(n_1686),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1573),
.Y(n_1810)
);

CKINVDCx5p33_ASAP7_75t_R g1811 ( 
.A(n_1686),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1453),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_R g1813 ( 
.A(n_1697),
.B(n_1182),
.Y(n_1813)
);

NOR2xp33_ASAP7_75t_R g1814 ( 
.A(n_1697),
.B(n_1182),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1573),
.Y(n_1815)
);

NOR2xp33_ASAP7_75t_L g1816 ( 
.A(n_1434),
.B(n_1402),
.Y(n_1816)
);

CKINVDCx16_ASAP7_75t_R g1817 ( 
.A(n_1531),
.Y(n_1817)
);

NOR2xp33_ASAP7_75t_L g1818 ( 
.A(n_1456),
.B(n_1402),
.Y(n_1818)
);

CKINVDCx5p33_ASAP7_75t_R g1819 ( 
.A(n_1686),
.Y(n_1819)
);

HB1xp67_ASAP7_75t_L g1820 ( 
.A(n_1648),
.Y(n_1820)
);

CKINVDCx5p33_ASAP7_75t_R g1821 ( 
.A(n_1618),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1573),
.Y(n_1822)
);

CKINVDCx5p33_ASAP7_75t_R g1823 ( 
.A(n_1620),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1455),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1577),
.Y(n_1825)
);

CKINVDCx20_ASAP7_75t_R g1826 ( 
.A(n_1528),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1455),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_1620),
.Y(n_1828)
);

INVx3_ASAP7_75t_L g1829 ( 
.A(n_1478),
.Y(n_1829)
);

NAND2xp33_ASAP7_75t_R g1830 ( 
.A(n_1528),
.B(n_1405),
.Y(n_1830)
);

CKINVDCx5p33_ASAP7_75t_R g1831 ( 
.A(n_1620),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1424),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_SL g1833 ( 
.A(n_1647),
.B(n_1405),
.Y(n_1833)
);

BUFx2_ASAP7_75t_L g1834 ( 
.A(n_1460),
.Y(n_1834)
);

CKINVDCx5p33_ASAP7_75t_R g1835 ( 
.A(n_1620),
.Y(n_1835)
);

CKINVDCx5p33_ASAP7_75t_R g1836 ( 
.A(n_1623),
.Y(n_1836)
);

CKINVDCx5p33_ASAP7_75t_R g1837 ( 
.A(n_1662),
.Y(n_1837)
);

CKINVDCx20_ASAP7_75t_R g1838 ( 
.A(n_1604),
.Y(n_1838)
);

NOR2xp33_ASAP7_75t_R g1839 ( 
.A(n_1697),
.B(n_1183),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1424),
.Y(n_1840)
);

CKINVDCx20_ASAP7_75t_R g1841 ( 
.A(n_1712),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1474),
.B(n_1003),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1577),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_SL g1844 ( 
.A(n_1647),
.B(n_1408),
.Y(n_1844)
);

CKINVDCx5p33_ASAP7_75t_R g1845 ( 
.A(n_1685),
.Y(n_1845)
);

CKINVDCx5p33_ASAP7_75t_R g1846 ( 
.A(n_1679),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1427),
.Y(n_1847)
);

CKINVDCx5p33_ASAP7_75t_R g1848 ( 
.A(n_1679),
.Y(n_1848)
);

CKINVDCx5p33_ASAP7_75t_R g1849 ( 
.A(n_1679),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1577),
.Y(n_1850)
);

CKINVDCx5p33_ASAP7_75t_R g1851 ( 
.A(n_1691),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1579),
.Y(n_1852)
);

CKINVDCx5p33_ASAP7_75t_R g1853 ( 
.A(n_1691),
.Y(n_1853)
);

NOR2xp67_ASAP7_75t_L g1854 ( 
.A(n_1483),
.B(n_1205),
.Y(n_1854)
);

CKINVDCx16_ASAP7_75t_R g1855 ( 
.A(n_1662),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1579),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1579),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1609),
.Y(n_1858)
);

INVxp67_ASAP7_75t_SL g1859 ( 
.A(n_1464),
.Y(n_1859)
);

INVx3_ASAP7_75t_L g1860 ( 
.A(n_1526),
.Y(n_1860)
);

HB1xp67_ASAP7_75t_L g1861 ( 
.A(n_1648),
.Y(n_1861)
);

BUFx6f_ASAP7_75t_L g1862 ( 
.A(n_1525),
.Y(n_1862)
);

CKINVDCx5p33_ASAP7_75t_R g1863 ( 
.A(n_1437),
.Y(n_1863)
);

NAND2xp33_ASAP7_75t_R g1864 ( 
.A(n_1652),
.B(n_1408),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1609),
.Y(n_1865)
);

INVx3_ASAP7_75t_L g1866 ( 
.A(n_1526),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1474),
.B(n_1003),
.Y(n_1867)
);

CKINVDCx20_ASAP7_75t_R g1868 ( 
.A(n_1673),
.Y(n_1868)
);

BUFx3_ASAP7_75t_L g1869 ( 
.A(n_1473),
.Y(n_1869)
);

CKINVDCx20_ASAP7_75t_R g1870 ( 
.A(n_1673),
.Y(n_1870)
);

NOR2x1p5_ASAP7_75t_L g1871 ( 
.A(n_1624),
.B(n_1055),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1507),
.B(n_1020),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1427),
.Y(n_1873)
);

NOR2x1p5_ASAP7_75t_L g1874 ( 
.A(n_1624),
.B(n_1628),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1564),
.Y(n_1875)
);

CKINVDCx16_ASAP7_75t_R g1876 ( 
.A(n_1684),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_R g1877 ( 
.A(n_1708),
.B(n_1183),
.Y(n_1877)
);

CKINVDCx5p33_ASAP7_75t_R g1878 ( 
.A(n_1437),
.Y(n_1878)
);

CKINVDCx5p33_ASAP7_75t_R g1879 ( 
.A(n_1650),
.Y(n_1879)
);

INVx1_ASAP7_75t_SL g1880 ( 
.A(n_1574),
.Y(n_1880)
);

CKINVDCx20_ASAP7_75t_R g1881 ( 
.A(n_1684),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1507),
.B(n_1020),
.Y(n_1882)
);

CKINVDCx16_ASAP7_75t_R g1883 ( 
.A(n_1703),
.Y(n_1883)
);

BUFx2_ASAP7_75t_L g1884 ( 
.A(n_1651),
.Y(n_1884)
);

CKINVDCx5p33_ASAP7_75t_R g1885 ( 
.A(n_1650),
.Y(n_1885)
);

CKINVDCx5p33_ASAP7_75t_R g1886 ( 
.A(n_1655),
.Y(n_1886)
);

CKINVDCx5p33_ASAP7_75t_R g1887 ( 
.A(n_1690),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1564),
.Y(n_1888)
);

CKINVDCx20_ASAP7_75t_R g1889 ( 
.A(n_1631),
.Y(n_1889)
);

CKINVDCx5p33_ASAP7_75t_R g1890 ( 
.A(n_1435),
.Y(n_1890)
);

NOR2xp33_ASAP7_75t_R g1891 ( 
.A(n_1708),
.B(n_1185),
.Y(n_1891)
);

CKINVDCx20_ASAP7_75t_R g1892 ( 
.A(n_1670),
.Y(n_1892)
);

INVx3_ASAP7_75t_L g1893 ( 
.A(n_1526),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1575),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1575),
.Y(n_1895)
);

CKINVDCx5p33_ASAP7_75t_R g1896 ( 
.A(n_1708),
.Y(n_1896)
);

NOR2xp33_ASAP7_75t_R g1897 ( 
.A(n_1693),
.B(n_1185),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1588),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1588),
.Y(n_1899)
);

CKINVDCx5p33_ASAP7_75t_R g1900 ( 
.A(n_1426),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1436),
.Y(n_1901)
);

CKINVDCx5p33_ASAP7_75t_R g1902 ( 
.A(n_1711),
.Y(n_1902)
);

CKINVDCx5p33_ASAP7_75t_R g1903 ( 
.A(n_1542),
.Y(n_1903)
);

CKINVDCx5p33_ASAP7_75t_R g1904 ( 
.A(n_1562),
.Y(n_1904)
);

BUFx10_ASAP7_75t_L g1905 ( 
.A(n_1657),
.Y(n_1905)
);

CKINVDCx5p33_ASAP7_75t_R g1906 ( 
.A(n_1522),
.Y(n_1906)
);

BUFx2_ASAP7_75t_L g1907 ( 
.A(n_1651),
.Y(n_1907)
);

HB1xp67_ASAP7_75t_L g1908 ( 
.A(n_1683),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1509),
.B(n_1043),
.Y(n_1909)
);

CKINVDCx5p33_ASAP7_75t_R g1910 ( 
.A(n_1572),
.Y(n_1910)
);

CKINVDCx5p33_ASAP7_75t_R g1911 ( 
.A(n_1497),
.Y(n_1911)
);

INVxp67_ASAP7_75t_L g1912 ( 
.A(n_1574),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1436),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1446),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1425),
.Y(n_1915)
);

CKINVDCx20_ASAP7_75t_R g1916 ( 
.A(n_1672),
.Y(n_1916)
);

CKINVDCx5p33_ASAP7_75t_R g1917 ( 
.A(n_1444),
.Y(n_1917)
);

INVxp67_ASAP7_75t_L g1918 ( 
.A(n_1683),
.Y(n_1918)
);

CKINVDCx20_ASAP7_75t_R g1919 ( 
.A(n_1705),
.Y(n_1919)
);

CKINVDCx5p33_ASAP7_75t_R g1920 ( 
.A(n_1617),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_1537),
.Y(n_1921)
);

CKINVDCx5p33_ASAP7_75t_R g1922 ( 
.A(n_1655),
.Y(n_1922)
);

CKINVDCx5p33_ASAP7_75t_R g1923 ( 
.A(n_1656),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1430),
.Y(n_1924)
);

HB1xp67_ASAP7_75t_L g1925 ( 
.A(n_1710),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1509),
.B(n_1043),
.Y(n_1926)
);

CKINVDCx20_ASAP7_75t_R g1927 ( 
.A(n_1463),
.Y(n_1927)
);

NOR2xp67_ASAP7_75t_L g1928 ( 
.A(n_1505),
.B(n_1420),
.Y(n_1928)
);

INVx8_ASAP7_75t_L g1929 ( 
.A(n_1698),
.Y(n_1929)
);

NOR2xp33_ASAP7_75t_L g1930 ( 
.A(n_1456),
.B(n_1420),
.Y(n_1930)
);

CKINVDCx5p33_ASAP7_75t_R g1931 ( 
.A(n_1656),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1446),
.Y(n_1932)
);

CKINVDCx5p33_ASAP7_75t_R g1933 ( 
.A(n_1664),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1448),
.B(n_998),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1555),
.B(n_1040),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1442),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1449),
.Y(n_1937)
);

CKINVDCx5p33_ASAP7_75t_R g1938 ( 
.A(n_1664),
.Y(n_1938)
);

CKINVDCx16_ASAP7_75t_R g1939 ( 
.A(n_1591),
.Y(n_1939)
);

CKINVDCx20_ASAP7_75t_R g1940 ( 
.A(n_1463),
.Y(n_1940)
);

INVx3_ASAP7_75t_L g1941 ( 
.A(n_1471),
.Y(n_1941)
);

CKINVDCx5p33_ASAP7_75t_R g1942 ( 
.A(n_1668),
.Y(n_1942)
);

CKINVDCx5p33_ASAP7_75t_R g1943 ( 
.A(n_1668),
.Y(n_1943)
);

CKINVDCx5p33_ASAP7_75t_R g1944 ( 
.A(n_1682),
.Y(n_1944)
);

NAND2xp33_ASAP7_75t_R g1945 ( 
.A(n_1652),
.B(n_1237),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_R g1946 ( 
.A(n_1695),
.B(n_1178),
.Y(n_1946)
);

CKINVDCx5p33_ASAP7_75t_R g1947 ( 
.A(n_1682),
.Y(n_1947)
);

CKINVDCx20_ASAP7_75t_R g1948 ( 
.A(n_1504),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1454),
.Y(n_1949)
);

CKINVDCx5p33_ASAP7_75t_R g1950 ( 
.A(n_1689),
.Y(n_1950)
);

BUFx2_ASAP7_75t_L g1951 ( 
.A(n_1640),
.Y(n_1951)
);

INVx3_ASAP7_75t_L g1952 ( 
.A(n_1471),
.Y(n_1952)
);

AND2x4_ASAP7_75t_L g1953 ( 
.A(n_1514),
.B(n_1076),
.Y(n_1953)
);

CKINVDCx5p33_ASAP7_75t_R g1954 ( 
.A(n_1689),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1457),
.Y(n_1955)
);

CKINVDCx5p33_ASAP7_75t_R g1956 ( 
.A(n_1661),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1459),
.Y(n_1957)
);

CKINVDCx5p33_ASAP7_75t_R g1958 ( 
.A(n_1667),
.Y(n_1958)
);

CKINVDCx5p33_ASAP7_75t_R g1959 ( 
.A(n_1669),
.Y(n_1959)
);

CKINVDCx5p33_ASAP7_75t_R g1960 ( 
.A(n_1674),
.Y(n_1960)
);

CKINVDCx5p33_ASAP7_75t_R g1961 ( 
.A(n_1675),
.Y(n_1961)
);

CKINVDCx5p33_ASAP7_75t_R g1962 ( 
.A(n_1676),
.Y(n_1962)
);

INVx2_ASAP7_75t_SL g1963 ( 
.A(n_1659),
.Y(n_1963)
);

CKINVDCx5p33_ASAP7_75t_R g1964 ( 
.A(n_1681),
.Y(n_1964)
);

CKINVDCx16_ASAP7_75t_R g1965 ( 
.A(n_1591),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1481),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1465),
.Y(n_1967)
);

CKINVDCx5p33_ASAP7_75t_R g1968 ( 
.A(n_1687),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_1694),
.Y(n_1969)
);

CKINVDCx5p33_ASAP7_75t_R g1970 ( 
.A(n_1694),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1469),
.Y(n_1971)
);

CKINVDCx5p33_ASAP7_75t_R g1972 ( 
.A(n_1700),
.Y(n_1972)
);

CKINVDCx5p33_ASAP7_75t_R g1973 ( 
.A(n_1700),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1472),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1475),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1481),
.Y(n_1976)
);

INVx3_ASAP7_75t_L g1977 ( 
.A(n_1471),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1479),
.Y(n_1978)
);

CKINVDCx5p33_ASAP7_75t_R g1979 ( 
.A(n_1701),
.Y(n_1979)
);

CKINVDCx5p33_ASAP7_75t_R g1980 ( 
.A(n_1701),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1482),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1448),
.B(n_998),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1484),
.Y(n_1983)
);

CKINVDCx5p33_ASAP7_75t_R g1984 ( 
.A(n_1706),
.Y(n_1984)
);

CKINVDCx5p33_ASAP7_75t_R g1985 ( 
.A(n_1706),
.Y(n_1985)
);

CKINVDCx5p33_ASAP7_75t_R g1986 ( 
.A(n_1707),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1491),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1485),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1485),
.Y(n_1989)
);

NOR2xp33_ASAP7_75t_R g1990 ( 
.A(n_1699),
.B(n_1178),
.Y(n_1990)
);

INVxp67_ASAP7_75t_L g1991 ( 
.A(n_1696),
.Y(n_1991)
);

CKINVDCx5p33_ASAP7_75t_R g1992 ( 
.A(n_1707),
.Y(n_1992)
);

CKINVDCx5p33_ASAP7_75t_R g1993 ( 
.A(n_1709),
.Y(n_1993)
);

CKINVDCx5p33_ASAP7_75t_R g1994 ( 
.A(n_1709),
.Y(n_1994)
);

CKINVDCx20_ASAP7_75t_R g1995 ( 
.A(n_1504),
.Y(n_1995)
);

AO21x2_ASAP7_75t_L g1996 ( 
.A1(n_1525),
.A2(n_1094),
.B(n_1093),
.Y(n_1996)
);

INVx3_ASAP7_75t_L g1997 ( 
.A(n_1471),
.Y(n_1997)
);

CKINVDCx5p33_ASAP7_75t_R g1998 ( 
.A(n_1506),
.Y(n_1998)
);

INVx2_ASAP7_75t_SL g1999 ( 
.A(n_1659),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1489),
.Y(n_2000)
);

BUFx10_ASAP7_75t_L g2001 ( 
.A(n_1657),
.Y(n_2001)
);

OA21x2_ASAP7_75t_L g2002 ( 
.A1(n_1592),
.A2(n_1098),
.B(n_929),
.Y(n_2002)
);

CKINVDCx5p33_ASAP7_75t_R g2003 ( 
.A(n_1702),
.Y(n_2003)
);

CKINVDCx5p33_ASAP7_75t_R g2004 ( 
.A(n_1628),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1489),
.Y(n_2005)
);

NOR2xp33_ASAP7_75t_R g2006 ( 
.A(n_1632),
.B(n_1118),
.Y(n_2006)
);

CKINVDCx5p33_ASAP7_75t_R g2007 ( 
.A(n_1633),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1966),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1966),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_SL g2010 ( 
.A(n_1771),
.B(n_1532),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1715),
.Y(n_2011)
);

INVx4_ASAP7_75t_SL g2012 ( 
.A(n_1963),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1934),
.B(n_1521),
.Y(n_2013)
);

INVx1_ASAP7_75t_SL g2014 ( 
.A(n_1880),
.Y(n_2014)
);

INVx1_ASAP7_75t_SL g2015 ( 
.A(n_1939),
.Y(n_2015)
);

BUFx6f_ASAP7_75t_L g2016 ( 
.A(n_1869),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1934),
.B(n_1982),
.Y(n_2017)
);

AOI22xp33_ASAP7_75t_L g2018 ( 
.A1(n_1963),
.A2(n_1999),
.B1(n_1476),
.B2(n_1816),
.Y(n_2018)
);

INVx4_ASAP7_75t_L g2019 ( 
.A(n_1803),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1976),
.Y(n_2020)
);

OR2x2_ASAP7_75t_L g2021 ( 
.A(n_1912),
.B(n_1640),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1982),
.B(n_1696),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1715),
.Y(n_2023)
);

NOR2xp33_ASAP7_75t_L g2024 ( 
.A(n_1991),
.B(n_1641),
.Y(n_2024)
);

AOI22xp33_ASAP7_75t_L g2025 ( 
.A1(n_1999),
.A2(n_1476),
.B1(n_1581),
.B2(n_1698),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1976),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1988),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1988),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1989),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1989),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1793),
.B(n_1580),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1717),
.Y(n_2032)
);

AOI22xp5_ASAP7_75t_L g2033 ( 
.A1(n_1918),
.A2(n_1698),
.B1(n_1443),
.B2(n_1476),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1842),
.B(n_1641),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_SL g2035 ( 
.A(n_1771),
.B(n_1776),
.Y(n_2035)
);

INVx3_ASAP7_75t_L g2036 ( 
.A(n_1869),
.Y(n_2036)
);

NOR2xp33_ASAP7_75t_L g2037 ( 
.A(n_1737),
.B(n_1644),
.Y(n_2037)
);

AOI22xp33_ASAP7_75t_L g2038 ( 
.A1(n_1858),
.A2(n_1476),
.B1(n_1581),
.B2(n_1698),
.Y(n_2038)
);

INVx1_ASAP7_75t_SL g2039 ( 
.A(n_1965),
.Y(n_2039)
);

BUFx3_ASAP7_75t_L g2040 ( 
.A(n_1756),
.Y(n_2040)
);

INVx5_ASAP7_75t_L g2041 ( 
.A(n_1929),
.Y(n_2041)
);

AOI22xp33_ASAP7_75t_L g2042 ( 
.A1(n_1865),
.A2(n_1476),
.B1(n_1698),
.B2(n_1671),
.Y(n_2042)
);

OR2x6_ASAP7_75t_L g2043 ( 
.A(n_1770),
.B(n_1644),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_2000),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_SL g2045 ( 
.A(n_1771),
.B(n_1532),
.Y(n_2045)
);

AND2x6_ASAP7_75t_L g2046 ( 
.A(n_1727),
.B(n_1633),
.Y(n_2046)
);

BUFx2_ASAP7_75t_L g2047 ( 
.A(n_1781),
.Y(n_2047)
);

BUFx8_ASAP7_75t_SL g2048 ( 
.A(n_1732),
.Y(n_2048)
);

AND2x4_ASAP7_75t_L g2049 ( 
.A(n_1874),
.B(n_1514),
.Y(n_2049)
);

OAI22xp33_ASAP7_75t_L g2050 ( 
.A1(n_1821),
.A2(n_1646),
.B1(n_1470),
.B2(n_1530),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1842),
.B(n_1867),
.Y(n_2051)
);

INVx4_ASAP7_75t_L g2052 ( 
.A(n_1803),
.Y(n_2052)
);

NOR2xp33_ASAP7_75t_L g2053 ( 
.A(n_1764),
.B(n_1646),
.Y(n_2053)
);

NAND2xp33_ASAP7_75t_L g2054 ( 
.A(n_1767),
.B(n_1698),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_1717),
.Y(n_2055)
);

AOI22xp33_ASAP7_75t_L g2056 ( 
.A1(n_1860),
.A2(n_1476),
.B1(n_1893),
.B2(n_1866),
.Y(n_2056)
);

NOR2xp33_ASAP7_75t_L g2057 ( 
.A(n_1798),
.B(n_1443),
.Y(n_2057)
);

NAND2xp33_ASAP7_75t_L g2058 ( 
.A(n_1767),
.B(n_1627),
.Y(n_2058)
);

INVx2_ASAP7_75t_SL g2059 ( 
.A(n_1823),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2000),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1722),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_1722),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_1867),
.B(n_1710),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_2005),
.Y(n_2064)
);

AOI22xp5_ASAP7_75t_L g2065 ( 
.A1(n_1818),
.A2(n_1462),
.B1(n_1678),
.B2(n_1663),
.Y(n_2065)
);

NOR2xp33_ASAP7_75t_L g2066 ( 
.A(n_1908),
.B(n_1637),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1935),
.B(n_1458),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1776),
.B(n_1458),
.Y(n_2068)
);

NOR2xp33_ASAP7_75t_L g2069 ( 
.A(n_1820),
.B(n_1710),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1776),
.B(n_1590),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_1829),
.B(n_1602),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_1829),
.B(n_1659),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_1829),
.B(n_1671),
.Y(n_2073)
);

CKINVDCx20_ASAP7_75t_R g2074 ( 
.A(n_1719),
.Y(n_2074)
);

AOI22xp33_ASAP7_75t_L g2075 ( 
.A1(n_1860),
.A2(n_1671),
.B1(n_801),
.B2(n_818),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2005),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1733),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1733),
.Y(n_2078)
);

NOR2xp33_ASAP7_75t_L g2079 ( 
.A(n_1861),
.B(n_1653),
.Y(n_2079)
);

AOI22xp5_ASAP7_75t_L g2080 ( 
.A1(n_1930),
.A2(n_1663),
.B1(n_1678),
.B2(n_1606),
.Y(n_2080)
);

INVxp67_ASAP7_75t_L g2081 ( 
.A(n_1951),
.Y(n_2081)
);

INVx5_ASAP7_75t_L g2082 ( 
.A(n_1929),
.Y(n_2082)
);

INVx2_ASAP7_75t_SL g2083 ( 
.A(n_1828),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_SL g2084 ( 
.A(n_1768),
.B(n_1532),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1953),
.B(n_1596),
.Y(n_2085)
);

INVx2_ASAP7_75t_SL g2086 ( 
.A(n_1835),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1800),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1800),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1812),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_1953),
.B(n_1596),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1812),
.Y(n_2091)
);

AO22x2_ASAP7_75t_L g2092 ( 
.A1(n_1833),
.A2(n_1634),
.B1(n_1649),
.B2(n_818),
.Y(n_2092)
);

BUFx6f_ASAP7_75t_L g2093 ( 
.A(n_1929),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1824),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_SL g2095 ( 
.A(n_1768),
.B(n_1532),
.Y(n_2095)
);

NAND2xp33_ASAP7_75t_L g2096 ( 
.A(n_1769),
.B(n_1627),
.Y(n_2096)
);

NOR2xp33_ASAP7_75t_L g2097 ( 
.A(n_1773),
.B(n_1634),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1824),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1827),
.Y(n_2099)
);

NOR2xp33_ASAP7_75t_L g2100 ( 
.A(n_1744),
.B(n_1634),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1953),
.B(n_1596),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1872),
.B(n_1429),
.Y(n_2102)
);

BUFx2_ASAP7_75t_L g2103 ( 
.A(n_1783),
.Y(n_2103)
);

INVx5_ASAP7_75t_L g2104 ( 
.A(n_1929),
.Y(n_2104)
);

NOR2xp33_ASAP7_75t_L g2105 ( 
.A(n_1884),
.B(n_1649),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1827),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_SL g2107 ( 
.A(n_1769),
.B(n_1541),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_1872),
.B(n_1440),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_1832),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_SL g2110 ( 
.A(n_1780),
.B(n_1541),
.Y(n_2110)
);

AOI22xp33_ASAP7_75t_L g2111 ( 
.A1(n_1860),
.A2(n_1893),
.B1(n_1866),
.B2(n_1725),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_1882),
.B(n_1626),
.Y(n_2112)
);

INVx3_ASAP7_75t_L g2113 ( 
.A(n_1941),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1832),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1840),
.Y(n_2115)
);

AOI22xp33_ASAP7_75t_L g2116 ( 
.A1(n_1866),
.A2(n_1027),
.B1(n_1547),
.B2(n_921),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1840),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1847),
.Y(n_2118)
);

INVx1_ASAP7_75t_SL g2119 ( 
.A(n_1831),
.Y(n_2119)
);

AND2x4_ASAP7_75t_L g2120 ( 
.A(n_1739),
.B(n_1601),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_1847),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1873),
.Y(n_2122)
);

BUFx3_ASAP7_75t_L g2123 ( 
.A(n_1831),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1873),
.Y(n_2124)
);

INVx3_ASAP7_75t_L g2125 ( 
.A(n_1941),
.Y(n_2125)
);

INVx5_ASAP7_75t_L g2126 ( 
.A(n_1862),
.Y(n_2126)
);

INVx3_ASAP7_75t_L g2127 ( 
.A(n_1941),
.Y(n_2127)
);

AND2x4_ASAP7_75t_L g2128 ( 
.A(n_1754),
.B(n_1755),
.Y(n_2128)
);

NOR2xp33_ASAP7_75t_L g2129 ( 
.A(n_1907),
.B(n_1649),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_SL g2130 ( 
.A(n_1780),
.B(n_1541),
.Y(n_2130)
);

AND2x2_ASAP7_75t_SL g2131 ( 
.A(n_1883),
.B(n_1639),
.Y(n_2131)
);

NOR2xp33_ASAP7_75t_L g2132 ( 
.A(n_1752),
.B(n_1663),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_1882),
.B(n_1438),
.Y(n_2133)
);

INVx4_ASAP7_75t_L g2134 ( 
.A(n_1785),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1901),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_1909),
.B(n_1541),
.Y(n_2136)
);

BUFx3_ASAP7_75t_L g2137 ( 
.A(n_1757),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_1909),
.B(n_1678),
.Y(n_2138)
);

BUFx4f_ASAP7_75t_L g2139 ( 
.A(n_1834),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1901),
.Y(n_2140)
);

INVx2_ASAP7_75t_SL g2141 ( 
.A(n_1969),
.Y(n_2141)
);

BUFx3_ASAP7_75t_L g2142 ( 
.A(n_1763),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_SL g2143 ( 
.A(n_1787),
.B(n_1466),
.Y(n_2143)
);

BUFx3_ASAP7_75t_L g2144 ( 
.A(n_1721),
.Y(n_2144)
);

OAI21xp33_ASAP7_75t_SL g2145 ( 
.A1(n_1915),
.A2(n_1936),
.B(n_1924),
.Y(n_2145)
);

CKINVDCx5p33_ASAP7_75t_R g2146 ( 
.A(n_1724),
.Y(n_2146)
);

BUFx6f_ASAP7_75t_SL g2147 ( 
.A(n_1905),
.Y(n_2147)
);

NAND3xp33_ASAP7_75t_L g2148 ( 
.A(n_1980),
.B(n_1045),
.C(n_1041),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_1913),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_SL g2150 ( 
.A(n_1788),
.B(n_1466),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_1926),
.B(n_1496),
.Y(n_2151)
);

CKINVDCx5p33_ASAP7_75t_R g2152 ( 
.A(n_1726),
.Y(n_2152)
);

INVx2_ASAP7_75t_SL g2153 ( 
.A(n_1970),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1913),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_1926),
.B(n_1500),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_1759),
.B(n_1601),
.Y(n_2156)
);

NOR2xp33_ASAP7_75t_L g2157 ( 
.A(n_1836),
.B(n_1630),
.Y(n_2157)
);

INVx4_ASAP7_75t_L g2158 ( 
.A(n_1790),
.Y(n_2158)
);

BUFx3_ASAP7_75t_L g2159 ( 
.A(n_1740),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1914),
.Y(n_2160)
);

AND3x2_ASAP7_75t_L g2161 ( 
.A(n_1730),
.B(n_944),
.C(n_943),
.Y(n_2161)
);

BUFx6f_ASAP7_75t_L g2162 ( 
.A(n_1905),
.Y(n_2162)
);

XOR2xp5_ASAP7_75t_R g2163 ( 
.A(n_1765),
.B(n_1128),
.Y(n_2163)
);

CKINVDCx5p33_ASAP7_75t_R g2164 ( 
.A(n_1714),
.Y(n_2164)
);

INVx5_ASAP7_75t_L g2165 ( 
.A(n_1862),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_SL g2166 ( 
.A(n_1794),
.B(n_1795),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1914),
.Y(n_2167)
);

NAND2xp33_ASAP7_75t_L g2168 ( 
.A(n_1797),
.B(n_1627),
.Y(n_2168)
);

OR2x2_ASAP7_75t_L g2169 ( 
.A(n_1718),
.B(n_1250),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_1932),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_1716),
.B(n_1502),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_1875),
.B(n_1503),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_1888),
.B(n_1510),
.Y(n_2173)
);

INVx3_ASAP7_75t_L g2174 ( 
.A(n_1952),
.Y(n_2174)
);

INVx4_ASAP7_75t_SL g2175 ( 
.A(n_1862),
.Y(n_2175)
);

AOI22xp5_ASAP7_75t_L g2176 ( 
.A1(n_1864),
.A2(n_1945),
.B1(n_1940),
.B2(n_1927),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1932),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_1937),
.Y(n_2178)
);

OR2x6_ASAP7_75t_L g2179 ( 
.A(n_1925),
.B(n_1473),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1949),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_SL g2181 ( 
.A(n_1799),
.B(n_1466),
.Y(n_2181)
);

INVx4_ASAP7_75t_L g2182 ( 
.A(n_1801),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_SL g2183 ( 
.A(n_1802),
.B(n_1806),
.Y(n_2183)
);

INVx5_ASAP7_75t_L g2184 ( 
.A(n_1862),
.Y(n_2184)
);

INVx4_ASAP7_75t_L g2185 ( 
.A(n_1807),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1955),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1957),
.Y(n_2187)
);

BUFx6f_ASAP7_75t_L g2188 ( 
.A(n_1905),
.Y(n_2188)
);

INVx3_ASAP7_75t_L g2189 ( 
.A(n_1952),
.Y(n_2189)
);

BUFx3_ASAP7_75t_L g2190 ( 
.A(n_1740),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_1894),
.B(n_1511),
.Y(n_2191)
);

BUFx6f_ASAP7_75t_L g2192 ( 
.A(n_2001),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1967),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_1895),
.B(n_1518),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_1971),
.Y(n_2195)
);

AND2x6_ASAP7_75t_L g2196 ( 
.A(n_1727),
.B(n_1639),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_SL g2197 ( 
.A(n_1809),
.B(n_1811),
.Y(n_2197)
);

INVxp33_ASAP7_75t_L g2198 ( 
.A(n_2006),
.Y(n_2198)
);

AND2x4_ASAP7_75t_L g2199 ( 
.A(n_1758),
.B(n_1606),
.Y(n_2199)
);

INVx3_ASAP7_75t_L g2200 ( 
.A(n_1952),
.Y(n_2200)
);

NAND3xp33_ASAP7_75t_L g2201 ( 
.A(n_1980),
.B(n_1045),
.C(n_1041),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_1898),
.B(n_1520),
.Y(n_2202)
);

AOI22xp33_ASAP7_75t_L g2203 ( 
.A1(n_1893),
.A2(n_1486),
.B1(n_1516),
.B2(n_1488),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1974),
.Y(n_2204)
);

OR2x2_ASAP7_75t_L g2205 ( 
.A(n_1746),
.B(n_1657),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_1975),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_1978),
.Y(n_2207)
);

AND2x6_ASAP7_75t_L g2208 ( 
.A(n_1727),
.B(n_1508),
.Y(n_2208)
);

NAND3xp33_ASAP7_75t_L g2209 ( 
.A(n_1984),
.B(n_1237),
.C(n_1090),
.Y(n_2209)
);

CKINVDCx20_ASAP7_75t_R g2210 ( 
.A(n_1751),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1981),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1983),
.Y(n_2212)
);

BUFx6f_ASAP7_75t_L g2213 ( 
.A(n_2001),
.Y(n_2213)
);

NOR2xp33_ASAP7_75t_L g2214 ( 
.A(n_1845),
.B(n_1523),
.Y(n_2214)
);

BUFx10_ASAP7_75t_L g2215 ( 
.A(n_1720),
.Y(n_2215)
);

BUFx2_ASAP7_75t_L g2216 ( 
.A(n_1784),
.Y(n_2216)
);

NOR2xp33_ASAP7_75t_L g2217 ( 
.A(n_1984),
.B(n_1524),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_1987),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_1899),
.B(n_1533),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_1766),
.B(n_1535),
.Y(n_2220)
);

OR2x2_ASAP7_75t_L g2221 ( 
.A(n_1855),
.B(n_1081),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_1774),
.Y(n_2222)
);

CKINVDCx5p33_ASAP7_75t_R g2223 ( 
.A(n_1713),
.Y(n_2223)
);

INVx5_ASAP7_75t_L g2224 ( 
.A(n_1862),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1777),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_SL g2226 ( 
.A(n_1819),
.B(n_1466),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_1791),
.Y(n_2227)
);

AOI22xp33_ASAP7_75t_SL g2228 ( 
.A1(n_1900),
.A2(n_1097),
.B1(n_1055),
.B2(n_742),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_1792),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_1759),
.B(n_1760),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1804),
.Y(n_2231)
);

BUFx6f_ASAP7_75t_L g2232 ( 
.A(n_2001),
.Y(n_2232)
);

BUFx6f_ASAP7_75t_L g2233 ( 
.A(n_1977),
.Y(n_2233)
);

NOR2xp33_ASAP7_75t_L g2234 ( 
.A(n_1985),
.B(n_1539),
.Y(n_2234)
);

INVx3_ASAP7_75t_L g2235 ( 
.A(n_1977),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_1805),
.B(n_1545),
.Y(n_2236)
);

CKINVDCx5p33_ASAP7_75t_R g2237 ( 
.A(n_1713),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_1808),
.B(n_1548),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1810),
.Y(n_2239)
);

BUFx3_ASAP7_75t_L g2240 ( 
.A(n_1743),
.Y(n_2240)
);

BUFx10_ASAP7_75t_L g2241 ( 
.A(n_1723),
.Y(n_2241)
);

BUFx2_ASAP7_75t_L g2242 ( 
.A(n_1826),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_1815),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_SL g2244 ( 
.A(n_1985),
.B(n_1513),
.Y(n_2244)
);

NOR2xp33_ASAP7_75t_L g2245 ( 
.A(n_1986),
.B(n_1551),
.Y(n_2245)
);

AND2x6_ASAP7_75t_L g2246 ( 
.A(n_1735),
.B(n_1822),
.Y(n_2246)
);

INVx4_ASAP7_75t_L g2247 ( 
.A(n_1760),
.Y(n_2247)
);

INVx4_ASAP7_75t_L g2248 ( 
.A(n_1761),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_1825),
.Y(n_2249)
);

NOR2xp33_ASAP7_75t_L g2250 ( 
.A(n_1986),
.B(n_1556),
.Y(n_2250)
);

INVx2_ASAP7_75t_L g2251 ( 
.A(n_1843),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_1850),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_1852),
.B(n_1558),
.Y(n_2253)
);

NOR2xp33_ASAP7_75t_L g2254 ( 
.A(n_1992),
.B(n_1993),
.Y(n_2254)
);

AOI22xp33_ASAP7_75t_L g2255 ( 
.A1(n_1906),
.A2(n_1488),
.B1(n_1516),
.B2(n_1486),
.Y(n_2255)
);

AOI22xp33_ASAP7_75t_L g2256 ( 
.A1(n_1906),
.A2(n_1488),
.B1(n_1516),
.B2(n_1486),
.Y(n_2256)
);

AND2x6_ASAP7_75t_L g2257 ( 
.A(n_1735),
.B(n_1606),
.Y(n_2257)
);

AOI22xp33_ASAP7_75t_L g2258 ( 
.A1(n_1900),
.A2(n_1488),
.B1(n_1516),
.B2(n_1486),
.Y(n_2258)
);

INVx2_ASAP7_75t_L g2259 ( 
.A(n_1856),
.Y(n_2259)
);

AND2x2_ASAP7_75t_L g2260 ( 
.A(n_1761),
.B(n_1433),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1857),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_1977),
.Y(n_2262)
);

AOI22xp33_ASAP7_75t_L g2263 ( 
.A1(n_1735),
.A2(n_1488),
.B1(n_1516),
.B2(n_1486),
.Y(n_2263)
);

AND2x2_ASAP7_75t_L g2264 ( 
.A(n_1762),
.B(n_1433),
.Y(n_2264)
);

NOR2xp33_ASAP7_75t_SL g2265 ( 
.A(n_1723),
.B(n_1184),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_1762),
.B(n_1433),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_1997),
.Y(n_2267)
);

OR2x2_ASAP7_75t_L g2268 ( 
.A(n_1876),
.B(n_1081),
.Y(n_2268)
);

AND2x6_ASAP7_75t_L g2269 ( 
.A(n_1997),
.B(n_1487),
.Y(n_2269)
);

AND2x4_ASAP7_75t_L g2270 ( 
.A(n_1741),
.B(n_1487),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_1997),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_1859),
.B(n_1567),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_2002),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1992),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_SL g2275 ( 
.A(n_1993),
.B(n_1513),
.Y(n_2275)
);

INVx4_ASAP7_75t_L g2276 ( 
.A(n_1748),
.Y(n_2276)
);

AND2x4_ASAP7_75t_L g2277 ( 
.A(n_1871),
.B(n_1487),
.Y(n_2277)
);

CKINVDCx5p33_ASAP7_75t_R g2278 ( 
.A(n_1728),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_2002),
.Y(n_2279)
);

BUFx6f_ASAP7_75t_L g2280 ( 
.A(n_1789),
.Y(n_2280)
);

OR2x2_ASAP7_75t_L g2281 ( 
.A(n_1844),
.B(n_1090),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_SL g2282 ( 
.A(n_1994),
.B(n_1513),
.Y(n_2282)
);

AND2x6_ASAP7_75t_L g2283 ( 
.A(n_1996),
.B(n_1519),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_1972),
.B(n_1973),
.Y(n_2284)
);

OR2x2_ASAP7_75t_L g2285 ( 
.A(n_1729),
.B(n_1096),
.Y(n_2285)
);

BUFx6f_ASAP7_75t_L g2286 ( 
.A(n_1789),
.Y(n_2286)
);

INVx3_ASAP7_75t_L g2287 ( 
.A(n_1996),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_1994),
.Y(n_2288)
);

NOR2xp33_ASAP7_75t_L g2289 ( 
.A(n_1979),
.B(n_1571),
.Y(n_2289)
);

AOI22xp33_ASAP7_75t_L g2290 ( 
.A1(n_1890),
.A2(n_1488),
.B1(n_1516),
.B2(n_1486),
.Y(n_2290)
);

INVx4_ASAP7_75t_L g2291 ( 
.A(n_1748),
.Y(n_2291)
);

BUFx6f_ASAP7_75t_L g2292 ( 
.A(n_1749),
.Y(n_2292)
);

BUFx8_ASAP7_75t_SL g2293 ( 
.A(n_1736),
.Y(n_2293)
);

INVx2_ASAP7_75t_L g2294 ( 
.A(n_2002),
.Y(n_2294)
);

INVx3_ASAP7_75t_L g2295 ( 
.A(n_1996),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_1896),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_1879),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_1885),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_SL g2299 ( 
.A(n_1886),
.B(n_1513),
.Y(n_2299)
);

BUFx3_ASAP7_75t_L g2300 ( 
.A(n_1743),
.Y(n_2300)
);

INVx3_ASAP7_75t_L g2301 ( 
.A(n_1896),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_1922),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_2031),
.B(n_2013),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2180),
.Y(n_2304)
);

NOR2xp33_ASAP7_75t_L g2305 ( 
.A(n_2157),
.B(n_1923),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_2011),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2186),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_2067),
.B(n_1931),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2187),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_2133),
.B(n_1933),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_2102),
.B(n_1938),
.Y(n_2311)
);

INVxp67_ASAP7_75t_L g2312 ( 
.A(n_2284),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2193),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_2023),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_2032),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_2055),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2108),
.B(n_1942),
.Y(n_2317)
);

BUFx6f_ASAP7_75t_L g2318 ( 
.A(n_2292),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_SL g2319 ( 
.A(n_2080),
.B(n_1943),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_2017),
.B(n_1944),
.Y(n_2320)
);

INVx2_ASAP7_75t_L g2321 ( 
.A(n_2061),
.Y(n_2321)
);

INVx2_ASAP7_75t_SL g2322 ( 
.A(n_2047),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2204),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2211),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_2051),
.B(n_1947),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2022),
.B(n_1950),
.Y(n_2326)
);

NOR2xp33_ASAP7_75t_L g2327 ( 
.A(n_2157),
.B(n_1954),
.Y(n_2327)
);

BUFx5_ASAP7_75t_L g2328 ( 
.A(n_2246),
.Y(n_2328)
);

AND2x2_ASAP7_75t_L g2329 ( 
.A(n_2034),
.B(n_1851),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_2062),
.Y(n_2330)
);

AND2x2_ASAP7_75t_L g2331 ( 
.A(n_2063),
.B(n_2138),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_2068),
.B(n_1846),
.Y(n_2332)
);

NOR2xp33_ASAP7_75t_L g2333 ( 
.A(n_2254),
.B(n_1292),
.Y(n_2333)
);

AND2x2_ASAP7_75t_L g2334 ( 
.A(n_2230),
.B(n_2254),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_2112),
.B(n_1848),
.Y(n_2335)
);

INVx3_ASAP7_75t_L g2336 ( 
.A(n_2016),
.Y(n_2336)
);

INVx2_ASAP7_75t_L g2337 ( 
.A(n_2098),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2136),
.B(n_1849),
.Y(n_2338)
);

AND2x2_ASAP7_75t_L g2339 ( 
.A(n_2037),
.B(n_1853),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_2109),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_2121),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_2037),
.B(n_2151),
.Y(n_2342)
);

INVx2_ASAP7_75t_SL g2343 ( 
.A(n_2139),
.Y(n_2343)
);

BUFx5_ASAP7_75t_L g2344 ( 
.A(n_2246),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2155),
.B(n_1928),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_2024),
.B(n_2007),
.Y(n_2346)
);

INVx2_ASAP7_75t_SL g2347 ( 
.A(n_2139),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_SL g2348 ( 
.A(n_2065),
.B(n_1956),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_SL g2349 ( 
.A(n_2050),
.B(n_1958),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2212),
.Y(n_2350)
);

NOR2xp33_ASAP7_75t_L g2351 ( 
.A(n_2014),
.B(n_1292),
.Y(n_2351)
);

NOR2xp33_ASAP7_75t_L g2352 ( 
.A(n_2214),
.B(n_1293),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2149),
.Y(n_2353)
);

NAND2xp33_ASAP7_75t_L g2354 ( 
.A(n_2292),
.B(n_2162),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_2170),
.Y(n_2355)
);

BUFx3_ASAP7_75t_L g2356 ( 
.A(n_2137),
.Y(n_2356)
);

INVx2_ASAP7_75t_L g2357 ( 
.A(n_2008),
.Y(n_2357)
);

NAND2xp33_ASAP7_75t_L g2358 ( 
.A(n_2292),
.B(n_1749),
.Y(n_2358)
);

INVx2_ASAP7_75t_L g2359 ( 
.A(n_2009),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2020),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_2024),
.B(n_2004),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_2057),
.B(n_2004),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_2057),
.B(n_2007),
.Y(n_2363)
);

INVx4_ASAP7_75t_L g2364 ( 
.A(n_2162),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_2053),
.B(n_2003),
.Y(n_2365)
);

BUFx5_ASAP7_75t_L g2366 ( 
.A(n_2246),
.Y(n_2366)
);

NOR2xp33_ASAP7_75t_L g2367 ( 
.A(n_2214),
.B(n_1293),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_2050),
.B(n_2003),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2097),
.B(n_1863),
.Y(n_2369)
);

NAND2xp33_ASAP7_75t_L g2370 ( 
.A(n_2292),
.B(n_2162),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2097),
.B(n_1878),
.Y(n_2371)
);

NOR2xp33_ASAP7_75t_L g2372 ( 
.A(n_2274),
.B(n_1296),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_SL g2373 ( 
.A(n_2297),
.B(n_1959),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_2026),
.Y(n_2374)
);

BUFx3_ASAP7_75t_L g2375 ( 
.A(n_2137),
.Y(n_2375)
);

NOR2xp33_ASAP7_75t_R g2376 ( 
.A(n_2164),
.B(n_1728),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2027),
.Y(n_2377)
);

NOR2xp67_ASAP7_75t_L g2378 ( 
.A(n_2134),
.B(n_1731),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2100),
.B(n_1515),
.Y(n_2379)
);

AND2x4_ASAP7_75t_L g2380 ( 
.A(n_2120),
.B(n_1750),
.Y(n_2380)
);

A2O1A1Ixp33_ASAP7_75t_L g2381 ( 
.A1(n_2100),
.A2(n_1854),
.B(n_1917),
.C(n_1921),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_2132),
.B(n_1515),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_SL g2383 ( 
.A(n_2298),
.B(n_1960),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_2028),
.Y(n_2384)
);

AOI221xp5_ASAP7_75t_L g2385 ( 
.A1(n_2228),
.A2(n_1917),
.B1(n_1921),
.B2(n_1910),
.C(n_1890),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2029),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2030),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_SL g2388 ( 
.A(n_2141),
.B(n_1961),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2132),
.B(n_2217),
.Y(n_2389)
);

NAND2xp33_ASAP7_75t_L g2390 ( 
.A(n_2162),
.B(n_1750),
.Y(n_2390)
);

BUFx6f_ASAP7_75t_SL g2391 ( 
.A(n_2215),
.Y(n_2391)
);

NAND2xp33_ASAP7_75t_L g2392 ( 
.A(n_2188),
.B(n_1753),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_2217),
.B(n_2234),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_SL g2394 ( 
.A(n_2153),
.B(n_1962),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_2234),
.B(n_1576),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_2245),
.B(n_2250),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_2245),
.B(n_1578),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_2053),
.B(n_1778),
.Y(n_2398)
);

INVx1_ASAP7_75t_SL g2399 ( 
.A(n_2015),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2044),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_2060),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_SL g2402 ( 
.A(n_2260),
.B(n_1964),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2064),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_SL g2404 ( 
.A(n_2264),
.B(n_1968),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_SL g2405 ( 
.A(n_2266),
.B(n_1813),
.Y(n_2405)
);

BUFx2_ASAP7_75t_L g2406 ( 
.A(n_2123),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_2076),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2077),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_2250),
.B(n_1582),
.Y(n_2409)
);

AND2x4_ASAP7_75t_L g2410 ( 
.A(n_2120),
.B(n_1753),
.Y(n_2410)
);

NOR2xp33_ASAP7_75t_SL g2411 ( 
.A(n_2223),
.B(n_1731),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2078),
.Y(n_2412)
);

OR2x2_ASAP7_75t_L g2413 ( 
.A(n_2021),
.B(n_1817),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_2087),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2088),
.Y(n_2415)
);

INVx2_ASAP7_75t_SL g2416 ( 
.A(n_2043),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_2069),
.B(n_1584),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2089),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_L g2419 ( 
.A(n_2069),
.B(n_1587),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2178),
.B(n_1593),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_2195),
.B(n_1595),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2206),
.B(n_1611),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_2207),
.B(n_1614),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2091),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_SL g2425 ( 
.A(n_2302),
.B(n_1814),
.Y(n_2425)
);

AOI22xp33_ASAP7_75t_L g2426 ( 
.A1(n_2128),
.A2(n_1920),
.B1(n_1911),
.B2(n_1902),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2218),
.B(n_2171),
.Y(n_2427)
);

BUFx5_ASAP7_75t_L g2428 ( 
.A(n_2246),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_L g2429 ( 
.A(n_2172),
.B(n_1619),
.Y(n_2429)
);

BUFx6f_ASAP7_75t_L g2430 ( 
.A(n_2016),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2173),
.B(n_1517),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2094),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_2191),
.B(n_1517),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_SL g2434 ( 
.A(n_2176),
.B(n_1839),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_2099),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2111),
.B(n_1498),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2111),
.B(n_1498),
.Y(n_2437)
);

AND2x2_ASAP7_75t_L g2438 ( 
.A(n_2105),
.B(n_1779),
.Y(n_2438)
);

INVx2_ASAP7_75t_L g2439 ( 
.A(n_2106),
.Y(n_2439)
);

INVx6_ASAP7_75t_L g2440 ( 
.A(n_2215),
.Y(n_2440)
);

BUFx12f_ASAP7_75t_L g2441 ( 
.A(n_2241),
.Y(n_2441)
);

AOI22xp5_ASAP7_75t_L g2442 ( 
.A1(n_2105),
.A2(n_1995),
.B1(n_1948),
.B2(n_1892),
.Y(n_2442)
);

INVxp67_ASAP7_75t_L g2443 ( 
.A(n_2079),
.Y(n_2443)
);

NOR2xp33_ASAP7_75t_L g2444 ( 
.A(n_2288),
.B(n_2119),
.Y(n_2444)
);

INVx2_ASAP7_75t_SL g2445 ( 
.A(n_2043),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2114),
.Y(n_2446)
);

NOR2xp33_ASAP7_75t_L g2447 ( 
.A(n_2081),
.B(n_1296),
.Y(n_2447)
);

OAI22xp5_ASAP7_75t_L g2448 ( 
.A1(n_2018),
.A2(n_1911),
.B1(n_1920),
.B2(n_1902),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2115),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2117),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2118),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_SL g2452 ( 
.A(n_2129),
.B(n_1877),
.Y(n_2452)
);

AOI22xp5_ASAP7_75t_L g2453 ( 
.A1(n_2129),
.A2(n_1916),
.B1(n_1919),
.B2(n_1889),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2085),
.B(n_1498),
.Y(n_2454)
);

INVx2_ASAP7_75t_L g2455 ( 
.A(n_2122),
.Y(n_2455)
);

NAND2x1_ASAP7_75t_L g2456 ( 
.A(n_2093),
.B(n_1445),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2124),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2135),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2140),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2090),
.B(n_1501),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_SL g2461 ( 
.A(n_2247),
.B(n_1891),
.Y(n_2461)
);

NOR2xp33_ASAP7_75t_L g2462 ( 
.A(n_2081),
.B(n_1304),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_L g2463 ( 
.A(n_2101),
.B(n_1501),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_L g2464 ( 
.A(n_2018),
.B(n_1501),
.Y(n_2464)
);

O2A1O1Ixp5_ASAP7_75t_L g2465 ( 
.A1(n_2084),
.A2(n_1568),
.B(n_1585),
.C(n_1552),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2056),
.B(n_2075),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_2056),
.B(n_1552),
.Y(n_2467)
);

INVx2_ASAP7_75t_SL g2468 ( 
.A(n_2043),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2154),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2160),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_L g2471 ( 
.A(n_2075),
.B(n_1552),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2033),
.B(n_1568),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2167),
.Y(n_2473)
);

AND2x2_ASAP7_75t_L g2474 ( 
.A(n_2156),
.B(n_1782),
.Y(n_2474)
);

BUFx3_ASAP7_75t_L g2475 ( 
.A(n_2142),
.Y(n_2475)
);

OR2x2_ASAP7_75t_L g2476 ( 
.A(n_2221),
.B(n_1736),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_2177),
.B(n_1568),
.Y(n_2477)
);

INVx2_ASAP7_75t_L g2478 ( 
.A(n_2222),
.Y(n_2478)
);

NOR2xp33_ASAP7_75t_L g2479 ( 
.A(n_2289),
.B(n_1304),
.Y(n_2479)
);

OR2x6_ASAP7_75t_L g2480 ( 
.A(n_2123),
.B(n_1473),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_L g2481 ( 
.A(n_2070),
.B(n_1585),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_SL g2482 ( 
.A(n_2247),
.B(n_2248),
.Y(n_2482)
);

AND2x4_ASAP7_75t_L g2483 ( 
.A(n_2199),
.B(n_1745),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_2225),
.B(n_1585),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2227),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2229),
.Y(n_2486)
);

CKINVDCx5p33_ASAP7_75t_R g2487 ( 
.A(n_2048),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_2231),
.B(n_1492),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_SL g2489 ( 
.A(n_2248),
.B(n_2301),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_2239),
.B(n_1492),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2252),
.B(n_1494),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_2243),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_SL g2493 ( 
.A(n_2301),
.B(n_1745),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_L g2494 ( 
.A(n_2261),
.B(n_1494),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2249),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2251),
.Y(n_2496)
);

NOR2xp33_ASAP7_75t_L g2497 ( 
.A(n_2289),
.B(n_1317),
.Y(n_2497)
);

NOR2xp33_ASAP7_75t_L g2498 ( 
.A(n_2166),
.B(n_1317),
.Y(n_2498)
);

BUFx6f_ASAP7_75t_L g2499 ( 
.A(n_2016),
.Y(n_2499)
);

AOI22xp5_ASAP7_75t_L g2500 ( 
.A1(n_2270),
.A2(n_1910),
.B1(n_1904),
.B2(n_1903),
.Y(n_2500)
);

NOR2x1p5_ASAP7_75t_L g2501 ( 
.A(n_2134),
.B(n_1747),
.Y(n_2501)
);

INVx2_ASAP7_75t_L g2502 ( 
.A(n_2259),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_L g2503 ( 
.A(n_2072),
.B(n_1512),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_2073),
.B(n_1512),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_SL g2505 ( 
.A(n_2158),
.B(n_1747),
.Y(n_2505)
);

NOR3xp33_ASAP7_75t_L g2506 ( 
.A(n_2166),
.B(n_1738),
.C(n_1796),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_SL g2507 ( 
.A(n_2158),
.B(n_1772),
.Y(n_2507)
);

AND2x6_ASAP7_75t_L g2508 ( 
.A(n_2093),
.B(n_2280),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2220),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2236),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2145),
.B(n_1527),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_SL g2512 ( 
.A(n_2182),
.B(n_1775),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2238),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2194),
.B(n_1527),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_L g2515 ( 
.A(n_2202),
.B(n_1529),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_2262),
.Y(n_2516)
);

BUFx8_ASAP7_75t_L g2517 ( 
.A(n_2103),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2253),
.Y(n_2518)
);

AND2x2_ASAP7_75t_L g2519 ( 
.A(n_2066),
.B(n_1734),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_2219),
.B(n_1529),
.Y(n_2520)
);

INVxp67_ASAP7_75t_L g2521 ( 
.A(n_2079),
.Y(n_2521)
);

INVxp33_ASAP7_75t_L g2522 ( 
.A(n_2268),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_2283),
.B(n_1538),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_SL g2524 ( 
.A(n_2182),
.B(n_1786),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2128),
.Y(n_2525)
);

AOI22xp33_ASAP7_75t_L g2526 ( 
.A1(n_2092),
.A2(n_1887),
.B1(n_1904),
.B2(n_1903),
.Y(n_2526)
);

NOR2xp33_ASAP7_75t_L g2527 ( 
.A(n_2183),
.B(n_1340),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_SL g2528 ( 
.A(n_2185),
.B(n_1734),
.Y(n_2528)
);

AO221x1_ASAP7_75t_L g2529 ( 
.A1(n_2092),
.A2(n_1534),
.B1(n_813),
.B2(n_989),
.C(n_992),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2283),
.B(n_1538),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_2283),
.B(n_2126),
.Y(n_2531)
);

NOR2xp33_ASAP7_75t_L g2532 ( 
.A(n_2183),
.B(n_1340),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_SL g2533 ( 
.A(n_2185),
.B(n_1517),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_2113),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2267),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_SL g2536 ( 
.A(n_2270),
.B(n_1517),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2113),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_L g2538 ( 
.A(n_2283),
.B(n_1544),
.Y(n_2538)
);

OR2x2_ASAP7_75t_L g2539 ( 
.A(n_2039),
.B(n_1738),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_SL g2540 ( 
.A(n_2197),
.B(n_1897),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_2283),
.B(n_1544),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_L g2542 ( 
.A(n_2126),
.B(n_1550),
.Y(n_2542)
);

AND2x4_ASAP7_75t_L g2543 ( 
.A(n_2483),
.B(n_2199),
.Y(n_2543)
);

AND2x2_ASAP7_75t_L g2544 ( 
.A(n_2365),
.B(n_2339),
.Y(n_2544)
);

NAND2xp5_ASAP7_75t_SL g2545 ( 
.A(n_2305),
.B(n_2059),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2304),
.Y(n_2546)
);

AND2x6_ASAP7_75t_L g2547 ( 
.A(n_2525),
.B(n_2188),
.Y(n_2547)
);

AND2x2_ASAP7_75t_L g2548 ( 
.A(n_2325),
.B(n_2334),
.Y(n_2548)
);

AOI22xp5_ASAP7_75t_L g2549 ( 
.A1(n_2352),
.A2(n_1187),
.B1(n_1195),
.B2(n_1184),
.Y(n_2549)
);

AO22x2_ASAP7_75t_L g2550 ( 
.A1(n_2349),
.A2(n_2281),
.B1(n_2244),
.B2(n_2275),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2303),
.B(n_2197),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_2303),
.B(n_2066),
.Y(n_2552)
);

INVx2_ASAP7_75t_SL g2553 ( 
.A(n_2356),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2307),
.Y(n_2554)
);

HB1xp67_ASAP7_75t_L g2555 ( 
.A(n_2322),
.Y(n_2555)
);

AOI22xp5_ASAP7_75t_L g2556 ( 
.A1(n_2367),
.A2(n_1195),
.B1(n_1203),
.B2(n_1187),
.Y(n_2556)
);

NAND2x1p5_ASAP7_75t_L g2557 ( 
.A(n_2318),
.B(n_2019),
.Y(n_2557)
);

INVx2_ASAP7_75t_L g2558 ( 
.A(n_2357),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2309),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2313),
.Y(n_2560)
);

INVx2_ASAP7_75t_L g2561 ( 
.A(n_2359),
.Y(n_2561)
);

AND2x2_ASAP7_75t_L g2562 ( 
.A(n_2329),
.B(n_2131),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2323),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2324),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_2342),
.B(n_2299),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2350),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2389),
.B(n_2299),
.Y(n_2567)
);

INVx2_ASAP7_75t_L g2568 ( 
.A(n_2374),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_L g2569 ( 
.A(n_2393),
.B(n_2296),
.Y(n_2569)
);

AOI22xp5_ASAP7_75t_L g2570 ( 
.A1(n_2327),
.A2(n_1203),
.B1(n_2265),
.B2(n_1365),
.Y(n_2570)
);

BUFx3_ASAP7_75t_L g2571 ( 
.A(n_2406),
.Y(n_2571)
);

AO22x2_ASAP7_75t_L g2572 ( 
.A1(n_2448),
.A2(n_2282),
.B1(n_2275),
.B2(n_2244),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_SL g2573 ( 
.A(n_2398),
.B(n_2083),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2485),
.Y(n_2574)
);

INVx3_ASAP7_75t_L g2575 ( 
.A(n_2318),
.Y(n_2575)
);

AO22x2_ASAP7_75t_L g2576 ( 
.A1(n_2396),
.A2(n_2282),
.B1(n_2285),
.B2(n_2095),
.Y(n_2576)
);

NOR2xp33_ASAP7_75t_L g2577 ( 
.A(n_2362),
.B(n_1128),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2509),
.B(n_2086),
.Y(n_2578)
);

AND2x4_ASAP7_75t_L g2579 ( 
.A(n_2483),
.B(n_2159),
.Y(n_2579)
);

NOR2xp33_ASAP7_75t_L g2580 ( 
.A(n_2363),
.B(n_1134),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2486),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_L g2582 ( 
.A(n_2510),
.B(n_2131),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_L g2583 ( 
.A(n_2513),
.B(n_2092),
.Y(n_2583)
);

INVx2_ASAP7_75t_L g2584 ( 
.A(n_2384),
.Y(n_2584)
);

AND2x2_ASAP7_75t_L g2585 ( 
.A(n_2331),
.B(n_2159),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_L g2586 ( 
.A(n_2518),
.B(n_2116),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2360),
.Y(n_2587)
);

AO22x2_ASAP7_75t_L g2588 ( 
.A1(n_2368),
.A2(n_2348),
.B1(n_2319),
.B2(n_2434),
.Y(n_2588)
);

NOR2xp33_ASAP7_75t_L g2589 ( 
.A(n_2311),
.B(n_1134),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2377),
.Y(n_2590)
);

OR2x2_ASAP7_75t_L g2591 ( 
.A(n_2311),
.B(n_2216),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2386),
.Y(n_2592)
);

AO22x2_ASAP7_75t_L g2593 ( 
.A1(n_2346),
.A2(n_2361),
.B1(n_2308),
.B2(n_2335),
.Y(n_2593)
);

CKINVDCx20_ASAP7_75t_R g2594 ( 
.A(n_2376),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_L g2595 ( 
.A(n_2310),
.B(n_2116),
.Y(n_2595)
);

BUFx6f_ASAP7_75t_L g2596 ( 
.A(n_2318),
.Y(n_2596)
);

INVx2_ASAP7_75t_L g2597 ( 
.A(n_2401),
.Y(n_2597)
);

NAND2x1p5_ASAP7_75t_L g2598 ( 
.A(n_2364),
.B(n_2019),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_L g2599 ( 
.A(n_2310),
.B(n_2276),
.Y(n_2599)
);

A2O1A1Ixp33_ASAP7_75t_L g2600 ( 
.A1(n_2345),
.A2(n_2054),
.B(n_2209),
.C(n_2038),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2387),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2400),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2403),
.Y(n_2603)
);

AO22x2_ASAP7_75t_L g2604 ( 
.A1(n_2308),
.A2(n_2095),
.B1(n_2107),
.B2(n_2084),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2408),
.Y(n_2605)
);

INVx2_ASAP7_75t_L g2606 ( 
.A(n_2407),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2412),
.Y(n_2607)
);

AO22x2_ASAP7_75t_L g2608 ( 
.A1(n_2335),
.A2(n_2110),
.B1(n_2130),
.B2(n_2107),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_2317),
.B(n_2276),
.Y(n_2609)
);

AO22x2_ASAP7_75t_L g2610 ( 
.A1(n_2317),
.A2(n_2130),
.B1(n_2110),
.B2(n_2148),
.Y(n_2610)
);

AO22x2_ASAP7_75t_L g2611 ( 
.A1(n_2332),
.A2(n_2201),
.B1(n_2295),
.B2(n_2287),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2415),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_2395),
.B(n_2291),
.Y(n_2613)
);

CKINVDCx20_ASAP7_75t_R g2614 ( 
.A(n_2487),
.Y(n_2614)
);

AOI22xp5_ASAP7_75t_L g2615 ( 
.A1(n_2479),
.A2(n_1365),
.B1(n_1369),
.B2(n_1353),
.Y(n_2615)
);

OAI221xp5_ASAP7_75t_L g2616 ( 
.A1(n_2385),
.A2(n_2228),
.B1(n_2169),
.B2(n_1887),
.C(n_978),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_2397),
.B(n_2291),
.Y(n_2617)
);

INVxp67_ASAP7_75t_L g2618 ( 
.A(n_2444),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2418),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2424),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_L g2621 ( 
.A(n_2409),
.B(n_2049),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2414),
.Y(n_2622)
);

AO22x2_ASAP7_75t_L g2623 ( 
.A1(n_2332),
.A2(n_2295),
.B1(n_2287),
.B2(n_2150),
.Y(n_2623)
);

AO22x2_ASAP7_75t_L g2624 ( 
.A1(n_2452),
.A2(n_2150),
.B1(n_2181),
.B2(n_2143),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2432),
.Y(n_2625)
);

BUFx6f_ASAP7_75t_L g2626 ( 
.A(n_2375),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2446),
.Y(n_2627)
);

AND2x2_ASAP7_75t_L g2628 ( 
.A(n_2438),
.B(n_2190),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2449),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2450),
.Y(n_2630)
);

NAND2x1p5_ASAP7_75t_L g2631 ( 
.A(n_2364),
.B(n_2052),
.Y(n_2631)
);

OAI21xp33_ASAP7_75t_L g2632 ( 
.A1(n_2497),
.A2(n_2198),
.B(n_1267),
.Y(n_2632)
);

NOR2xp33_ASAP7_75t_L g2633 ( 
.A(n_2369),
.B(n_1139),
.Y(n_2633)
);

AO22x2_ASAP7_75t_L g2634 ( 
.A1(n_2519),
.A2(n_2181),
.B1(n_2226),
.B2(n_2143),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2451),
.Y(n_2635)
);

AO22x2_ASAP7_75t_L g2636 ( 
.A1(n_2338),
.A2(n_2226),
.B1(n_2012),
.B2(n_2205),
.Y(n_2636)
);

A2O1A1Ixp33_ASAP7_75t_L g2637 ( 
.A1(n_2381),
.A2(n_2038),
.B(n_2071),
.C(n_2025),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2457),
.Y(n_2638)
);

AND2x2_ASAP7_75t_L g2639 ( 
.A(n_2474),
.B(n_2190),
.Y(n_2639)
);

AO22x2_ASAP7_75t_L g2640 ( 
.A1(n_2338),
.A2(n_2012),
.B1(n_2279),
.B2(n_2273),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_L g2641 ( 
.A(n_2427),
.B(n_2049),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2435),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_L g2643 ( 
.A(n_2443),
.B(n_2240),
.Y(n_2643)
);

AND2x4_ASAP7_75t_L g2644 ( 
.A(n_2380),
.B(n_2240),
.Y(n_2644)
);

AO22x2_ASAP7_75t_L g2645 ( 
.A1(n_2529),
.A2(n_2012),
.B1(n_2294),
.B2(n_2175),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2458),
.Y(n_2646)
);

BUFx8_ASAP7_75t_L g2647 ( 
.A(n_2391),
.Y(n_2647)
);

OAI22xp5_ASAP7_75t_L g2648 ( 
.A1(n_2526),
.A2(n_2025),
.B1(n_2042),
.B2(n_2179),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2469),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_L g2650 ( 
.A(n_2521),
.B(n_2300),
.Y(n_2650)
);

INVx2_ASAP7_75t_SL g2651 ( 
.A(n_2475),
.Y(n_2651)
);

AO22x2_ASAP7_75t_L g2652 ( 
.A1(n_2540),
.A2(n_2175),
.B1(n_2052),
.B2(n_2163),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2470),
.Y(n_2653)
);

AND2x4_ASAP7_75t_L g2654 ( 
.A(n_2380),
.B(n_2300),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_L g2655 ( 
.A(n_2417),
.B(n_2272),
.Y(n_2655)
);

BUFx3_ASAP7_75t_L g2656 ( 
.A(n_2440),
.Y(n_2656)
);

AND2x4_ASAP7_75t_L g2657 ( 
.A(n_2410),
.B(n_2179),
.Y(n_2657)
);

INVxp67_ASAP7_75t_L g2658 ( 
.A(n_2413),
.Y(n_2658)
);

HB1xp67_ASAP7_75t_L g2659 ( 
.A(n_2399),
.Y(n_2659)
);

CKINVDCx5p33_ASAP7_75t_R g2660 ( 
.A(n_2391),
.Y(n_2660)
);

BUFx8_ASAP7_75t_L g2661 ( 
.A(n_2441),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2473),
.Y(n_2662)
);

NAND2x1p5_ASAP7_75t_L g2663 ( 
.A(n_2430),
.B(n_2188),
.Y(n_2663)
);

AND2x4_ASAP7_75t_L g2664 ( 
.A(n_2410),
.B(n_2179),
.Y(n_2664)
);

AO22x2_ASAP7_75t_L g2665 ( 
.A1(n_2371),
.A2(n_2175),
.B1(n_2277),
.B2(n_2161),
.Y(n_2665)
);

OR2x6_ASAP7_75t_L g2666 ( 
.A(n_2440),
.B(n_2142),
.Y(n_2666)
);

AOI22xp5_ASAP7_75t_L g2667 ( 
.A1(n_2333),
.A2(n_1369),
.B1(n_1375),
.B2(n_1353),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_L g2668 ( 
.A(n_2419),
.B(n_2382),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2439),
.Y(n_2669)
);

INVx3_ASAP7_75t_L g2670 ( 
.A(n_2440),
.Y(n_2670)
);

AOI22xp5_ASAP7_75t_L g2671 ( 
.A1(n_2498),
.A2(n_1387),
.B1(n_1395),
.B2(n_1375),
.Y(n_2671)
);

INVx2_ASAP7_75t_SL g2672 ( 
.A(n_2343),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_L g2673 ( 
.A(n_2320),
.B(n_2161),
.Y(n_2673)
);

INVxp67_ASAP7_75t_L g2674 ( 
.A(n_2351),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2455),
.Y(n_2675)
);

OAI221xp5_ASAP7_75t_L g2676 ( 
.A1(n_2326),
.A2(n_1022),
.B1(n_1830),
.B2(n_1998),
.C(n_1837),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2459),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2495),
.Y(n_2678)
);

NOR2xp33_ASAP7_75t_L g2679 ( 
.A(n_2326),
.B(n_2320),
.Y(n_2679)
);

NOR2xp67_ASAP7_75t_L g2680 ( 
.A(n_2312),
.B(n_2237),
.Y(n_2680)
);

NOR2xp33_ASAP7_75t_L g2681 ( 
.A(n_2447),
.B(n_1139),
.Y(n_2681)
);

BUFx8_ASAP7_75t_L g2682 ( 
.A(n_2347),
.Y(n_2682)
);

AO22x2_ASAP7_75t_L g2683 ( 
.A1(n_2466),
.A2(n_2277),
.B1(n_2144),
.B2(n_1083),
.Y(n_2683)
);

AO22x2_ASAP7_75t_L g2684 ( 
.A1(n_2466),
.A2(n_2144),
.B1(n_728),
.B2(n_2271),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2496),
.Y(n_2685)
);

INVxp67_ASAP7_75t_L g2686 ( 
.A(n_2411),
.Y(n_2686)
);

AOI22xp5_ASAP7_75t_SL g2687 ( 
.A1(n_2372),
.A2(n_1162),
.B1(n_1169),
.B2(n_1156),
.Y(n_2687)
);

AOI22xp5_ASAP7_75t_L g2688 ( 
.A1(n_2527),
.A2(n_1395),
.B1(n_1396),
.B2(n_1387),
.Y(n_2688)
);

AOI22xp33_ASAP7_75t_L g2689 ( 
.A1(n_2506),
.A2(n_1998),
.B1(n_1519),
.B2(n_1742),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2488),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2488),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2490),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2429),
.B(n_2278),
.Y(n_2693)
);

AOI22xp5_ASAP7_75t_L g2694 ( 
.A1(n_2532),
.A2(n_2462),
.B1(n_1399),
.B2(n_1412),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2490),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2491),
.Y(n_2696)
);

AND2x4_ASAP7_75t_L g2697 ( 
.A(n_2501),
.B(n_2188),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2491),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2494),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2494),
.Y(n_2700)
);

AND2x4_ASAP7_75t_L g2701 ( 
.A(n_2416),
.B(n_2192),
.Y(n_2701)
);

NAND2xp33_ASAP7_75t_L g2702 ( 
.A(n_2508),
.B(n_2192),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2306),
.Y(n_2703)
);

AO22x2_ASAP7_75t_L g2704 ( 
.A1(n_2445),
.A2(n_2010),
.B1(n_2045),
.B2(n_1097),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_L g2705 ( 
.A(n_2379),
.B(n_2192),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_L g2706 ( 
.A(n_2514),
.B(n_2192),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2314),
.Y(n_2707)
);

AOI22xp5_ASAP7_75t_L g2708 ( 
.A1(n_2453),
.A2(n_1399),
.B1(n_1412),
.B2(n_1396),
.Y(n_2708)
);

CKINVDCx5p33_ASAP7_75t_R g2709 ( 
.A(n_2517),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_2514),
.B(n_2213),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2315),
.Y(n_2711)
);

AO22x2_ASAP7_75t_L g2712 ( 
.A1(n_2468),
.A2(n_2045),
.B1(n_2010),
.B2(n_2040),
.Y(n_2712)
);

AND2x2_ASAP7_75t_L g2713 ( 
.A(n_2426),
.B(n_2198),
.Y(n_2713)
);

OAI221xp5_ASAP7_75t_L g2714 ( 
.A1(n_2500),
.A2(n_1837),
.B1(n_1096),
.B2(n_1107),
.C(n_1106),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2316),
.Y(n_2715)
);

BUFx8_ASAP7_75t_L g2716 ( 
.A(n_2539),
.Y(n_2716)
);

HB1xp67_ASAP7_75t_L g2717 ( 
.A(n_2480),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2321),
.Y(n_2718)
);

INVxp67_ASAP7_75t_L g2719 ( 
.A(n_2373),
.Y(n_2719)
);

AO22x2_ASAP7_75t_L g2720 ( 
.A1(n_2471),
.A2(n_2035),
.B1(n_2127),
.B2(n_2125),
.Y(n_2720)
);

INVx2_ASAP7_75t_L g2721 ( 
.A(n_2330),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2337),
.Y(n_2722)
);

BUFx8_ASAP7_75t_L g2723 ( 
.A(n_2476),
.Y(n_2723)
);

AO22x2_ASAP7_75t_L g2724 ( 
.A1(n_2471),
.A2(n_2035),
.B1(n_2127),
.B2(n_2125),
.Y(n_2724)
);

AO22x2_ASAP7_75t_L g2725 ( 
.A1(n_2472),
.A2(n_2174),
.B1(n_2200),
.B2(n_2189),
.Y(n_2725)
);

BUFx3_ASAP7_75t_L g2726 ( 
.A(n_2517),
.Y(n_2726)
);

INVx2_ASAP7_75t_L g2727 ( 
.A(n_2340),
.Y(n_2727)
);

AND2x2_ASAP7_75t_L g2728 ( 
.A(n_2442),
.B(n_2242),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2341),
.Y(n_2729)
);

AND2x4_ASAP7_75t_L g2730 ( 
.A(n_2480),
.B(n_2213),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2353),
.Y(n_2731)
);

CKINVDCx20_ASAP7_75t_R g2732 ( 
.A(n_2388),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2355),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2478),
.Y(n_2734)
);

AND2x4_ASAP7_75t_L g2735 ( 
.A(n_2480),
.B(n_2213),
.Y(n_2735)
);

OAI221xp5_ASAP7_75t_L g2736 ( 
.A1(n_2383),
.A2(n_1100),
.B1(n_1108),
.B2(n_1107),
.C(n_1106),
.Y(n_2736)
);

AND2x2_ASAP7_75t_L g2737 ( 
.A(n_2544),
.B(n_2492),
.Y(n_2737)
);

AND2x2_ASAP7_75t_SL g2738 ( 
.A(n_2702),
.B(n_2354),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_L g2739 ( 
.A(n_2552),
.B(n_2515),
.Y(n_2739)
);

AND2x2_ASAP7_75t_L g2740 ( 
.A(n_2548),
.B(n_2502),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_L g2741 ( 
.A(n_2679),
.B(n_2515),
.Y(n_2741)
);

AOI21xp5_ASAP7_75t_L g2742 ( 
.A1(n_2655),
.A2(n_2165),
.B(n_2126),
.Y(n_2742)
);

INVx5_ASAP7_75t_L g2743 ( 
.A(n_2547),
.Y(n_2743)
);

BUFx2_ASAP7_75t_L g2744 ( 
.A(n_2659),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_L g2745 ( 
.A(n_2551),
.B(n_2520),
.Y(n_2745)
);

OAI22xp5_ASAP7_75t_L g2746 ( 
.A1(n_2618),
.A2(n_2394),
.B1(n_2378),
.B2(n_2522),
.Y(n_2746)
);

AOI21xp5_ASAP7_75t_L g2747 ( 
.A1(n_2668),
.A2(n_2165),
.B(n_2126),
.Y(n_2747)
);

INVx2_ASAP7_75t_L g2748 ( 
.A(n_2558),
.Y(n_2748)
);

AOI21xp5_ASAP7_75t_L g2749 ( 
.A1(n_2637),
.A2(n_2184),
.B(n_2165),
.Y(n_2749)
);

AND2x2_ASAP7_75t_L g2750 ( 
.A(n_2562),
.B(n_1519),
.Y(n_2750)
);

NOR2xp67_ASAP7_75t_L g2751 ( 
.A(n_2670),
.B(n_2146),
.Y(n_2751)
);

AOI21xp5_ASAP7_75t_L g2752 ( 
.A1(n_2600),
.A2(n_2184),
.B(n_2165),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_2693),
.B(n_2520),
.Y(n_2753)
);

BUFx6f_ASAP7_75t_L g2754 ( 
.A(n_2656),
.Y(n_2754)
);

INVx2_ASAP7_75t_L g2755 ( 
.A(n_2561),
.Y(n_2755)
);

AOI21xp5_ASAP7_75t_L g2756 ( 
.A1(n_2613),
.A2(n_2224),
.B(n_2184),
.Y(n_2756)
);

A2O1A1Ixp33_ASAP7_75t_L g2757 ( 
.A1(n_2595),
.A2(n_2425),
.B(n_2370),
.C(n_2405),
.Y(n_2757)
);

AO22x1_ASAP7_75t_L g2758 ( 
.A1(n_2723),
.A2(n_2152),
.B1(n_1108),
.B2(n_1110),
.Y(n_2758)
);

AOI21xp5_ASAP7_75t_L g2759 ( 
.A1(n_2617),
.A2(n_2224),
.B(n_2184),
.Y(n_2759)
);

A2O1A1Ixp33_ASAP7_75t_L g2760 ( 
.A1(n_2586),
.A2(n_2420),
.B(n_2422),
.C(n_2421),
.Y(n_2760)
);

BUFx6f_ASAP7_75t_L g2761 ( 
.A(n_2596),
.Y(n_2761)
);

AOI21xp5_ASAP7_75t_L g2762 ( 
.A1(n_2565),
.A2(n_2224),
.B(n_2096),
.Y(n_2762)
);

OAI21xp5_ASAP7_75t_L g2763 ( 
.A1(n_2567),
.A2(n_2472),
.B(n_2465),
.Y(n_2763)
);

AOI21xp5_ASAP7_75t_L g2764 ( 
.A1(n_2648),
.A2(n_2224),
.B(n_2058),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2568),
.Y(n_2765)
);

NOR3xp33_ASAP7_75t_L g2766 ( 
.A(n_2632),
.B(n_2404),
.C(n_2402),
.Y(n_2766)
);

AOI21xp5_ASAP7_75t_L g2767 ( 
.A1(n_2706),
.A2(n_2168),
.B(n_2531),
.Y(n_2767)
);

OAI21xp5_ASAP7_75t_L g2768 ( 
.A1(n_2583),
.A2(n_2464),
.B(n_2511),
.Y(n_2768)
);

AOI21xp5_ASAP7_75t_L g2769 ( 
.A1(n_2710),
.A2(n_2531),
.B(n_2042),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2569),
.B(n_2493),
.Y(n_2770)
);

NOR2xp33_ASAP7_75t_SL g2771 ( 
.A(n_2616),
.B(n_1742),
.Y(n_2771)
);

INVx2_ASAP7_75t_L g2772 ( 
.A(n_2584),
.Y(n_2772)
);

A2O1A1Ixp33_ASAP7_75t_L g2773 ( 
.A1(n_2599),
.A2(n_2423),
.B(n_2461),
.C(n_2358),
.Y(n_2773)
);

O2A1O1Ixp33_ASAP7_75t_L g2774 ( 
.A1(n_2676),
.A2(n_2714),
.B(n_2609),
.C(n_2736),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2546),
.Y(n_2775)
);

AOI22xp5_ASAP7_75t_L g2776 ( 
.A1(n_2633),
.A2(n_1162),
.B1(n_1169),
.B2(n_1156),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_L g2777 ( 
.A(n_2621),
.B(n_2505),
.Y(n_2777)
);

AO21x1_ASAP7_75t_L g2778 ( 
.A1(n_2705),
.A2(n_2511),
.B(n_2464),
.Y(n_2778)
);

AOI22xp5_ASAP7_75t_L g2779 ( 
.A1(n_2577),
.A2(n_1177),
.B1(n_1423),
.B2(n_1419),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_L g2780 ( 
.A(n_2580),
.B(n_2528),
.Y(n_2780)
);

AOI21xp5_ASAP7_75t_L g2781 ( 
.A1(n_2588),
.A2(n_2481),
.B(n_2503),
.Y(n_2781)
);

BUFx6f_ASAP7_75t_L g2782 ( 
.A(n_2596),
.Y(n_2782)
);

AOI221xp5_ASAP7_75t_L g2783 ( 
.A1(n_2588),
.A2(n_1534),
.B1(n_1110),
.B2(n_1100),
.C(n_928),
.Y(n_2783)
);

OAI22xp5_ASAP7_75t_L g2784 ( 
.A1(n_2582),
.A2(n_2437),
.B1(n_2436),
.B2(n_2467),
.Y(n_2784)
);

BUFx3_ASAP7_75t_L g2785 ( 
.A(n_2626),
.Y(n_2785)
);

AOI33xp33_ASAP7_75t_L g2786 ( 
.A1(n_2694),
.A2(n_1086),
.A3(n_1089),
.B1(n_1087),
.B2(n_1082),
.B3(n_1078),
.Y(n_2786)
);

NOR2xp67_ASAP7_75t_SL g2787 ( 
.A(n_2726),
.B(n_2507),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2554),
.Y(n_2788)
);

OAI21x1_ASAP7_75t_L g2789 ( 
.A1(n_2690),
.A2(n_2504),
.B(n_2503),
.Y(n_2789)
);

AOI21xp5_ASAP7_75t_L g2790 ( 
.A1(n_2593),
.A2(n_2481),
.B(n_2504),
.Y(n_2790)
);

AOI21xp5_ASAP7_75t_L g2791 ( 
.A1(n_2593),
.A2(n_2530),
.B(n_2523),
.Y(n_2791)
);

BUFx6f_ASAP7_75t_L g2792 ( 
.A(n_2626),
.Y(n_2792)
);

AOI21xp5_ASAP7_75t_L g2793 ( 
.A1(n_2608),
.A2(n_2530),
.B(n_2523),
.Y(n_2793)
);

AOI21xp5_ASAP7_75t_L g2794 ( 
.A1(n_2608),
.A2(n_2541),
.B(n_2538),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_2589),
.B(n_2512),
.Y(n_2795)
);

NOR2x1_ASAP7_75t_L g2796 ( 
.A(n_2545),
.B(n_2524),
.Y(n_2796)
);

AOI21xp5_ASAP7_75t_L g2797 ( 
.A1(n_2604),
.A2(n_2541),
.B(n_2538),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2559),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_2674),
.B(n_2431),
.Y(n_2799)
);

AOI21xp5_ASAP7_75t_L g2800 ( 
.A1(n_2604),
.A2(n_2392),
.B(n_2390),
.Y(n_2800)
);

AOI221xp5_ASAP7_75t_L g2801 ( 
.A1(n_2684),
.A2(n_1423),
.B1(n_1419),
.B2(n_1990),
.C(n_1946),
.Y(n_2801)
);

NOR2xp33_ASAP7_75t_L g2802 ( 
.A(n_2681),
.B(n_1177),
.Y(n_2802)
);

AOI21xp5_ASAP7_75t_L g2803 ( 
.A1(n_2691),
.A2(n_2437),
.B(n_2436),
.Y(n_2803)
);

CKINVDCx8_ASAP7_75t_R g2804 ( 
.A(n_2709),
.Y(n_2804)
);

CKINVDCx20_ASAP7_75t_R g2805 ( 
.A(n_2614),
.Y(n_2805)
);

AOI21xp5_ASAP7_75t_L g2806 ( 
.A1(n_2692),
.A2(n_2433),
.B(n_2454),
.Y(n_2806)
);

INVx2_ASAP7_75t_L g2807 ( 
.A(n_2597),
.Y(n_2807)
);

OAI22xp5_ASAP7_75t_L g2808 ( 
.A1(n_2689),
.A2(n_2467),
.B1(n_2484),
.B2(n_2482),
.Y(n_2808)
);

OAI21xp5_ASAP7_75t_L g2809 ( 
.A1(n_2695),
.A2(n_2460),
.B(n_2454),
.Y(n_2809)
);

AOI21xp5_ASAP7_75t_L g2810 ( 
.A1(n_2696),
.A2(n_2463),
.B(n_2460),
.Y(n_2810)
);

AOI21xp5_ASAP7_75t_L g2811 ( 
.A1(n_2698),
.A2(n_2463),
.B(n_2082),
.Y(n_2811)
);

NAND2x1p5_ASAP7_75t_L g2812 ( 
.A(n_2730),
.B(n_2213),
.Y(n_2812)
);

AO21x1_ASAP7_75t_L g2813 ( 
.A1(n_2673),
.A2(n_2533),
.B(n_2542),
.Y(n_2813)
);

OAI22xp5_ASAP7_75t_L g2814 ( 
.A1(n_2699),
.A2(n_2484),
.B1(n_2489),
.B2(n_2255),
.Y(n_2814)
);

INVx2_ASAP7_75t_L g2815 ( 
.A(n_2606),
.Y(n_2815)
);

O2A1O1Ixp5_ASAP7_75t_L g2816 ( 
.A1(n_2573),
.A2(n_2536),
.B(n_2542),
.C(n_2477),
.Y(n_2816)
);

BUFx3_ASAP7_75t_L g2817 ( 
.A(n_2571),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_2578),
.B(n_2241),
.Y(n_2818)
);

AOI21xp5_ASAP7_75t_L g2819 ( 
.A1(n_2700),
.A2(n_2082),
.B(n_2041),
.Y(n_2819)
);

OAI22xp5_ASAP7_75t_L g2820 ( 
.A1(n_2570),
.A2(n_1841),
.B1(n_1742),
.B2(n_1868),
.Y(n_2820)
);

OAI22xp33_ASAP7_75t_L g2821 ( 
.A1(n_2615),
.A2(n_1239),
.B1(n_1246),
.B2(n_1233),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2560),
.Y(n_2822)
);

INVx2_ASAP7_75t_L g2823 ( 
.A(n_2622),
.Y(n_2823)
);

AOI22xp5_ASAP7_75t_L g2824 ( 
.A1(n_2549),
.A2(n_1870),
.B1(n_1881),
.B2(n_1838),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2563),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2564),
.Y(n_2826)
);

OAI21xp5_ASAP7_75t_L g2827 ( 
.A1(n_2641),
.A2(n_2477),
.B(n_2208),
.Y(n_2827)
);

OAI21xp5_ASAP7_75t_L g2828 ( 
.A1(n_2703),
.A2(n_2208),
.B(n_2535),
.Y(n_2828)
);

AOI21xp5_ASAP7_75t_L g2829 ( 
.A1(n_2720),
.A2(n_2082),
.B(n_2041),
.Y(n_2829)
);

AOI21xp5_ASAP7_75t_L g2830 ( 
.A1(n_2720),
.A2(n_2082),
.B(n_2041),
.Y(n_2830)
);

AOI22xp5_ASAP7_75t_L g2831 ( 
.A1(n_2556),
.A2(n_1239),
.B1(n_1246),
.B2(n_1233),
.Y(n_2831)
);

AOI21xp5_ASAP7_75t_L g2832 ( 
.A1(n_2724),
.A2(n_2104),
.B(n_2041),
.Y(n_2832)
);

OAI22xp5_ASAP7_75t_L g2833 ( 
.A1(n_2671),
.A2(n_2147),
.B1(n_2256),
.B2(n_2255),
.Y(n_2833)
);

OAI22xp5_ASAP7_75t_L g2834 ( 
.A1(n_2688),
.A2(n_2147),
.B1(n_2256),
.B2(n_2232),
.Y(n_2834)
);

AOI21xp5_ASAP7_75t_L g2835 ( 
.A1(n_2724),
.A2(n_2104),
.B(n_2610),
.Y(n_2835)
);

AOI21x1_ASAP7_75t_L g2836 ( 
.A1(n_2645),
.A2(n_1625),
.B(n_2456),
.Y(n_2836)
);

OAI21xp5_ASAP7_75t_L g2837 ( 
.A1(n_2707),
.A2(n_2208),
.B(n_2196),
.Y(n_2837)
);

O2A1O1Ixp33_ASAP7_75t_L g2838 ( 
.A1(n_2719),
.A2(n_1089),
.B(n_1087),
.C(n_1114),
.Y(n_2838)
);

HB1xp67_ASAP7_75t_L g2839 ( 
.A(n_2555),
.Y(n_2839)
);

AOI21xp5_ASAP7_75t_L g2840 ( 
.A1(n_2610),
.A2(n_2104),
.B(n_2280),
.Y(n_2840)
);

CKINVDCx20_ASAP7_75t_R g2841 ( 
.A(n_2594),
.Y(n_2841)
);

OAI21xp5_ASAP7_75t_L g2842 ( 
.A1(n_2711),
.A2(n_2208),
.B(n_2196),
.Y(n_2842)
);

NOR2xp33_ASAP7_75t_L g2843 ( 
.A(n_2667),
.B(n_2210),
.Y(n_2843)
);

HB1xp67_ASAP7_75t_L g2844 ( 
.A(n_2585),
.Y(n_2844)
);

A2O1A1Ixp33_ASAP7_75t_L g2845 ( 
.A1(n_2713),
.A2(n_2516),
.B(n_2290),
.C(n_2258),
.Y(n_2845)
);

NOR3xp33_ASAP7_75t_L g2846 ( 
.A(n_2686),
.B(n_1080),
.C(n_1077),
.Y(n_2846)
);

AOI22xp5_ASAP7_75t_L g2847 ( 
.A1(n_2732),
.A2(n_1251),
.B1(n_2074),
.B2(n_1215),
.Y(n_2847)
);

OR2x2_ASAP7_75t_L g2848 ( 
.A(n_2591),
.B(n_2336),
.Y(n_2848)
);

AO21x1_ASAP7_75t_L g2849 ( 
.A1(n_2587),
.A2(n_2534),
.B(n_2537),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_L g2850 ( 
.A(n_2628),
.B(n_2336),
.Y(n_2850)
);

OAI22xp5_ASAP7_75t_L g2851 ( 
.A1(n_2643),
.A2(n_2232),
.B1(n_2104),
.B2(n_2258),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_L g2852 ( 
.A(n_2639),
.B(n_1473),
.Y(n_2852)
);

AOI21xp5_ASAP7_75t_L g2853 ( 
.A1(n_2572),
.A2(n_2286),
.B(n_2280),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_L g2854 ( 
.A(n_2658),
.B(n_1565),
.Y(n_2854)
);

A2O1A1Ixp33_ASAP7_75t_L g2855 ( 
.A1(n_2687),
.A2(n_2290),
.B(n_2036),
.C(n_1598),
.Y(n_2855)
);

AOI21xp5_ASAP7_75t_L g2856 ( 
.A1(n_2572),
.A2(n_2286),
.B(n_2280),
.Y(n_2856)
);

INVx2_ASAP7_75t_SL g2857 ( 
.A(n_2666),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_L g2858 ( 
.A(n_2650),
.B(n_1565),
.Y(n_2858)
);

AND2x4_ASAP7_75t_L g2859 ( 
.A(n_2657),
.B(n_2430),
.Y(n_2859)
);

OAI21xp33_ASAP7_75t_L g2860 ( 
.A1(n_2708),
.A2(n_1251),
.B(n_1215),
.Y(n_2860)
);

AOI21xp5_ASAP7_75t_L g2861 ( 
.A1(n_2624),
.A2(n_2286),
.B(n_2093),
.Y(n_2861)
);

AOI21xp5_ASAP7_75t_L g2862 ( 
.A1(n_2624),
.A2(n_2286),
.B(n_2093),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_L g2863 ( 
.A(n_2728),
.B(n_1565),
.Y(n_2863)
);

A2O1A1Ixp33_ASAP7_75t_L g2864 ( 
.A1(n_2590),
.A2(n_2036),
.B(n_1598),
.C(n_1594),
.Y(n_2864)
);

AND2x2_ASAP7_75t_L g2865 ( 
.A(n_2579),
.B(n_2430),
.Y(n_2865)
);

OAI21xp33_ASAP7_75t_L g2866 ( 
.A1(n_2684),
.A2(n_1217),
.B(n_1211),
.Y(n_2866)
);

HB1xp67_ASAP7_75t_L g2867 ( 
.A(n_2553),
.Y(n_2867)
);

OAI21xp5_ASAP7_75t_L g2868 ( 
.A1(n_2715),
.A2(n_2208),
.B(n_2196),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_SL g2869 ( 
.A(n_2680),
.B(n_2232),
.Y(n_2869)
);

BUFx3_ASAP7_75t_L g2870 ( 
.A(n_2666),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2566),
.Y(n_2871)
);

AOI21xp5_ASAP7_75t_L g2872 ( 
.A1(n_2623),
.A2(n_2263),
.B(n_2203),
.Y(n_2872)
);

A2O1A1Ixp33_ASAP7_75t_L g2873 ( 
.A1(n_2592),
.A2(n_1594),
.B(n_2232),
.C(n_1559),
.Y(n_2873)
);

AND2x2_ASAP7_75t_L g2874 ( 
.A(n_2579),
.B(n_2499),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_SL g2875 ( 
.A(n_2716),
.B(n_2499),
.Y(n_2875)
);

INVx2_ASAP7_75t_L g2876 ( 
.A(n_2642),
.Y(n_2876)
);

A2O1A1Ixp33_ASAP7_75t_L g2877 ( 
.A1(n_2601),
.A2(n_1559),
.B(n_1563),
.C(n_1550),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_L g2878 ( 
.A(n_2644),
.B(n_1565),
.Y(n_2878)
);

AND2x2_ASAP7_75t_L g2879 ( 
.A(n_2543),
.B(n_2499),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_L g2880 ( 
.A(n_2644),
.B(n_2016),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2654),
.B(n_1563),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2574),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2654),
.B(n_2657),
.Y(n_2883)
);

AOI22xp5_ASAP7_75t_L g2884 ( 
.A1(n_2652),
.A2(n_1217),
.B1(n_2269),
.B2(n_2257),
.Y(n_2884)
);

AND2x2_ASAP7_75t_SL g2885 ( 
.A(n_2697),
.B(n_2293),
.Y(n_2885)
);

AOI21xp5_ASAP7_75t_L g2886 ( 
.A1(n_2623),
.A2(n_2263),
.B(n_2203),
.Y(n_2886)
);

AOI21xp5_ASAP7_75t_L g2887 ( 
.A1(n_2634),
.A2(n_2189),
.B(n_2174),
.Y(n_2887)
);

NOR2xp33_ASAP7_75t_L g2888 ( 
.A(n_2543),
.B(n_2048),
.Y(n_2888)
);

BUFx2_ASAP7_75t_L g2889 ( 
.A(n_2716),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2581),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_L g2891 ( 
.A(n_2664),
.B(n_1566),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_SL g2892 ( 
.A(n_2664),
.B(n_2328),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_L g2893 ( 
.A(n_2669),
.B(n_1566),
.Y(n_2893)
);

OAI21xp5_ASAP7_75t_L g2894 ( 
.A1(n_2718),
.A2(n_2196),
.B(n_2046),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_L g2895 ( 
.A(n_2675),
.B(n_2677),
.Y(n_2895)
);

AOI21xp5_ASAP7_75t_L g2896 ( 
.A1(n_2634),
.A2(n_2235),
.B(n_2200),
.Y(n_2896)
);

CKINVDCx10_ASAP7_75t_R g2897 ( 
.A(n_2661),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_L g2898 ( 
.A(n_2734),
.B(n_1569),
.Y(n_2898)
);

AOI21xp5_ASAP7_75t_L g2899 ( 
.A1(n_2576),
.A2(n_2235),
.B(n_2233),
.Y(n_2899)
);

NOR2xp67_ASAP7_75t_L g2900 ( 
.A(n_2651),
.B(n_2233),
.Y(n_2900)
);

NAND2xp5_ASAP7_75t_L g2901 ( 
.A(n_2678),
.B(n_1569),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_2721),
.Y(n_2902)
);

O2A1O1Ixp33_ASAP7_75t_L g2903 ( 
.A1(n_2717),
.A2(n_1586),
.B(n_1589),
.C(n_1583),
.Y(n_2903)
);

INVx2_ASAP7_75t_L g2904 ( 
.A(n_2727),
.Y(n_2904)
);

AOI21xp5_ASAP7_75t_L g2905 ( 
.A1(n_2576),
.A2(n_2233),
.B(n_2328),
.Y(n_2905)
);

INVxp33_ASAP7_75t_L g2906 ( 
.A(n_2701),
.Y(n_2906)
);

AOI21xp5_ASAP7_75t_L g2907 ( 
.A1(n_2550),
.A2(n_2233),
.B(n_2328),
.Y(n_2907)
);

AOI21xp5_ASAP7_75t_L g2908 ( 
.A1(n_2550),
.A2(n_2344),
.B(n_2328),
.Y(n_2908)
);

NAND2xp5_ASAP7_75t_L g2909 ( 
.A(n_2685),
.B(n_1583),
.Y(n_2909)
);

OAI22xp5_ASAP7_75t_L g2910 ( 
.A1(n_2602),
.A2(n_583),
.B1(n_651),
.B2(n_478),
.Y(n_2910)
);

AOI21xp5_ASAP7_75t_L g2911 ( 
.A1(n_2725),
.A2(n_2344),
.B(n_2328),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_L g2912 ( 
.A(n_2722),
.B(n_1586),
.Y(n_2912)
);

NOR2xp33_ASAP7_75t_L g2913 ( 
.A(n_2672),
.B(n_2293),
.Y(n_2913)
);

BUFx4f_ASAP7_75t_L g2914 ( 
.A(n_2697),
.Y(n_2914)
);

CKINVDCx6p67_ASAP7_75t_R g2915 ( 
.A(n_2701),
.Y(n_2915)
);

INVx2_ASAP7_75t_L g2916 ( 
.A(n_2603),
.Y(n_2916)
);

A2O1A1Ixp33_ASAP7_75t_L g2917 ( 
.A1(n_2605),
.A2(n_1589),
.B(n_461),
.C(n_464),
.Y(n_2917)
);

AND2x2_ASAP7_75t_L g2918 ( 
.A(n_2683),
.B(n_456),
.Y(n_2918)
);

AOI21xp5_ASAP7_75t_L g2919 ( 
.A1(n_2725),
.A2(n_2344),
.B(n_2328),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_L g2920 ( 
.A(n_2729),
.B(n_2269),
.Y(n_2920)
);

INVx2_ASAP7_75t_L g2921 ( 
.A(n_2607),
.Y(n_2921)
);

INVx4_ASAP7_75t_L g2922 ( 
.A(n_2547),
.Y(n_2922)
);

INVx3_ASAP7_75t_L g2923 ( 
.A(n_2547),
.Y(n_2923)
);

NAND2x1p5_ASAP7_75t_L g2924 ( 
.A(n_2730),
.B(n_2735),
.Y(n_2924)
);

AOI21x1_ASAP7_75t_L g2925 ( 
.A1(n_2645),
.A2(n_2611),
.B(n_2636),
.Y(n_2925)
);

INVx4_ASAP7_75t_L g2926 ( 
.A(n_2575),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2612),
.Y(n_2927)
);

O2A1O1Ixp33_ASAP7_75t_L g2928 ( 
.A1(n_2774),
.A2(n_2619),
.B(n_2625),
.C(n_2620),
.Y(n_2928)
);

AOI21x1_ASAP7_75t_L g2929 ( 
.A1(n_2840),
.A2(n_2611),
.B(n_2683),
.Y(n_2929)
);

NOR3xp33_ASAP7_75t_SL g2930 ( 
.A(n_2866),
.B(n_2660),
.C(n_583),
.Y(n_2930)
);

HB1xp67_ASAP7_75t_L g2931 ( 
.A(n_2848),
.Y(n_2931)
);

NOR2xp33_ASAP7_75t_L g2932 ( 
.A(n_2802),
.B(n_2731),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_L g2933 ( 
.A(n_2753),
.B(n_2627),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_L g2934 ( 
.A(n_2741),
.B(n_2629),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_L g2935 ( 
.A(n_2770),
.B(n_2630),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2775),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_SL g2937 ( 
.A(n_2771),
.B(n_2735),
.Y(n_2937)
);

INVx3_ASAP7_75t_L g2938 ( 
.A(n_2922),
.Y(n_2938)
);

AOI21xp5_ASAP7_75t_L g2939 ( 
.A1(n_2738),
.A2(n_2636),
.B(n_2712),
.Y(n_2939)
);

AOI21xp5_ASAP7_75t_L g2940 ( 
.A1(n_2790),
.A2(n_2712),
.B(n_2640),
.Y(n_2940)
);

NOR2x1_ASAP7_75t_L g2941 ( 
.A(n_2796),
.B(n_2635),
.Y(n_2941)
);

AOI22xp5_ASAP7_75t_L g2942 ( 
.A1(n_2771),
.A2(n_2652),
.B1(n_2665),
.B2(n_2704),
.Y(n_2942)
);

OAI22xp5_ASAP7_75t_L g2943 ( 
.A1(n_2779),
.A2(n_2665),
.B1(n_2638),
.B2(n_2649),
.Y(n_2943)
);

BUFx4f_ASAP7_75t_L g2944 ( 
.A(n_2792),
.Y(n_2944)
);

O2A1O1Ixp33_ASAP7_75t_L g2945 ( 
.A1(n_2757),
.A2(n_2646),
.B(n_2662),
.C(n_2653),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_L g2946 ( 
.A(n_2739),
.B(n_2745),
.Y(n_2946)
);

NAND2x1p5_ASAP7_75t_L g2947 ( 
.A(n_2743),
.B(n_2733),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_SL g2948 ( 
.A(n_2795),
.B(n_2557),
.Y(n_2948)
);

INVx1_ASAP7_75t_SL g2949 ( 
.A(n_2744),
.Y(n_2949)
);

NOR2xp33_ASAP7_75t_L g2950 ( 
.A(n_2776),
.B(n_2682),
.Y(n_2950)
);

CKINVDCx5p33_ASAP7_75t_R g2951 ( 
.A(n_2897),
.Y(n_2951)
);

NAND2xp5_ASAP7_75t_SL g2952 ( 
.A(n_2766),
.B(n_2598),
.Y(n_2952)
);

NOR2xp33_ASAP7_75t_R g2953 ( 
.A(n_2805),
.B(n_2647),
.Y(n_2953)
);

AOI21xp5_ASAP7_75t_L g2954 ( 
.A1(n_2781),
.A2(n_2640),
.B(n_2704),
.Y(n_2954)
);

BUFx3_ASAP7_75t_L g2955 ( 
.A(n_2792),
.Y(n_2955)
);

AOI21xp5_ASAP7_75t_L g2956 ( 
.A1(n_2829),
.A2(n_2663),
.B(n_2631),
.Y(n_2956)
);

O2A1O1Ixp5_ASAP7_75t_L g2957 ( 
.A1(n_2813),
.A2(n_2800),
.B(n_2791),
.C(n_2835),
.Y(n_2957)
);

NAND2x1p5_ASAP7_75t_L g2958 ( 
.A(n_2743),
.B(n_2508),
.Y(n_2958)
);

BUFx3_ASAP7_75t_L g2959 ( 
.A(n_2792),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_SL g2960 ( 
.A(n_2780),
.B(n_2647),
.Y(n_2960)
);

OR2x2_ASAP7_75t_L g2961 ( 
.A(n_2844),
.B(n_1600),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_L g2962 ( 
.A(n_2777),
.B(n_2682),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_2916),
.Y(n_2963)
);

AND2x4_ASAP7_75t_L g2964 ( 
.A(n_2870),
.B(n_2508),
.Y(n_2964)
);

O2A1O1Ixp33_ASAP7_75t_SL g2965 ( 
.A1(n_2773),
.A2(n_1616),
.B(n_1098),
.C(n_2508),
.Y(n_2965)
);

AOI21x1_ASAP7_75t_L g2966 ( 
.A1(n_2836),
.A2(n_929),
.B(n_922),
.Y(n_2966)
);

AOI21xp5_ASAP7_75t_L g2967 ( 
.A1(n_2830),
.A2(n_2366),
.B(n_2344),
.Y(n_2967)
);

BUFx12f_ASAP7_75t_L g2968 ( 
.A(n_2754),
.Y(n_2968)
);

BUFx12f_ASAP7_75t_L g2969 ( 
.A(n_2754),
.Y(n_2969)
);

OAI22xp5_ASAP7_75t_L g2970 ( 
.A1(n_2801),
.A2(n_651),
.B1(n_652),
.B2(n_478),
.Y(n_2970)
);

NOR3xp33_ASAP7_75t_L g2971 ( 
.A(n_2783),
.B(n_658),
.C(n_652),
.Y(n_2971)
);

NAND3xp33_ASAP7_75t_L g2972 ( 
.A(n_2786),
.B(n_661),
.C(n_658),
.Y(n_2972)
);

NOR2xp33_ASAP7_75t_R g2973 ( 
.A(n_2841),
.B(n_2508),
.Y(n_2973)
);

AOI21xp5_ASAP7_75t_L g2974 ( 
.A1(n_2832),
.A2(n_2366),
.B(n_2344),
.Y(n_2974)
);

AOI21x1_ASAP7_75t_L g2975 ( 
.A1(n_2853),
.A2(n_933),
.B(n_922),
.Y(n_2975)
);

INVx5_ASAP7_75t_L g2976 ( 
.A(n_2743),
.Y(n_2976)
);

AO31x2_ASAP7_75t_L g2977 ( 
.A1(n_2778),
.A2(n_971),
.A3(n_977),
.B(n_933),
.Y(n_2977)
);

AOI21xp5_ASAP7_75t_L g2978 ( 
.A1(n_2742),
.A2(n_2749),
.B(n_2752),
.Y(n_2978)
);

NOR3xp33_ASAP7_75t_SL g2979 ( 
.A(n_2821),
.B(n_662),
.C(n_661),
.Y(n_2979)
);

OAI22xp5_ASAP7_75t_L g2980 ( 
.A1(n_2831),
.A2(n_2884),
.B1(n_2818),
.B2(n_2860),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2788),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2798),
.Y(n_2982)
);

INVxp67_ASAP7_75t_SL g2983 ( 
.A(n_2839),
.Y(n_2983)
);

BUFx3_ASAP7_75t_L g2984 ( 
.A(n_2785),
.Y(n_2984)
);

BUFx3_ASAP7_75t_L g2985 ( 
.A(n_2754),
.Y(n_2985)
);

AOI21xp5_ASAP7_75t_L g2986 ( 
.A1(n_2747),
.A2(n_2366),
.B(n_2344),
.Y(n_2986)
);

INVx2_ASAP7_75t_L g2987 ( 
.A(n_2921),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_SL g2988 ( 
.A(n_2746),
.B(n_2366),
.Y(n_2988)
);

O2A1O1Ixp33_ASAP7_75t_SL g2989 ( 
.A1(n_2855),
.A2(n_2869),
.B(n_2875),
.C(n_2917),
.Y(n_2989)
);

AOI22xp33_ASAP7_75t_L g2990 ( 
.A1(n_2918),
.A2(n_2257),
.B1(n_2269),
.B2(n_2196),
.Y(n_2990)
);

BUFx6f_ASAP7_75t_L g2991 ( 
.A(n_2817),
.Y(n_2991)
);

HB1xp67_ASAP7_75t_L g2992 ( 
.A(n_2822),
.Y(n_2992)
);

INVx2_ASAP7_75t_L g2993 ( 
.A(n_2748),
.Y(n_2993)
);

O2A1O1Ixp5_ASAP7_75t_L g2994 ( 
.A1(n_2908),
.A2(n_2366),
.B(n_2428),
.C(n_1477),
.Y(n_2994)
);

A2O1A1Ixp33_ASAP7_75t_L g2995 ( 
.A1(n_2838),
.A2(n_461),
.B(n_464),
.C(n_456),
.Y(n_2995)
);

O2A1O1Ixp33_ASAP7_75t_L g2996 ( 
.A1(n_2833),
.A2(n_887),
.B(n_664),
.C(n_665),
.Y(n_2996)
);

O2A1O1Ixp5_ASAP7_75t_L g2997 ( 
.A1(n_2828),
.A2(n_2366),
.B(n_2428),
.C(n_1477),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2825),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2799),
.B(n_662),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2826),
.Y(n_3000)
);

NOR2xp33_ASAP7_75t_R g3001 ( 
.A(n_2804),
.B(n_2046),
.Y(n_3001)
);

O2A1O1Ixp33_ASAP7_75t_L g3002 ( 
.A1(n_2834),
.A2(n_665),
.B(n_666),
.C(n_664),
.Y(n_3002)
);

OAI21x1_ASAP7_75t_L g3003 ( 
.A1(n_2911),
.A2(n_1477),
.B(n_1450),
.Y(n_3003)
);

AOI21xp5_ASAP7_75t_L g3004 ( 
.A1(n_2760),
.A2(n_2428),
.B(n_2257),
.Y(n_3004)
);

OAI21xp33_ASAP7_75t_SL g3005 ( 
.A1(n_2828),
.A2(n_2809),
.B(n_2789),
.Y(n_3005)
);

BUFx3_ASAP7_75t_L g3006 ( 
.A(n_2761),
.Y(n_3006)
);

BUFx8_ASAP7_75t_L g3007 ( 
.A(n_2889),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2871),
.Y(n_3008)
);

OAI22xp5_ASAP7_75t_L g3009 ( 
.A1(n_2824),
.A2(n_670),
.B1(n_672),
.B2(n_666),
.Y(n_3009)
);

INVx3_ASAP7_75t_L g3010 ( 
.A(n_2922),
.Y(n_3010)
);

INVx2_ASAP7_75t_L g3011 ( 
.A(n_2755),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2882),
.Y(n_3012)
);

OAI22xp5_ASAP7_75t_L g3013 ( 
.A1(n_2743),
.A2(n_672),
.B1(n_673),
.B2(n_670),
.Y(n_3013)
);

NAND2xp5_ASAP7_75t_L g3014 ( 
.A(n_2737),
.B(n_673),
.Y(n_3014)
);

OAI22xp5_ASAP7_75t_L g3015 ( 
.A1(n_2863),
.A2(n_2847),
.B1(n_2820),
.B2(n_2914),
.Y(n_3015)
);

O2A1O1Ixp33_ASAP7_75t_L g3016 ( 
.A1(n_2808),
.A2(n_681),
.B(n_684),
.C(n_674),
.Y(n_3016)
);

OAI22xp5_ASAP7_75t_L g3017 ( 
.A1(n_2890),
.A2(n_681),
.B1(n_684),
.B2(n_674),
.Y(n_3017)
);

OAI21x1_ASAP7_75t_L g3018 ( 
.A1(n_2919),
.A2(n_1450),
.B(n_1428),
.Y(n_3018)
);

NOR2xp67_ASAP7_75t_L g3019 ( 
.A(n_2751),
.B(n_246),
.Y(n_3019)
);

NOR2xp33_ASAP7_75t_L g3020 ( 
.A(n_2883),
.B(n_479),
.Y(n_3020)
);

AOI21xp5_ASAP7_75t_L g3021 ( 
.A1(n_2811),
.A2(n_2428),
.B(n_2257),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2927),
.Y(n_3022)
);

INVx2_ASAP7_75t_SL g3023 ( 
.A(n_2761),
.Y(n_3023)
);

AOI21xp5_ASAP7_75t_L g3024 ( 
.A1(n_2856),
.A2(n_2806),
.B(n_2819),
.Y(n_3024)
);

OAI22xp5_ASAP7_75t_L g3025 ( 
.A1(n_2914),
.A2(n_748),
.B1(n_752),
.B2(n_739),
.Y(n_3025)
);

AOI21x1_ASAP7_75t_L g3026 ( 
.A1(n_2905),
.A2(n_977),
.B(n_971),
.Y(n_3026)
);

AOI21xp5_ASAP7_75t_L g3027 ( 
.A1(n_2764),
.A2(n_2428),
.B(n_2257),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2895),
.Y(n_3028)
);

O2A1O1Ixp5_ASAP7_75t_L g3029 ( 
.A1(n_2793),
.A2(n_2428),
.B(n_1010),
.C(n_1046),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2765),
.Y(n_3030)
);

BUFx6f_ASAP7_75t_L g3031 ( 
.A(n_2761),
.Y(n_3031)
);

INVx3_ASAP7_75t_L g3032 ( 
.A(n_2859),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_2740),
.B(n_739),
.Y(n_3033)
);

AOI21xp5_ASAP7_75t_L g3034 ( 
.A1(n_2861),
.A2(n_1464),
.B(n_2246),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2850),
.B(n_748),
.Y(n_3035)
);

INVx2_ASAP7_75t_L g3036 ( 
.A(n_2772),
.Y(n_3036)
);

INVx2_ASAP7_75t_L g3037 ( 
.A(n_2807),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2815),
.Y(n_3038)
);

NOR2xp33_ASAP7_75t_R g3039 ( 
.A(n_2915),
.B(n_2046),
.Y(n_3039)
);

INVxp67_ASAP7_75t_L g3040 ( 
.A(n_2867),
.Y(n_3040)
);

OAI22xp5_ASAP7_75t_L g3041 ( 
.A1(n_2843),
.A2(n_480),
.B1(n_585),
.B2(n_479),
.Y(n_3041)
);

AND2x4_ASAP7_75t_L g3042 ( 
.A(n_2857),
.B(n_2046),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_L g3043 ( 
.A(n_2823),
.B(n_480),
.Y(n_3043)
);

AND2x4_ASAP7_75t_L g3044 ( 
.A(n_2859),
.B(n_2046),
.Y(n_3044)
);

AND2x2_ASAP7_75t_SL g3045 ( 
.A(n_2885),
.B(n_815),
.Y(n_3045)
);

AO22x1_ASAP7_75t_L g3046 ( 
.A1(n_2906),
.A2(n_649),
.B1(n_656),
.B2(n_585),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2876),
.Y(n_3047)
);

INVx2_ASAP7_75t_L g3048 ( 
.A(n_2902),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2904),
.B(n_649),
.Y(n_3049)
);

OAI22xp5_ASAP7_75t_L g3050 ( 
.A1(n_2845),
.A2(n_660),
.B1(n_663),
.B2(n_656),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_SL g3051 ( 
.A(n_2808),
.B(n_1615),
.Y(n_3051)
);

AOI21xp5_ASAP7_75t_L g3052 ( 
.A1(n_2862),
.A2(n_1464),
.B(n_1597),
.Y(n_3052)
);

NOR2xp33_ASAP7_75t_L g3053 ( 
.A(n_2880),
.B(n_660),
.Y(n_3053)
);

BUFx3_ASAP7_75t_L g3054 ( 
.A(n_2782),
.Y(n_3054)
);

AND2x2_ASAP7_75t_L g3055 ( 
.A(n_2750),
.B(n_663),
.Y(n_3055)
);

OAI21xp33_ASAP7_75t_L g3056 ( 
.A1(n_2910),
.A2(n_677),
.B(n_671),
.Y(n_3056)
);

INVx1_ASAP7_75t_SL g3057 ( 
.A(n_2891),
.Y(n_3057)
);

NOR2xp33_ASAP7_75t_L g3058 ( 
.A(n_2852),
.B(n_671),
.Y(n_3058)
);

NOR2xp33_ASAP7_75t_L g3059 ( 
.A(n_2865),
.B(n_677),
.Y(n_3059)
);

AO32x2_ASAP7_75t_L g3060 ( 
.A1(n_2784),
.A2(n_990),
.A3(n_7),
.B1(n_4),
.B2(n_5),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2849),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_L g3062 ( 
.A(n_2858),
.B(n_678),
.Y(n_3062)
);

NOR2xp33_ASAP7_75t_R g3063 ( 
.A(n_2874),
.B(n_678),
.Y(n_3063)
);

AO21x1_ASAP7_75t_L g3064 ( 
.A1(n_2887),
.A2(n_1023),
.B(n_1010),
.Y(n_3064)
);

AOI22xp33_ASAP7_75t_L g3065 ( 
.A1(n_2846),
.A2(n_2269),
.B1(n_744),
.B2(n_749),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2901),
.Y(n_3066)
);

CKINVDCx5p33_ASAP7_75t_R g3067 ( 
.A(n_2913),
.Y(n_3067)
);

OR2x2_ASAP7_75t_L g3068 ( 
.A(n_2784),
.B(n_1023),
.Y(n_3068)
);

HB1xp67_ASAP7_75t_L g3069 ( 
.A(n_2924),
.Y(n_3069)
);

A2O1A1Ixp33_ASAP7_75t_L g3070 ( 
.A1(n_2794),
.A2(n_744),
.B(n_749),
.C(n_683),
.Y(n_3070)
);

OR2x6_ASAP7_75t_L g3071 ( 
.A(n_2907),
.B(n_1615),
.Y(n_3071)
);

NOR2x1_ASAP7_75t_L g3072 ( 
.A(n_2923),
.B(n_2900),
.Y(n_3072)
);

NOR2xp67_ASAP7_75t_L g3073 ( 
.A(n_2881),
.B(n_2854),
.Y(n_3073)
);

AND2x2_ASAP7_75t_L g3074 ( 
.A(n_2879),
.B(n_683),
.Y(n_3074)
);

INVx4_ASAP7_75t_L g3075 ( 
.A(n_2782),
.Y(n_3075)
);

INVx2_ASAP7_75t_L g3076 ( 
.A(n_2893),
.Y(n_3076)
);

INVx1_ASAP7_75t_SL g3077 ( 
.A(n_2892),
.Y(n_3077)
);

INVx2_ASAP7_75t_L g3078 ( 
.A(n_2898),
.Y(n_3078)
);

NAND2xp5_ASAP7_75t_SL g3079 ( 
.A(n_2816),
.B(n_1615),
.Y(n_3079)
);

NAND2xp33_ASAP7_75t_SL g3080 ( 
.A(n_2787),
.B(n_567),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2909),
.B(n_575),
.Y(n_3081)
);

INVx3_ASAP7_75t_L g3082 ( 
.A(n_2923),
.Y(n_3082)
);

NOR2xp67_ASAP7_75t_L g3083 ( 
.A(n_2888),
.B(n_249),
.Y(n_3083)
);

AND2x4_ASAP7_75t_L g3084 ( 
.A(n_2926),
.B(n_2269),
.Y(n_3084)
);

NAND2xp5_ASAP7_75t_SL g3085 ( 
.A(n_2827),
.B(n_1615),
.Y(n_3085)
);

OAI21xp33_ASAP7_75t_L g3086 ( 
.A1(n_2910),
.A2(n_591),
.B(n_580),
.Y(n_3086)
);

INVx4_ASAP7_75t_L g3087 ( 
.A(n_2782),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_2809),
.B(n_597),
.Y(n_3088)
);

BUFx8_ASAP7_75t_SL g3089 ( 
.A(n_2878),
.Y(n_3089)
);

CKINVDCx20_ASAP7_75t_R g3090 ( 
.A(n_2926),
.Y(n_3090)
);

BUFx6f_ASAP7_75t_L g3091 ( 
.A(n_2924),
.Y(n_3091)
);

BUFx6f_ASAP7_75t_L g3092 ( 
.A(n_2812),
.Y(n_3092)
);

AND2x2_ASAP7_75t_L g3093 ( 
.A(n_2812),
.B(n_598),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_2912),
.Y(n_3094)
);

NOR2xp33_ASAP7_75t_L g3095 ( 
.A(n_2758),
.B(n_606),
.Y(n_3095)
);

AND2x4_ASAP7_75t_L g3096 ( 
.A(n_2920),
.B(n_250),
.Y(n_3096)
);

O2A1O1Ixp33_ASAP7_75t_L g3097 ( 
.A1(n_2873),
.A2(n_2814),
.B(n_2827),
.C(n_2851),
.Y(n_3097)
);

NOR2xp33_ASAP7_75t_L g3098 ( 
.A(n_2903),
.B(n_611),
.Y(n_3098)
);

BUFx3_ASAP7_75t_L g3099 ( 
.A(n_2814),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_L g3100 ( 
.A(n_2803),
.B(n_612),
.Y(n_3100)
);

NOR2xp33_ASAP7_75t_L g3101 ( 
.A(n_2768),
.B(n_615),
.Y(n_3101)
);

OAI22xp5_ASAP7_75t_L g3102 ( 
.A1(n_2864),
.A2(n_620),
.B1(n_623),
.B2(n_618),
.Y(n_3102)
);

AOI21xp5_ASAP7_75t_L g3103 ( 
.A1(n_2810),
.A2(n_1464),
.B(n_1597),
.Y(n_3103)
);

NOR2x1_ASAP7_75t_L g3104 ( 
.A(n_2899),
.B(n_1046),
.Y(n_3104)
);

AOI21xp5_ASAP7_75t_L g3105 ( 
.A1(n_2756),
.A2(n_1599),
.B(n_1597),
.Y(n_3105)
);

INVx2_ASAP7_75t_L g3106 ( 
.A(n_2925),
.Y(n_3106)
);

A2O1A1Ixp33_ASAP7_75t_SL g3107 ( 
.A1(n_2837),
.A2(n_2868),
.B(n_2842),
.C(n_2763),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_L g3108 ( 
.A(n_2768),
.B(n_627),
.Y(n_3108)
);

OAI21x1_ASAP7_75t_L g3109 ( 
.A1(n_2896),
.A2(n_1450),
.B(n_1428),
.Y(n_3109)
);

O2A1O1Ixp33_ASAP7_75t_L g3110 ( 
.A1(n_2877),
.A2(n_1063),
.B(n_1103),
.C(n_1102),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_2763),
.Y(n_3111)
);

OAI21xp33_ASAP7_75t_SL g3112 ( 
.A1(n_2894),
.A2(n_1102),
.B(n_1063),
.Y(n_3112)
);

INVx3_ASAP7_75t_L g3113 ( 
.A(n_2837),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_SL g3114 ( 
.A(n_2759),
.B(n_990),
.Y(n_3114)
);

INVx2_ASAP7_75t_L g3115 ( 
.A(n_2894),
.Y(n_3115)
);

O2A1O1Ixp5_ASAP7_75t_SL g3116 ( 
.A1(n_2842),
.A2(n_1428),
.B(n_990),
.C(n_692),
.Y(n_3116)
);

NOR2x1_ASAP7_75t_SL g3117 ( 
.A(n_2797),
.B(n_1597),
.Y(n_3117)
);

O2A1O1Ixp33_ASAP7_75t_L g3118 ( 
.A1(n_2868),
.A2(n_1103),
.B(n_10),
.C(n_8),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_L g3119 ( 
.A(n_2769),
.B(n_2767),
.Y(n_3119)
);

NOR2xp33_ASAP7_75t_L g3120 ( 
.A(n_2762),
.B(n_630),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_L g3121 ( 
.A(n_2872),
.B(n_694),
.Y(n_3121)
);

AOI221xp5_ASAP7_75t_L g3122 ( 
.A1(n_2886),
.A2(n_736),
.B1(n_738),
.B2(n_735),
.C(n_715),
.Y(n_3122)
);

OAI22x1_ASAP7_75t_L g3123 ( 
.A1(n_2884),
.A2(n_12),
.B1(n_8),
.B2(n_9),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_2753),
.B(n_9),
.Y(n_3124)
);

INVx3_ASAP7_75t_L g3125 ( 
.A(n_2922),
.Y(n_3125)
);

INVx2_ASAP7_75t_L g3126 ( 
.A(n_2916),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_2775),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_L g3128 ( 
.A(n_2753),
.B(n_12),
.Y(n_3128)
);

NOR2xp33_ASAP7_75t_L g3129 ( 
.A(n_2962),
.B(n_13),
.Y(n_3129)
);

AND2x4_ASAP7_75t_L g3130 ( 
.A(n_2983),
.B(n_254),
.Y(n_3130)
);

BUFx3_ASAP7_75t_L g3131 ( 
.A(n_2968),
.Y(n_3131)
);

HB1xp67_ASAP7_75t_L g3132 ( 
.A(n_2931),
.Y(n_3132)
);

INVx1_ASAP7_75t_SL g3133 ( 
.A(n_2949),
.Y(n_3133)
);

AND2x4_ASAP7_75t_L g3134 ( 
.A(n_2949),
.B(n_2936),
.Y(n_3134)
);

BUFx6f_ASAP7_75t_L g3135 ( 
.A(n_2991),
.Y(n_3135)
);

OAI21xp33_ASAP7_75t_L g3136 ( 
.A1(n_3101),
.A2(n_1599),
.B(n_1597),
.Y(n_3136)
);

BUFx6f_ASAP7_75t_L g3137 ( 
.A(n_2991),
.Y(n_3137)
);

AOI22xp5_ASAP7_75t_L g3138 ( 
.A1(n_2971),
.A2(n_1627),
.B1(n_1603),
.B2(n_1605),
.Y(n_3138)
);

AOI21xp5_ASAP7_75t_L g3139 ( 
.A1(n_3051),
.A2(n_1603),
.B(n_1599),
.Y(n_3139)
);

CKINVDCx20_ASAP7_75t_R g3140 ( 
.A(n_2951),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_2981),
.Y(n_3141)
);

INVx4_ASAP7_75t_L g3142 ( 
.A(n_2938),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_2982),
.Y(n_3143)
);

OAI22xp5_ASAP7_75t_L g3144 ( 
.A1(n_2979),
.A2(n_1603),
.B1(n_1605),
.B2(n_1599),
.Y(n_3144)
);

AOI21xp5_ASAP7_75t_L g3145 ( 
.A1(n_2965),
.A2(n_1603),
.B(n_1599),
.Y(n_3145)
);

INVx3_ASAP7_75t_L g3146 ( 
.A(n_3091),
.Y(n_3146)
);

INVx3_ASAP7_75t_L g3147 ( 
.A(n_3091),
.Y(n_3147)
);

OR2x6_ASAP7_75t_L g3148 ( 
.A(n_2937),
.B(n_1603),
.Y(n_3148)
);

AOI22xp5_ASAP7_75t_L g3149 ( 
.A1(n_2980),
.A2(n_1627),
.B1(n_1610),
.B2(n_1613),
.Y(n_3149)
);

INVx1_ASAP7_75t_SL g3150 ( 
.A(n_3090),
.Y(n_3150)
);

INVx1_ASAP7_75t_SL g3151 ( 
.A(n_2984),
.Y(n_3151)
);

BUFx6f_ASAP7_75t_L g3152 ( 
.A(n_2991),
.Y(n_3152)
);

INVxp67_ASAP7_75t_SL g3153 ( 
.A(n_2992),
.Y(n_3153)
);

BUFx12f_ASAP7_75t_L g3154 ( 
.A(n_3007),
.Y(n_3154)
);

AOI21xp5_ASAP7_75t_L g3155 ( 
.A1(n_3024),
.A2(n_1610),
.B(n_1605),
.Y(n_3155)
);

BUFx6f_ASAP7_75t_L g3156 ( 
.A(n_3031),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_2998),
.Y(n_3157)
);

CKINVDCx6p67_ASAP7_75t_R g3158 ( 
.A(n_2969),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_SL g3159 ( 
.A(n_2946),
.B(n_1605),
.Y(n_3159)
);

INVx2_ASAP7_75t_L g3160 ( 
.A(n_2963),
.Y(n_3160)
);

INVx3_ASAP7_75t_L g3161 ( 
.A(n_3091),
.Y(n_3161)
);

INVx2_ASAP7_75t_SL g3162 ( 
.A(n_2985),
.Y(n_3162)
);

INVx2_ASAP7_75t_L g3163 ( 
.A(n_2987),
.Y(n_3163)
);

BUFx2_ASAP7_75t_L g3164 ( 
.A(n_3069),
.Y(n_3164)
);

BUFx3_ASAP7_75t_L g3165 ( 
.A(n_2955),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_3000),
.Y(n_3166)
);

BUFx3_ASAP7_75t_L g3167 ( 
.A(n_2959),
.Y(n_3167)
);

AND2x4_ASAP7_75t_L g3168 ( 
.A(n_3008),
.B(n_258),
.Y(n_3168)
);

BUFx6f_ASAP7_75t_L g3169 ( 
.A(n_3031),
.Y(n_3169)
);

NOR2xp33_ASAP7_75t_L g3170 ( 
.A(n_2932),
.B(n_13),
.Y(n_3170)
);

BUFx2_ASAP7_75t_L g3171 ( 
.A(n_3089),
.Y(n_3171)
);

BUFx6f_ASAP7_75t_L g3172 ( 
.A(n_3031),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_3012),
.Y(n_3173)
);

BUFx2_ASAP7_75t_L g3174 ( 
.A(n_2973),
.Y(n_3174)
);

INVx1_ASAP7_75t_SL g3175 ( 
.A(n_3063),
.Y(n_3175)
);

BUFx2_ASAP7_75t_L g3176 ( 
.A(n_3040),
.Y(n_3176)
);

BUFx6f_ASAP7_75t_L g3177 ( 
.A(n_2944),
.Y(n_3177)
);

INVxp67_ASAP7_75t_L g3178 ( 
.A(n_3014),
.Y(n_3178)
);

NAND2xp5_ASAP7_75t_L g3179 ( 
.A(n_3057),
.B(n_3028),
.Y(n_3179)
);

AOI22xp5_ASAP7_75t_L g3180 ( 
.A1(n_3015),
.A2(n_1627),
.B1(n_1610),
.B2(n_1613),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_3022),
.Y(n_3181)
);

INVx4_ASAP7_75t_L g3182 ( 
.A(n_2938),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_3127),
.Y(n_3183)
);

INVx2_ASAP7_75t_L g3184 ( 
.A(n_3126),
.Y(n_3184)
);

INVx3_ASAP7_75t_L g3185 ( 
.A(n_3092),
.Y(n_3185)
);

INVx2_ASAP7_75t_L g3186 ( 
.A(n_3030),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_3061),
.Y(n_3187)
);

CKINVDCx5p33_ASAP7_75t_R g3188 ( 
.A(n_2953),
.Y(n_3188)
);

BUFx2_ASAP7_75t_L g3189 ( 
.A(n_3092),
.Y(n_3189)
);

AND2x2_ASAP7_75t_L g3190 ( 
.A(n_3057),
.B(n_14),
.Y(n_3190)
);

CKINVDCx8_ASAP7_75t_R g3191 ( 
.A(n_3067),
.Y(n_3191)
);

INVx2_ASAP7_75t_L g3192 ( 
.A(n_3038),
.Y(n_3192)
);

BUFx2_ASAP7_75t_L g3193 ( 
.A(n_3092),
.Y(n_3193)
);

INVx2_ASAP7_75t_L g3194 ( 
.A(n_3047),
.Y(n_3194)
);

OR2x6_ASAP7_75t_L g3195 ( 
.A(n_2939),
.B(n_1605),
.Y(n_3195)
);

AOI22xp5_ASAP7_75t_L g3196 ( 
.A1(n_2960),
.A2(n_1613),
.B1(n_1610),
.B2(n_1495),
.Y(n_3196)
);

BUFx4_ASAP7_75t_SL g3197 ( 
.A(n_3006),
.Y(n_3197)
);

BUFx12f_ASAP7_75t_L g3198 ( 
.A(n_3007),
.Y(n_3198)
);

INVx1_ASAP7_75t_SL g3199 ( 
.A(n_3054),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_L g3200 ( 
.A(n_2933),
.B(n_14),
.Y(n_3200)
);

INVx2_ASAP7_75t_L g3201 ( 
.A(n_2993),
.Y(n_3201)
);

AOI22xp33_ASAP7_75t_SL g3202 ( 
.A1(n_3099),
.A2(n_819),
.B1(n_836),
.B2(n_816),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_3111),
.Y(n_3203)
);

BUFx3_ASAP7_75t_L g3204 ( 
.A(n_2944),
.Y(n_3204)
);

OR2x6_ASAP7_75t_L g3205 ( 
.A(n_2952),
.B(n_1610),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_3106),
.Y(n_3206)
);

AOI22xp33_ASAP7_75t_L g3207 ( 
.A1(n_3123),
.A2(n_1613),
.B1(n_1495),
.B2(n_1557),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_3119),
.Y(n_3208)
);

INVx5_ASAP7_75t_L g3209 ( 
.A(n_2976),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_2929),
.Y(n_3210)
);

INVx2_ASAP7_75t_SL g3211 ( 
.A(n_3023),
.Y(n_3211)
);

HAxp5_ASAP7_75t_L g3212 ( 
.A(n_2970),
.B(n_15),
.CON(n_3212),
.SN(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_3011),
.Y(n_3213)
);

AOI222xp33_ASAP7_75t_L g3214 ( 
.A1(n_2970),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.C1(n_19),
.C2(n_20),
.Y(n_3214)
);

O2A1O1Ixp33_ASAP7_75t_L g3215 ( 
.A1(n_3016),
.A2(n_21),
.B(n_17),
.C(n_20),
.Y(n_3215)
);

AND2x2_ASAP7_75t_L g3216 ( 
.A(n_3077),
.B(n_21),
.Y(n_3216)
);

BUFx2_ASAP7_75t_L g3217 ( 
.A(n_3032),
.Y(n_3217)
);

BUFx2_ASAP7_75t_L g3218 ( 
.A(n_3032),
.Y(n_3218)
);

BUFx12f_ASAP7_75t_L g3219 ( 
.A(n_3045),
.Y(n_3219)
);

HB1xp67_ASAP7_75t_L g3220 ( 
.A(n_3077),
.Y(n_3220)
);

NOR2xp33_ASAP7_75t_L g3221 ( 
.A(n_3020),
.B(n_22),
.Y(n_3221)
);

BUFx2_ASAP7_75t_L g3222 ( 
.A(n_3075),
.Y(n_3222)
);

HB1xp67_ASAP7_75t_L g3223 ( 
.A(n_2941),
.Y(n_3223)
);

BUFx2_ASAP7_75t_L g3224 ( 
.A(n_3075),
.Y(n_3224)
);

NOR2xp33_ASAP7_75t_L g3225 ( 
.A(n_3059),
.B(n_3095),
.Y(n_3225)
);

INVx6_ASAP7_75t_SL g3226 ( 
.A(n_2964),
.Y(n_3226)
);

AND2x4_ASAP7_75t_L g3227 ( 
.A(n_3010),
.B(n_259),
.Y(n_3227)
);

AND2x4_ASAP7_75t_L g3228 ( 
.A(n_3010),
.B(n_268),
.Y(n_3228)
);

OR2x2_ASAP7_75t_L g3229 ( 
.A(n_2935),
.B(n_2961),
.Y(n_3229)
);

BUFx2_ASAP7_75t_L g3230 ( 
.A(n_3087),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_3036),
.Y(n_3231)
);

BUFx6f_ASAP7_75t_L g3232 ( 
.A(n_3087),
.Y(n_3232)
);

INVx2_ASAP7_75t_L g3233 ( 
.A(n_3037),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_3048),
.Y(n_3234)
);

BUFx2_ASAP7_75t_L g3235 ( 
.A(n_3125),
.Y(n_3235)
);

OAI22xp5_ASAP7_75t_L g3236 ( 
.A1(n_2930),
.A2(n_1613),
.B1(n_1554),
.B2(n_1557),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_L g3237 ( 
.A(n_2934),
.B(n_22),
.Y(n_3237)
);

INVx3_ASAP7_75t_L g3238 ( 
.A(n_2947),
.Y(n_3238)
);

INVx3_ASAP7_75t_SL g3239 ( 
.A(n_3074),
.Y(n_3239)
);

AOI22xp5_ASAP7_75t_L g3240 ( 
.A1(n_2972),
.A2(n_2950),
.B1(n_3080),
.B2(n_2943),
.Y(n_3240)
);

CKINVDCx11_ASAP7_75t_R g3241 ( 
.A(n_2964),
.Y(n_3241)
);

AND2x4_ASAP7_75t_L g3242 ( 
.A(n_3125),
.B(n_269),
.Y(n_3242)
);

NAND2xp33_ASAP7_75t_L g3243 ( 
.A(n_3056),
.B(n_1561),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_2957),
.Y(n_3244)
);

INVx2_ASAP7_75t_L g3245 ( 
.A(n_3076),
.Y(n_3245)
);

BUFx3_ASAP7_75t_L g3246 ( 
.A(n_3082),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_L g3247 ( 
.A(n_3066),
.B(n_24),
.Y(n_3247)
);

BUFx6f_ASAP7_75t_L g3248 ( 
.A(n_2976),
.Y(n_3248)
);

INVx3_ASAP7_75t_L g3249 ( 
.A(n_2947),
.Y(n_3249)
);

INVx2_ASAP7_75t_SL g3250 ( 
.A(n_3082),
.Y(n_3250)
);

INVx3_ASAP7_75t_L g3251 ( 
.A(n_2976),
.Y(n_3251)
);

INVx1_ASAP7_75t_SL g3252 ( 
.A(n_3033),
.Y(n_3252)
);

BUFx2_ASAP7_75t_L g3253 ( 
.A(n_3072),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_2940),
.Y(n_3254)
);

AOI22xp33_ASAP7_75t_L g3255 ( 
.A1(n_2972),
.A2(n_1495),
.B1(n_1557),
.B2(n_1554),
.Y(n_3255)
);

INVx5_ASAP7_75t_L g3256 ( 
.A(n_3071),
.Y(n_3256)
);

BUFx3_ASAP7_75t_L g3257 ( 
.A(n_2958),
.Y(n_3257)
);

AND2x2_ASAP7_75t_L g3258 ( 
.A(n_3113),
.B(n_24),
.Y(n_3258)
);

INVx3_ASAP7_75t_L g3259 ( 
.A(n_2958),
.Y(n_3259)
);

AND2x2_ASAP7_75t_L g3260 ( 
.A(n_3113),
.B(n_25),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_3060),
.Y(n_3261)
);

INVx2_ASAP7_75t_SL g3262 ( 
.A(n_3039),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_3060),
.Y(n_3263)
);

AND2x4_ASAP7_75t_L g3264 ( 
.A(n_3073),
.B(n_270),
.Y(n_3264)
);

INVx2_ASAP7_75t_L g3265 ( 
.A(n_3078),
.Y(n_3265)
);

CKINVDCx5p33_ASAP7_75t_R g3266 ( 
.A(n_3001),
.Y(n_3266)
);

BUFx3_ASAP7_75t_L g3267 ( 
.A(n_3044),
.Y(n_3267)
);

INVx5_ASAP7_75t_L g3268 ( 
.A(n_3071),
.Y(n_3268)
);

AND2x4_ASAP7_75t_L g3269 ( 
.A(n_2942),
.B(n_271),
.Y(n_3269)
);

AOI21xp5_ASAP7_75t_L g3270 ( 
.A1(n_3004),
.A2(n_2978),
.B(n_3100),
.Y(n_3270)
);

AND2x4_ASAP7_75t_L g3271 ( 
.A(n_2942),
.B(n_272),
.Y(n_3271)
);

CKINVDCx5p33_ASAP7_75t_R g3272 ( 
.A(n_3035),
.Y(n_3272)
);

OR2x6_ASAP7_75t_SL g3273 ( 
.A(n_3121),
.B(n_28),
.Y(n_3273)
);

INVx2_ASAP7_75t_L g3274 ( 
.A(n_3094),
.Y(n_3274)
);

BUFx3_ASAP7_75t_L g3275 ( 
.A(n_3044),
.Y(n_3275)
);

INVx1_ASAP7_75t_L g3276 ( 
.A(n_3060),
.Y(n_3276)
);

AND2x4_ASAP7_75t_L g3277 ( 
.A(n_3042),
.B(n_275),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_3071),
.Y(n_3278)
);

BUFx6f_ASAP7_75t_L g3279 ( 
.A(n_3042),
.Y(n_3279)
);

INVx3_ASAP7_75t_L g3280 ( 
.A(n_3084),
.Y(n_3280)
);

AO32x1_ASAP7_75t_L g3281 ( 
.A1(n_3050),
.A2(n_31),
.A3(n_28),
.B1(n_29),
.B2(n_32),
.Y(n_3281)
);

BUFx6f_ASAP7_75t_L g3282 ( 
.A(n_3084),
.Y(n_3282)
);

AOI22xp33_ASAP7_75t_L g3283 ( 
.A1(n_3098),
.A2(n_1495),
.B1(n_1557),
.B2(n_1554),
.Y(n_3283)
);

INVx1_ASAP7_75t_SL g3284 ( 
.A(n_3093),
.Y(n_3284)
);

NOR2xp67_ASAP7_75t_SL g3285 ( 
.A(n_2956),
.B(n_1495),
.Y(n_3285)
);

CKINVDCx5p33_ASAP7_75t_R g3286 ( 
.A(n_3055),
.Y(n_3286)
);

INVx2_ASAP7_75t_L g3287 ( 
.A(n_3115),
.Y(n_3287)
);

NAND3xp33_ASAP7_75t_L g3288 ( 
.A(n_3108),
.B(n_1557),
.C(n_1554),
.Y(n_3288)
);

NOR2xp33_ASAP7_75t_R g3289 ( 
.A(n_3058),
.B(n_276),
.Y(n_3289)
);

OR2x2_ASAP7_75t_L g3290 ( 
.A(n_3124),
.B(n_3128),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_L g3291 ( 
.A(n_3053),
.B(n_31),
.Y(n_3291)
);

AND2x4_ASAP7_75t_L g3292 ( 
.A(n_2948),
.B(n_278),
.Y(n_3292)
);

AND2x4_ASAP7_75t_SL g3293 ( 
.A(n_3096),
.B(n_1471),
.Y(n_3293)
);

NOR2xp33_ASAP7_75t_L g3294 ( 
.A(n_2999),
.B(n_33),
.Y(n_3294)
);

INVx3_ASAP7_75t_L g3295 ( 
.A(n_3096),
.Y(n_3295)
);

BUFx3_ASAP7_75t_L g3296 ( 
.A(n_3043),
.Y(n_3296)
);

INVx2_ASAP7_75t_L g3297 ( 
.A(n_2977),
.Y(n_3297)
);

NAND3xp33_ASAP7_75t_L g3298 ( 
.A(n_3122),
.B(n_3050),
.C(n_3120),
.Y(n_3298)
);

INVx2_ASAP7_75t_L g3299 ( 
.A(n_2977),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_2928),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_2945),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_2977),
.Y(n_3302)
);

OR2x2_ASAP7_75t_L g3303 ( 
.A(n_3085),
.B(n_3068),
.Y(n_3303)
);

OR2x6_ASAP7_75t_L g3304 ( 
.A(n_2988),
.B(n_816),
.Y(n_3304)
);

OAI22xp5_ASAP7_75t_SL g3305 ( 
.A1(n_3009),
.A2(n_36),
.B1(n_33),
.B2(n_34),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_L g3306 ( 
.A(n_3088),
.B(n_34),
.Y(n_3306)
);

INVx3_ASAP7_75t_L g3307 ( 
.A(n_3109),
.Y(n_3307)
);

INVx8_ASAP7_75t_L g3308 ( 
.A(n_3083),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_2954),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_3005),
.Y(n_3310)
);

BUFx3_ASAP7_75t_L g3311 ( 
.A(n_3049),
.Y(n_3311)
);

INVx1_ASAP7_75t_L g3312 ( 
.A(n_3005),
.Y(n_3312)
);

BUFx6f_ASAP7_75t_L g3313 ( 
.A(n_3062),
.Y(n_3313)
);

INVx3_ASAP7_75t_L g3314 ( 
.A(n_3018),
.Y(n_3314)
);

INVx2_ASAP7_75t_SL g3315 ( 
.A(n_3081),
.Y(n_3315)
);

OAI222xp33_ASAP7_75t_L g3316 ( 
.A1(n_3002),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.C1(n_41),
.C2(n_42),
.Y(n_3316)
);

CKINVDCx5p33_ASAP7_75t_R g3317 ( 
.A(n_3025),
.Y(n_3317)
);

AOI221xp5_ASAP7_75t_L g3318 ( 
.A1(n_3056),
.A2(n_1561),
.B1(n_1560),
.B2(n_1554),
.C(n_867),
.Y(n_3318)
);

NOR2xp33_ASAP7_75t_L g3319 ( 
.A(n_3041),
.B(n_37),
.Y(n_3319)
);

INVx6_ASAP7_75t_L g3320 ( 
.A(n_3019),
.Y(n_3320)
);

OR2x2_ASAP7_75t_L g3321 ( 
.A(n_3107),
.B(n_816),
.Y(n_3321)
);

INVx1_ASAP7_75t_SL g3322 ( 
.A(n_3046),
.Y(n_3322)
);

AOI21xp5_ASAP7_75t_L g3323 ( 
.A1(n_3079),
.A2(n_1561),
.B(n_1560),
.Y(n_3323)
);

AOI21xp5_ASAP7_75t_L g3324 ( 
.A1(n_3118),
.A2(n_1561),
.B(n_1560),
.Y(n_3324)
);

INVxp67_ASAP7_75t_L g3325 ( 
.A(n_3013),
.Y(n_3325)
);

AOI22xp5_ASAP7_75t_L g3326 ( 
.A1(n_3086),
.A2(n_2989),
.B1(n_3114),
.B2(n_3065),
.Y(n_3326)
);

INVx2_ASAP7_75t_SL g3327 ( 
.A(n_3104),
.Y(n_3327)
);

AND2x4_ASAP7_75t_L g3328 ( 
.A(n_3021),
.B(n_279),
.Y(n_3328)
);

AOI22xp33_ASAP7_75t_L g3329 ( 
.A1(n_3086),
.A2(n_1561),
.B1(n_1560),
.B2(n_836),
.Y(n_3329)
);

BUFx6f_ASAP7_75t_L g3330 ( 
.A(n_3003),
.Y(n_3330)
);

NAND2xp33_ASAP7_75t_SL g3331 ( 
.A(n_3013),
.B(n_819),
.Y(n_3331)
);

BUFx3_ASAP7_75t_L g3332 ( 
.A(n_3017),
.Y(n_3332)
);

AOI22xp33_ASAP7_75t_L g3333 ( 
.A1(n_2990),
.A2(n_1560),
.B1(n_836),
.B2(n_857),
.Y(n_3333)
);

O2A1O1Ixp33_ASAP7_75t_L g3334 ( 
.A1(n_2996),
.A2(n_41),
.B(n_39),
.C(n_40),
.Y(n_3334)
);

CKINVDCx5p33_ASAP7_75t_R g3335 ( 
.A(n_3017),
.Y(n_3335)
);

INVx2_ASAP7_75t_SL g3336 ( 
.A(n_3102),
.Y(n_3336)
);

OR2x6_ASAP7_75t_L g3337 ( 
.A(n_3097),
.B(n_819),
.Y(n_3337)
);

HB1xp67_ASAP7_75t_L g3338 ( 
.A(n_2975),
.Y(n_3338)
);

BUFx6f_ASAP7_75t_L g3339 ( 
.A(n_3026),
.Y(n_3339)
);

INVx6_ASAP7_75t_L g3340 ( 
.A(n_2995),
.Y(n_3340)
);

BUFx2_ASAP7_75t_L g3341 ( 
.A(n_3112),
.Y(n_3341)
);

AND2x6_ASAP7_75t_L g3342 ( 
.A(n_3269),
.B(n_3117),
.Y(n_3342)
);

INVx2_ASAP7_75t_L g3343 ( 
.A(n_3134),
.Y(n_3343)
);

BUFx3_ASAP7_75t_L g3344 ( 
.A(n_3154),
.Y(n_3344)
);

OAI21x1_ASAP7_75t_L g3345 ( 
.A1(n_3270),
.A2(n_2994),
.B(n_3052),
.Y(n_3345)
);

BUFx3_ASAP7_75t_L g3346 ( 
.A(n_3198),
.Y(n_3346)
);

INVx2_ASAP7_75t_SL g3347 ( 
.A(n_3135),
.Y(n_3347)
);

AND2x2_ASAP7_75t_L g3348 ( 
.A(n_3132),
.B(n_3034),
.Y(n_3348)
);

INVx2_ASAP7_75t_L g3349 ( 
.A(n_3134),
.Y(n_3349)
);

BUFx6f_ASAP7_75t_L g3350 ( 
.A(n_3135),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_3141),
.Y(n_3351)
);

NOR2xp33_ASAP7_75t_L g3352 ( 
.A(n_3225),
.B(n_3070),
.Y(n_3352)
);

OA21x2_ASAP7_75t_L g3353 ( 
.A1(n_3244),
.A2(n_3105),
.B(n_3029),
.Y(n_3353)
);

BUFx3_ASAP7_75t_L g3354 ( 
.A(n_3140),
.Y(n_3354)
);

O2A1O1Ixp33_ASAP7_75t_L g3355 ( 
.A1(n_3316),
.A2(n_3334),
.B(n_3215),
.C(n_3212),
.Y(n_3355)
);

OR2x6_ASAP7_75t_L g3356 ( 
.A(n_3195),
.B(n_3027),
.Y(n_3356)
);

INVx5_ASAP7_75t_L g3357 ( 
.A(n_3248),
.Y(n_3357)
);

NAND2xp5_ASAP7_75t_L g3358 ( 
.A(n_3208),
.B(n_3112),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_L g3359 ( 
.A(n_3208),
.B(n_3064),
.Y(n_3359)
);

INVx3_ASAP7_75t_L g3360 ( 
.A(n_3146),
.Y(n_3360)
);

AOI22xp33_ASAP7_75t_L g3361 ( 
.A1(n_3298),
.A2(n_2986),
.B1(n_2974),
.B2(n_2967),
.Y(n_3361)
);

AO22x1_ASAP7_75t_L g3362 ( 
.A1(n_3170),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_3362)
);

BUFx12f_ASAP7_75t_L g3363 ( 
.A(n_3188),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_3141),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_3143),
.Y(n_3365)
);

BUFx12f_ASAP7_75t_L g3366 ( 
.A(n_3286),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_3143),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_L g3368 ( 
.A(n_3179),
.B(n_3103),
.Y(n_3368)
);

NOR2xp67_ASAP7_75t_SL g3369 ( 
.A(n_3191),
.B(n_819),
.Y(n_3369)
);

INVx1_ASAP7_75t_SL g3370 ( 
.A(n_3133),
.Y(n_3370)
);

BUFx6f_ASAP7_75t_L g3371 ( 
.A(n_3135),
.Y(n_3371)
);

BUFx3_ASAP7_75t_L g3372 ( 
.A(n_3137),
.Y(n_3372)
);

INVx2_ASAP7_75t_L g3373 ( 
.A(n_3157),
.Y(n_3373)
);

BUFx3_ASAP7_75t_L g3374 ( 
.A(n_3137),
.Y(n_3374)
);

AOI21xp5_ASAP7_75t_L g3375 ( 
.A1(n_3243),
.A2(n_2997),
.B(n_3110),
.Y(n_3375)
);

INVx1_ASAP7_75t_SL g3376 ( 
.A(n_3164),
.Y(n_3376)
);

INVx4_ASAP7_75t_L g3377 ( 
.A(n_3137),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_3166),
.Y(n_3378)
);

INVx2_ASAP7_75t_L g3379 ( 
.A(n_3186),
.Y(n_3379)
);

INVx2_ASAP7_75t_L g3380 ( 
.A(n_3192),
.Y(n_3380)
);

INVx3_ASAP7_75t_SL g3381 ( 
.A(n_3158),
.Y(n_3381)
);

INVx1_ASAP7_75t_L g3382 ( 
.A(n_3166),
.Y(n_3382)
);

INVxp67_ASAP7_75t_L g3383 ( 
.A(n_3176),
.Y(n_3383)
);

INVx2_ASAP7_75t_L g3384 ( 
.A(n_3194),
.Y(n_3384)
);

AOI21xp5_ASAP7_75t_L g3385 ( 
.A1(n_3136),
.A2(n_3116),
.B(n_2966),
.Y(n_3385)
);

INVx4_ASAP7_75t_L g3386 ( 
.A(n_3152),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_3173),
.Y(n_3387)
);

NOR2xp33_ASAP7_75t_L g3388 ( 
.A(n_3313),
.B(n_46),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_L g3389 ( 
.A(n_3153),
.B(n_3220),
.Y(n_3389)
);

BUFx3_ASAP7_75t_L g3390 ( 
.A(n_3152),
.Y(n_3390)
);

BUFx6f_ASAP7_75t_L g3391 ( 
.A(n_3152),
.Y(n_3391)
);

INVx2_ASAP7_75t_L g3392 ( 
.A(n_3173),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_L g3393 ( 
.A(n_3229),
.B(n_46),
.Y(n_3393)
);

AND2x2_ASAP7_75t_L g3394 ( 
.A(n_3284),
.B(n_47),
.Y(n_3394)
);

CKINVDCx5p33_ASAP7_75t_R g3395 ( 
.A(n_3197),
.Y(n_3395)
);

OAI22xp5_ASAP7_75t_SL g3396 ( 
.A1(n_3335),
.A2(n_51),
.B1(n_48),
.B2(n_50),
.Y(n_3396)
);

O2A1O1Ixp33_ASAP7_75t_SL g3397 ( 
.A1(n_3221),
.A2(n_3291),
.B(n_3306),
.C(n_3322),
.Y(n_3397)
);

AND2x2_ASAP7_75t_L g3398 ( 
.A(n_3239),
.B(n_52),
.Y(n_3398)
);

AOI21xp33_ASAP7_75t_SL g3399 ( 
.A1(n_3308),
.A2(n_53),
.B(n_54),
.Y(n_3399)
);

AOI21xp5_ASAP7_75t_L g3400 ( 
.A1(n_3324),
.A2(n_1461),
.B(n_1451),
.Y(n_3400)
);

OA21x2_ASAP7_75t_L g3401 ( 
.A1(n_3244),
.A2(n_54),
.B(n_55),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_3203),
.B(n_55),
.Y(n_3402)
);

OAI21x1_ASAP7_75t_L g3403 ( 
.A1(n_3155),
.A2(n_284),
.B(n_282),
.Y(n_3403)
);

O2A1O1Ixp5_ASAP7_75t_L g3404 ( 
.A1(n_3319),
.A2(n_59),
.B(n_57),
.C(n_58),
.Y(n_3404)
);

O2A1O1Ixp33_ASAP7_75t_L g3405 ( 
.A1(n_3214),
.A2(n_62),
.B(n_57),
.C(n_61),
.Y(n_3405)
);

INVxp67_ASAP7_75t_L g3406 ( 
.A(n_3313),
.Y(n_3406)
);

CKINVDCx5p33_ASAP7_75t_R g3407 ( 
.A(n_3171),
.Y(n_3407)
);

AND2x2_ASAP7_75t_L g3408 ( 
.A(n_3217),
.B(n_61),
.Y(n_3408)
);

INVx1_ASAP7_75t_L g3409 ( 
.A(n_3181),
.Y(n_3409)
);

AOI21xp5_ASAP7_75t_L g3410 ( 
.A1(n_3331),
.A2(n_1461),
.B(n_1451),
.Y(n_3410)
);

INVx3_ASAP7_75t_L g3411 ( 
.A(n_3146),
.Y(n_3411)
);

NAND2xp5_ASAP7_75t_L g3412 ( 
.A(n_3203),
.B(n_65),
.Y(n_3412)
);

AOI21xp33_ASAP7_75t_SL g3413 ( 
.A1(n_3308),
.A2(n_67),
.B(n_68),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_L g3414 ( 
.A(n_3274),
.B(n_3245),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_SL g3415 ( 
.A(n_3240),
.B(n_819),
.Y(n_3415)
);

AOI21xp5_ASAP7_75t_L g3416 ( 
.A1(n_3318),
.A2(n_1461),
.B(n_1451),
.Y(n_3416)
);

INVx1_ASAP7_75t_L g3417 ( 
.A(n_3181),
.Y(n_3417)
);

A2O1A1Ixp33_ASAP7_75t_L g3418 ( 
.A1(n_3326),
.A2(n_3271),
.B(n_3269),
.C(n_3294),
.Y(n_3418)
);

BUFx2_ASAP7_75t_L g3419 ( 
.A(n_3189),
.Y(n_3419)
);

OAI22xp5_ASAP7_75t_L g3420 ( 
.A1(n_3273),
.A2(n_70),
.B1(n_67),
.B2(n_69),
.Y(n_3420)
);

OAI22xp5_ASAP7_75t_L g3421 ( 
.A1(n_3332),
.A2(n_74),
.B1(n_71),
.B2(n_73),
.Y(n_3421)
);

NAND2xp5_ASAP7_75t_L g3422 ( 
.A(n_3265),
.B(n_73),
.Y(n_3422)
);

AOI21xp5_ASAP7_75t_L g3423 ( 
.A1(n_3145),
.A2(n_1461),
.B(n_1451),
.Y(n_3423)
);

OR2x2_ASAP7_75t_L g3424 ( 
.A(n_3183),
.B(n_75),
.Y(n_3424)
);

INVx2_ASAP7_75t_L g3425 ( 
.A(n_3183),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_3206),
.Y(n_3426)
);

AND2x4_ASAP7_75t_L g3427 ( 
.A(n_3278),
.B(n_75),
.Y(n_3427)
);

AND2x2_ASAP7_75t_L g3428 ( 
.A(n_3218),
.B(n_3150),
.Y(n_3428)
);

INVxp67_ASAP7_75t_SL g3429 ( 
.A(n_3223),
.Y(n_3429)
);

INVx1_ASAP7_75t_SL g3430 ( 
.A(n_3253),
.Y(n_3430)
);

AND2x2_ASAP7_75t_L g3431 ( 
.A(n_3193),
.B(n_76),
.Y(n_3431)
);

OAI21xp33_ASAP7_75t_L g3432 ( 
.A1(n_3301),
.A2(n_76),
.B(n_77),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_L g3433 ( 
.A(n_3213),
.B(n_78),
.Y(n_3433)
);

OAI22xp5_ASAP7_75t_L g3434 ( 
.A1(n_3305),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_3434)
);

AOI22xp33_ASAP7_75t_L g3435 ( 
.A1(n_3340),
.A2(n_857),
.B1(n_867),
.B2(n_836),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_SL g3436 ( 
.A(n_3313),
.B(n_836),
.Y(n_3436)
);

AOI21xp5_ASAP7_75t_L g3437 ( 
.A1(n_3288),
.A2(n_1461),
.B(n_1451),
.Y(n_3437)
);

INVx2_ASAP7_75t_L g3438 ( 
.A(n_3213),
.Y(n_3438)
);

INVx1_ASAP7_75t_SL g3439 ( 
.A(n_3235),
.Y(n_3439)
);

INVx3_ASAP7_75t_L g3440 ( 
.A(n_3147),
.Y(n_3440)
);

BUFx12f_ASAP7_75t_L g3441 ( 
.A(n_3272),
.Y(n_3441)
);

AOI21xp33_ASAP7_75t_SL g3442 ( 
.A1(n_3317),
.A2(n_81),
.B(n_82),
.Y(n_3442)
);

INVxp67_ASAP7_75t_SL g3443 ( 
.A(n_3187),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_L g3444 ( 
.A(n_3231),
.B(n_83),
.Y(n_3444)
);

OAI22xp5_ASAP7_75t_L g3445 ( 
.A1(n_3325),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_3445)
);

OR2x2_ASAP7_75t_L g3446 ( 
.A(n_3254),
.B(n_84),
.Y(n_3446)
);

BUFx3_ASAP7_75t_L g3447 ( 
.A(n_3165),
.Y(n_3447)
);

INVxp67_ASAP7_75t_L g3448 ( 
.A(n_3296),
.Y(n_3448)
);

AOI21xp5_ASAP7_75t_L g3449 ( 
.A1(n_3337),
.A2(n_3281),
.B(n_3300),
.Y(n_3449)
);

INVx2_ASAP7_75t_SL g3450 ( 
.A(n_3167),
.Y(n_3450)
);

INVx1_ASAP7_75t_L g3451 ( 
.A(n_3206),
.Y(n_3451)
);

NAND2x1p5_ASAP7_75t_L g3452 ( 
.A(n_3209),
.B(n_857),
.Y(n_3452)
);

NOR2xp33_ASAP7_75t_L g3453 ( 
.A(n_3315),
.B(n_85),
.Y(n_3453)
);

NAND2x1p5_ASAP7_75t_L g3454 ( 
.A(n_3209),
.B(n_857),
.Y(n_3454)
);

CKINVDCx5p33_ASAP7_75t_R g3455 ( 
.A(n_3219),
.Y(n_3455)
);

AND2x2_ASAP7_75t_L g3456 ( 
.A(n_3151),
.B(n_87),
.Y(n_3456)
);

AND2x4_ASAP7_75t_L g3457 ( 
.A(n_3278),
.B(n_88),
.Y(n_3457)
);

INVx2_ASAP7_75t_L g3458 ( 
.A(n_3231),
.Y(n_3458)
);

A2O1A1Ixp33_ASAP7_75t_SL g3459 ( 
.A1(n_3254),
.A2(n_93),
.B(n_91),
.C(n_92),
.Y(n_3459)
);

INVx2_ASAP7_75t_SL g3460 ( 
.A(n_3162),
.Y(n_3460)
);

BUFx3_ASAP7_75t_L g3461 ( 
.A(n_3131),
.Y(n_3461)
);

INVx3_ASAP7_75t_L g3462 ( 
.A(n_3147),
.Y(n_3462)
);

OR2x6_ASAP7_75t_L g3463 ( 
.A(n_3195),
.B(n_857),
.Y(n_3463)
);

INVx2_ASAP7_75t_L g3464 ( 
.A(n_3234),
.Y(n_3464)
);

INVx6_ASAP7_75t_L g3465 ( 
.A(n_3177),
.Y(n_3465)
);

INVx1_ASAP7_75t_SL g3466 ( 
.A(n_3222),
.Y(n_3466)
);

OAI22xp5_ASAP7_75t_L g3467 ( 
.A1(n_3271),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_3467)
);

NAND2xp33_ASAP7_75t_L g3468 ( 
.A(n_3289),
.B(n_867),
.Y(n_3468)
);

OAI22xp5_ASAP7_75t_L g3469 ( 
.A1(n_3207),
.A2(n_94),
.B1(n_96),
.B2(n_98),
.Y(n_3469)
);

OR2x6_ASAP7_75t_L g3470 ( 
.A(n_3309),
.B(n_867),
.Y(n_3470)
);

OAI21xp5_ASAP7_75t_L g3471 ( 
.A1(n_3336),
.A2(n_99),
.B(n_100),
.Y(n_3471)
);

OAI22xp5_ASAP7_75t_SL g3472 ( 
.A1(n_3337),
.A2(n_99),
.B1(n_101),
.B2(n_103),
.Y(n_3472)
);

AND2x4_ASAP7_75t_L g3473 ( 
.A(n_3238),
.B(n_101),
.Y(n_3473)
);

INVxp67_ASAP7_75t_SL g3474 ( 
.A(n_3187),
.Y(n_3474)
);

OAI21xp5_ASAP7_75t_L g3475 ( 
.A1(n_3149),
.A2(n_104),
.B(n_105),
.Y(n_3475)
);

INVx4_ASAP7_75t_L g3476 ( 
.A(n_3232),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_L g3477 ( 
.A(n_3261),
.B(n_106),
.Y(n_3477)
);

AND2x2_ASAP7_75t_L g3478 ( 
.A(n_3199),
.B(n_106),
.Y(n_3478)
);

AOI22xp33_ASAP7_75t_L g3479 ( 
.A1(n_3340),
.A2(n_867),
.B1(n_108),
.B2(n_109),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_L g3480 ( 
.A(n_3234),
.B(n_3160),
.Y(n_3480)
);

NAND2x1p5_ASAP7_75t_L g3481 ( 
.A(n_3209),
.B(n_1431),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_3163),
.Y(n_3482)
);

AND2x2_ASAP7_75t_L g3483 ( 
.A(n_3280),
.B(n_107),
.Y(n_3483)
);

AND2x4_ASAP7_75t_L g3484 ( 
.A(n_3238),
.B(n_108),
.Y(n_3484)
);

NOR2xp67_ASAP7_75t_SL g3485 ( 
.A(n_3320),
.B(n_3311),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3184),
.Y(n_3486)
);

INVx2_ASAP7_75t_L g3487 ( 
.A(n_3201),
.Y(n_3487)
);

INVx2_ASAP7_75t_L g3488 ( 
.A(n_3233),
.Y(n_3488)
);

AOI21xp5_ASAP7_75t_L g3489 ( 
.A1(n_3281),
.A2(n_1431),
.B(n_110),
.Y(n_3489)
);

NOR2xp67_ASAP7_75t_SL g3490 ( 
.A(n_3320),
.B(n_1431),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_L g3491 ( 
.A(n_3261),
.B(n_112),
.Y(n_3491)
);

AND2x2_ASAP7_75t_L g3492 ( 
.A(n_3280),
.B(n_114),
.Y(n_3492)
);

AND2x4_ASAP7_75t_L g3493 ( 
.A(n_3249),
.B(n_114),
.Y(n_3493)
);

BUFx2_ASAP7_75t_SL g3494 ( 
.A(n_3211),
.Y(n_3494)
);

A2O1A1Ixp33_ASAP7_75t_L g3495 ( 
.A1(n_3292),
.A2(n_115),
.B(n_116),
.C(n_117),
.Y(n_3495)
);

BUFx6f_ASAP7_75t_L g3496 ( 
.A(n_3232),
.Y(n_3496)
);

INVx1_ASAP7_75t_L g3497 ( 
.A(n_3309),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_3210),
.Y(n_3498)
);

AOI221xp5_ASAP7_75t_L g3499 ( 
.A1(n_3263),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.C(n_119),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_L g3500 ( 
.A(n_3290),
.B(n_3252),
.Y(n_3500)
);

AND2x2_ASAP7_75t_L g3501 ( 
.A(n_3161),
.B(n_120),
.Y(n_3501)
);

INVx1_ASAP7_75t_L g3502 ( 
.A(n_3210),
.Y(n_3502)
);

AOI21xp5_ASAP7_75t_L g3503 ( 
.A1(n_3281),
.A2(n_1431),
.B(n_120),
.Y(n_3503)
);

INVx2_ASAP7_75t_L g3504 ( 
.A(n_3287),
.Y(n_3504)
);

INVx1_ASAP7_75t_L g3505 ( 
.A(n_3263),
.Y(n_3505)
);

OR2x2_ASAP7_75t_L g3506 ( 
.A(n_3310),
.B(n_3312),
.Y(n_3506)
);

A2O1A1Ixp33_ASAP7_75t_L g3507 ( 
.A1(n_3292),
.A2(n_121),
.B(n_123),
.C(n_124),
.Y(n_3507)
);

INVxp67_ASAP7_75t_L g3508 ( 
.A(n_3224),
.Y(n_3508)
);

BUFx12f_ASAP7_75t_L g3509 ( 
.A(n_3177),
.Y(n_3509)
);

CKINVDCx5p33_ASAP7_75t_R g3510 ( 
.A(n_3241),
.Y(n_3510)
);

CKINVDCx11_ASAP7_75t_R g3511 ( 
.A(n_3175),
.Y(n_3511)
);

INVx6_ASAP7_75t_L g3512 ( 
.A(n_3357),
.Y(n_3512)
);

INVx2_ASAP7_75t_L g3513 ( 
.A(n_3506),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_3351),
.Y(n_3514)
);

BUFx6f_ASAP7_75t_L g3515 ( 
.A(n_3496),
.Y(n_3515)
);

OAI21xp5_ASAP7_75t_L g3516 ( 
.A1(n_3355),
.A2(n_3180),
.B(n_3283),
.Y(n_3516)
);

OAI22xp33_ASAP7_75t_L g3517 ( 
.A1(n_3467),
.A2(n_3148),
.B1(n_3295),
.B2(n_3205),
.Y(n_3517)
);

INVx4_ASAP7_75t_L g3518 ( 
.A(n_3381),
.Y(n_3518)
);

OAI22xp5_ASAP7_75t_L g3519 ( 
.A1(n_3418),
.A2(n_3276),
.B1(n_3178),
.B2(n_3148),
.Y(n_3519)
);

CKINVDCx11_ASAP7_75t_R g3520 ( 
.A(n_3511),
.Y(n_3520)
);

AOI22xp33_ASAP7_75t_L g3521 ( 
.A1(n_3352),
.A2(n_3396),
.B1(n_3432),
.B2(n_3415),
.Y(n_3521)
);

CKINVDCx11_ASAP7_75t_R g3522 ( 
.A(n_3363),
.Y(n_3522)
);

INVx2_ASAP7_75t_L g3523 ( 
.A(n_3438),
.Y(n_3523)
);

AOI22xp33_ASAP7_75t_SL g3524 ( 
.A1(n_3396),
.A2(n_3276),
.B1(n_3129),
.B2(n_3341),
.Y(n_3524)
);

AOI22xp33_ASAP7_75t_SL g3525 ( 
.A1(n_3420),
.A2(n_3190),
.B1(n_3216),
.B2(n_3258),
.Y(n_3525)
);

OAI22x1_ASAP7_75t_L g3526 ( 
.A1(n_3430),
.A2(n_3310),
.B1(n_3312),
.B2(n_3295),
.Y(n_3526)
);

BUFx8_ASAP7_75t_L g3527 ( 
.A(n_3398),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_L g3528 ( 
.A(n_3429),
.B(n_3302),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_3364),
.Y(n_3529)
);

AOI22xp33_ASAP7_75t_L g3530 ( 
.A1(n_3432),
.A2(n_3328),
.B1(n_3264),
.B2(n_3327),
.Y(n_3530)
);

AOI22xp33_ASAP7_75t_L g3531 ( 
.A1(n_3434),
.A2(n_3328),
.B1(n_3264),
.B2(n_3275),
.Y(n_3531)
);

INVx3_ASAP7_75t_L g3532 ( 
.A(n_3360),
.Y(n_3532)
);

CKINVDCx5p33_ASAP7_75t_R g3533 ( 
.A(n_3354),
.Y(n_3533)
);

BUFx12f_ASAP7_75t_L g3534 ( 
.A(n_3395),
.Y(n_3534)
);

INVx8_ASAP7_75t_L g3535 ( 
.A(n_3509),
.Y(n_3535)
);

INVx1_ASAP7_75t_SL g3536 ( 
.A(n_3370),
.Y(n_3536)
);

AOI22xp33_ASAP7_75t_L g3537 ( 
.A1(n_3434),
.A2(n_3267),
.B1(n_3282),
.B2(n_3279),
.Y(n_3537)
);

CKINVDCx5p33_ASAP7_75t_R g3538 ( 
.A(n_3407),
.Y(n_3538)
);

INVx4_ASAP7_75t_L g3539 ( 
.A(n_3510),
.Y(n_3539)
);

CKINVDCx20_ASAP7_75t_R g3540 ( 
.A(n_3455),
.Y(n_3540)
);

CKINVDCx6p67_ASAP7_75t_R g3541 ( 
.A(n_3441),
.Y(n_3541)
);

BUFx2_ASAP7_75t_L g3542 ( 
.A(n_3419),
.Y(n_3542)
);

CKINVDCx5p33_ASAP7_75t_R g3543 ( 
.A(n_3366),
.Y(n_3543)
);

INVx2_ASAP7_75t_L g3544 ( 
.A(n_3458),
.Y(n_3544)
);

OAI22xp33_ASAP7_75t_L g3545 ( 
.A1(n_3467),
.A2(n_3205),
.B1(n_3196),
.B2(n_3256),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_3365),
.Y(n_3546)
);

AOI22xp33_ASAP7_75t_L g3547 ( 
.A1(n_3342),
.A2(n_3282),
.B1(n_3279),
.B2(n_3168),
.Y(n_3547)
);

INVx6_ASAP7_75t_L g3548 ( 
.A(n_3357),
.Y(n_3548)
);

INVx1_ASAP7_75t_L g3549 ( 
.A(n_3367),
.Y(n_3549)
);

INVx2_ASAP7_75t_L g3550 ( 
.A(n_3464),
.Y(n_3550)
);

AOI22xp33_ASAP7_75t_L g3551 ( 
.A1(n_3342),
.A2(n_3282),
.B1(n_3279),
.B2(n_3168),
.Y(n_3551)
);

BUFx2_ASAP7_75t_L g3552 ( 
.A(n_3508),
.Y(n_3552)
);

AOI22xp33_ASAP7_75t_L g3553 ( 
.A1(n_3342),
.A2(n_3260),
.B1(n_3130),
.B2(n_3257),
.Y(n_3553)
);

INVx1_ASAP7_75t_SL g3554 ( 
.A(n_3370),
.Y(n_3554)
);

AOI22xp33_ASAP7_75t_L g3555 ( 
.A1(n_3342),
.A2(n_3130),
.B1(n_3277),
.B2(n_3304),
.Y(n_3555)
);

BUFx2_ASAP7_75t_L g3556 ( 
.A(n_3406),
.Y(n_3556)
);

BUFx4f_ASAP7_75t_SL g3557 ( 
.A(n_3344),
.Y(n_3557)
);

AOI22xp33_ASAP7_75t_L g3558 ( 
.A1(n_3420),
.A2(n_3277),
.B1(n_3304),
.B2(n_3174),
.Y(n_3558)
);

INVx2_ASAP7_75t_L g3559 ( 
.A(n_3392),
.Y(n_3559)
);

BUFx12f_ASAP7_75t_L g3560 ( 
.A(n_3346),
.Y(n_3560)
);

INVx1_ASAP7_75t_L g3561 ( 
.A(n_3378),
.Y(n_3561)
);

AOI22xp33_ASAP7_75t_SL g3562 ( 
.A1(n_3471),
.A2(n_3237),
.B1(n_3200),
.B2(n_3256),
.Y(n_3562)
);

OAI22xp33_ASAP7_75t_L g3563 ( 
.A1(n_3475),
.A2(n_3268),
.B1(n_3256),
.B2(n_3303),
.Y(n_3563)
);

INVx1_ASAP7_75t_L g3564 ( 
.A(n_3382),
.Y(n_3564)
);

INVx2_ASAP7_75t_L g3565 ( 
.A(n_3425),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_3387),
.Y(n_3566)
);

INVx2_ASAP7_75t_L g3567 ( 
.A(n_3373),
.Y(n_3567)
);

AOI22xp33_ASAP7_75t_L g3568 ( 
.A1(n_3475),
.A2(n_3255),
.B1(n_3293),
.B2(n_3249),
.Y(n_3568)
);

AOI22xp33_ASAP7_75t_L g3569 ( 
.A1(n_3499),
.A2(n_3138),
.B1(n_3228),
.B2(n_3227),
.Y(n_3569)
);

INVx6_ASAP7_75t_L g3570 ( 
.A(n_3357),
.Y(n_3570)
);

CKINVDCx5p33_ASAP7_75t_R g3571 ( 
.A(n_3447),
.Y(n_3571)
);

OAI22xp5_ASAP7_75t_L g3572 ( 
.A1(n_3472),
.A2(n_3202),
.B1(n_3329),
.B2(n_3247),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_3497),
.B(n_3297),
.Y(n_3573)
);

INVx2_ASAP7_75t_L g3574 ( 
.A(n_3409),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_3417),
.Y(n_3575)
);

AOI22xp33_ASAP7_75t_L g3576 ( 
.A1(n_3471),
.A2(n_3227),
.B1(n_3242),
.B2(n_3228),
.Y(n_3576)
);

CKINVDCx6p67_ASAP7_75t_R g3577 ( 
.A(n_3461),
.Y(n_3577)
);

OAI22xp33_ASAP7_75t_L g3578 ( 
.A1(n_3442),
.A2(n_3268),
.B1(n_3259),
.B2(n_3248),
.Y(n_3578)
);

OAI22xp5_ASAP7_75t_L g3579 ( 
.A1(n_3472),
.A2(n_3507),
.B1(n_3495),
.B2(n_3405),
.Y(n_3579)
);

BUFx12f_ASAP7_75t_L g3580 ( 
.A(n_3456),
.Y(n_3580)
);

AOI22xp33_ASAP7_75t_L g3581 ( 
.A1(n_3421),
.A2(n_3242),
.B1(n_3259),
.B2(n_3285),
.Y(n_3581)
);

INVx2_ASAP7_75t_L g3582 ( 
.A(n_3439),
.Y(n_3582)
);

INVx3_ASAP7_75t_L g3583 ( 
.A(n_3360),
.Y(n_3583)
);

AOI22xp5_ASAP7_75t_L g3584 ( 
.A1(n_3468),
.A2(n_3262),
.B1(n_3159),
.B2(n_3236),
.Y(n_3584)
);

AOI22xp33_ASAP7_75t_L g3585 ( 
.A1(n_3421),
.A2(n_3445),
.B1(n_3485),
.B2(n_3479),
.Y(n_3585)
);

INVxp67_ASAP7_75t_SL g3586 ( 
.A(n_3443),
.Y(n_3586)
);

AOI22xp33_ASAP7_75t_L g3587 ( 
.A1(n_3445),
.A2(n_3226),
.B1(n_3144),
.B2(n_3339),
.Y(n_3587)
);

NAND2x1p5_ASAP7_75t_L g3588 ( 
.A(n_3490),
.B(n_3268),
.Y(n_3588)
);

INVx1_ASAP7_75t_L g3589 ( 
.A(n_3498),
.Y(n_3589)
);

INVx1_ASAP7_75t_L g3590 ( 
.A(n_3502),
.Y(n_3590)
);

NAND2xp5_ASAP7_75t_L g3591 ( 
.A(n_3505),
.B(n_3474),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_L g3592 ( 
.A(n_3482),
.B(n_3299),
.Y(n_3592)
);

INVx1_ASAP7_75t_L g3593 ( 
.A(n_3426),
.Y(n_3593)
);

INVx1_ASAP7_75t_SL g3594 ( 
.A(n_3494),
.Y(n_3594)
);

OAI22xp5_ASAP7_75t_L g3595 ( 
.A1(n_3442),
.A2(n_3226),
.B1(n_3333),
.B2(n_3266),
.Y(n_3595)
);

BUFx6f_ASAP7_75t_L g3596 ( 
.A(n_3496),
.Y(n_3596)
);

OAI21xp33_ASAP7_75t_L g3597 ( 
.A1(n_3449),
.A2(n_3321),
.B(n_3246),
.Y(n_3597)
);

BUFx2_ASAP7_75t_L g3598 ( 
.A(n_3466),
.Y(n_3598)
);

BUFx6f_ASAP7_75t_L g3599 ( 
.A(n_3496),
.Y(n_3599)
);

INVx6_ASAP7_75t_L g3600 ( 
.A(n_3476),
.Y(n_3600)
);

AND2x2_ASAP7_75t_L g3601 ( 
.A(n_3376),
.B(n_3161),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_3451),
.Y(n_3602)
);

BUFx8_ASAP7_75t_SL g3603 ( 
.A(n_3473),
.Y(n_3603)
);

BUFx10_ASAP7_75t_L g3604 ( 
.A(n_3388),
.Y(n_3604)
);

NAND2xp5_ASAP7_75t_L g3605 ( 
.A(n_3486),
.B(n_3338),
.Y(n_3605)
);

INVx1_ASAP7_75t_SL g3606 ( 
.A(n_3500),
.Y(n_3606)
);

AOI22xp33_ASAP7_75t_L g3607 ( 
.A1(n_3469),
.A2(n_3339),
.B1(n_3230),
.B2(n_3185),
.Y(n_3607)
);

BUFx3_ASAP7_75t_L g3608 ( 
.A(n_3450),
.Y(n_3608)
);

BUFx2_ASAP7_75t_SL g3609 ( 
.A(n_3460),
.Y(n_3609)
);

AOI22xp33_ASAP7_75t_L g3610 ( 
.A1(n_3469),
.A2(n_3339),
.B1(n_3185),
.B2(n_3330),
.Y(n_3610)
);

NAND2xp5_ASAP7_75t_L g3611 ( 
.A(n_3379),
.B(n_3314),
.Y(n_3611)
);

NAND2xp5_ASAP7_75t_L g3612 ( 
.A(n_3380),
.B(n_3314),
.Y(n_3612)
);

HB1xp67_ASAP7_75t_L g3613 ( 
.A(n_3376),
.Y(n_3613)
);

CKINVDCx11_ASAP7_75t_R g3614 ( 
.A(n_3350),
.Y(n_3614)
);

INVx3_ASAP7_75t_SL g3615 ( 
.A(n_3427),
.Y(n_3615)
);

INVx1_ASAP7_75t_L g3616 ( 
.A(n_3480),
.Y(n_3616)
);

INVx8_ASAP7_75t_L g3617 ( 
.A(n_3473),
.Y(n_3617)
);

CKINVDCx11_ASAP7_75t_R g3618 ( 
.A(n_3350),
.Y(n_3618)
);

CKINVDCx20_ASAP7_75t_R g3619 ( 
.A(n_3428),
.Y(n_3619)
);

BUFx8_ASAP7_75t_L g3620 ( 
.A(n_3478),
.Y(n_3620)
);

AOI22xp33_ASAP7_75t_L g3621 ( 
.A1(n_3448),
.A2(n_3330),
.B1(n_3250),
.B2(n_3182),
.Y(n_3621)
);

CKINVDCx11_ASAP7_75t_R g3622 ( 
.A(n_3350),
.Y(n_3622)
);

AOI22xp33_ASAP7_75t_L g3623 ( 
.A1(n_3348),
.A2(n_3343),
.B1(n_3349),
.B2(n_3356),
.Y(n_3623)
);

BUFx4f_ASAP7_75t_SL g3624 ( 
.A(n_3372),
.Y(n_3624)
);

INVx1_ASAP7_75t_L g3625 ( 
.A(n_3384),
.Y(n_3625)
);

AND2x2_ASAP7_75t_L g3626 ( 
.A(n_3439),
.B(n_3251),
.Y(n_3626)
);

CKINVDCx6p67_ASAP7_75t_R g3627 ( 
.A(n_3374),
.Y(n_3627)
);

INVx1_ASAP7_75t_L g3628 ( 
.A(n_3487),
.Y(n_3628)
);

INVx2_ASAP7_75t_L g3629 ( 
.A(n_3466),
.Y(n_3629)
);

CKINVDCx20_ASAP7_75t_R g3630 ( 
.A(n_3383),
.Y(n_3630)
);

CKINVDCx20_ASAP7_75t_R g3631 ( 
.A(n_3390),
.Y(n_3631)
);

INVx1_ASAP7_75t_SL g3632 ( 
.A(n_3430),
.Y(n_3632)
);

CKINVDCx5p33_ASAP7_75t_R g3633 ( 
.A(n_3371),
.Y(n_3633)
);

AOI22xp33_ASAP7_75t_SL g3634 ( 
.A1(n_3401),
.A2(n_3248),
.B1(n_3251),
.B2(n_3177),
.Y(n_3634)
);

AOI22xp33_ASAP7_75t_L g3635 ( 
.A1(n_3356),
.A2(n_3330),
.B1(n_3142),
.B2(n_3182),
.Y(n_3635)
);

AOI22xp33_ASAP7_75t_SL g3636 ( 
.A1(n_3401),
.A2(n_3204),
.B1(n_3142),
.B2(n_3139),
.Y(n_3636)
);

AOI22xp33_ASAP7_75t_L g3637 ( 
.A1(n_3356),
.A2(n_3427),
.B1(n_3457),
.B2(n_3453),
.Y(n_3637)
);

BUFx2_ASAP7_75t_L g3638 ( 
.A(n_3411),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3488),
.Y(n_3639)
);

INVx4_ASAP7_75t_L g3640 ( 
.A(n_3371),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3414),
.Y(n_3641)
);

OAI22xp5_ASAP7_75t_L g3642 ( 
.A1(n_3399),
.A2(n_3323),
.B1(n_3172),
.B2(n_3169),
.Y(n_3642)
);

AOI22xp33_ASAP7_75t_L g3643 ( 
.A1(n_3457),
.A2(n_3232),
.B1(n_3307),
.B2(n_3172),
.Y(n_3643)
);

BUFx12f_ASAP7_75t_L g3644 ( 
.A(n_3394),
.Y(n_3644)
);

INVx2_ASAP7_75t_L g3645 ( 
.A(n_3411),
.Y(n_3645)
);

INVx2_ASAP7_75t_L g3646 ( 
.A(n_3440),
.Y(n_3646)
);

INVx2_ASAP7_75t_L g3647 ( 
.A(n_3589),
.Y(n_3647)
);

OA21x2_ASAP7_75t_L g3648 ( 
.A1(n_3597),
.A2(n_3491),
.B(n_3477),
.Y(n_3648)
);

INVx2_ASAP7_75t_L g3649 ( 
.A(n_3590),
.Y(n_3649)
);

BUFx3_ASAP7_75t_L g3650 ( 
.A(n_3520),
.Y(n_3650)
);

OAI21xp5_ASAP7_75t_L g3651 ( 
.A1(n_3524),
.A2(n_3404),
.B(n_3397),
.Y(n_3651)
);

HB1xp67_ASAP7_75t_L g3652 ( 
.A(n_3613),
.Y(n_3652)
);

INVx2_ASAP7_75t_L g3653 ( 
.A(n_3574),
.Y(n_3653)
);

INVx1_ASAP7_75t_L g3654 ( 
.A(n_3605),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_3605),
.Y(n_3655)
);

INVx1_ASAP7_75t_L g3656 ( 
.A(n_3514),
.Y(n_3656)
);

INVx3_ASAP7_75t_L g3657 ( 
.A(n_3512),
.Y(n_3657)
);

INVx1_ASAP7_75t_L g3658 ( 
.A(n_3529),
.Y(n_3658)
);

INVx2_ASAP7_75t_L g3659 ( 
.A(n_3546),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_3549),
.Y(n_3660)
);

HB1xp67_ASAP7_75t_L g3661 ( 
.A(n_3598),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_L g3662 ( 
.A(n_3606),
.B(n_3389),
.Y(n_3662)
);

INVx2_ASAP7_75t_L g3663 ( 
.A(n_3561),
.Y(n_3663)
);

BUFx2_ASAP7_75t_L g3664 ( 
.A(n_3512),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_L g3665 ( 
.A(n_3536),
.B(n_3477),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_3564),
.Y(n_3666)
);

INVx1_ASAP7_75t_L g3667 ( 
.A(n_3566),
.Y(n_3667)
);

AND2x4_ASAP7_75t_L g3668 ( 
.A(n_3586),
.B(n_3440),
.Y(n_3668)
);

INVxp67_ASAP7_75t_SL g3669 ( 
.A(n_3526),
.Y(n_3669)
);

INVx3_ASAP7_75t_L g3670 ( 
.A(n_3512),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3575),
.Y(n_3671)
);

INVx1_ASAP7_75t_L g3672 ( 
.A(n_3586),
.Y(n_3672)
);

INVx2_ASAP7_75t_L g3673 ( 
.A(n_3611),
.Y(n_3673)
);

AND2x2_ASAP7_75t_L g3674 ( 
.A(n_3542),
.B(n_3462),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_3591),
.Y(n_3675)
);

OR2x6_ASAP7_75t_L g3676 ( 
.A(n_3588),
.B(n_3470),
.Y(n_3676)
);

NOR2xp33_ASAP7_75t_L g3677 ( 
.A(n_3518),
.B(n_3393),
.Y(n_3677)
);

AND2x2_ASAP7_75t_L g3678 ( 
.A(n_3626),
.B(n_3462),
.Y(n_3678)
);

BUFx2_ASAP7_75t_L g3679 ( 
.A(n_3548),
.Y(n_3679)
);

AOI21x1_ASAP7_75t_L g3680 ( 
.A1(n_3528),
.A2(n_3491),
.B(n_3611),
.Y(n_3680)
);

OAI22xp5_ASAP7_75t_L g3681 ( 
.A1(n_3524),
.A2(n_3463),
.B1(n_3446),
.B2(n_3412),
.Y(n_3681)
);

HB1xp67_ASAP7_75t_L g3682 ( 
.A(n_3528),
.Y(n_3682)
);

OAI22xp33_ASAP7_75t_L g3683 ( 
.A1(n_3579),
.A2(n_3463),
.B1(n_3470),
.B2(n_3358),
.Y(n_3683)
);

INVx2_ASAP7_75t_L g3684 ( 
.A(n_3612),
.Y(n_3684)
);

BUFx3_ASAP7_75t_L g3685 ( 
.A(n_3534),
.Y(n_3685)
);

INVx2_ASAP7_75t_L g3686 ( 
.A(n_3612),
.Y(n_3686)
);

NAND2x1_ASAP7_75t_L g3687 ( 
.A(n_3548),
.B(n_3470),
.Y(n_3687)
);

OAI21xp5_ASAP7_75t_L g3688 ( 
.A1(n_3579),
.A2(n_3413),
.B(n_3399),
.Y(n_3688)
);

AOI21x1_ASAP7_75t_L g3689 ( 
.A1(n_3519),
.A2(n_3412),
.B(n_3402),
.Y(n_3689)
);

OAI21xp5_ASAP7_75t_L g3690 ( 
.A1(n_3519),
.A2(n_3413),
.B(n_3402),
.Y(n_3690)
);

AND2x4_ASAP7_75t_L g3691 ( 
.A(n_3532),
.B(n_3504),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_3593),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_3602),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3591),
.Y(n_3694)
);

OAI221xp5_ASAP7_75t_SL g3695 ( 
.A1(n_3521),
.A2(n_3361),
.B1(n_3424),
.B2(n_3362),
.C(n_3408),
.Y(n_3695)
);

AOI22xp5_ASAP7_75t_L g3696 ( 
.A1(n_3595),
.A2(n_3369),
.B1(n_3493),
.B2(n_3484),
.Y(n_3696)
);

INVx2_ASAP7_75t_L g3697 ( 
.A(n_3513),
.Y(n_3697)
);

OAI21xp5_ASAP7_75t_L g3698 ( 
.A1(n_3562),
.A2(n_3368),
.B(n_3422),
.Y(n_3698)
);

INVx2_ASAP7_75t_L g3699 ( 
.A(n_3523),
.Y(n_3699)
);

AND2x4_ASAP7_75t_L g3700 ( 
.A(n_3532),
.B(n_3476),
.Y(n_3700)
);

INVx2_ASAP7_75t_L g3701 ( 
.A(n_3544),
.Y(n_3701)
);

INVx1_ASAP7_75t_L g3702 ( 
.A(n_3616),
.Y(n_3702)
);

INVxp67_ASAP7_75t_L g3703 ( 
.A(n_3552),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_3641),
.Y(n_3704)
);

NAND2x1p5_ASAP7_75t_L g3705 ( 
.A(n_3554),
.B(n_3345),
.Y(n_3705)
);

AOI22xp33_ASAP7_75t_SL g3706 ( 
.A1(n_3516),
.A2(n_3484),
.B1(n_3493),
.B2(n_3431),
.Y(n_3706)
);

INVx1_ASAP7_75t_L g3707 ( 
.A(n_3592),
.Y(n_3707)
);

INVx3_ASAP7_75t_L g3708 ( 
.A(n_3548),
.Y(n_3708)
);

AOI21xp33_ASAP7_75t_SL g3709 ( 
.A1(n_3535),
.A2(n_3444),
.B(n_3433),
.Y(n_3709)
);

INVx1_ASAP7_75t_L g3710 ( 
.A(n_3592),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_L g3711 ( 
.A(n_3632),
.B(n_3359),
.Y(n_3711)
);

AND2x2_ASAP7_75t_L g3712 ( 
.A(n_3601),
.B(n_3347),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_L g3713 ( 
.A(n_3582),
.B(n_3483),
.Y(n_3713)
);

AND2x2_ASAP7_75t_L g3714 ( 
.A(n_3556),
.B(n_3377),
.Y(n_3714)
);

INVx2_ASAP7_75t_L g3715 ( 
.A(n_3550),
.Y(n_3715)
);

INVx2_ASAP7_75t_SL g3716 ( 
.A(n_3570),
.Y(n_3716)
);

INVx2_ASAP7_75t_L g3717 ( 
.A(n_3559),
.Y(n_3717)
);

OAI22xp5_ASAP7_75t_L g3718 ( 
.A1(n_3585),
.A2(n_3463),
.B1(n_3465),
.B2(n_3377),
.Y(n_3718)
);

INVx1_ASAP7_75t_L g3719 ( 
.A(n_3625),
.Y(n_3719)
);

CKINVDCx20_ASAP7_75t_R g3720 ( 
.A(n_3540),
.Y(n_3720)
);

BUFx2_ASAP7_75t_L g3721 ( 
.A(n_3570),
.Y(n_3721)
);

INVx1_ASAP7_75t_L g3722 ( 
.A(n_3628),
.Y(n_3722)
);

INVx2_ASAP7_75t_L g3723 ( 
.A(n_3565),
.Y(n_3723)
);

INVx2_ASAP7_75t_L g3724 ( 
.A(n_3573),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3639),
.Y(n_3725)
);

AOI22xp33_ASAP7_75t_L g3726 ( 
.A1(n_3516),
.A2(n_3465),
.B1(n_3385),
.B2(n_3436),
.Y(n_3726)
);

INVx2_ASAP7_75t_L g3727 ( 
.A(n_3573),
.Y(n_3727)
);

INVx2_ASAP7_75t_L g3728 ( 
.A(n_3567),
.Y(n_3728)
);

AO21x1_ASAP7_75t_L g3729 ( 
.A1(n_3578),
.A2(n_3503),
.B(n_3489),
.Y(n_3729)
);

INVx3_ASAP7_75t_L g3730 ( 
.A(n_3570),
.Y(n_3730)
);

CKINVDCx5p33_ASAP7_75t_R g3731 ( 
.A(n_3522),
.Y(n_3731)
);

INVx1_ASAP7_75t_L g3732 ( 
.A(n_3629),
.Y(n_3732)
);

INVx2_ASAP7_75t_L g3733 ( 
.A(n_3583),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_3638),
.Y(n_3734)
);

OAI21x1_ASAP7_75t_L g3735 ( 
.A1(n_3635),
.A2(n_3423),
.B(n_3307),
.Y(n_3735)
);

INVx2_ASAP7_75t_SL g3736 ( 
.A(n_3600),
.Y(n_3736)
);

INVx1_ASAP7_75t_L g3737 ( 
.A(n_3645),
.Y(n_3737)
);

HB1xp67_ASAP7_75t_L g3738 ( 
.A(n_3646),
.Y(n_3738)
);

AND2x4_ASAP7_75t_L g3739 ( 
.A(n_3583),
.B(n_3386),
.Y(n_3739)
);

AND2x2_ASAP7_75t_L g3740 ( 
.A(n_3623),
.B(n_3386),
.Y(n_3740)
);

INVx4_ASAP7_75t_L g3741 ( 
.A(n_3518),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3609),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_L g3743 ( 
.A(n_3562),
.B(n_3492),
.Y(n_3743)
);

AND2x2_ASAP7_75t_L g3744 ( 
.A(n_3594),
.B(n_3371),
.Y(n_3744)
);

BUFx3_ASAP7_75t_L g3745 ( 
.A(n_3603),
.Y(n_3745)
);

HB1xp67_ASAP7_75t_L g3746 ( 
.A(n_3619),
.Y(n_3746)
);

BUFx3_ASAP7_75t_L g3747 ( 
.A(n_3560),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3600),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3600),
.Y(n_3749)
);

HB1xp67_ASAP7_75t_L g3750 ( 
.A(n_3608),
.Y(n_3750)
);

INVx1_ASAP7_75t_L g3751 ( 
.A(n_3515),
.Y(n_3751)
);

HB1xp67_ASAP7_75t_L g3752 ( 
.A(n_3515),
.Y(n_3752)
);

CKINVDCx20_ASAP7_75t_R g3753 ( 
.A(n_3557),
.Y(n_3753)
);

BUFx3_ASAP7_75t_L g3754 ( 
.A(n_3577),
.Y(n_3754)
);

INVx2_ASAP7_75t_L g3755 ( 
.A(n_3640),
.Y(n_3755)
);

AOI22xp5_ASAP7_75t_L g3756 ( 
.A1(n_3595),
.A2(n_3501),
.B1(n_3391),
.B2(n_3403),
.Y(n_3756)
);

BUFx3_ASAP7_75t_L g3757 ( 
.A(n_3535),
.Y(n_3757)
);

INVx2_ASAP7_75t_L g3758 ( 
.A(n_3640),
.Y(n_3758)
);

INVx1_ASAP7_75t_L g3759 ( 
.A(n_3634),
.Y(n_3759)
);

INVx2_ASAP7_75t_L g3760 ( 
.A(n_3515),
.Y(n_3760)
);

AO21x1_ASAP7_75t_SL g3761 ( 
.A1(n_3610),
.A2(n_3435),
.B(n_3459),
.Y(n_3761)
);

INVx2_ASAP7_75t_L g3762 ( 
.A(n_3596),
.Y(n_3762)
);

OR2x2_ASAP7_75t_L g3763 ( 
.A(n_3634),
.B(n_3353),
.Y(n_3763)
);

AOI222xp33_ASAP7_75t_L g3764 ( 
.A1(n_3572),
.A2(n_121),
.B1(n_124),
.B2(n_125),
.C1(n_127),
.C2(n_128),
.Y(n_3764)
);

INVx2_ASAP7_75t_L g3765 ( 
.A(n_3596),
.Y(n_3765)
);

OAI21x1_ASAP7_75t_L g3766 ( 
.A1(n_3588),
.A2(n_3353),
.B(n_3400),
.Y(n_3766)
);

INVx1_ASAP7_75t_L g3767 ( 
.A(n_3596),
.Y(n_3767)
);

OAI22xp33_ASAP7_75t_L g3768 ( 
.A1(n_3545),
.A2(n_3375),
.B1(n_3391),
.B2(n_3416),
.Y(n_3768)
);

INVx1_ASAP7_75t_L g3769 ( 
.A(n_3599),
.Y(n_3769)
);

INVx2_ASAP7_75t_L g3770 ( 
.A(n_3599),
.Y(n_3770)
);

BUFx4f_ASAP7_75t_L g3771 ( 
.A(n_3541),
.Y(n_3771)
);

INVx2_ASAP7_75t_L g3772 ( 
.A(n_3599),
.Y(n_3772)
);

INVx1_ASAP7_75t_L g3773 ( 
.A(n_3647),
.Y(n_3773)
);

INVx1_ASAP7_75t_L g3774 ( 
.A(n_3647),
.Y(n_3774)
);

INVx2_ASAP7_75t_L g3775 ( 
.A(n_3649),
.Y(n_3775)
);

OAI21x1_ASAP7_75t_L g3776 ( 
.A1(n_3705),
.A2(n_3621),
.B(n_3643),
.Y(n_3776)
);

NAND2xp5_ASAP7_75t_L g3777 ( 
.A(n_3698),
.B(n_3525),
.Y(n_3777)
);

INVx2_ASAP7_75t_L g3778 ( 
.A(n_3649),
.Y(n_3778)
);

CKINVDCx20_ASAP7_75t_R g3779 ( 
.A(n_3720),
.Y(n_3779)
);

BUFx2_ASAP7_75t_L g3780 ( 
.A(n_3741),
.Y(n_3780)
);

INVx2_ASAP7_75t_L g3781 ( 
.A(n_3659),
.Y(n_3781)
);

AND2x4_ASAP7_75t_L g3782 ( 
.A(n_3664),
.B(n_3637),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_3659),
.Y(n_3783)
);

AOI22xp33_ASAP7_75t_L g3784 ( 
.A1(n_3651),
.A2(n_3563),
.B1(n_3572),
.B2(n_3604),
.Y(n_3784)
);

CKINVDCx6p67_ASAP7_75t_R g3785 ( 
.A(n_3650),
.Y(n_3785)
);

INVx2_ASAP7_75t_L g3786 ( 
.A(n_3663),
.Y(n_3786)
);

AND2x2_ASAP7_75t_L g3787 ( 
.A(n_3657),
.B(n_3627),
.Y(n_3787)
);

INVx2_ASAP7_75t_L g3788 ( 
.A(n_3663),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3656),
.Y(n_3789)
);

BUFx12f_ASAP7_75t_SL g3790 ( 
.A(n_3741),
.Y(n_3790)
);

NAND2xp5_ASAP7_75t_L g3791 ( 
.A(n_3648),
.B(n_3525),
.Y(n_3791)
);

OAI21x1_ASAP7_75t_L g3792 ( 
.A1(n_3705),
.A2(n_3553),
.B(n_3642),
.Y(n_3792)
);

INVx3_ASAP7_75t_L g3793 ( 
.A(n_3741),
.Y(n_3793)
);

INVx2_ASAP7_75t_L g3794 ( 
.A(n_3653),
.Y(n_3794)
);

OAI21x1_ASAP7_75t_L g3795 ( 
.A1(n_3705),
.A2(n_3642),
.B(n_3551),
.Y(n_3795)
);

AO21x2_ASAP7_75t_L g3796 ( 
.A1(n_3759),
.A2(n_3763),
.B(n_3690),
.Y(n_3796)
);

AND2x2_ASAP7_75t_L g3797 ( 
.A(n_3657),
.B(n_3615),
.Y(n_3797)
);

AND2x2_ASAP7_75t_L g3798 ( 
.A(n_3657),
.B(n_3615),
.Y(n_3798)
);

INVx1_ASAP7_75t_L g3799 ( 
.A(n_3658),
.Y(n_3799)
);

AO21x2_ASAP7_75t_L g3800 ( 
.A1(n_3759),
.A2(n_3437),
.B(n_3517),
.Y(n_3800)
);

NAND2xp5_ASAP7_75t_L g3801 ( 
.A(n_3648),
.B(n_3636),
.Y(n_3801)
);

OR2x2_ASAP7_75t_L g3802 ( 
.A(n_3682),
.B(n_3636),
.Y(n_3802)
);

HB1xp67_ASAP7_75t_L g3803 ( 
.A(n_3652),
.Y(n_3803)
);

INVx1_ASAP7_75t_L g3804 ( 
.A(n_3660),
.Y(n_3804)
);

INVx1_ASAP7_75t_L g3805 ( 
.A(n_3666),
.Y(n_3805)
);

HB1xp67_ASAP7_75t_L g3806 ( 
.A(n_3661),
.Y(n_3806)
);

HB1xp67_ASAP7_75t_L g3807 ( 
.A(n_3672),
.Y(n_3807)
);

OR2x2_ASAP7_75t_L g3808 ( 
.A(n_3675),
.B(n_3654),
.Y(n_3808)
);

INVx2_ASAP7_75t_L g3809 ( 
.A(n_3653),
.Y(n_3809)
);

INVx2_ASAP7_75t_L g3810 ( 
.A(n_3699),
.Y(n_3810)
);

AO21x2_ASAP7_75t_L g3811 ( 
.A1(n_3763),
.A2(n_3410),
.B(n_3584),
.Y(n_3811)
);

INVx2_ASAP7_75t_L g3812 ( 
.A(n_3699),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3667),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_3671),
.Y(n_3814)
);

INVx2_ASAP7_75t_L g3815 ( 
.A(n_3701),
.Y(n_3815)
);

OA21x2_ASAP7_75t_L g3816 ( 
.A1(n_3735),
.A2(n_3607),
.B(n_3587),
.Y(n_3816)
);

BUFx2_ASAP7_75t_L g3817 ( 
.A(n_3664),
.Y(n_3817)
);

AND2x2_ASAP7_75t_L g3818 ( 
.A(n_3670),
.B(n_3708),
.Y(n_3818)
);

AND2x2_ASAP7_75t_L g3819 ( 
.A(n_3670),
.B(n_3708),
.Y(n_3819)
);

INVx3_ASAP7_75t_L g3820 ( 
.A(n_3670),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_3692),
.Y(n_3821)
);

OAI21x1_ASAP7_75t_L g3822 ( 
.A1(n_3680),
.A2(n_3547),
.B(n_3530),
.Y(n_3822)
);

OAI21x1_ASAP7_75t_L g3823 ( 
.A1(n_3680),
.A2(n_3555),
.B(n_3581),
.Y(n_3823)
);

INVx1_ASAP7_75t_SL g3824 ( 
.A(n_3679),
.Y(n_3824)
);

INVx1_ASAP7_75t_L g3825 ( 
.A(n_3693),
.Y(n_3825)
);

INVx1_ASAP7_75t_L g3826 ( 
.A(n_3672),
.Y(n_3826)
);

INVx2_ASAP7_75t_SL g3827 ( 
.A(n_3757),
.Y(n_3827)
);

INVx3_ASAP7_75t_L g3828 ( 
.A(n_3708),
.Y(n_3828)
);

INVx2_ASAP7_75t_L g3829 ( 
.A(n_3701),
.Y(n_3829)
);

INVx2_ASAP7_75t_L g3830 ( 
.A(n_3715),
.Y(n_3830)
);

AND2x2_ASAP7_75t_L g3831 ( 
.A(n_3730),
.B(n_3604),
.Y(n_3831)
);

INVx2_ASAP7_75t_L g3832 ( 
.A(n_3715),
.Y(n_3832)
);

AND2x2_ASAP7_75t_L g3833 ( 
.A(n_3730),
.B(n_3633),
.Y(n_3833)
);

INVx1_ASAP7_75t_L g3834 ( 
.A(n_3719),
.Y(n_3834)
);

INVx2_ASAP7_75t_L g3835 ( 
.A(n_3717),
.Y(n_3835)
);

INVx2_ASAP7_75t_L g3836 ( 
.A(n_3717),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_L g3837 ( 
.A(n_3648),
.B(n_3630),
.Y(n_3837)
);

OR2x2_ASAP7_75t_L g3838 ( 
.A(n_3675),
.B(n_3655),
.Y(n_3838)
);

OAI21x1_ASAP7_75t_SL g3839 ( 
.A1(n_3688),
.A2(n_3539),
.B(n_3576),
.Y(n_3839)
);

INVx1_ASAP7_75t_L g3840 ( 
.A(n_3722),
.Y(n_3840)
);

INVx2_ASAP7_75t_L g3841 ( 
.A(n_3723),
.Y(n_3841)
);

NAND2xp5_ASAP7_75t_L g3842 ( 
.A(n_3703),
.B(n_3617),
.Y(n_3842)
);

AND2x2_ASAP7_75t_L g3843 ( 
.A(n_3730),
.B(n_3614),
.Y(n_3843)
);

INVx1_ASAP7_75t_L g3844 ( 
.A(n_3725),
.Y(n_3844)
);

OAI21x1_ASAP7_75t_L g3845 ( 
.A1(n_3735),
.A2(n_3537),
.B(n_3531),
.Y(n_3845)
);

INVx1_ASAP7_75t_L g3846 ( 
.A(n_3704),
.Y(n_3846)
);

OAI21x1_ASAP7_75t_L g3847 ( 
.A1(n_3689),
.A2(n_3558),
.B(n_3481),
.Y(n_3847)
);

INVx2_ASAP7_75t_L g3848 ( 
.A(n_3723),
.Y(n_3848)
);

INVx1_ASAP7_75t_L g3849 ( 
.A(n_3702),
.Y(n_3849)
);

INVx1_ASAP7_75t_L g3850 ( 
.A(n_3728),
.Y(n_3850)
);

INVxp33_ASAP7_75t_L g3851 ( 
.A(n_3650),
.Y(n_3851)
);

HB1xp67_ASAP7_75t_L g3852 ( 
.A(n_3694),
.Y(n_3852)
);

INVx1_ASAP7_75t_L g3853 ( 
.A(n_3728),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_3707),
.Y(n_3854)
);

NOR2xp33_ASAP7_75t_L g3855 ( 
.A(n_3731),
.B(n_3539),
.Y(n_3855)
);

INVx3_ASAP7_75t_L g3856 ( 
.A(n_3668),
.Y(n_3856)
);

INVx2_ASAP7_75t_L g3857 ( 
.A(n_3668),
.Y(n_3857)
);

INVx2_ASAP7_75t_L g3858 ( 
.A(n_3668),
.Y(n_3858)
);

BUFx6f_ASAP7_75t_L g3859 ( 
.A(n_3771),
.Y(n_3859)
);

INVx1_ASAP7_75t_L g3860 ( 
.A(n_3710),
.Y(n_3860)
);

AND2x2_ASAP7_75t_L g3861 ( 
.A(n_3679),
.B(n_3618),
.Y(n_3861)
);

INVx1_ASAP7_75t_L g3862 ( 
.A(n_3724),
.Y(n_3862)
);

AO21x2_ASAP7_75t_L g3863 ( 
.A1(n_3689),
.A2(n_3622),
.B(n_3620),
.Y(n_3863)
);

BUFx8_ASAP7_75t_L g3864 ( 
.A(n_3747),
.Y(n_3864)
);

INVx1_ASAP7_75t_L g3865 ( 
.A(n_3724),
.Y(n_3865)
);

NAND2xp5_ASAP7_75t_L g3866 ( 
.A(n_3681),
.B(n_3711),
.Y(n_3866)
);

HB1xp67_ASAP7_75t_L g3867 ( 
.A(n_3697),
.Y(n_3867)
);

INVx1_ASAP7_75t_L g3868 ( 
.A(n_3727),
.Y(n_3868)
);

INVx2_ASAP7_75t_L g3869 ( 
.A(n_3727),
.Y(n_3869)
);

INVx1_ASAP7_75t_L g3870 ( 
.A(n_3697),
.Y(n_3870)
);

CKINVDCx20_ASAP7_75t_R g3871 ( 
.A(n_3720),
.Y(n_3871)
);

OR2x2_ASAP7_75t_L g3872 ( 
.A(n_3673),
.B(n_3617),
.Y(n_3872)
);

INVx2_ASAP7_75t_L g3873 ( 
.A(n_3673),
.Y(n_3873)
);

INVx2_ASAP7_75t_L g3874 ( 
.A(n_3684),
.Y(n_3874)
);

HB1xp67_ASAP7_75t_L g3875 ( 
.A(n_3721),
.Y(n_3875)
);

INVx2_ASAP7_75t_SL g3876 ( 
.A(n_3757),
.Y(n_3876)
);

INVx2_ASAP7_75t_L g3877 ( 
.A(n_3684),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_3686),
.Y(n_3878)
);

INVx1_ASAP7_75t_L g3879 ( 
.A(n_3686),
.Y(n_3879)
);

INVx1_ASAP7_75t_L g3880 ( 
.A(n_3732),
.Y(n_3880)
);

INVx2_ASAP7_75t_L g3881 ( 
.A(n_3733),
.Y(n_3881)
);

INVx2_ASAP7_75t_L g3882 ( 
.A(n_3733),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_3738),
.Y(n_3883)
);

INVx2_ASAP7_75t_L g3884 ( 
.A(n_3737),
.Y(n_3884)
);

INVx2_ASAP7_75t_L g3885 ( 
.A(n_3691),
.Y(n_3885)
);

AND2x4_ASAP7_75t_SL g3886 ( 
.A(n_3746),
.B(n_3631),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_3752),
.Y(n_3887)
);

OA21x2_ASAP7_75t_L g3888 ( 
.A1(n_3766),
.A2(n_3568),
.B(n_3569),
.Y(n_3888)
);

OR2x2_ASAP7_75t_L g3889 ( 
.A(n_3669),
.B(n_3617),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3760),
.Y(n_3890)
);

AO21x2_ASAP7_75t_L g3891 ( 
.A1(n_3729),
.A2(n_3620),
.B(n_3454),
.Y(n_3891)
);

AND2x2_ASAP7_75t_L g3892 ( 
.A(n_3721),
.B(n_3571),
.Y(n_3892)
);

NAND2xp33_ASAP7_75t_R g3893 ( 
.A(n_3731),
.B(n_3543),
.Y(n_3893)
);

INVx2_ASAP7_75t_L g3894 ( 
.A(n_3691),
.Y(n_3894)
);

INVx2_ASAP7_75t_L g3895 ( 
.A(n_3691),
.Y(n_3895)
);

A2O1A1Ixp33_ASAP7_75t_L g3896 ( 
.A1(n_3784),
.A2(n_3695),
.B(n_3771),
.C(n_3745),
.Y(n_3896)
);

OAI22xp5_ASAP7_75t_L g3897 ( 
.A1(n_3777),
.A2(n_3696),
.B1(n_3683),
.B2(n_3768),
.Y(n_3897)
);

NAND2xp5_ASAP7_75t_L g3898 ( 
.A(n_3796),
.B(n_3743),
.Y(n_3898)
);

AOI22xp5_ASAP7_75t_L g3899 ( 
.A1(n_3796),
.A2(n_3764),
.B1(n_3729),
.B2(n_3718),
.Y(n_3899)
);

OAI21xp5_ASAP7_75t_L g3900 ( 
.A1(n_3791),
.A2(n_3756),
.B(n_3706),
.Y(n_3900)
);

INVx1_ASAP7_75t_L g3901 ( 
.A(n_3807),
.Y(n_3901)
);

OAI21xp5_ASAP7_75t_L g3902 ( 
.A1(n_3823),
.A2(n_3740),
.B(n_3677),
.Y(n_3902)
);

NAND2xp5_ASAP7_75t_L g3903 ( 
.A(n_3796),
.B(n_3709),
.Y(n_3903)
);

AND2x2_ASAP7_75t_L g3904 ( 
.A(n_3861),
.B(n_3716),
.Y(n_3904)
);

OAI21xp5_ASAP7_75t_L g3905 ( 
.A1(n_3823),
.A2(n_3740),
.B(n_3771),
.Y(n_3905)
);

OAI211xp5_ASAP7_75t_SL g3906 ( 
.A1(n_3801),
.A2(n_3866),
.B(n_3837),
.C(n_3802),
.Y(n_3906)
);

INVx3_ASAP7_75t_L g3907 ( 
.A(n_3785),
.Y(n_3907)
);

NAND2xp5_ASAP7_75t_L g3908 ( 
.A(n_3887),
.B(n_3755),
.Y(n_3908)
);

NAND3xp33_ASAP7_75t_L g3909 ( 
.A(n_3802),
.B(n_3726),
.C(n_3755),
.Y(n_3909)
);

NAND2xp5_ASAP7_75t_L g3910 ( 
.A(n_3887),
.B(n_3758),
.Y(n_3910)
);

INVx2_ASAP7_75t_L g3911 ( 
.A(n_3856),
.Y(n_3911)
);

AOI22xp33_ASAP7_75t_SL g3912 ( 
.A1(n_3839),
.A2(n_3754),
.B1(n_3745),
.B2(n_3742),
.Y(n_3912)
);

BUFx12f_ASAP7_75t_L g3913 ( 
.A(n_3864),
.Y(n_3913)
);

AOI22xp5_ASAP7_75t_L g3914 ( 
.A1(n_3863),
.A2(n_3716),
.B1(n_3676),
.B2(n_3748),
.Y(n_3914)
);

INVx1_ASAP7_75t_L g3915 ( 
.A(n_3789),
.Y(n_3915)
);

INVx4_ASAP7_75t_L g3916 ( 
.A(n_3859),
.Y(n_3916)
);

AND2x2_ASAP7_75t_L g3917 ( 
.A(n_3861),
.B(n_3749),
.Y(n_3917)
);

AO32x2_ASAP7_75t_L g3918 ( 
.A1(n_3827),
.A2(n_3736),
.A3(n_3665),
.B1(n_3750),
.B2(n_3758),
.Y(n_3918)
);

NOR2xp33_ASAP7_75t_L g3919 ( 
.A(n_3851),
.B(n_3747),
.Y(n_3919)
);

A2O1A1Ixp33_ASAP7_75t_L g3920 ( 
.A1(n_3845),
.A2(n_3754),
.B(n_3687),
.C(n_3685),
.Y(n_3920)
);

INVx3_ASAP7_75t_L g3921 ( 
.A(n_3785),
.Y(n_3921)
);

AND2x4_ASAP7_75t_L g3922 ( 
.A(n_3797),
.B(n_3736),
.Y(n_3922)
);

AND2x2_ASAP7_75t_L g3923 ( 
.A(n_3843),
.B(n_3714),
.Y(n_3923)
);

INVx1_ASAP7_75t_SL g3924 ( 
.A(n_3886),
.Y(n_3924)
);

AND2x2_ASAP7_75t_L g3925 ( 
.A(n_3843),
.B(n_3714),
.Y(n_3925)
);

OR2x2_ASAP7_75t_L g3926 ( 
.A(n_3803),
.B(n_3662),
.Y(n_3926)
);

AO21x2_ASAP7_75t_L g3927 ( 
.A1(n_3863),
.A2(n_3762),
.B(n_3760),
.Y(n_3927)
);

AND2x2_ASAP7_75t_L g3928 ( 
.A(n_3787),
.B(n_3700),
.Y(n_3928)
);

AOI22xp5_ASAP7_75t_L g3929 ( 
.A1(n_3863),
.A2(n_3891),
.B1(n_3782),
.B2(n_3798),
.Y(n_3929)
);

A2O1A1Ixp33_ASAP7_75t_L g3930 ( 
.A1(n_3845),
.A2(n_3687),
.B(n_3685),
.C(n_3535),
.Y(n_3930)
);

OR2x2_ASAP7_75t_L g3931 ( 
.A(n_3806),
.B(n_3713),
.Y(n_3931)
);

AND2x2_ASAP7_75t_L g3932 ( 
.A(n_3787),
.B(n_3700),
.Y(n_3932)
);

AND2x4_ASAP7_75t_L g3933 ( 
.A(n_3797),
.B(n_3744),
.Y(n_3933)
);

INVx2_ASAP7_75t_L g3934 ( 
.A(n_3856),
.Y(n_3934)
);

O2A1O1Ixp33_ASAP7_75t_L g3935 ( 
.A1(n_3891),
.A2(n_3751),
.B(n_3767),
.C(n_3769),
.Y(n_3935)
);

OR2x2_ASAP7_75t_L g3936 ( 
.A(n_3889),
.B(n_3734),
.Y(n_3936)
);

OA21x2_ASAP7_75t_L g3937 ( 
.A1(n_3792),
.A2(n_3772),
.B(n_3765),
.Y(n_3937)
);

OR2x6_ASAP7_75t_L g3938 ( 
.A(n_3859),
.B(n_3580),
.Y(n_3938)
);

INVx4_ASAP7_75t_L g3939 ( 
.A(n_3859),
.Y(n_3939)
);

AND2x2_ASAP7_75t_L g3940 ( 
.A(n_3892),
.B(n_3798),
.Y(n_3940)
);

AND2x2_ASAP7_75t_L g3941 ( 
.A(n_3892),
.B(n_3833),
.Y(n_3941)
);

A2O1A1Ixp33_ASAP7_75t_L g3942 ( 
.A1(n_3847),
.A2(n_3753),
.B(n_3766),
.C(n_3744),
.Y(n_3942)
);

O2A1O1Ixp33_ASAP7_75t_SL g3943 ( 
.A1(n_3889),
.A2(n_3753),
.B(n_3770),
.C(n_3765),
.Y(n_3943)
);

AND2x2_ASAP7_75t_L g3944 ( 
.A(n_3833),
.B(n_3831),
.Y(n_3944)
);

AND2x4_ASAP7_75t_L g3945 ( 
.A(n_3831),
.B(n_3827),
.Y(n_3945)
);

HB1xp67_ASAP7_75t_L g3946 ( 
.A(n_3817),
.Y(n_3946)
);

AND2x4_ASAP7_75t_SL g3947 ( 
.A(n_3859),
.B(n_3674),
.Y(n_3947)
);

INVx1_ASAP7_75t_L g3948 ( 
.A(n_3789),
.Y(n_3948)
);

OR2x2_ASAP7_75t_L g3949 ( 
.A(n_3872),
.B(n_3883),
.Y(n_3949)
);

A2O1A1Ixp33_ASAP7_75t_L g3950 ( 
.A1(n_3847),
.A2(n_3700),
.B(n_3761),
.C(n_3739),
.Y(n_3950)
);

AND2x2_ASAP7_75t_L g3951 ( 
.A(n_3818),
.B(n_3674),
.Y(n_3951)
);

NAND2xp5_ASAP7_75t_L g3952 ( 
.A(n_3876),
.B(n_3824),
.Y(n_3952)
);

NAND2xp5_ASAP7_75t_L g3953 ( 
.A(n_3876),
.B(n_3762),
.Y(n_3953)
);

INVx3_ASAP7_75t_L g3954 ( 
.A(n_3886),
.Y(n_3954)
);

AOI21xp5_ASAP7_75t_L g3955 ( 
.A1(n_3891),
.A2(n_3676),
.B(n_3538),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_L g3956 ( 
.A(n_3824),
.B(n_3770),
.Y(n_3956)
);

AND2x2_ASAP7_75t_L g3957 ( 
.A(n_3818),
.B(n_3739),
.Y(n_3957)
);

NAND2xp33_ASAP7_75t_L g3958 ( 
.A(n_3859),
.B(n_3533),
.Y(n_3958)
);

INVx1_ASAP7_75t_L g3959 ( 
.A(n_3799),
.Y(n_3959)
);

AND2x2_ASAP7_75t_L g3960 ( 
.A(n_3819),
.B(n_3739),
.Y(n_3960)
);

OAI22xp5_ASAP7_75t_L g3961 ( 
.A1(n_3888),
.A2(n_3676),
.B1(n_3772),
.B2(n_3624),
.Y(n_3961)
);

AO32x2_ASAP7_75t_L g3962 ( 
.A1(n_3875),
.A2(n_3761),
.A3(n_3644),
.B1(n_3527),
.B2(n_3712),
.Y(n_3962)
);

AO32x1_ASAP7_75t_L g3963 ( 
.A1(n_3819),
.A2(n_3712),
.A3(n_3678),
.B1(n_3676),
.B2(n_3527),
.Y(n_3963)
);

AOI22xp5_ASAP7_75t_L g3964 ( 
.A1(n_3782),
.A2(n_3678),
.B1(n_3391),
.B2(n_3452),
.Y(n_3964)
);

NAND2xp5_ASAP7_75t_L g3965 ( 
.A(n_3782),
.B(n_3172),
.Y(n_3965)
);

INVx1_ASAP7_75t_L g3966 ( 
.A(n_3799),
.Y(n_3966)
);

INVx2_ASAP7_75t_L g3967 ( 
.A(n_3856),
.Y(n_3967)
);

A2O1A1Ixp33_ASAP7_75t_L g3968 ( 
.A1(n_3822),
.A2(n_3169),
.B(n_3156),
.C(n_130),
.Y(n_3968)
);

OAI21xp5_ASAP7_75t_L g3969 ( 
.A1(n_3822),
.A2(n_128),
.B(n_129),
.Y(n_3969)
);

NOR2xp33_ASAP7_75t_L g3970 ( 
.A(n_3886),
.B(n_131),
.Y(n_3970)
);

AND2x2_ASAP7_75t_L g3971 ( 
.A(n_3782),
.B(n_3156),
.Y(n_3971)
);

INVx1_ASAP7_75t_L g3972 ( 
.A(n_3804),
.Y(n_3972)
);

HB1xp67_ASAP7_75t_L g3973 ( 
.A(n_3817),
.Y(n_3973)
);

AOI22xp33_ASAP7_75t_L g3974 ( 
.A1(n_3839),
.A2(n_3169),
.B1(n_3156),
.B2(n_135),
.Y(n_3974)
);

CKINVDCx20_ASAP7_75t_R g3975 ( 
.A(n_3779),
.Y(n_3975)
);

O2A1O1Ixp33_ASAP7_75t_SL g3976 ( 
.A1(n_3855),
.A2(n_132),
.B(n_134),
.C(n_136),
.Y(n_3976)
);

OA21x2_ASAP7_75t_L g3977 ( 
.A1(n_3792),
.A2(n_134),
.B(n_136),
.Y(n_3977)
);

AND2x2_ASAP7_75t_L g3978 ( 
.A(n_3857),
.B(n_137),
.Y(n_3978)
);

BUFx3_ASAP7_75t_L g3979 ( 
.A(n_3864),
.Y(n_3979)
);

AND2x2_ASAP7_75t_L g3980 ( 
.A(n_3857),
.B(n_138),
.Y(n_3980)
);

AND2x2_ASAP7_75t_L g3981 ( 
.A(n_3858),
.B(n_3885),
.Y(n_3981)
);

OAI21xp5_ASAP7_75t_L g3982 ( 
.A1(n_3795),
.A2(n_139),
.B(n_141),
.Y(n_3982)
);

NAND2x1p5_ASAP7_75t_L g3983 ( 
.A(n_3795),
.B(n_3820),
.Y(n_3983)
);

AND2x2_ASAP7_75t_L g3984 ( 
.A(n_3858),
.B(n_141),
.Y(n_3984)
);

OR2x2_ASAP7_75t_L g3985 ( 
.A(n_3872),
.B(n_143),
.Y(n_3985)
);

INVx2_ASAP7_75t_L g3986 ( 
.A(n_3856),
.Y(n_3986)
);

NAND2xp5_ASAP7_75t_L g3987 ( 
.A(n_3883),
.B(n_143),
.Y(n_3987)
);

AND2x2_ASAP7_75t_L g3988 ( 
.A(n_3885),
.B(n_144),
.Y(n_3988)
);

BUFx3_ASAP7_75t_L g3989 ( 
.A(n_3864),
.Y(n_3989)
);

AND2x2_ASAP7_75t_L g3990 ( 
.A(n_3894),
.B(n_145),
.Y(n_3990)
);

AOI221xp5_ASAP7_75t_L g3991 ( 
.A1(n_3811),
.A2(n_147),
.B1(n_150),
.B2(n_151),
.C(n_154),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_3804),
.Y(n_3992)
);

NOR2x1_ASAP7_75t_SL g3993 ( 
.A(n_3811),
.B(n_151),
.Y(n_3993)
);

AOI211xp5_ASAP7_75t_L g3994 ( 
.A1(n_3776),
.A2(n_155),
.B(n_156),
.C(n_157),
.Y(n_3994)
);

AND2x4_ASAP7_75t_L g3995 ( 
.A(n_3793),
.B(n_156),
.Y(n_3995)
);

BUFx2_ASAP7_75t_L g3996 ( 
.A(n_3790),
.Y(n_3996)
);

AOI22xp5_ASAP7_75t_L g3997 ( 
.A1(n_3888),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_3997)
);

BUFx6f_ASAP7_75t_L g3998 ( 
.A(n_3780),
.Y(n_3998)
);

AND2x2_ASAP7_75t_L g3999 ( 
.A(n_3894),
.B(n_3780),
.Y(n_3999)
);

AND2x2_ASAP7_75t_L g4000 ( 
.A(n_3895),
.B(n_160),
.Y(n_4000)
);

INVx2_ASAP7_75t_L g4001 ( 
.A(n_3820),
.Y(n_4001)
);

AOI221xp5_ASAP7_75t_L g4002 ( 
.A1(n_3811),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.C(n_165),
.Y(n_4002)
);

INVx1_ASAP7_75t_L g4003 ( 
.A(n_3805),
.Y(n_4003)
);

AND2x4_ASAP7_75t_SL g4004 ( 
.A(n_3871),
.B(n_162),
.Y(n_4004)
);

HB1xp67_ASAP7_75t_L g4005 ( 
.A(n_3852),
.Y(n_4005)
);

NAND2xp5_ASAP7_75t_L g4006 ( 
.A(n_3890),
.B(n_163),
.Y(n_4006)
);

OR2x6_ASAP7_75t_L g4007 ( 
.A(n_3793),
.B(n_165),
.Y(n_4007)
);

NOR2xp33_ASAP7_75t_L g4008 ( 
.A(n_3864),
.B(n_167),
.Y(n_4008)
);

AND2x2_ASAP7_75t_L g4009 ( 
.A(n_3895),
.B(n_168),
.Y(n_4009)
);

AND2x2_ASAP7_75t_L g4010 ( 
.A(n_3895),
.B(n_168),
.Y(n_4010)
);

AND2x4_ASAP7_75t_L g4011 ( 
.A(n_3793),
.B(n_170),
.Y(n_4011)
);

AO32x2_ASAP7_75t_L g4012 ( 
.A1(n_3790),
.A2(n_170),
.A3(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_4012)
);

AND2x4_ASAP7_75t_L g4013 ( 
.A(n_3793),
.B(n_171),
.Y(n_4013)
);

INVx3_ASAP7_75t_L g4014 ( 
.A(n_3820),
.Y(n_4014)
);

INVx1_ASAP7_75t_L g4015 ( 
.A(n_3946),
.Y(n_4015)
);

NAND2x1_ASAP7_75t_L g4016 ( 
.A(n_3954),
.B(n_3820),
.Y(n_4016)
);

BUFx3_ASAP7_75t_L g4017 ( 
.A(n_3913),
.Y(n_4017)
);

INVx2_ASAP7_75t_L g4018 ( 
.A(n_3998),
.Y(n_4018)
);

INVx2_ASAP7_75t_L g4019 ( 
.A(n_3998),
.Y(n_4019)
);

NAND2xp5_ASAP7_75t_L g4020 ( 
.A(n_3924),
.B(n_3890),
.Y(n_4020)
);

INVx2_ASAP7_75t_L g4021 ( 
.A(n_3998),
.Y(n_4021)
);

INVx1_ASAP7_75t_L g4022 ( 
.A(n_3973),
.Y(n_4022)
);

NAND2xp5_ASAP7_75t_SL g4023 ( 
.A(n_3954),
.B(n_3994),
.Y(n_4023)
);

AND2x2_ASAP7_75t_L g4024 ( 
.A(n_3941),
.B(n_3828),
.Y(n_4024)
);

NOR2xp33_ASAP7_75t_L g4025 ( 
.A(n_3907),
.B(n_3842),
.Y(n_4025)
);

AND2x2_ASAP7_75t_L g4026 ( 
.A(n_3940),
.B(n_3828),
.Y(n_4026)
);

INVx1_ASAP7_75t_L g4027 ( 
.A(n_3915),
.Y(n_4027)
);

INVx2_ASAP7_75t_L g4028 ( 
.A(n_4014),
.Y(n_4028)
);

INVx1_ASAP7_75t_L g4029 ( 
.A(n_3915),
.Y(n_4029)
);

INVx3_ASAP7_75t_L g4030 ( 
.A(n_3907),
.Y(n_4030)
);

INVx3_ASAP7_75t_L g4031 ( 
.A(n_3921),
.Y(n_4031)
);

AND2x2_ASAP7_75t_L g4032 ( 
.A(n_3904),
.B(n_3923),
.Y(n_4032)
);

INVx2_ASAP7_75t_L g4033 ( 
.A(n_4014),
.Y(n_4033)
);

NAND2xp5_ASAP7_75t_L g4034 ( 
.A(n_3997),
.B(n_4000),
.Y(n_4034)
);

AND2x2_ASAP7_75t_L g4035 ( 
.A(n_3925),
.B(n_3828),
.Y(n_4035)
);

AND2x2_ASAP7_75t_L g4036 ( 
.A(n_3944),
.B(n_3828),
.Y(n_4036)
);

INVx3_ASAP7_75t_L g4037 ( 
.A(n_3921),
.Y(n_4037)
);

OAI222xp33_ASAP7_75t_L g4038 ( 
.A1(n_3899),
.A2(n_3808),
.B1(n_3838),
.B2(n_3826),
.C1(n_3860),
.C2(n_3854),
.Y(n_4038)
);

INVx1_ASAP7_75t_L g4039 ( 
.A(n_3948),
.Y(n_4039)
);

HB1xp67_ASAP7_75t_L g4040 ( 
.A(n_4005),
.Y(n_4040)
);

INVx1_ASAP7_75t_L g4041 ( 
.A(n_3948),
.Y(n_4041)
);

INVx1_ASAP7_75t_L g4042 ( 
.A(n_3966),
.Y(n_4042)
);

NOR2xp33_ASAP7_75t_L g4043 ( 
.A(n_3979),
.B(n_3888),
.Y(n_4043)
);

BUFx3_ASAP7_75t_L g4044 ( 
.A(n_3989),
.Y(n_4044)
);

OR2x2_ASAP7_75t_L g4045 ( 
.A(n_3901),
.B(n_3808),
.Y(n_4045)
);

OR2x2_ASAP7_75t_L g4046 ( 
.A(n_3901),
.B(n_3838),
.Y(n_4046)
);

AND2x2_ASAP7_75t_L g4047 ( 
.A(n_3928),
.B(n_3776),
.Y(n_4047)
);

OAI21x1_ASAP7_75t_L g4048 ( 
.A1(n_3983),
.A2(n_3935),
.B(n_3955),
.Y(n_4048)
);

INVx2_ASAP7_75t_L g4049 ( 
.A(n_3918),
.Y(n_4049)
);

HB1xp67_ASAP7_75t_L g4050 ( 
.A(n_3952),
.Y(n_4050)
);

OR2x2_ASAP7_75t_L g4051 ( 
.A(n_3926),
.B(n_3854),
.Y(n_4051)
);

INVx2_ASAP7_75t_L g4052 ( 
.A(n_3918),
.Y(n_4052)
);

HB1xp67_ASAP7_75t_L g4053 ( 
.A(n_4007),
.Y(n_4053)
);

INVx1_ASAP7_75t_L g4054 ( 
.A(n_3966),
.Y(n_4054)
);

AND2x2_ASAP7_75t_L g4055 ( 
.A(n_3932),
.B(n_3933),
.Y(n_4055)
);

INVx1_ASAP7_75t_L g4056 ( 
.A(n_3992),
.Y(n_4056)
);

AND2x2_ASAP7_75t_L g4057 ( 
.A(n_3933),
.B(n_3800),
.Y(n_4057)
);

AND2x2_ASAP7_75t_L g4058 ( 
.A(n_3947),
.B(n_3800),
.Y(n_4058)
);

INVx2_ASAP7_75t_L g4059 ( 
.A(n_3918),
.Y(n_4059)
);

OR2x2_ASAP7_75t_L g4060 ( 
.A(n_3956),
.B(n_3860),
.Y(n_4060)
);

AND2x2_ASAP7_75t_L g4061 ( 
.A(n_3957),
.B(n_3800),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_3992),
.Y(n_4062)
);

INVx2_ASAP7_75t_L g4063 ( 
.A(n_3993),
.Y(n_4063)
);

AND2x2_ASAP7_75t_L g4064 ( 
.A(n_3960),
.B(n_3867),
.Y(n_4064)
);

AND2x4_ASAP7_75t_L g4065 ( 
.A(n_3993),
.B(n_3826),
.Y(n_4065)
);

AOI33xp33_ASAP7_75t_L g4066 ( 
.A1(n_3912),
.A2(n_3849),
.A3(n_3846),
.B1(n_3814),
.B2(n_3805),
.B3(n_3813),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_L g4067 ( 
.A(n_4009),
.B(n_3846),
.Y(n_4067)
);

INVx2_ASAP7_75t_L g4068 ( 
.A(n_3911),
.Y(n_4068)
);

AND2x2_ASAP7_75t_L g4069 ( 
.A(n_3962),
.B(n_3881),
.Y(n_4069)
);

AND2x2_ASAP7_75t_L g4070 ( 
.A(n_3962),
.B(n_3881),
.Y(n_4070)
);

AND2x4_ASAP7_75t_SL g4071 ( 
.A(n_3938),
.B(n_3849),
.Y(n_4071)
);

AND2x2_ASAP7_75t_L g4072 ( 
.A(n_3962),
.B(n_3882),
.Y(n_4072)
);

INVxp67_ASAP7_75t_L g4073 ( 
.A(n_3919),
.Y(n_4073)
);

INVx2_ASAP7_75t_L g4074 ( 
.A(n_3934),
.Y(n_4074)
);

OR2x2_ASAP7_75t_L g4075 ( 
.A(n_3931),
.B(n_3949),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_3959),
.Y(n_4076)
);

INVx1_ASAP7_75t_L g4077 ( 
.A(n_3972),
.Y(n_4077)
);

OAI22xp33_ASAP7_75t_L g4078 ( 
.A1(n_3929),
.A2(n_3888),
.B1(n_3816),
.B2(n_3880),
.Y(n_4078)
);

HB1xp67_ASAP7_75t_L g4079 ( 
.A(n_4007),
.Y(n_4079)
);

OR2x2_ASAP7_75t_L g4080 ( 
.A(n_3936),
.B(n_3870),
.Y(n_4080)
);

INVx3_ASAP7_75t_L g4081 ( 
.A(n_3977),
.Y(n_4081)
);

NAND2xp5_ASAP7_75t_L g4082 ( 
.A(n_4010),
.B(n_3813),
.Y(n_4082)
);

OR2x2_ASAP7_75t_L g4083 ( 
.A(n_3908),
.B(n_3870),
.Y(n_4083)
);

NOR2xp33_ASAP7_75t_L g4084 ( 
.A(n_3938),
.B(n_3816),
.Y(n_4084)
);

AND2x2_ASAP7_75t_L g4085 ( 
.A(n_3996),
.B(n_3882),
.Y(n_4085)
);

INVx2_ASAP7_75t_L g4086 ( 
.A(n_3967),
.Y(n_4086)
);

OAI21xp5_ASAP7_75t_L g4087 ( 
.A1(n_3896),
.A2(n_3816),
.B(n_3880),
.Y(n_4087)
);

INVx2_ASAP7_75t_L g4088 ( 
.A(n_3986),
.Y(n_4088)
);

INVx2_ASAP7_75t_L g4089 ( 
.A(n_3945),
.Y(n_4089)
);

INVx2_ASAP7_75t_L g4090 ( 
.A(n_3945),
.Y(n_4090)
);

AND2x2_ASAP7_75t_L g4091 ( 
.A(n_3951),
.B(n_3816),
.Y(n_4091)
);

AND2x2_ASAP7_75t_L g4092 ( 
.A(n_3922),
.B(n_3884),
.Y(n_4092)
);

INVxp67_ASAP7_75t_R g4093 ( 
.A(n_3978),
.Y(n_4093)
);

INVx1_ASAP7_75t_L g4094 ( 
.A(n_4003),
.Y(n_4094)
);

INVx2_ASAP7_75t_L g4095 ( 
.A(n_3927),
.Y(n_4095)
);

AOI22xp33_ASAP7_75t_L g4096 ( 
.A1(n_3906),
.A2(n_3884),
.B1(n_3850),
.B2(n_3853),
.Y(n_4096)
);

INVx1_ASAP7_75t_L g4097 ( 
.A(n_4012),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_L g4098 ( 
.A(n_3980),
.B(n_3814),
.Y(n_4098)
);

AND2x2_ASAP7_75t_L g4099 ( 
.A(n_3922),
.B(n_3794),
.Y(n_4099)
);

CKINVDCx20_ASAP7_75t_R g4100 ( 
.A(n_3975),
.Y(n_4100)
);

INVx3_ASAP7_75t_L g4101 ( 
.A(n_3977),
.Y(n_4101)
);

INVx1_ASAP7_75t_L g4102 ( 
.A(n_4012),
.Y(n_4102)
);

AO31x2_ASAP7_75t_L g4103 ( 
.A1(n_3898),
.A2(n_3786),
.A3(n_3775),
.B(n_3788),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_4012),
.Y(n_4104)
);

INVx2_ASAP7_75t_L g4105 ( 
.A(n_3917),
.Y(n_4105)
);

AND2x2_ASAP7_75t_L g4106 ( 
.A(n_3971),
.B(n_3794),
.Y(n_4106)
);

OR2x2_ASAP7_75t_L g4107 ( 
.A(n_3910),
.B(n_3953),
.Y(n_4107)
);

OAI211xp5_ASAP7_75t_L g4108 ( 
.A1(n_4087),
.A2(n_4002),
.B(n_3991),
.C(n_3903),
.Y(n_4108)
);

AND2x2_ASAP7_75t_L g4109 ( 
.A(n_4032),
.B(n_3916),
.Y(n_4109)
);

NAND2xp5_ASAP7_75t_L g4110 ( 
.A(n_4097),
.B(n_4102),
.Y(n_4110)
);

OAI221xp5_ASAP7_75t_SL g4111 ( 
.A1(n_4066),
.A2(n_4078),
.B1(n_3974),
.B2(n_4102),
.C(n_4097),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_L g4112 ( 
.A(n_4104),
.B(n_3995),
.Y(n_4112)
);

NAND3xp33_ASAP7_75t_L g4113 ( 
.A(n_4104),
.B(n_3969),
.C(n_4043),
.Y(n_4113)
);

NAND3xp33_ASAP7_75t_L g4114 ( 
.A(n_4081),
.B(n_3968),
.C(n_3982),
.Y(n_4114)
);

NAND3xp33_ASAP7_75t_L g4115 ( 
.A(n_4081),
.B(n_3909),
.C(n_3902),
.Y(n_4115)
);

AOI221xp5_ASAP7_75t_L g4116 ( 
.A1(n_4038),
.A2(n_3900),
.B1(n_3897),
.B2(n_3905),
.C(n_3943),
.Y(n_4116)
);

AOI22xp5_ASAP7_75t_L g4117 ( 
.A1(n_4023),
.A2(n_3914),
.B1(n_3961),
.B2(n_3958),
.Y(n_4117)
);

AOI221xp5_ASAP7_75t_L g4118 ( 
.A1(n_4040),
.A2(n_3976),
.B1(n_3942),
.B2(n_3920),
.C(n_3950),
.Y(n_4118)
);

NAND2xp5_ASAP7_75t_L g4119 ( 
.A(n_4053),
.B(n_3995),
.Y(n_4119)
);

OA211x2_ASAP7_75t_L g4120 ( 
.A1(n_4016),
.A2(n_4084),
.B(n_4025),
.C(n_4073),
.Y(n_4120)
);

AND2x2_ASAP7_75t_L g4121 ( 
.A(n_4032),
.B(n_3916),
.Y(n_4121)
);

NAND2xp5_ASAP7_75t_L g4122 ( 
.A(n_4079),
.B(n_4011),
.Y(n_4122)
);

NAND3xp33_ASAP7_75t_L g4123 ( 
.A(n_4081),
.B(n_4101),
.C(n_4063),
.Y(n_4123)
);

AOI22xp33_ASAP7_75t_L g4124 ( 
.A1(n_4034),
.A2(n_4008),
.B1(n_3970),
.B2(n_3939),
.Y(n_4124)
);

OAI22xp5_ASAP7_75t_L g4125 ( 
.A1(n_4081),
.A2(n_3930),
.B1(n_3964),
.B2(n_3965),
.Y(n_4125)
);

NAND2xp5_ASAP7_75t_L g4126 ( 
.A(n_4089),
.B(n_4013),
.Y(n_4126)
);

OAI221xp5_ASAP7_75t_SL g4127 ( 
.A1(n_4101),
.A2(n_3987),
.B1(n_3985),
.B2(n_4006),
.C(n_3999),
.Y(n_4127)
);

INVx2_ASAP7_75t_L g4128 ( 
.A(n_4065),
.Y(n_4128)
);

NAND4xp25_ASAP7_75t_L g4129 ( 
.A(n_4044),
.B(n_3939),
.C(n_3981),
.D(n_3893),
.Y(n_4129)
);

NAND2xp5_ASAP7_75t_L g4130 ( 
.A(n_4089),
.B(n_4011),
.Y(n_4130)
);

NAND2xp5_ASAP7_75t_L g4131 ( 
.A(n_4090),
.B(n_4013),
.Y(n_4131)
);

AOI221xp5_ASAP7_75t_L g4132 ( 
.A1(n_4101),
.A2(n_4001),
.B1(n_3984),
.B2(n_3990),
.C(n_3988),
.Y(n_4132)
);

OAI21xp5_ASAP7_75t_L g4133 ( 
.A1(n_4048),
.A2(n_4065),
.B(n_4101),
.Y(n_4133)
);

AND2x4_ASAP7_75t_SL g4134 ( 
.A(n_4030),
.B(n_3775),
.Y(n_4134)
);

AND2x2_ASAP7_75t_L g4135 ( 
.A(n_4093),
.B(n_4004),
.Y(n_4135)
);

AOI22xp33_ASAP7_75t_L g4136 ( 
.A1(n_4065),
.A2(n_3937),
.B1(n_3835),
.B2(n_3832),
.Y(n_4136)
);

AND2x2_ASAP7_75t_L g4137 ( 
.A(n_4093),
.B(n_3937),
.Y(n_4137)
);

AOI221xp5_ASAP7_75t_L g4138 ( 
.A1(n_4050),
.A2(n_4022),
.B1(n_4015),
.B2(n_4049),
.C(n_4059),
.Y(n_4138)
);

NAND3xp33_ASAP7_75t_L g4139 ( 
.A(n_4063),
.B(n_3853),
.C(n_3850),
.Y(n_4139)
);

OAI21xp5_ASAP7_75t_L g4140 ( 
.A1(n_4048),
.A2(n_3840),
.B(n_3834),
.Y(n_4140)
);

AND2x2_ASAP7_75t_L g4141 ( 
.A(n_4055),
.B(n_3809),
.Y(n_4141)
);

AND2x2_ASAP7_75t_L g4142 ( 
.A(n_4055),
.B(n_3809),
.Y(n_4142)
);

AND2x2_ASAP7_75t_L g4143 ( 
.A(n_4026),
.B(n_3810),
.Y(n_4143)
);

AND2x2_ASAP7_75t_L g4144 ( 
.A(n_4026),
.B(n_3810),
.Y(n_4144)
);

NAND3xp33_ASAP7_75t_L g4145 ( 
.A(n_4095),
.B(n_3840),
.C(n_3834),
.Y(n_4145)
);

AND2x2_ASAP7_75t_L g4146 ( 
.A(n_4044),
.B(n_3821),
.Y(n_4146)
);

NAND3xp33_ASAP7_75t_L g4147 ( 
.A(n_4095),
.B(n_3844),
.C(n_3825),
.Y(n_4147)
);

AND2x2_ASAP7_75t_L g4148 ( 
.A(n_4035),
.B(n_3812),
.Y(n_4148)
);

INVx1_ASAP7_75t_L g4149 ( 
.A(n_4015),
.Y(n_4149)
);

NAND2xp5_ASAP7_75t_SL g4150 ( 
.A(n_4065),
.B(n_3844),
.Y(n_4150)
);

AND2x2_ASAP7_75t_L g4151 ( 
.A(n_4035),
.B(n_3812),
.Y(n_4151)
);

NAND2xp5_ASAP7_75t_L g4152 ( 
.A(n_4090),
.B(n_3821),
.Y(n_4152)
);

AND2x2_ASAP7_75t_L g4153 ( 
.A(n_4044),
.B(n_3825),
.Y(n_4153)
);

NOR2xp67_ASAP7_75t_L g4154 ( 
.A(n_4030),
.B(n_3778),
.Y(n_4154)
);

OAI21xp5_ASAP7_75t_SL g4155 ( 
.A1(n_4071),
.A2(n_3963),
.B(n_3879),
.Y(n_4155)
);

NAND2xp5_ASAP7_75t_L g4156 ( 
.A(n_4105),
.B(n_3815),
.Y(n_4156)
);

NAND2xp5_ASAP7_75t_L g4157 ( 
.A(n_4105),
.B(n_3815),
.Y(n_4157)
);

AND2x2_ASAP7_75t_L g4158 ( 
.A(n_4024),
.B(n_3829),
.Y(n_4158)
);

AND2x2_ASAP7_75t_L g4159 ( 
.A(n_4024),
.B(n_3829),
.Y(n_4159)
);

INVxp67_ASAP7_75t_L g4160 ( 
.A(n_4030),
.Y(n_4160)
);

OAI221xp5_ASAP7_75t_L g4161 ( 
.A1(n_4017),
.A2(n_3963),
.B1(n_3879),
.B2(n_3878),
.C(n_3865),
.Y(n_4161)
);

OAI33xp33_ASAP7_75t_L g4162 ( 
.A1(n_4110),
.A2(n_4022),
.A3(n_4059),
.B1(n_4049),
.B2(n_4052),
.B3(n_4094),
.Y(n_4162)
);

AND2x2_ASAP7_75t_L g4163 ( 
.A(n_4135),
.B(n_4017),
.Y(n_4163)
);

INVx5_ASAP7_75t_L g4164 ( 
.A(n_4128),
.Y(n_4164)
);

OR2x2_ASAP7_75t_L g4165 ( 
.A(n_4112),
.B(n_4075),
.Y(n_4165)
);

INVx1_ASAP7_75t_L g4166 ( 
.A(n_4128),
.Y(n_4166)
);

NAND2xp5_ASAP7_75t_L g4167 ( 
.A(n_4124),
.B(n_4018),
.Y(n_4167)
);

AND2x2_ASAP7_75t_L g4168 ( 
.A(n_4109),
.B(n_4017),
.Y(n_4168)
);

INVx1_ASAP7_75t_L g4169 ( 
.A(n_4123),
.Y(n_4169)
);

NAND2xp5_ASAP7_75t_L g4170 ( 
.A(n_4124),
.B(n_4018),
.Y(n_4170)
);

AND2x2_ASAP7_75t_L g4171 ( 
.A(n_4109),
.B(n_4030),
.Y(n_4171)
);

INVx4_ASAP7_75t_L g4172 ( 
.A(n_4146),
.Y(n_4172)
);

OAI21xp5_ASAP7_75t_L g4173 ( 
.A1(n_4115),
.A2(n_4058),
.B(n_4052),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_4150),
.Y(n_4174)
);

BUFx3_ASAP7_75t_L g4175 ( 
.A(n_4121),
.Y(n_4175)
);

AND2x2_ASAP7_75t_L g4176 ( 
.A(n_4141),
.B(n_4031),
.Y(n_4176)
);

AND2x2_ASAP7_75t_L g4177 ( 
.A(n_4141),
.B(n_4031),
.Y(n_4177)
);

OR2x2_ASAP7_75t_L g4178 ( 
.A(n_4149),
.B(n_4075),
.Y(n_4178)
);

NOR2xp33_ASAP7_75t_L g4179 ( 
.A(n_4129),
.B(n_4100),
.Y(n_4179)
);

INVx2_ASAP7_75t_L g4180 ( 
.A(n_4134),
.Y(n_4180)
);

INVx2_ASAP7_75t_L g4181 ( 
.A(n_4134),
.Y(n_4181)
);

BUFx2_ASAP7_75t_L g4182 ( 
.A(n_4133),
.Y(n_4182)
);

INVx3_ASAP7_75t_L g4183 ( 
.A(n_4137),
.Y(n_4183)
);

AND2x2_ASAP7_75t_L g4184 ( 
.A(n_4142),
.B(n_4031),
.Y(n_4184)
);

OR2x2_ASAP7_75t_L g4185 ( 
.A(n_4150),
.B(n_4045),
.Y(n_4185)
);

AND2x2_ASAP7_75t_L g4186 ( 
.A(n_4142),
.B(n_4031),
.Y(n_4186)
);

O2A1O1Ixp5_ASAP7_75t_L g4187 ( 
.A1(n_4111),
.A2(n_4108),
.B(n_4140),
.C(n_4114),
.Y(n_4187)
);

AO31x2_ASAP7_75t_L g4188 ( 
.A1(n_4125),
.A2(n_4019),
.A3(n_4021),
.B(n_4027),
.Y(n_4188)
);

INVx1_ASAP7_75t_L g4189 ( 
.A(n_4119),
.Y(n_4189)
);

AND2x2_ASAP7_75t_L g4190 ( 
.A(n_4143),
.B(n_4037),
.Y(n_4190)
);

AND2x4_ASAP7_75t_SL g4191 ( 
.A(n_4153),
.B(n_4037),
.Y(n_4191)
);

BUFx2_ASAP7_75t_L g4192 ( 
.A(n_4160),
.Y(n_4192)
);

AO21x2_ASAP7_75t_L g4193 ( 
.A1(n_4145),
.A2(n_4147),
.B(n_4113),
.Y(n_4193)
);

NAND5xp2_ASAP7_75t_L g4194 ( 
.A(n_4116),
.B(n_4047),
.C(n_4069),
.D(n_4070),
.E(n_4072),
.Y(n_4194)
);

INVx1_ASAP7_75t_L g4195 ( 
.A(n_4122),
.Y(n_4195)
);

INVx1_ASAP7_75t_L g4196 ( 
.A(n_4152),
.Y(n_4196)
);

AOI22xp5_ASAP7_75t_L g4197 ( 
.A1(n_4118),
.A2(n_4064),
.B1(n_4036),
.B2(n_4047),
.Y(n_4197)
);

AND2x2_ASAP7_75t_L g4198 ( 
.A(n_4143),
.B(n_4037),
.Y(n_4198)
);

AOI21xp5_ASAP7_75t_L g4199 ( 
.A1(n_4138),
.A2(n_3963),
.B(n_4071),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_4156),
.Y(n_4200)
);

NOR2xp33_ASAP7_75t_R g4201 ( 
.A(n_4126),
.B(n_4037),
.Y(n_4201)
);

OAI33xp33_ASAP7_75t_L g4202 ( 
.A1(n_4130),
.A2(n_4077),
.A3(n_4076),
.B1(n_4094),
.B2(n_4021),
.B3(n_4019),
.Y(n_4202)
);

AOI221xp5_ASAP7_75t_L g4203 ( 
.A1(n_4127),
.A2(n_4072),
.B1(n_4070),
.B2(n_4069),
.C(n_4058),
.Y(n_4203)
);

INVx2_ASAP7_75t_L g4204 ( 
.A(n_4144),
.Y(n_4204)
);

AND2x2_ASAP7_75t_SL g4205 ( 
.A(n_4117),
.B(n_4071),
.Y(n_4205)
);

AOI21xp5_ASAP7_75t_L g4206 ( 
.A1(n_4155),
.A2(n_4016),
.B(n_4067),
.Y(n_4206)
);

BUFx2_ASAP7_75t_L g4207 ( 
.A(n_4131),
.Y(n_4207)
);

AND2x2_ASAP7_75t_L g4208 ( 
.A(n_4144),
.B(n_4036),
.Y(n_4208)
);

AND2x2_ASAP7_75t_L g4209 ( 
.A(n_4158),
.B(n_4064),
.Y(n_4209)
);

AND2x2_ASAP7_75t_L g4210 ( 
.A(n_4158),
.B(n_4085),
.Y(n_4210)
);

INVx2_ASAP7_75t_L g4211 ( 
.A(n_4148),
.Y(n_4211)
);

NAND2xp5_ASAP7_75t_L g4212 ( 
.A(n_4132),
.B(n_4085),
.Y(n_4212)
);

OAI21xp33_ASAP7_75t_L g4213 ( 
.A1(n_4157),
.A2(n_4020),
.B(n_4107),
.Y(n_4213)
);

AND2x2_ASAP7_75t_L g4214 ( 
.A(n_4168),
.B(n_4092),
.Y(n_4214)
);

NOR2xp33_ASAP7_75t_L g4215 ( 
.A(n_4168),
.B(n_4082),
.Y(n_4215)
);

AND2x2_ASAP7_75t_L g4216 ( 
.A(n_4163),
.B(n_4092),
.Y(n_4216)
);

AND2x2_ASAP7_75t_L g4217 ( 
.A(n_4163),
.B(n_4099),
.Y(n_4217)
);

INVxp67_ASAP7_75t_SL g4218 ( 
.A(n_4185),
.Y(n_4218)
);

INVx1_ASAP7_75t_L g4219 ( 
.A(n_4185),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_4178),
.Y(n_4220)
);

AND2x2_ASAP7_75t_L g4221 ( 
.A(n_4209),
.B(n_4099),
.Y(n_4221)
);

AND2x2_ASAP7_75t_L g4222 ( 
.A(n_4209),
.B(n_4106),
.Y(n_4222)
);

INVx2_ASAP7_75t_L g4223 ( 
.A(n_4164),
.Y(n_4223)
);

INVx1_ASAP7_75t_L g4224 ( 
.A(n_4178),
.Y(n_4224)
);

AND2x2_ASAP7_75t_L g4225 ( 
.A(n_4171),
.B(n_4106),
.Y(n_4225)
);

INVx1_ASAP7_75t_L g4226 ( 
.A(n_4204),
.Y(n_4226)
);

OR2x2_ASAP7_75t_L g4227 ( 
.A(n_4193),
.B(n_4045),
.Y(n_4227)
);

INVx1_ASAP7_75t_L g4228 ( 
.A(n_4204),
.Y(n_4228)
);

NAND2xp5_ASAP7_75t_L g4229 ( 
.A(n_4171),
.B(n_4098),
.Y(n_4229)
);

NAND2xp5_ASAP7_75t_L g4230 ( 
.A(n_4210),
.B(n_4148),
.Y(n_4230)
);

HB1xp67_ASAP7_75t_L g4231 ( 
.A(n_4164),
.Y(n_4231)
);

AND2x2_ASAP7_75t_L g4232 ( 
.A(n_4210),
.B(n_4151),
.Y(n_4232)
);

INVx3_ASAP7_75t_L g4233 ( 
.A(n_4188),
.Y(n_4233)
);

INVx1_ASAP7_75t_L g4234 ( 
.A(n_4211),
.Y(n_4234)
);

INVx1_ASAP7_75t_L g4235 ( 
.A(n_4211),
.Y(n_4235)
);

AND2x4_ASAP7_75t_L g4236 ( 
.A(n_4164),
.B(n_4154),
.Y(n_4236)
);

OR2x2_ASAP7_75t_L g4237 ( 
.A(n_4193),
.B(n_4046),
.Y(n_4237)
);

AOI22xp33_ASAP7_75t_L g4238 ( 
.A1(n_4194),
.A2(n_4120),
.B1(n_4061),
.B2(n_4091),
.Y(n_4238)
);

AND2x2_ASAP7_75t_L g4239 ( 
.A(n_4208),
.B(n_4151),
.Y(n_4239)
);

AND2x2_ASAP7_75t_L g4240 ( 
.A(n_4208),
.B(n_4159),
.Y(n_4240)
);

INVx2_ASAP7_75t_L g4241 ( 
.A(n_4164),
.Y(n_4241)
);

INVx1_ASAP7_75t_L g4242 ( 
.A(n_4193),
.Y(n_4242)
);

OR2x2_ASAP7_75t_L g4243 ( 
.A(n_4165),
.B(n_4046),
.Y(n_4243)
);

INVx1_ASAP7_75t_L g4244 ( 
.A(n_4166),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_4164),
.Y(n_4245)
);

INVx2_ASAP7_75t_L g4246 ( 
.A(n_4191),
.Y(n_4246)
);

INVx1_ASAP7_75t_L g4247 ( 
.A(n_4190),
.Y(n_4247)
);

INVx2_ASAP7_75t_L g4248 ( 
.A(n_4191),
.Y(n_4248)
);

INVx1_ASAP7_75t_L g4249 ( 
.A(n_4190),
.Y(n_4249)
);

NAND2xp5_ASAP7_75t_L g4250 ( 
.A(n_4176),
.B(n_4107),
.Y(n_4250)
);

OR2x2_ASAP7_75t_L g4251 ( 
.A(n_4165),
.B(n_4169),
.Y(n_4251)
);

INVx2_ASAP7_75t_L g4252 ( 
.A(n_4198),
.Y(n_4252)
);

HB1xp67_ASAP7_75t_L g4253 ( 
.A(n_4231),
.Y(n_4253)
);

INVx2_ASAP7_75t_L g4254 ( 
.A(n_4233),
.Y(n_4254)
);

AND2x2_ASAP7_75t_L g4255 ( 
.A(n_4217),
.B(n_4176),
.Y(n_4255)
);

OR2x2_ASAP7_75t_L g4256 ( 
.A(n_4227),
.B(n_4173),
.Y(n_4256)
);

INVx1_ASAP7_75t_L g4257 ( 
.A(n_4233),
.Y(n_4257)
);

AND2x4_ASAP7_75t_SL g4258 ( 
.A(n_4217),
.B(n_4172),
.Y(n_4258)
);

AND2x2_ASAP7_75t_L g4259 ( 
.A(n_4216),
.B(n_4214),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_4220),
.Y(n_4260)
);

INVx1_ASAP7_75t_L g4261 ( 
.A(n_4233),
.Y(n_4261)
);

HB1xp67_ASAP7_75t_L g4262 ( 
.A(n_4236),
.Y(n_4262)
);

INVx1_ASAP7_75t_L g4263 ( 
.A(n_4233),
.Y(n_4263)
);

INVx2_ASAP7_75t_L g4264 ( 
.A(n_4236),
.Y(n_4264)
);

NAND2xp5_ASAP7_75t_L g4265 ( 
.A(n_4216),
.B(n_4192),
.Y(n_4265)
);

INVx2_ASAP7_75t_L g4266 ( 
.A(n_4236),
.Y(n_4266)
);

OR2x2_ASAP7_75t_L g4267 ( 
.A(n_4227),
.B(n_4237),
.Y(n_4267)
);

HB1xp67_ASAP7_75t_L g4268 ( 
.A(n_4236),
.Y(n_4268)
);

OR2x2_ASAP7_75t_L g4269 ( 
.A(n_4237),
.B(n_4183),
.Y(n_4269)
);

OR2x2_ASAP7_75t_L g4270 ( 
.A(n_4243),
.B(n_4183),
.Y(n_4270)
);

INVx1_ASAP7_75t_L g4271 ( 
.A(n_4220),
.Y(n_4271)
);

AND2x2_ASAP7_75t_L g4272 ( 
.A(n_4214),
.B(n_4177),
.Y(n_4272)
);

AND2x2_ASAP7_75t_L g4273 ( 
.A(n_4221),
.B(n_4177),
.Y(n_4273)
);

INVx1_ASAP7_75t_L g4274 ( 
.A(n_4224),
.Y(n_4274)
);

INVx3_ASAP7_75t_L g4275 ( 
.A(n_4223),
.Y(n_4275)
);

INVx2_ASAP7_75t_L g4276 ( 
.A(n_4223),
.Y(n_4276)
);

AND2x2_ASAP7_75t_L g4277 ( 
.A(n_4221),
.B(n_4184),
.Y(n_4277)
);

INVx1_ASAP7_75t_L g4278 ( 
.A(n_4224),
.Y(n_4278)
);

AOI22xp5_ASAP7_75t_L g4279 ( 
.A1(n_4256),
.A2(n_4182),
.B1(n_4238),
.B2(n_4218),
.Y(n_4279)
);

INVx2_ASAP7_75t_SL g4280 ( 
.A(n_4258),
.Y(n_4280)
);

INVx2_ASAP7_75t_L g4281 ( 
.A(n_4270),
.Y(n_4281)
);

AOI32xp33_ASAP7_75t_L g4282 ( 
.A1(n_4256),
.A2(n_4242),
.A3(n_4219),
.B1(n_4174),
.B2(n_4170),
.Y(n_4282)
);

XNOR2x2_ASAP7_75t_L g4283 ( 
.A(n_4267),
.B(n_4242),
.Y(n_4283)
);

O2A1O1Ixp33_ASAP7_75t_L g4284 ( 
.A1(n_4267),
.A2(n_4187),
.B(n_4219),
.C(n_4199),
.Y(n_4284)
);

INVx2_ASAP7_75t_L g4285 ( 
.A(n_4270),
.Y(n_4285)
);

INVx1_ASAP7_75t_L g4286 ( 
.A(n_4269),
.Y(n_4286)
);

O2A1O1Ixp5_ASAP7_75t_L g4287 ( 
.A1(n_4269),
.A2(n_4162),
.B(n_4172),
.C(n_4212),
.Y(n_4287)
);

NOR2xp33_ASAP7_75t_L g4288 ( 
.A(n_4265),
.B(n_4175),
.Y(n_4288)
);

OR2x2_ASAP7_75t_L g4289 ( 
.A(n_4259),
.B(n_4243),
.Y(n_4289)
);

NAND2xp5_ASAP7_75t_L g4290 ( 
.A(n_4259),
.B(n_4232),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_4262),
.Y(n_4291)
);

INVx1_ASAP7_75t_L g4292 ( 
.A(n_4268),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_4273),
.Y(n_4293)
);

INVx1_ASAP7_75t_L g4294 ( 
.A(n_4273),
.Y(n_4294)
);

INVx1_ASAP7_75t_L g4295 ( 
.A(n_4277),
.Y(n_4295)
);

INVx1_ASAP7_75t_L g4296 ( 
.A(n_4277),
.Y(n_4296)
);

NAND2x1p5_ASAP7_75t_L g4297 ( 
.A(n_4255),
.B(n_4175),
.Y(n_4297)
);

OAI32xp33_ASAP7_75t_L g4298 ( 
.A1(n_4278),
.A2(n_4251),
.A3(n_4167),
.B1(n_4246),
.B2(n_4248),
.Y(n_4298)
);

OR2x2_ASAP7_75t_L g4299 ( 
.A(n_4289),
.B(n_4230),
.Y(n_4299)
);

OAI22xp5_ASAP7_75t_L g4300 ( 
.A1(n_4279),
.A2(n_4197),
.B1(n_4203),
.B2(n_4205),
.Y(n_4300)
);

XNOR2xp5_ASAP7_75t_L g4301 ( 
.A(n_4279),
.B(n_4205),
.Y(n_4301)
);

XOR2x2_ASAP7_75t_L g4302 ( 
.A(n_4297),
.B(n_4179),
.Y(n_4302)
);

INVx1_ASAP7_75t_SL g4303 ( 
.A(n_4290),
.Y(n_4303)
);

INVxp67_ASAP7_75t_SL g4304 ( 
.A(n_4283),
.Y(n_4304)
);

INVx1_ASAP7_75t_L g4305 ( 
.A(n_4291),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_4292),
.Y(n_4306)
);

AND2x4_ASAP7_75t_L g4307 ( 
.A(n_4281),
.B(n_4258),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_4286),
.Y(n_4308)
);

NOR2xp33_ASAP7_75t_L g4309 ( 
.A(n_4280),
.B(n_4172),
.Y(n_4309)
);

NOR2xp33_ASAP7_75t_L g4310 ( 
.A(n_4298),
.B(n_4207),
.Y(n_4310)
);

INVx2_ASAP7_75t_L g4311 ( 
.A(n_4285),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_4293),
.Y(n_4312)
);

XOR2x2_ASAP7_75t_L g4313 ( 
.A(n_4288),
.B(n_4255),
.Y(n_4313)
);

OR2x2_ASAP7_75t_L g4314 ( 
.A(n_4294),
.B(n_4252),
.Y(n_4314)
);

NAND2xp5_ASAP7_75t_L g4315 ( 
.A(n_4295),
.B(n_4272),
.Y(n_4315)
);

INVxp67_ASAP7_75t_L g4316 ( 
.A(n_4309),
.Y(n_4316)
);

CKINVDCx16_ASAP7_75t_R g4317 ( 
.A(n_4301),
.Y(n_4317)
);

INVx4_ASAP7_75t_L g4318 ( 
.A(n_4307),
.Y(n_4318)
);

INVx1_ASAP7_75t_L g4319 ( 
.A(n_4307),
.Y(n_4319)
);

INVx1_ASAP7_75t_SL g4320 ( 
.A(n_4314),
.Y(n_4320)
);

NAND2xp5_ASAP7_75t_L g4321 ( 
.A(n_4304),
.B(n_4272),
.Y(n_4321)
);

NAND2xp5_ASAP7_75t_L g4322 ( 
.A(n_4310),
.B(n_4247),
.Y(n_4322)
);

NAND2xp5_ASAP7_75t_L g4323 ( 
.A(n_4311),
.B(n_4247),
.Y(n_4323)
);

HB1xp67_ASAP7_75t_L g4324 ( 
.A(n_4313),
.Y(n_4324)
);

NOR2x1_ASAP7_75t_L g4325 ( 
.A(n_4299),
.B(n_4275),
.Y(n_4325)
);

AND2x2_ASAP7_75t_L g4326 ( 
.A(n_4303),
.B(n_4296),
.Y(n_4326)
);

INVx1_ASAP7_75t_SL g4327 ( 
.A(n_4315),
.Y(n_4327)
);

INVx1_ASAP7_75t_L g4328 ( 
.A(n_4325),
.Y(n_4328)
);

AND2x2_ASAP7_75t_SL g4329 ( 
.A(n_4318),
.B(n_4251),
.Y(n_4329)
);

OAI221xp5_ASAP7_75t_L g4330 ( 
.A1(n_4321),
.A2(n_4282),
.B1(n_4284),
.B2(n_4300),
.C(n_4287),
.Y(n_4330)
);

OAI21xp5_ASAP7_75t_L g4331 ( 
.A1(n_4316),
.A2(n_4248),
.B(n_4246),
.Y(n_4331)
);

INVx2_ASAP7_75t_L g4332 ( 
.A(n_4318),
.Y(n_4332)
);

NAND2xp5_ASAP7_75t_L g4333 ( 
.A(n_4319),
.B(n_4249),
.Y(n_4333)
);

AND2x2_ASAP7_75t_SL g4334 ( 
.A(n_4317),
.B(n_4278),
.Y(n_4334)
);

INVx1_ASAP7_75t_L g4335 ( 
.A(n_4326),
.Y(n_4335)
);

NAND3xp33_ASAP7_75t_SL g4336 ( 
.A(n_4330),
.B(n_4282),
.C(n_4320),
.Y(n_4336)
);

AND2x2_ASAP7_75t_L g4337 ( 
.A(n_4329),
.B(n_4215),
.Y(n_4337)
);

OR2x2_ASAP7_75t_L g4338 ( 
.A(n_4332),
.B(n_4252),
.Y(n_4338)
);

NAND3xp33_ASAP7_75t_SL g4339 ( 
.A(n_4328),
.B(n_4327),
.C(n_4308),
.Y(n_4339)
);

INVx1_ASAP7_75t_L g4340 ( 
.A(n_4334),
.Y(n_4340)
);

OAI32xp33_ASAP7_75t_L g4341 ( 
.A1(n_4333),
.A2(n_4249),
.A3(n_4322),
.B1(n_4306),
.B2(n_4305),
.Y(n_4341)
);

AOI21xp33_ASAP7_75t_SL g4342 ( 
.A1(n_4328),
.A2(n_4253),
.B(n_4260),
.Y(n_4342)
);

INVx1_ASAP7_75t_L g4343 ( 
.A(n_4331),
.Y(n_4343)
);

INVx1_ASAP7_75t_L g4344 ( 
.A(n_4335),
.Y(n_4344)
);

INVx2_ASAP7_75t_L g4345 ( 
.A(n_4329),
.Y(n_4345)
);

INVx1_ASAP7_75t_L g4346 ( 
.A(n_4329),
.Y(n_4346)
);

INVx1_ASAP7_75t_L g4347 ( 
.A(n_4329),
.Y(n_4347)
);

NAND2xp5_ASAP7_75t_L g4348 ( 
.A(n_4329),
.B(n_4271),
.Y(n_4348)
);

AOI21xp5_ASAP7_75t_L g4349 ( 
.A1(n_4348),
.A2(n_4302),
.B(n_4324),
.Y(n_4349)
);

AOI22xp33_ASAP7_75t_L g4350 ( 
.A1(n_4336),
.A2(n_4180),
.B1(n_4181),
.B2(n_4183),
.Y(n_4350)
);

NAND2xp5_ASAP7_75t_L g4351 ( 
.A(n_4337),
.B(n_4274),
.Y(n_4351)
);

NAND2xp5_ASAP7_75t_L g4352 ( 
.A(n_4346),
.B(n_4226),
.Y(n_4352)
);

INVx1_ASAP7_75t_L g4353 ( 
.A(n_4338),
.Y(n_4353)
);

NAND2xp5_ASAP7_75t_L g4354 ( 
.A(n_4347),
.B(n_4226),
.Y(n_4354)
);

OR2x2_ASAP7_75t_L g4355 ( 
.A(n_4345),
.B(n_4250),
.Y(n_4355)
);

NAND2xp5_ASAP7_75t_L g4356 ( 
.A(n_4342),
.B(n_4228),
.Y(n_4356)
);

OR2x2_ASAP7_75t_L g4357 ( 
.A(n_4340),
.B(n_4229),
.Y(n_4357)
);

NAND2xp5_ASAP7_75t_L g4358 ( 
.A(n_4342),
.B(n_4228),
.Y(n_4358)
);

INVx1_ASAP7_75t_L g4359 ( 
.A(n_4343),
.Y(n_4359)
);

AND2x2_ASAP7_75t_L g4360 ( 
.A(n_4344),
.B(n_4189),
.Y(n_4360)
);

NAND2xp5_ASAP7_75t_L g4361 ( 
.A(n_4341),
.B(n_4234),
.Y(n_4361)
);

INVx1_ASAP7_75t_L g4362 ( 
.A(n_4339),
.Y(n_4362)
);

NAND2xp5_ASAP7_75t_L g4363 ( 
.A(n_4337),
.B(n_4234),
.Y(n_4363)
);

INVx1_ASAP7_75t_L g4364 ( 
.A(n_4337),
.Y(n_4364)
);

INVx1_ASAP7_75t_L g4365 ( 
.A(n_4337),
.Y(n_4365)
);

AND2x4_ASAP7_75t_L g4366 ( 
.A(n_4345),
.B(n_4264),
.Y(n_4366)
);

INVx1_ASAP7_75t_L g4367 ( 
.A(n_4337),
.Y(n_4367)
);

INVx1_ASAP7_75t_L g4368 ( 
.A(n_4337),
.Y(n_4368)
);

AND2x2_ASAP7_75t_L g4369 ( 
.A(n_4337),
.B(n_4195),
.Y(n_4369)
);

AND2x2_ASAP7_75t_L g4370 ( 
.A(n_4337),
.B(n_4232),
.Y(n_4370)
);

OAI322xp33_ASAP7_75t_L g4371 ( 
.A1(n_4361),
.A2(n_4312),
.A3(n_4323),
.B1(n_4245),
.B2(n_4266),
.C1(n_4264),
.C2(n_4276),
.Y(n_4371)
);

HB1xp67_ASAP7_75t_L g4372 ( 
.A(n_4370),
.Y(n_4372)
);

AOI221xp5_ASAP7_75t_L g4373 ( 
.A1(n_4350),
.A2(n_4235),
.B1(n_4244),
.B2(n_4245),
.C(n_4266),
.Y(n_4373)
);

OAI22xp5_ASAP7_75t_SL g4374 ( 
.A1(n_4362),
.A2(n_4276),
.B1(n_4275),
.B2(n_4257),
.Y(n_4374)
);

INVx1_ASAP7_75t_L g4375 ( 
.A(n_4356),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_4358),
.Y(n_4376)
);

OAI22xp33_ASAP7_75t_L g4377 ( 
.A1(n_4355),
.A2(n_4180),
.B1(n_4181),
.B2(n_4235),
.Y(n_4377)
);

AND4x1_ASAP7_75t_L g4378 ( 
.A(n_4349),
.B(n_4257),
.C(n_4263),
.D(n_4261),
.Y(n_4378)
);

INVx1_ASAP7_75t_SL g4379 ( 
.A(n_4366),
.Y(n_4379)
);

OAI22xp5_ASAP7_75t_L g4380 ( 
.A1(n_4357),
.A2(n_4200),
.B1(n_4196),
.B2(n_4244),
.Y(n_4380)
);

AOI22xp5_ASAP7_75t_SL g4381 ( 
.A1(n_4366),
.A2(n_4275),
.B1(n_4263),
.B2(n_4261),
.Y(n_4381)
);

HB1xp67_ASAP7_75t_L g4382 ( 
.A(n_4363),
.Y(n_4382)
);

AOI221xp5_ASAP7_75t_L g4383 ( 
.A1(n_4359),
.A2(n_4353),
.B1(n_4352),
.B2(n_4354),
.C(n_4365),
.Y(n_4383)
);

OAI322xp33_ASAP7_75t_L g4384 ( 
.A1(n_4351),
.A2(n_4241),
.A3(n_4254),
.B1(n_4206),
.B2(n_4225),
.C1(n_4239),
.C2(n_4240),
.Y(n_4384)
);

OAI22xp5_ASAP7_75t_L g4385 ( 
.A1(n_4364),
.A2(n_4241),
.B1(n_4225),
.B2(n_4239),
.Y(n_4385)
);

AOI22xp5_ASAP7_75t_L g4386 ( 
.A1(n_4367),
.A2(n_4240),
.B1(n_4202),
.B2(n_4222),
.Y(n_4386)
);

OAI322xp33_ASAP7_75t_L g4387 ( 
.A1(n_4368),
.A2(n_4254),
.A3(n_4198),
.B1(n_4186),
.B2(n_4184),
.C1(n_4222),
.C2(n_4188),
.Y(n_4387)
);

OAI322xp33_ASAP7_75t_L g4388 ( 
.A1(n_4360),
.A2(n_4186),
.A3(n_4188),
.B1(n_4201),
.B2(n_4139),
.C1(n_4039),
.C2(n_4041),
.Y(n_4388)
);

OAI22xp5_ASAP7_75t_L g4389 ( 
.A1(n_4369),
.A2(n_4161),
.B1(n_4136),
.B2(n_4213),
.Y(n_4389)
);

INVx1_ASAP7_75t_L g4390 ( 
.A(n_4370),
.Y(n_4390)
);

INVx1_ASAP7_75t_L g4391 ( 
.A(n_4370),
.Y(n_4391)
);

INVx1_ASAP7_75t_L g4392 ( 
.A(n_4370),
.Y(n_4392)
);

INVx1_ASAP7_75t_L g4393 ( 
.A(n_4370),
.Y(n_4393)
);

NAND4xp25_ASAP7_75t_SL g4394 ( 
.A(n_4350),
.B(n_4136),
.C(n_4201),
.D(n_4057),
.Y(n_4394)
);

AOI22xp5_ASAP7_75t_L g4395 ( 
.A1(n_4370),
.A2(n_4077),
.B1(n_4076),
.B2(n_4074),
.Y(n_4395)
);

OAI22xp5_ASAP7_75t_L g4396 ( 
.A1(n_4350),
.A2(n_4068),
.B1(n_4074),
.B2(n_4088),
.Y(n_4396)
);

AOI22xp5_ASAP7_75t_L g4397 ( 
.A1(n_4389),
.A2(n_4068),
.B1(n_4086),
.B2(n_4088),
.Y(n_4397)
);

OAI21xp33_ASAP7_75t_L g4398 ( 
.A1(n_4386),
.A2(n_4086),
.B(n_4033),
.Y(n_4398)
);

NAND3xp33_ASAP7_75t_SL g4399 ( 
.A(n_4379),
.B(n_4057),
.C(n_4061),
.Y(n_4399)
);

NAND4xp25_ASAP7_75t_SL g4400 ( 
.A(n_4383),
.B(n_4188),
.C(n_4054),
.D(n_4056),
.Y(n_4400)
);

INVx1_ASAP7_75t_L g4401 ( 
.A(n_4381),
.Y(n_4401)
);

INVx1_ASAP7_75t_L g4402 ( 
.A(n_4374),
.Y(n_4402)
);

NOR2x1_ASAP7_75t_L g4403 ( 
.A(n_4371),
.B(n_4390),
.Y(n_4403)
);

INVx1_ASAP7_75t_L g4404 ( 
.A(n_4384),
.Y(n_4404)
);

INVx1_ASAP7_75t_L g4405 ( 
.A(n_4387),
.Y(n_4405)
);

OAI21xp33_ASAP7_75t_L g4406 ( 
.A1(n_4391),
.A2(n_4033),
.B(n_4028),
.Y(n_4406)
);

NOR3xp33_ASAP7_75t_L g4407 ( 
.A(n_4392),
.B(n_4029),
.C(n_4027),
.Y(n_4407)
);

INVx1_ASAP7_75t_L g4408 ( 
.A(n_4372),
.Y(n_4408)
);

NOR3x1_ASAP7_75t_L g4409 ( 
.A(n_4385),
.B(n_4039),
.C(n_4029),
.Y(n_4409)
);

INVx1_ASAP7_75t_L g4410 ( 
.A(n_4393),
.Y(n_4410)
);

NAND2xp5_ASAP7_75t_SL g4411 ( 
.A(n_4377),
.B(n_4028),
.Y(n_4411)
);

OAI21xp33_ASAP7_75t_L g4412 ( 
.A1(n_4394),
.A2(n_4042),
.B(n_4041),
.Y(n_4412)
);

NAND2xp5_ASAP7_75t_SL g4413 ( 
.A(n_4373),
.B(n_4042),
.Y(n_4413)
);

AOI22xp5_ASAP7_75t_L g4414 ( 
.A1(n_4396),
.A2(n_4054),
.B1(n_4056),
.B2(n_4062),
.Y(n_4414)
);

AOI22xp5_ASAP7_75t_L g4415 ( 
.A1(n_4380),
.A2(n_4062),
.B1(n_4091),
.B2(n_4096),
.Y(n_4415)
);

AND2x2_ASAP7_75t_L g4416 ( 
.A(n_4382),
.B(n_4395),
.Y(n_4416)
);

AND2x2_ASAP7_75t_L g4417 ( 
.A(n_4378),
.B(n_4051),
.Y(n_4417)
);

INVx2_ASAP7_75t_L g4418 ( 
.A(n_4375),
.Y(n_4418)
);

NOR3xp33_ASAP7_75t_SL g4419 ( 
.A(n_4376),
.B(n_4103),
.C(n_173),
.Y(n_4419)
);

INVx1_ASAP7_75t_L g4420 ( 
.A(n_4388),
.Y(n_4420)
);

NAND4xp25_ASAP7_75t_L g4421 ( 
.A(n_4403),
.B(n_4408),
.C(n_4410),
.D(n_4404),
.Y(n_4421)
);

INVx2_ASAP7_75t_L g4422 ( 
.A(n_4417),
.Y(n_4422)
);

OAI322xp33_ASAP7_75t_L g4423 ( 
.A1(n_4405),
.A2(n_4060),
.A3(n_4083),
.B1(n_4051),
.B2(n_4080),
.C1(n_4103),
.C2(n_3848),
.Y(n_4423)
);

OAI322xp33_ASAP7_75t_L g4424 ( 
.A1(n_4411),
.A2(n_4060),
.A3(n_4083),
.B1(n_4080),
.B2(n_4103),
.C1(n_3848),
.C2(n_3835),
.Y(n_4424)
);

NAND2xp5_ASAP7_75t_SL g4425 ( 
.A(n_4406),
.B(n_3869),
.Y(n_4425)
);

NOR2x1p5_ASAP7_75t_SL g4426 ( 
.A(n_4420),
.B(n_4103),
.Y(n_4426)
);

INVx1_ASAP7_75t_L g4427 ( 
.A(n_4409),
.Y(n_4427)
);

NAND3xp33_ASAP7_75t_L g4428 ( 
.A(n_4402),
.B(n_3878),
.C(n_3832),
.Y(n_4428)
);

NAND4xp75_ASAP7_75t_L g4429 ( 
.A(n_4401),
.B(n_174),
.C(n_175),
.D(n_177),
.Y(n_4429)
);

NAND4xp75_ASAP7_75t_L g4430 ( 
.A(n_4416),
.B(n_174),
.C(n_179),
.D(n_180),
.Y(n_4430)
);

AOI211xp5_ASAP7_75t_L g4431 ( 
.A1(n_4400),
.A2(n_4103),
.B(n_182),
.C(n_183),
.Y(n_4431)
);

NOR2x1p5_ASAP7_75t_SL g4432 ( 
.A(n_4418),
.B(n_4419),
.Y(n_4432)
);

NAND2xp5_ASAP7_75t_SL g4433 ( 
.A(n_4397),
.B(n_3869),
.Y(n_4433)
);

NAND5xp2_ASAP7_75t_L g4434 ( 
.A(n_4398),
.B(n_179),
.C(n_182),
.D(n_184),
.E(n_185),
.Y(n_4434)
);

NAND3xp33_ASAP7_75t_L g4435 ( 
.A(n_4413),
.B(n_3836),
.C(n_3830),
.Y(n_4435)
);

OR2x2_ASAP7_75t_L g4436 ( 
.A(n_4415),
.B(n_3830),
.Y(n_4436)
);

NOR3xp33_ASAP7_75t_L g4437 ( 
.A(n_4399),
.B(n_184),
.C(n_187),
.Y(n_4437)
);

NAND3xp33_ASAP7_75t_L g4438 ( 
.A(n_4421),
.B(n_4407),
.C(n_4412),
.Y(n_4438)
);

NOR4xp25_ASAP7_75t_L g4439 ( 
.A(n_4427),
.B(n_4414),
.C(n_3773),
.D(n_3774),
.Y(n_4439)
);

NOR3x1_ASAP7_75t_L g4440 ( 
.A(n_4429),
.B(n_4430),
.C(n_4428),
.Y(n_4440)
);

NOR2x1_ASAP7_75t_L g4441 ( 
.A(n_4422),
.B(n_187),
.Y(n_4441)
);

NOR4xp25_ASAP7_75t_L g4442 ( 
.A(n_4423),
.B(n_3773),
.C(n_3774),
.D(n_3783),
.Y(n_4442)
);

NAND2xp5_ASAP7_75t_L g4443 ( 
.A(n_4437),
.B(n_3836),
.Y(n_4443)
);

OAI211xp5_ASAP7_75t_SL g4444 ( 
.A1(n_4431),
.A2(n_188),
.B(n_189),
.C(n_190),
.Y(n_4444)
);

NOR3xp33_ASAP7_75t_L g4445 ( 
.A(n_4434),
.B(n_188),
.C(n_190),
.Y(n_4445)
);

NOR2x1_ASAP7_75t_L g4446 ( 
.A(n_4424),
.B(n_4425),
.Y(n_4446)
);

NOR3xp33_ASAP7_75t_L g4447 ( 
.A(n_4432),
.B(n_191),
.C(n_192),
.Y(n_4447)
);

AOI211xp5_ASAP7_75t_L g4448 ( 
.A1(n_4436),
.A2(n_191),
.B(n_192),
.C(n_193),
.Y(n_4448)
);

NOR2x1p5_ASAP7_75t_SL g4449 ( 
.A(n_4426),
.B(n_3841),
.Y(n_4449)
);

OAI211xp5_ASAP7_75t_L g4450 ( 
.A1(n_4433),
.A2(n_193),
.B(n_196),
.C(n_197),
.Y(n_4450)
);

AO22x1_ASAP7_75t_L g4451 ( 
.A1(n_4435),
.A2(n_3841),
.B1(n_3781),
.B2(n_3786),
.Y(n_4451)
);

NAND2xp5_ASAP7_75t_L g4452 ( 
.A(n_4437),
.B(n_3869),
.Y(n_4452)
);

AOI21xp33_ASAP7_75t_SL g4453 ( 
.A1(n_4447),
.A2(n_196),
.B(n_198),
.Y(n_4453)
);

OAI21xp33_ASAP7_75t_SL g4454 ( 
.A1(n_4441),
.A2(n_3783),
.B(n_3862),
.Y(n_4454)
);

NAND4xp25_ASAP7_75t_L g4455 ( 
.A(n_4445),
.B(n_198),
.C(n_199),
.D(n_200),
.Y(n_4455)
);

OA22x2_ASAP7_75t_L g4456 ( 
.A1(n_4450),
.A2(n_3778),
.B1(n_3781),
.B2(n_3788),
.Y(n_4456)
);

NAND3xp33_ASAP7_75t_SL g4457 ( 
.A(n_4448),
.B(n_199),
.C(n_200),
.Y(n_4457)
);

OAI22x1_ASAP7_75t_L g4458 ( 
.A1(n_4438),
.A2(n_3877),
.B1(n_3874),
.B2(n_3873),
.Y(n_4458)
);

AOI211xp5_ASAP7_75t_SL g4459 ( 
.A1(n_4444),
.A2(n_201),
.B(n_202),
.C(n_203),
.Y(n_4459)
);

O2A1O1Ixp5_ASAP7_75t_L g4460 ( 
.A1(n_4452),
.A2(n_3877),
.B(n_3874),
.C(n_3873),
.Y(n_4460)
);

AOI22xp5_ASAP7_75t_L g4461 ( 
.A1(n_4443),
.A2(n_4446),
.B1(n_4439),
.B2(n_4442),
.Y(n_4461)
);

OAI211xp5_ASAP7_75t_L g4462 ( 
.A1(n_4440),
.A2(n_4449),
.B(n_4451),
.C(n_204),
.Y(n_4462)
);

BUFx2_ASAP7_75t_L g4463 ( 
.A(n_4441),
.Y(n_4463)
);

OAI22xp33_ASAP7_75t_L g4464 ( 
.A1(n_4443),
.A2(n_3868),
.B1(n_3865),
.B2(n_3862),
.Y(n_4464)
);

O2A1O1Ixp33_ASAP7_75t_L g4465 ( 
.A1(n_4447),
.A2(n_201),
.B(n_203),
.C(n_205),
.Y(n_4465)
);

OAI21xp33_ASAP7_75t_L g4466 ( 
.A1(n_4445),
.A2(n_3868),
.B(n_207),
.Y(n_4466)
);

OAI22xp5_ASAP7_75t_L g4467 ( 
.A1(n_4438),
.A2(n_205),
.B1(n_207),
.B2(n_208),
.Y(n_4467)
);

OAI211xp5_ASAP7_75t_SL g4468 ( 
.A1(n_4446),
.A2(n_211),
.B(n_212),
.C(n_213),
.Y(n_4468)
);

AOI221xp5_ASAP7_75t_L g4469 ( 
.A1(n_4439),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.C(n_215),
.Y(n_4469)
);

OAI221xp5_ASAP7_75t_SL g4470 ( 
.A1(n_4445),
.A2(n_214),
.B1(n_215),
.B2(n_217),
.C(n_218),
.Y(n_4470)
);

AO22x1_ASAP7_75t_L g4471 ( 
.A1(n_4463),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_4471)
);

INVx1_ASAP7_75t_L g4472 ( 
.A(n_4465),
.Y(n_4472)
);

AOI22xp5_ASAP7_75t_L g4473 ( 
.A1(n_4455),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_4473)
);

INVx2_ASAP7_75t_L g4474 ( 
.A(n_4458),
.Y(n_4474)
);

INVx1_ASAP7_75t_L g4475 ( 
.A(n_4468),
.Y(n_4475)
);

NAND2xp5_ASAP7_75t_L g4476 ( 
.A(n_4469),
.B(n_223),
.Y(n_4476)
);

INVx2_ASAP7_75t_L g4477 ( 
.A(n_4456),
.Y(n_4477)
);

INVx1_ASAP7_75t_L g4478 ( 
.A(n_4457),
.Y(n_4478)
);

AOI22xp5_ASAP7_75t_L g4479 ( 
.A1(n_4466),
.A2(n_224),
.B1(n_230),
.B2(n_231),
.Y(n_4479)
);

AND2x4_ASAP7_75t_L g4480 ( 
.A(n_4461),
.B(n_224),
.Y(n_4480)
);

CKINVDCx20_ASAP7_75t_R g4481 ( 
.A(n_4467),
.Y(n_4481)
);

OR2x2_ASAP7_75t_L g4482 ( 
.A(n_4470),
.B(n_4453),
.Y(n_4482)
);

NAND2xp5_ASAP7_75t_L g4483 ( 
.A(n_4459),
.B(n_231),
.Y(n_4483)
);

INVx2_ASAP7_75t_L g4484 ( 
.A(n_4460),
.Y(n_4484)
);

INVx1_ASAP7_75t_L g4485 ( 
.A(n_4462),
.Y(n_4485)
);

INVx1_ASAP7_75t_L g4486 ( 
.A(n_4454),
.Y(n_4486)
);

INVx1_ASAP7_75t_L g4487 ( 
.A(n_4464),
.Y(n_4487)
);

NOR4xp75_ASAP7_75t_SL g4488 ( 
.A(n_4483),
.B(n_232),
.C(n_233),
.D(n_234),
.Y(n_4488)
);

AND2x2_ASAP7_75t_L g4489 ( 
.A(n_4480),
.B(n_234),
.Y(n_4489)
);

OAI22xp5_ASAP7_75t_L g4490 ( 
.A1(n_4473),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.Y(n_4490)
);

NOR2x1_ASAP7_75t_L g4491 ( 
.A(n_4486),
.B(n_235),
.Y(n_4491)
);

AND3x4_ASAP7_75t_L g4492 ( 
.A(n_4477),
.B(n_4474),
.C(n_4484),
.Y(n_4492)
);

NAND2xp5_ASAP7_75t_L g4493 ( 
.A(n_4479),
.B(n_236),
.Y(n_4493)
);

NOR2x1_ASAP7_75t_L g4494 ( 
.A(n_4478),
.B(n_238),
.Y(n_4494)
);

NOR2xp33_ASAP7_75t_R g4495 ( 
.A(n_4481),
.B(n_239),
.Y(n_4495)
);

NAND2xp5_ASAP7_75t_L g4496 ( 
.A(n_4475),
.B(n_240),
.Y(n_4496)
);

NOR2xp33_ASAP7_75t_R g4497 ( 
.A(n_4485),
.B(n_241),
.Y(n_4497)
);

NAND3xp33_ASAP7_75t_L g4498 ( 
.A(n_4487),
.B(n_1431),
.C(n_287),
.Y(n_4498)
);

OAI221xp5_ASAP7_75t_L g4499 ( 
.A1(n_4496),
.A2(n_4476),
.B1(n_4472),
.B2(n_4482),
.C(n_4471),
.Y(n_4499)
);

NAND4xp75_ASAP7_75t_L g4500 ( 
.A(n_4491),
.B(n_286),
.C(n_292),
.D(n_294),
.Y(n_4500)
);

INVx1_ASAP7_75t_L g4501 ( 
.A(n_4494),
.Y(n_4501)
);

O2A1O1Ixp33_ASAP7_75t_L g4502 ( 
.A1(n_4490),
.A2(n_295),
.B(n_296),
.C(n_301),
.Y(n_4502)
);

NOR2x1_ASAP7_75t_SL g4503 ( 
.A(n_4489),
.B(n_303),
.Y(n_4503)
);

NOR3xp33_ASAP7_75t_L g4504 ( 
.A(n_4493),
.B(n_306),
.C(n_309),
.Y(n_4504)
);

INVx1_ASAP7_75t_L g4505 ( 
.A(n_4503),
.Y(n_4505)
);

OAI22xp5_ASAP7_75t_L g4506 ( 
.A1(n_4499),
.A2(n_4492),
.B1(n_4498),
.B2(n_4501),
.Y(n_4506)
);

INVx1_ASAP7_75t_L g4507 ( 
.A(n_4500),
.Y(n_4507)
);

OAI21xp5_ASAP7_75t_L g4508 ( 
.A1(n_4506),
.A2(n_4502),
.B(n_4504),
.Y(n_4508)
);

AOI22xp5_ASAP7_75t_L g4509 ( 
.A1(n_4507),
.A2(n_4488),
.B1(n_4497),
.B2(n_4495),
.Y(n_4509)
);

OAI22xp5_ASAP7_75t_L g4510 ( 
.A1(n_4509),
.A2(n_4505),
.B1(n_4508),
.B2(n_314),
.Y(n_4510)
);

OAI211xp5_ASAP7_75t_SL g4511 ( 
.A1(n_4510),
.A2(n_311),
.B(n_313),
.C(n_317),
.Y(n_4511)
);

BUFx2_ASAP7_75t_L g4512 ( 
.A(n_4511),
.Y(n_4512)
);

INVx2_ASAP7_75t_L g4513 ( 
.A(n_4512),
.Y(n_4513)
);

OAI21xp5_ASAP7_75t_L g4514 ( 
.A1(n_4513),
.A2(n_319),
.B(n_321),
.Y(n_4514)
);

NAND2xp5_ASAP7_75t_L g4515 ( 
.A(n_4514),
.B(n_322),
.Y(n_4515)
);

AOI21xp5_ASAP7_75t_L g4516 ( 
.A1(n_4515),
.A2(n_324),
.B(n_330),
.Y(n_4516)
);

NAND3xp33_ASAP7_75t_L g4517 ( 
.A(n_4516),
.B(n_332),
.C(n_334),
.Y(n_4517)
);

AOI222xp33_ASAP7_75t_L g4518 ( 
.A1(n_4517),
.A2(n_1445),
.B1(n_340),
.B2(n_342),
.C1(n_343),
.C2(n_344),
.Y(n_4518)
);

BUFx2_ASAP7_75t_L g4519 ( 
.A(n_4518),
.Y(n_4519)
);

AOI221xp5_ASAP7_75t_L g4520 ( 
.A1(n_4519),
.A2(n_335),
.B1(n_346),
.B2(n_354),
.C(n_355),
.Y(n_4520)
);

AOI22xp5_ASAP7_75t_L g4521 ( 
.A1(n_4519),
.A2(n_1445),
.B1(n_357),
.B2(n_360),
.Y(n_4521)
);

AOI22xp33_ASAP7_75t_L g4522 ( 
.A1(n_4521),
.A2(n_1445),
.B1(n_361),
.B2(n_367),
.Y(n_4522)
);

AOI21xp33_ASAP7_75t_SL g4523 ( 
.A1(n_4520),
.A2(n_356),
.B(n_370),
.Y(n_4523)
);

AOI211xp5_ASAP7_75t_L g4524 ( 
.A1(n_4523),
.A2(n_4522),
.B(n_376),
.C(n_377),
.Y(n_4524)
);


endmodule