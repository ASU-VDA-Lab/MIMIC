module real_aes_2144_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_746;
wire n_153;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_0), .B(n_472), .Y(n_486) );
AOI222xp33_ASAP7_75t_L g102 ( .A1(n_1), .A2(n_103), .B1(n_759), .B2(n_770), .C1(n_786), .C2(n_788), .Y(n_102) );
AOI22xp5_ASAP7_75t_SL g775 ( .A1(n_1), .A2(n_776), .B1(n_779), .B2(n_780), .Y(n_775) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_1), .Y(n_780) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_2), .A2(n_471), .B(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_3), .B(n_766), .Y(n_765) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_4), .B(n_255), .Y(n_497) );
INVx1_ASAP7_75t_L g129 ( .A(n_5), .Y(n_129) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_6), .B(n_148), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_7), .B(n_255), .Y(n_526) );
INVx1_ASAP7_75t_L g157 ( .A(n_8), .Y(n_157) );
CKINVDCx16_ASAP7_75t_R g766 ( .A(n_9), .Y(n_766) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_10), .Y(n_174) );
NAND2xp33_ASAP7_75t_L g567 ( .A(n_11), .B(n_252), .Y(n_567) );
INVx2_ASAP7_75t_L g118 ( .A(n_12), .Y(n_118) );
AOI221x1_ASAP7_75t_L g470 ( .A1(n_13), .A2(n_26), .B1(n_471), .B2(n_472), .C(n_473), .Y(n_470) );
CKINVDCx16_ASAP7_75t_R g453 ( .A(n_14), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_15), .B(n_472), .Y(n_563) );
INVx1_ASAP7_75t_L g253 ( .A(n_16), .Y(n_253) );
AO21x2_ASAP7_75t_L g561 ( .A1(n_17), .A2(n_154), .B(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_18), .B(n_200), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_19), .B(n_255), .Y(n_550) );
AO21x1_ASAP7_75t_L g492 ( .A1(n_20), .A2(n_472), .B(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g457 ( .A(n_21), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_22), .Y(n_785) );
INVx1_ASAP7_75t_L g250 ( .A(n_23), .Y(n_250) );
INVx1_ASAP7_75t_SL g215 ( .A(n_24), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_25), .B(n_135), .Y(n_236) );
AOI33xp33_ASAP7_75t_L g186 ( .A1(n_27), .A2(n_56), .A3(n_124), .B1(n_133), .B2(n_187), .B3(n_188), .Y(n_186) );
NAND2x1_ASAP7_75t_L g484 ( .A(n_28), .B(n_255), .Y(n_484) );
NAND2x1_ASAP7_75t_L g525 ( .A(n_29), .B(n_252), .Y(n_525) );
INVx1_ASAP7_75t_L g166 ( .A(n_30), .Y(n_166) );
OA21x2_ASAP7_75t_L g117 ( .A1(n_31), .A2(n_88), .B(n_118), .Y(n_117) );
OR2x2_ASAP7_75t_L g149 ( .A(n_31), .B(n_88), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_32), .B(n_143), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_33), .B(n_252), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_34), .A2(n_93), .B1(n_747), .B2(n_748), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_34), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_35), .B(n_255), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_36), .B(n_252), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_37), .A2(n_471), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g123 ( .A(n_38), .Y(n_123) );
AND2x2_ASAP7_75t_L g141 ( .A(n_38), .B(n_129), .Y(n_141) );
AND2x2_ASAP7_75t_L g147 ( .A(n_38), .B(n_126), .Y(n_147) );
OR2x6_ASAP7_75t_L g455 ( .A(n_39), .B(n_456), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_40), .A2(n_745), .B1(n_750), .B2(n_755), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g169 ( .A(n_41), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g776 ( .A1(n_42), .A2(n_53), .B1(n_777), .B2(n_778), .Y(n_776) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_42), .Y(n_777) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_43), .B(n_472), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_44), .B(n_143), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g229 ( .A1(n_45), .A2(n_116), .B1(n_148), .B2(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_46), .B(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_47), .B(n_135), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_48), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_49), .B(n_252), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_50), .B(n_154), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_51), .B(n_135), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_52), .A2(n_471), .B(n_524), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_53), .Y(n_778) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_54), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_55), .B(n_252), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_57), .B(n_135), .Y(n_198) );
INVx1_ASAP7_75t_L g128 ( .A(n_58), .Y(n_128) );
INVx1_ASAP7_75t_L g137 ( .A(n_58), .Y(n_137) );
AND2x2_ASAP7_75t_L g199 ( .A(n_59), .B(n_200), .Y(n_199) );
AOI221xp5_ASAP7_75t_L g155 ( .A1(n_60), .A2(n_76), .B1(n_121), .B2(n_143), .C(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_61), .B(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_62), .B(n_255), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_63), .B(n_116), .Y(n_176) );
AOI21xp5_ASAP7_75t_SL g120 ( .A1(n_64), .A2(n_121), .B(n_130), .Y(n_120) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_65), .A2(n_471), .B(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g247 ( .A(n_66), .Y(n_247) );
AO21x1_ASAP7_75t_L g494 ( .A1(n_67), .A2(n_471), .B(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_68), .B(n_472), .Y(n_515) );
INVx1_ASAP7_75t_L g197 ( .A(n_69), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_70), .B(n_472), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_71), .A2(n_121), .B(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g508 ( .A(n_72), .B(n_201), .Y(n_508) );
INVx1_ASAP7_75t_L g126 ( .A(n_73), .Y(n_126) );
INVx1_ASAP7_75t_L g139 ( .A(n_73), .Y(n_139) );
AND2x2_ASAP7_75t_L g528 ( .A(n_74), .B(n_115), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_75), .B(n_143), .Y(n_189) );
AND2x2_ASAP7_75t_L g217 ( .A(n_77), .B(n_115), .Y(n_217) );
INVx1_ASAP7_75t_L g248 ( .A(n_78), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_79), .A2(n_121), .B(n_214), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_80), .A2(n_121), .B(n_181), .C(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g458 ( .A(n_81), .Y(n_458) );
AND2x2_ASAP7_75t_L g513 ( .A(n_82), .B(n_115), .Y(n_513) );
AND2x2_ASAP7_75t_SL g114 ( .A(n_83), .B(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_84), .B(n_472), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_85), .A2(n_121), .B1(n_184), .B2(n_185), .Y(n_183) );
XNOR2xp5_ASAP7_75t_L g745 ( .A(n_86), .B(n_746), .Y(n_745) );
AND2x2_ASAP7_75t_L g493 ( .A(n_87), .B(n_148), .Y(n_493) );
AND2x2_ASAP7_75t_L g487 ( .A(n_89), .B(n_115), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_90), .B(n_252), .Y(n_551) );
INVx1_ASAP7_75t_L g131 ( .A(n_91), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_92), .B(n_255), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_93), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_94), .B(n_252), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_95), .A2(n_471), .B(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g190 ( .A(n_96), .B(n_115), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_97), .B(n_255), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g163 ( .A1(n_98), .A2(n_164), .B(n_165), .C(n_168), .Y(n_163) );
BUFx2_ASAP7_75t_L g767 ( .A(n_99), .Y(n_767) );
BUFx2_ASAP7_75t_SL g792 ( .A(n_99), .Y(n_792) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_100), .A2(n_471), .B(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_101), .B(n_135), .Y(n_134) );
OAI21xp5_ASAP7_75t_SL g103 ( .A1(n_104), .A2(n_745), .B(n_749), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OAI22xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_450), .B1(n_459), .B2(n_463), .Y(n_105) );
INVx2_ASAP7_75t_L g754 ( .A(n_106), .Y(n_754) );
BUFx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
NAND3x1_ASAP7_75t_L g107 ( .A(n_108), .B(n_340), .C(n_405), .Y(n_107) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_294), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_239), .B(n_267), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_202), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_150), .Y(n_111) );
AOI21xp33_ASAP7_75t_L g341 ( .A1(n_112), .A2(n_342), .B(n_353), .Y(n_341) );
AND2x2_ASAP7_75t_SL g376 ( .A(n_112), .B(n_283), .Y(n_376) );
AND2x2_ASAP7_75t_L g391 ( .A(n_112), .B(n_392), .Y(n_391) );
OR2x6_ASAP7_75t_L g401 ( .A(n_112), .B(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g403 ( .A(n_112), .B(n_393), .Y(n_403) );
BUFx6f_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g277 ( .A(n_113), .Y(n_277) );
AND2x2_ASAP7_75t_L g290 ( .A(n_113), .B(n_291), .Y(n_290) );
INVx4_ASAP7_75t_L g309 ( .A(n_113), .Y(n_309) );
AND2x2_ASAP7_75t_L g312 ( .A(n_113), .B(n_228), .Y(n_312) );
NOR2x1_ASAP7_75t_SL g315 ( .A(n_113), .B(n_243), .Y(n_315) );
AND2x4_ASAP7_75t_L g327 ( .A(n_113), .B(n_325), .Y(n_327) );
OR2x2_ASAP7_75t_L g337 ( .A(n_113), .B(n_209), .Y(n_337) );
NAND2xp5_ASAP7_75t_SL g354 ( .A(n_113), .B(n_349), .Y(n_354) );
OR2x6_ASAP7_75t_L g113 ( .A(n_114), .B(n_119), .Y(n_113) );
OAI22xp5_ASAP7_75t_L g162 ( .A1(n_115), .A2(n_163), .B1(n_169), .B2(n_170), .Y(n_162) );
INVx3_ASAP7_75t_L g170 ( .A(n_115), .Y(n_170) );
INVx4_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_116), .B(n_173), .Y(n_172) );
INVx3_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
BUFx4f_ASAP7_75t_L g154 ( .A(n_117), .Y(n_154) );
AND2x4_ASAP7_75t_L g148 ( .A(n_118), .B(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_SL g201 ( .A(n_118), .B(n_149), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_142), .B(n_148), .Y(n_119) );
INVxp67_ASAP7_75t_L g175 ( .A(n_121), .Y(n_175) );
AND2x4_ASAP7_75t_L g121 ( .A(n_122), .B(n_127), .Y(n_121) );
NOR2x1p5_ASAP7_75t_L g122 ( .A(n_123), .B(n_124), .Y(n_122) );
INVx1_ASAP7_75t_L g188 ( .A(n_124), .Y(n_188) );
INVx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OR2x6_ASAP7_75t_L g132 ( .A(n_125), .B(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x6_ASAP7_75t_L g252 ( .A(n_126), .B(n_136), .Y(n_252) );
AND2x6_ASAP7_75t_L g471 ( .A(n_127), .B(n_147), .Y(n_471) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
INVx2_ASAP7_75t_L g133 ( .A(n_128), .Y(n_133) );
AND2x4_ASAP7_75t_L g255 ( .A(n_128), .B(n_138), .Y(n_255) );
HB1xp67_ASAP7_75t_L g145 ( .A(n_129), .Y(n_145) );
O2A1O1Ixp33_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_132), .B(n_134), .C(n_140), .Y(n_130) );
O2A1O1Ixp33_ASAP7_75t_SL g156 ( .A1(n_132), .A2(n_140), .B(n_157), .C(n_158), .Y(n_156) );
INVxp67_ASAP7_75t_L g164 ( .A(n_132), .Y(n_164) );
O2A1O1Ixp33_ASAP7_75t_L g196 ( .A1(n_132), .A2(n_140), .B(n_197), .C(n_198), .Y(n_196) );
O2A1O1Ixp33_ASAP7_75t_SL g214 ( .A1(n_132), .A2(n_140), .B(n_215), .C(n_216), .Y(n_214) );
INVx2_ASAP7_75t_L g238 ( .A(n_132), .Y(n_238) );
OAI22xp5_ASAP7_75t_L g246 ( .A1(n_132), .A2(n_167), .B1(n_247), .B2(n_248), .Y(n_246) );
AND2x2_ASAP7_75t_L g144 ( .A(n_133), .B(n_145), .Y(n_144) );
INVxp33_ASAP7_75t_L g187 ( .A(n_133), .Y(n_187) );
INVx1_ASAP7_75t_L g167 ( .A(n_135), .Y(n_167) );
AND2x4_ASAP7_75t_L g472 ( .A(n_135), .B(n_141), .Y(n_472) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_138), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g184 ( .A(n_140), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_140), .A2(n_236), .B(n_237), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_140), .B(n_148), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_140), .A2(n_474), .B(n_475), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_140), .A2(n_484), .B(n_485), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_140), .A2(n_496), .B(n_497), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_140), .A2(n_505), .B(n_506), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_140), .A2(n_518), .B(n_519), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_140), .A2(n_525), .B(n_526), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_140), .A2(n_550), .B(n_551), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_140), .A2(n_566), .B(n_567), .Y(n_565) );
INVx5_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
HB1xp67_ASAP7_75t_L g168 ( .A(n_141), .Y(n_168) );
INVx1_ASAP7_75t_L g177 ( .A(n_143), .Y(n_177) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_146), .Y(n_143) );
INVx1_ASAP7_75t_L g231 ( .A(n_144), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_146), .Y(n_232) );
BUFx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_148), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_SL g546 ( .A(n_148), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_148), .A2(n_563), .B(n_564), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g377 ( .A1(n_150), .A2(n_283), .B1(n_378), .B2(n_379), .Y(n_377) );
INVx1_ASAP7_75t_SL g421 ( .A(n_150), .Y(n_421) );
AND2x2_ASAP7_75t_L g150 ( .A(n_151), .B(n_178), .Y(n_150) );
INVx2_ASAP7_75t_L g352 ( .A(n_151), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_151), .B(n_298), .Y(n_424) );
AND2x2_ASAP7_75t_L g151 ( .A(n_152), .B(n_160), .Y(n_151) );
BUFx3_ASAP7_75t_L g270 ( .A(n_152), .Y(n_270) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g263 ( .A(n_153), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_153), .B(n_180), .Y(n_285) );
AND2x4_ASAP7_75t_L g302 ( .A(n_153), .B(n_303), .Y(n_302) );
INVxp67_ASAP7_75t_L g318 ( .A(n_153), .Y(n_318) );
INVx2_ASAP7_75t_L g375 ( .A(n_153), .Y(n_375) );
OA21x2_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_155), .B(n_159), .Y(n_153) );
INVx2_ASAP7_75t_SL g181 ( .A(n_154), .Y(n_181) );
AND2x2_ASAP7_75t_L g293 ( .A(n_160), .B(n_259), .Y(n_293) );
NOR2xp67_ASAP7_75t_L g339 ( .A(n_160), .B(n_262), .Y(n_339) );
AND2x2_ASAP7_75t_L g358 ( .A(n_160), .B(n_262), .Y(n_358) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g220 ( .A(n_161), .Y(n_220) );
INVx1_ASAP7_75t_L g301 ( .A(n_161), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_161), .B(n_192), .Y(n_320) );
AND2x4_ASAP7_75t_L g374 ( .A(n_161), .B(n_375), .Y(n_374) );
OR2x2_ASAP7_75t_L g161 ( .A(n_162), .B(n_171), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
AO21x2_ASAP7_75t_L g192 ( .A1(n_170), .A2(n_193), .B(n_199), .Y(n_192) );
AO21x2_ASAP7_75t_L g262 ( .A1(n_170), .A2(n_193), .B(n_199), .Y(n_262) );
AO21x2_ASAP7_75t_L g480 ( .A1(n_170), .A2(n_481), .B(n_487), .Y(n_480) );
AO21x2_ASAP7_75t_L g501 ( .A1(n_170), .A2(n_502), .B(n_508), .Y(n_501) );
AO21x2_ASAP7_75t_L g535 ( .A1(n_170), .A2(n_502), .B(n_508), .Y(n_535) );
AO21x2_ASAP7_75t_L g539 ( .A1(n_170), .A2(n_481), .B(n_487), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_175), .B1(n_176), .B2(n_177), .Y(n_171) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g333 ( .A(n_178), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_178), .B(n_391), .Y(n_390) );
AND2x4_ASAP7_75t_L g178 ( .A(n_179), .B(n_191), .Y(n_178) );
AND2x2_ASAP7_75t_L g317 ( .A(n_179), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g357 ( .A(n_179), .Y(n_357) );
AND2x2_ASAP7_75t_L g362 ( .A(n_179), .B(n_262), .Y(n_362) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_180), .B(n_192), .Y(n_222) );
AO21x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_190), .Y(n_180) );
AO21x2_ASAP7_75t_L g259 ( .A1(n_181), .A2(n_182), .B(n_190), .Y(n_259) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_183), .B(n_189), .Y(n_182) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx3_ASAP7_75t_L g298 ( .A(n_191), .Y(n_298) );
NAND2x1p5_ASAP7_75t_L g416 ( .A(n_191), .B(n_270), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_191), .B(n_220), .Y(n_437) );
INVx3_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_192), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_200), .Y(n_210) );
OA21x2_ASAP7_75t_L g469 ( .A1(n_200), .A2(n_470), .B(n_476), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_200), .A2(n_515), .B(n_516), .Y(n_514) );
OA21x2_ASAP7_75t_L g615 ( .A1(n_200), .A2(n_470), .B(n_476), .Y(n_615) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
OAI21xp33_ASAP7_75t_SL g202 ( .A1(n_203), .A2(n_218), .B(n_223), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
HB1xp67_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_205), .B(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g275 ( .A(n_206), .Y(n_275) );
AND2x2_ASAP7_75t_L g289 ( .A(n_206), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g323 ( .A(n_206), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g389 ( .A(n_206), .B(n_307), .Y(n_389) );
NOR3xp33_ASAP7_75t_L g435 ( .A(n_206), .B(n_436), .C(n_437), .Y(n_435) );
INVx3_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_207), .Y(n_266) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g282 ( .A(n_209), .Y(n_282) );
AND2x2_ASAP7_75t_L g288 ( .A(n_209), .B(n_243), .Y(n_288) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_209), .Y(n_299) );
AND2x2_ASAP7_75t_L g344 ( .A(n_209), .B(n_242), .Y(n_344) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_209), .Y(n_367) );
INVx1_ASAP7_75t_L g384 ( .A(n_209), .Y(n_384) );
AO21x2_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_217), .Y(n_209) );
AO21x2_ASAP7_75t_L g521 ( .A1(n_210), .A2(n_522), .B(n_528), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
INVx1_ASAP7_75t_L g426 ( .A(n_218), .Y(n_426) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_221), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_219), .B(n_297), .Y(n_398) );
INVx1_ASAP7_75t_SL g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g260 ( .A(n_220), .B(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AOI211x1_ASAP7_75t_L g294 ( .A1(n_224), .A2(n_295), .B(n_304), .C(n_321), .Y(n_294) );
INVx2_ASAP7_75t_SL g224 ( .A(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_SL g287 ( .A(n_225), .B(n_288), .Y(n_287) );
AND2x4_ASAP7_75t_L g347 ( .A(n_225), .B(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g283 ( .A(n_227), .B(n_242), .Y(n_283) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x4_ASAP7_75t_L g241 ( .A(n_228), .B(n_242), .Y(n_241) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_228), .Y(n_308) );
INVx1_ASAP7_75t_L g325 ( .A(n_228), .Y(n_325) );
AND2x2_ASAP7_75t_L g393 ( .A(n_228), .B(n_243), .Y(n_393) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_234), .Y(n_228) );
NOR3xp33_ASAP7_75t_L g230 ( .A(n_231), .B(n_232), .C(n_233), .Y(n_230) );
OAI21xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_257), .B(n_264), .Y(n_239) );
NOR2x1_ASAP7_75t_L g412 ( .A(n_240), .B(n_309), .Y(n_412) );
INVx2_ASAP7_75t_L g444 ( .A(n_240), .Y(n_444) );
INVx4_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g276 ( .A(n_241), .B(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g349 ( .A(n_242), .Y(n_349) );
INVx3_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g291 ( .A(n_243), .Y(n_291) );
AND2x4_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
OAI21xp5_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_249), .B(n_256), .Y(n_245) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_251), .B1(n_253), .B2(n_254), .Y(n_249) );
INVxp67_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVxp67_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_260), .Y(n_257) );
OR2x2_ASAP7_75t_L g351 ( .A(n_258), .B(n_352), .Y(n_351) );
NAND2x1_ASAP7_75t_SL g373 ( .A(n_258), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x4_ASAP7_75t_L g273 ( .A(n_259), .B(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g303 ( .A(n_259), .Y(n_303) );
INVx1_ASAP7_75t_L g427 ( .A(n_260), .Y(n_427) );
AND2x2_ASAP7_75t_L g292 ( .A(n_261), .B(n_293), .Y(n_292) );
NOR2x1_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
INVx2_ASAP7_75t_L g274 ( .A(n_262), .Y(n_274) );
INVxp33_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g331 ( .A(n_266), .B(n_324), .Y(n_331) );
OAI211xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_271), .B(n_278), .C(n_286), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g355 ( .A(n_269), .B(n_356), .Y(n_355) );
NOR2xp67_ASAP7_75t_SL g360 ( .A(n_269), .B(n_361), .Y(n_360) );
INVx3_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_270), .B(n_357), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_272), .B(n_276), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
AND2x2_ASAP7_75t_L g404 ( .A(n_273), .B(n_374), .Y(n_404) );
AOI222xp33_ASAP7_75t_L g422 ( .A1(n_276), .A2(n_423), .B1(n_425), .B2(n_428), .C1(n_429), .C2(n_432), .Y(n_422) );
INVx1_ASAP7_75t_L g386 ( .A(n_277), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_284), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
BUFx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_282), .Y(n_313) );
AND2x4_ASAP7_75t_SL g348 ( .A(n_282), .B(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g402 ( .A(n_283), .Y(n_402) );
AND2x2_ASAP7_75t_L g447 ( .A(n_283), .B(n_299), .Y(n_447) );
AND2x2_ASAP7_75t_L g328 ( .A(n_284), .B(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g441 ( .A(n_285), .B(n_320), .Y(n_441) );
OAI21xp33_ASAP7_75t_SL g286 ( .A1(n_287), .A2(n_289), .B(n_292), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g408 ( .A1(n_287), .A2(n_307), .B(n_348), .Y(n_408) );
AND2x2_ASAP7_75t_L g432 ( .A(n_288), .B(n_309), .Y(n_432) );
NOR2xp33_ASAP7_75t_SL g442 ( .A(n_288), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g380 ( .A(n_291), .Y(n_380) );
NOR2x1_ASAP7_75t_L g385 ( .A(n_291), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g415 ( .A(n_293), .Y(n_415) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_300), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
AND2x2_ASAP7_75t_L g418 ( .A(n_298), .B(n_302), .Y(n_418) );
BUFx2_ASAP7_75t_L g306 ( .A(n_299), .Y(n_306) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx1_ASAP7_75t_L g329 ( .A(n_301), .Y(n_329) );
INVx2_ASAP7_75t_L g335 ( .A(n_301), .Y(n_335) );
AND2x2_ASAP7_75t_L g371 ( .A(n_301), .B(n_362), .Y(n_371) );
AND2x4_ASAP7_75t_L g338 ( .A(n_302), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g378 ( .A(n_302), .B(n_335), .Y(n_378) );
AND2x2_ASAP7_75t_L g429 ( .A(n_302), .B(n_430), .Y(n_429) );
AOI31xp33_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_310), .A3(n_314), .B(n_316), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
AND2x2_ASAP7_75t_L g326 ( .A(n_306), .B(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_SL g307 ( .A(n_308), .B(n_309), .Y(n_307) );
AND2x4_ASAP7_75t_L g324 ( .A(n_309), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_312), .A2(n_364), .B1(n_395), .B2(n_398), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_312), .B(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g449 ( .A(n_312), .B(n_365), .Y(n_449) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g364 ( .A(n_315), .B(n_365), .Y(n_364) );
NAND2x1p5_ASAP7_75t_L g316 ( .A(n_317), .B(n_319), .Y(n_316) );
AND2x2_ASAP7_75t_L g387 ( .A(n_317), .B(n_358), .Y(n_387) );
INVx1_ASAP7_75t_L g397 ( .A(n_319), .Y(n_397) );
INVx2_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_322), .B(n_330), .Y(n_321) );
OAI21xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_326), .B(n_328), .Y(n_322) );
INVx1_ASAP7_75t_L g420 ( .A(n_323), .Y(n_420) );
AND2x2_ASAP7_75t_L g428 ( .A(n_324), .B(n_380), .Y(n_428) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_324), .Y(n_434) );
AND2x2_ASAP7_75t_L g379 ( .A(n_327), .B(n_380), .Y(n_379) );
AOI22xp33_ASAP7_75t_SL g330 ( .A1(n_331), .A2(n_332), .B1(n_336), .B2(n_338), .Y(n_330) );
NOR2xp33_ASAP7_75t_SL g332 ( .A(n_333), .B(n_334), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g445 ( .A1(n_333), .A2(n_352), .B1(n_446), .B2(n_448), .Y(n_445) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx2_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g345 ( .A(n_338), .Y(n_345) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_368), .Y(n_340) );
OAI21xp33_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_345), .B(n_346), .Y(n_342) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
OAI21xp33_ASAP7_75t_L g346 ( .A1(n_344), .A2(n_347), .B(n_350), .Y(n_346) );
AOI22xp33_ASAP7_75t_SL g370 ( .A1(n_347), .A2(n_371), .B1(n_372), .B2(n_376), .Y(n_370) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_355), .B1(n_359), .B2(n_363), .Y(n_353) );
INVx1_ASAP7_75t_L g388 ( .A(n_356), .Y(n_388) );
NAND2x1p5_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NOR2xp67_ASAP7_75t_L g368 ( .A(n_369), .B(n_381), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_370), .B(n_377), .Y(n_369) );
INVx2_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
NAND2xp33_ASAP7_75t_SL g423 ( .A(n_373), .B(n_424), .Y(n_423) );
INVx3_ASAP7_75t_L g396 ( .A(n_374), .Y(n_396) );
INVx3_ASAP7_75t_L g410 ( .A(n_378), .Y(n_410) );
INVxp67_ASAP7_75t_L g439 ( .A(n_379), .Y(n_439) );
NAND4xp25_ASAP7_75t_L g381 ( .A(n_382), .B(n_390), .C(n_394), .D(n_399), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_387), .B1(n_388), .B2(n_389), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
AND2x2_ASAP7_75t_L g392 ( .A(n_384), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g440 ( .A(n_388), .Y(n_440) );
NAND2xp33_ASAP7_75t_SL g395 ( .A(n_396), .B(n_397), .Y(n_395) );
OAI21xp33_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_403), .B(n_404), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AND3x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_422), .C(n_433), .Y(n_405) );
AOI221x1_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_409), .B1(n_411), .B2(n_413), .C(n_419), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NAND2xp33_ASAP7_75t_SL g413 ( .A(n_414), .B(n_417), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
NAND2xp33_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AOI211xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_435), .B(n_438), .C(n_445), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_440), .B1(n_441), .B2(n_442), .Y(n_438) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
CKINVDCx5p33_ASAP7_75t_R g753 ( .A(n_451), .Y(n_753) );
CKINVDCx11_ASAP7_75t_R g451 ( .A(n_452), .Y(n_451) );
OR2x6_ASAP7_75t_SL g452 ( .A(n_453), .B(n_454), .Y(n_452) );
AND2x6_ASAP7_75t_SL g462 ( .A(n_453), .B(n_455), .Y(n_462) );
OR2x2_ASAP7_75t_L g758 ( .A(n_453), .B(n_455), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_453), .B(n_454), .Y(n_769) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
CKINVDCx6p67_ASAP7_75t_R g459 ( .A(n_460), .Y(n_459) );
CKINVDCx11_ASAP7_75t_R g751 ( .A(n_460), .Y(n_751) );
INVx3_ASAP7_75t_SL g460 ( .A(n_461), .Y(n_460) );
CKINVDCx5p33_ASAP7_75t_R g461 ( .A(n_462), .Y(n_461) );
INVx3_ASAP7_75t_L g752 ( .A(n_463), .Y(n_752) );
XNOR2x2_ASAP7_75t_SL g774 ( .A(n_463), .B(n_775), .Y(n_774) );
NAND4xp75_ASAP7_75t_L g463 ( .A(n_464), .B(n_655), .C(n_695), .D(n_724), .Y(n_463) );
NOR2x1_ASAP7_75t_L g464 ( .A(n_465), .B(n_617), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_574), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_509), .B(n_529), .Y(n_466) );
AND2x2_ASAP7_75t_SL g467 ( .A(n_468), .B(n_477), .Y(n_467) );
AND2x4_ASAP7_75t_L g573 ( .A(n_468), .B(n_534), .Y(n_573) );
INVx1_ASAP7_75t_SL g626 ( .A(n_468), .Y(n_626) );
AOI21xp33_ASAP7_75t_L g661 ( .A1(n_468), .A2(n_662), .B(n_665), .Y(n_661) );
A2O1A1Ixp33_ASAP7_75t_SL g665 ( .A1(n_468), .A2(n_666), .B(n_667), .C(n_668), .Y(n_665) );
NAND2x1_ASAP7_75t_L g706 ( .A(n_468), .B(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_468), .B(n_667), .Y(n_728) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g532 ( .A(n_469), .Y(n_532) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_469), .Y(n_605) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_488), .Y(n_477) );
AND2x2_ASAP7_75t_L g597 ( .A(n_478), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g678 ( .A(n_478), .B(n_534), .Y(n_678) );
INVx1_ASAP7_75t_L g738 ( .A(n_478), .Y(n_738) );
BUFx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g582 ( .A(n_479), .B(n_500), .Y(n_582) );
AND2x2_ASAP7_75t_L g707 ( .A(n_479), .B(n_501), .Y(n_707) );
AND2x2_ASAP7_75t_L g712 ( .A(n_479), .B(n_672), .Y(n_712) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVxp67_ASAP7_75t_L g588 ( .A(n_480), .Y(n_588) );
BUFx3_ASAP7_75t_L g621 ( .A(n_480), .Y(n_621) );
AND2x2_ASAP7_75t_L g667 ( .A(n_480), .B(n_501), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_482), .B(n_486), .Y(n_481) );
AND2x2_ASAP7_75t_L g652 ( .A(n_488), .B(n_531), .Y(n_652) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_500), .Y(n_488) );
AND2x4_ASAP7_75t_L g534 ( .A(n_489), .B(n_535), .Y(n_534) );
OR2x2_ASAP7_75t_L g644 ( .A(n_489), .B(n_628), .Y(n_644) );
AND2x2_ASAP7_75t_SL g687 ( .A(n_489), .B(n_615), .Y(n_687) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx2_ASAP7_75t_L g623 ( .A(n_490), .Y(n_623) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g584 ( .A(n_491), .Y(n_584) );
OAI21x1_ASAP7_75t_SL g491 ( .A1(n_492), .A2(n_494), .B(n_498), .Y(n_491) );
INVx1_ASAP7_75t_L g499 ( .A(n_493), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_500), .B(n_584), .Y(n_587) );
AND2x2_ASAP7_75t_L g672 ( .A(n_500), .B(n_615), .Y(n_672) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g669 ( .A(n_501), .B(n_532), .Y(n_669) );
AND2x2_ASAP7_75t_L g689 ( .A(n_501), .B(n_615), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_503), .B(n_507), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_509), .B(n_578), .Y(n_607) );
AOI221xp5_ASAP7_75t_L g700 ( .A1(n_509), .A2(n_701), .B1(n_702), .B2(n_703), .C(n_705), .Y(n_700) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
OAI332xp33_ASAP7_75t_L g734 ( .A1(n_510), .A2(n_594), .A3(n_601), .B1(n_660), .B2(n_735), .B3(n_736), .C1(n_737), .C2(n_739), .Y(n_734) );
NAND2x1p5_ASAP7_75t_L g510 ( .A(n_511), .B(n_520), .Y(n_510) );
AND2x2_ASAP7_75t_L g540 ( .A(n_511), .B(n_521), .Y(n_540) );
AND2x2_ASAP7_75t_L g557 ( .A(n_511), .B(n_558), .Y(n_557) );
INVx4_ASAP7_75t_L g569 ( .A(n_511), .Y(n_569) );
AND2x2_ASAP7_75t_SL g629 ( .A(n_511), .B(n_570), .Y(n_629) );
INVx5_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NOR2x1_ASAP7_75t_SL g591 ( .A(n_512), .B(n_558), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_512), .B(n_520), .Y(n_595) );
AND2x2_ASAP7_75t_L g602 ( .A(n_512), .B(n_521), .Y(n_602) );
BUFx2_ASAP7_75t_L g637 ( .A(n_512), .Y(n_637) );
AND2x2_ASAP7_75t_L g692 ( .A(n_512), .B(n_561), .Y(n_692) );
OR2x6_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
OR2x2_ASAP7_75t_L g560 ( .A(n_520), .B(n_561), .Y(n_560) );
AND2x4_ASAP7_75t_L g570 ( .A(n_520), .B(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g610 ( .A(n_520), .Y(n_610) );
AND2x2_ASAP7_75t_L g680 ( .A(n_520), .B(n_579), .Y(n_680) );
AND2x2_ASAP7_75t_L g693 ( .A(n_520), .B(n_694), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_520), .B(n_694), .Y(n_711) );
INVx4_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_521), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_527), .Y(n_522) );
OAI32xp33_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_536), .A3(n_541), .B1(n_555), .B2(n_572), .Y(n_529) );
INVx2_ASAP7_75t_L g638 ( .A(n_530), .Y(n_638) );
OR2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_533), .Y(n_530) );
INVx1_ASAP7_75t_L g649 ( .A(n_531), .Y(n_649) );
BUFx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x4_ASAP7_75t_L g583 ( .A(n_532), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g716 ( .A(n_532), .B(n_621), .Y(n_716) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g628 ( .A(n_535), .Y(n_628) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_540), .Y(n_537) );
INVx2_ASAP7_75t_L g616 ( .A(n_538), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_538), .B(n_659), .Y(n_658) );
BUFx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x4_ASAP7_75t_SL g627 ( .A(n_539), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g704 ( .A(n_539), .Y(n_704) );
AND2x2_ASAP7_75t_L g722 ( .A(n_539), .B(n_584), .Y(n_722) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NOR2xp67_ASAP7_75t_SL g666 ( .A(n_542), .B(n_595), .Y(n_666) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_543), .B(n_577), .Y(n_664) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g740 ( .A(n_544), .B(n_610), .Y(n_740) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g571 ( .A(n_545), .Y(n_571) );
INVx2_ASAP7_75t_L g612 ( .A(n_545), .Y(n_612) );
AO21x2_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_547), .B(n_553), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_546), .B(n_554), .Y(n_553) );
AO21x2_ASAP7_75t_L g558 ( .A1(n_546), .A2(n_547), .B(n_553), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_552), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_556), .B(n_568), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_556), .B(n_614), .Y(n_699) );
AND2x4_ASAP7_75t_L g556 ( .A(n_557), .B(n_559), .Y(n_556) );
AND3x2_ASAP7_75t_L g654 ( .A(n_557), .B(n_601), .C(n_610), .Y(n_654) );
AND2x2_ASAP7_75t_L g578 ( .A(n_558), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_558), .B(n_561), .Y(n_635) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OR2x2_ASAP7_75t_L g589 ( .A(n_560), .B(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g579 ( .A(n_561), .Y(n_579) );
INVx1_ASAP7_75t_L g594 ( .A(n_561), .Y(n_594) );
BUFx3_ASAP7_75t_L g601 ( .A(n_561), .Y(n_601) );
AND2x2_ASAP7_75t_L g611 ( .A(n_561), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
AND2x4_ASAP7_75t_L g620 ( .A(n_569), .B(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_569), .B(n_579), .Y(n_663) );
AND2x2_ASAP7_75t_L g619 ( .A(n_570), .B(n_594), .Y(n_619) );
INVx2_ASAP7_75t_L g646 ( .A(n_570), .Y(n_646) );
INVx1_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
AOI211xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_580), .B(n_585), .C(n_606), .Y(n_574) );
OAI21xp5_ASAP7_75t_L g726 ( .A1(n_575), .A2(n_702), .B(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_578), .B(n_637), .Y(n_636) );
AOI211xp5_ASAP7_75t_SL g656 ( .A1(n_578), .A2(n_657), .B(n_661), .C(n_670), .Y(n_656) );
AND2x2_ASAP7_75t_L g642 ( .A(n_579), .B(n_602), .Y(n_642) );
OR2x2_ASAP7_75t_L g645 ( .A(n_579), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g732 ( .A(n_582), .B(n_687), .Y(n_732) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_583), .B(n_628), .Y(n_641) );
AOI221xp5_ASAP7_75t_L g697 ( .A1(n_583), .A2(n_609), .B1(n_689), .B2(n_692), .C(n_698), .Y(n_697) );
AND2x4_ASAP7_75t_L g614 ( .A(n_584), .B(n_615), .Y(n_614) );
OR2x2_ASAP7_75t_L g660 ( .A(n_584), .B(n_615), .Y(n_660) );
OAI221xp5_ASAP7_75t_SL g585 ( .A1(n_586), .A2(n_589), .B1(n_592), .B2(n_596), .C(n_599), .Y(n_585) );
AND2x2_ASAP7_75t_L g731 ( .A(n_586), .B(n_732), .Y(n_731) );
OR2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx1_ASAP7_75t_L g598 ( .A(n_587), .Y(n_598) );
INVx1_ASAP7_75t_L g684 ( .A(n_588), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_589), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g603 ( .A(n_591), .B(n_594), .Y(n_603) );
AND2x2_ASAP7_75t_L g679 ( .A(n_591), .B(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g604 ( .A(n_598), .B(n_605), .Y(n_604) );
OAI21xp5_ASAP7_75t_SL g599 ( .A1(n_600), .A2(n_603), .B(n_604), .Y(n_599) );
INVx1_ASAP7_75t_L g723 ( .A(n_600), .Y(n_723) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
AND2x2_ASAP7_75t_L g702 ( .A(n_601), .B(n_629), .Y(n_702) );
AND2x2_ASAP7_75t_SL g675 ( .A(n_602), .B(n_611), .Y(n_675) );
AOI21xp33_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_608), .B(n_613), .Y(n_606) );
OAI22xp33_ASAP7_75t_L g643 ( .A1(n_607), .A2(n_641), .B1(n_644), .B2(n_645), .Y(n_643) );
INVx1_ASAP7_75t_L g713 ( .A(n_607), .Y(n_713) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx1_ASAP7_75t_L g633 ( .A(n_610), .Y(n_633) );
INVx1_ASAP7_75t_L g694 ( .A(n_612), .Y(n_694) );
NAND2xp5_ASAP7_75t_SL g613 ( .A(n_614), .B(n_616), .Y(n_613) );
NAND2xp5_ASAP7_75t_SL g735 ( .A(n_614), .B(n_684), .Y(n_735) );
AND2x2_ASAP7_75t_L g703 ( .A(n_615), .B(n_704), .Y(n_703) );
OAI211xp5_ASAP7_75t_L g696 ( .A1(n_616), .A2(n_697), .B(n_700), .C(n_708), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_639), .Y(n_617) );
AOI322xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_620), .A3(n_622), .B1(n_624), .B2(n_629), .C1(n_630), .C2(n_638), .Y(n_618) );
CKINVDCx16_ASAP7_75t_R g736 ( .A(n_620), .Y(n_736) );
AND2x2_ASAP7_75t_L g686 ( .A(n_621), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_SL g720 ( .A(n_621), .Y(n_720) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NOR2xp33_ASAP7_75t_SL g671 ( .A(n_623), .B(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_SL g677 ( .A(n_623), .B(n_669), .Y(n_677) );
AND2x2_ASAP7_75t_L g701 ( .A(n_623), .B(n_667), .Y(n_701) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
INVx1_ASAP7_75t_L g673 ( .A(n_627), .Y(n_673) );
NAND2xp33_ASAP7_75t_SL g630 ( .A(n_631), .B(n_636), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AOI221xp5_ASAP7_75t_SL g676 ( .A1(n_632), .A2(n_677), .B1(n_678), .B2(n_679), .C(n_681), .Y(n_676) );
AND2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
INVxp67_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g743 ( .A(n_635), .Y(n_743) );
AOI211xp5_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_642), .B(n_643), .C(n_647), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_SL g718 ( .A(n_642), .Y(n_718) );
INVx1_ASAP7_75t_L g650 ( .A(n_644), .Y(n_650) );
OR2x2_ASAP7_75t_L g737 ( .A(n_644), .B(n_738), .Y(n_737) );
INVx2_ASAP7_75t_SL g733 ( .A(n_645), .Y(n_733) );
AOI21xp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_651), .B(n_653), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_649), .B(n_667), .Y(n_744) );
INVx1_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_676), .Y(n_655) );
INVx1_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_659), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
OR2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
OR2x2_ASAP7_75t_L g710 ( .A(n_663), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AOI21xp33_ASAP7_75t_SL g670 ( .A1(n_671), .A2(n_673), .B(n_674), .Y(n_670) );
INVx2_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
AOI31xp33_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_685), .A3(n_688), .B(n_690), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_687), .B(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
AND2x4_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AOI221xp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_712), .B1(n_713), .B2(n_714), .C(n_717), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVxp67_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_719), .B1(n_721), .B2(n_723), .Y(n_717) );
CKINVDCx16_ASAP7_75t_R g721 ( .A(n_722), .Y(n_721) );
NOR3xp33_ASAP7_75t_L g724 ( .A(n_725), .B(n_734), .C(n_741), .Y(n_724) );
NAND2xp5_ASAP7_75t_SL g725 ( .A(n_726), .B(n_729), .Y(n_725) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_733), .Y(n_729) );
INVxp67_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g741 ( .A(n_742), .B(n_744), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
OAI22x1_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_752), .B1(n_753), .B2(n_754), .Y(n_750) );
CKINVDCx5p33_ASAP7_75t_R g755 ( .A(n_756), .Y(n_755) );
CKINVDCx5p33_ASAP7_75t_R g756 ( .A(n_757), .Y(n_756) );
INVx3_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_SL g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_L g761 ( .A(n_762), .B(n_768), .Y(n_761) );
INVxp67_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
NAND2xp5_ASAP7_75t_SL g763 ( .A(n_764), .B(n_767), .Y(n_763) );
INVx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
OR2x2_ASAP7_75t_SL g787 ( .A(n_765), .B(n_767), .Y(n_787) );
AOI21xp5_ASAP7_75t_L g789 ( .A1(n_765), .A2(n_790), .B(n_793), .Y(n_789) );
BUFx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
BUFx3_ASAP7_75t_L g773 ( .A(n_769), .Y(n_773) );
BUFx2_ASAP7_75t_L g794 ( .A(n_769), .Y(n_794) );
INVxp67_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
AOI21xp5_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_774), .B(n_781), .Y(n_771) );
HB1xp67_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_773), .Y(n_784) );
INVx1_ASAP7_75t_L g779 ( .A(n_776), .Y(n_779) );
NOR2xp33_ASAP7_75t_SL g781 ( .A(n_782), .B(n_785), .Y(n_781) );
INVx1_ASAP7_75t_SL g782 ( .A(n_783), .Y(n_782) );
BUFx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_SL g788 ( .A(n_789), .Y(n_788) );
CKINVDCx11_ASAP7_75t_R g790 ( .A(n_791), .Y(n_790) );
CKINVDCx8_ASAP7_75t_R g791 ( .A(n_792), .Y(n_791) );
INVx2_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
endmodule