module real_aes_617_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_531, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_531;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_417;
wire n_363;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_0), .A2(n_178), .B1(n_179), .B2(n_182), .Y(n_177) );
INVx1_ASAP7_75t_L g182 ( .A(n_0), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_1), .B(n_223), .Y(n_249) );
AO22x2_ASAP7_75t_L g88 ( .A1(n_2), .A2(n_55), .B1(n_89), .B2(n_90), .Y(n_88) );
INVx1_ASAP7_75t_L g195 ( .A(n_3), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_4), .B(n_208), .Y(n_274) );
NAND2xp33_ASAP7_75t_SL g316 ( .A(n_5), .B(n_214), .Y(n_316) );
INVx1_ASAP7_75t_L g309 ( .A(n_6), .Y(n_309) );
AO22x2_ASAP7_75t_L g92 ( .A1(n_7), .A2(n_16), .B1(n_89), .B2(n_93), .Y(n_92) );
AND2x2_ASAP7_75t_L g272 ( .A(n_8), .B(n_231), .Y(n_272) );
INVx2_ASAP7_75t_L g229 ( .A(n_9), .Y(n_229) );
AOI221x1_ASAP7_75t_L g311 ( .A1(n_10), .A2(n_216), .B1(n_312), .B2(n_314), .C(n_315), .Y(n_311) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_11), .B(n_208), .Y(n_207) );
AOI22xp33_ASAP7_75t_L g119 ( .A1(n_12), .A2(n_33), .B1(n_120), .B2(n_127), .Y(n_119) );
AOI221xp5_ASAP7_75t_SL g238 ( .A1(n_13), .A2(n_30), .B1(n_208), .B2(n_216), .C(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_14), .B(n_223), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_15), .A2(n_216), .B(n_276), .Y(n_275) );
OAI221xp5_ASAP7_75t_L g187 ( .A1(n_16), .A2(n_55), .B1(n_57), .B2(n_188), .C(n_190), .Y(n_187) );
OA21x2_ASAP7_75t_L g228 ( .A1(n_17), .A2(n_71), .B(n_229), .Y(n_228) );
OR2x2_ASAP7_75t_L g232 ( .A(n_17), .B(n_71), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g179 ( .A1(n_18), .A2(n_22), .B1(n_180), .B2(n_181), .Y(n_179) );
INVxp67_ASAP7_75t_L g180 ( .A(n_18), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_19), .B(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g298 ( .A(n_20), .B(n_237), .Y(n_298) );
AOI22xp33_ASAP7_75t_L g146 ( .A1(n_21), .A2(n_37), .B1(n_147), .B2(n_151), .Y(n_146) );
INVx1_ASAP7_75t_L g181 ( .A(n_22), .Y(n_181) );
INVx3_ASAP7_75t_L g89 ( .A(n_23), .Y(n_89) );
AOI22xp33_ASAP7_75t_L g138 ( .A1(n_24), .A2(n_61), .B1(n_139), .B2(n_142), .Y(n_138) );
AOI222xp33_ASAP7_75t_L g155 ( .A1(n_25), .A2(n_43), .B1(n_51), .B2(n_156), .C1(n_159), .C2(n_163), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_26), .A2(n_216), .B(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_27), .B(n_225), .Y(n_240) );
INVx1_ASAP7_75t_SL g97 ( .A(n_28), .Y(n_97) );
INVx1_ASAP7_75t_L g197 ( .A(n_29), .Y(n_197) );
AND2x2_ASAP7_75t_L g214 ( .A(n_29), .B(n_195), .Y(n_214) );
AND2x2_ASAP7_75t_L g217 ( .A(n_29), .B(n_218), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_31), .A2(n_64), .B1(n_216), .B2(n_265), .Y(n_264) );
AOI22xp5_ASAP7_75t_L g512 ( .A1(n_31), .A2(n_81), .B1(n_82), .B2(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_31), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_32), .B(n_223), .Y(n_296) );
AO22x2_ASAP7_75t_L g100 ( .A1(n_34), .A2(n_57), .B1(n_89), .B2(n_101), .Y(n_100) );
AOI22xp5_ASAP7_75t_L g170 ( .A1(n_35), .A2(n_171), .B1(n_172), .B2(n_173), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_35), .Y(n_171) );
AND2x2_ASAP7_75t_L g252 ( .A(n_36), .B(n_237), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_38), .B(n_237), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g84 ( .A1(n_39), .A2(n_60), .B1(n_85), .B2(n_102), .Y(n_84) );
INVx1_ASAP7_75t_L g211 ( .A(n_40), .Y(n_211) );
INVx1_ASAP7_75t_L g220 ( .A(n_40), .Y(n_220) );
INVx1_ASAP7_75t_L g172 ( .A(n_41), .Y(n_172) );
INVx1_ASAP7_75t_L g98 ( .A(n_42), .Y(n_98) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_44), .B(n_208), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g130 ( .A1(n_45), .A2(n_70), .B1(n_131), .B2(n_134), .Y(n_130) );
AND2x2_ASAP7_75t_L g289 ( .A(n_46), .B(n_237), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_47), .B(n_225), .Y(n_250) );
AND2x2_ASAP7_75t_SL g230 ( .A(n_48), .B(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_49), .B(n_223), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_50), .A2(n_216), .B(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_52), .B(n_225), .Y(n_278) );
AND2x2_ASAP7_75t_SL g269 ( .A(n_53), .B(n_227), .Y(n_269) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_54), .A2(n_81), .B1(n_82), .B2(n_167), .Y(n_80) );
INVx1_ASAP7_75t_L g167 ( .A(n_54), .Y(n_167) );
INVxp33_ASAP7_75t_L g192 ( .A(n_55), .Y(n_192) );
INVx1_ASAP7_75t_L g213 ( .A(n_56), .Y(n_213) );
INVx1_ASAP7_75t_L g218 ( .A(n_56), .Y(n_218) );
INVxp67_ASAP7_75t_L g191 ( .A(n_57), .Y(n_191) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_58), .A2(n_81), .B1(n_82), .B2(n_522), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_58), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g107 ( .A1(n_59), .A2(n_68), .B1(n_108), .B2(n_114), .Y(n_107) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_62), .A2(n_65), .B1(n_208), .B2(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_63), .B(n_208), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_66), .B(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_67), .B(n_223), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_69), .A2(n_216), .B(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_72), .B(n_225), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_73), .B(n_208), .Y(n_251) );
INVxp67_ASAP7_75t_L g313 ( .A(n_74), .Y(n_313) );
OAI22xp5_ASAP7_75t_SL g175 ( .A1(n_75), .A2(n_176), .B1(n_177), .B2(n_183), .Y(n_175) );
INVx1_ASAP7_75t_L g183 ( .A(n_75), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_75), .B(n_225), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_76), .A2(n_216), .B(n_221), .Y(n_215) );
BUFx2_ASAP7_75t_SL g189 ( .A(n_77), .Y(n_189) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_184), .B1(n_198), .B2(n_510), .C(n_511), .Y(n_78) );
XOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_168), .Y(n_79) );
INVx1_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NAND4xp75_ASAP7_75t_SL g82 ( .A(n_83), .B(n_118), .C(n_137), .D(n_155), .Y(n_82) );
AND2x2_ASAP7_75t_L g83 ( .A(n_84), .B(n_107), .Y(n_83) );
BUFx6f_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
AND2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_94), .Y(n_86) );
AND2x4_ASAP7_75t_L g129 ( .A(n_87), .B(n_126), .Y(n_129) );
AND2x2_ASAP7_75t_L g150 ( .A(n_87), .B(n_112), .Y(n_150) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_91), .Y(n_87) );
INVx2_ASAP7_75t_L g111 ( .A(n_88), .Y(n_111) );
AND2x2_ASAP7_75t_L g145 ( .A(n_88), .B(n_92), .Y(n_145) );
INVx1_ASAP7_75t_L g90 ( .A(n_89), .Y(n_90) );
INVx2_ASAP7_75t_L g93 ( .A(n_89), .Y(n_93) );
OAI22x1_ASAP7_75t_L g95 ( .A1(n_89), .A2(n_96), .B1(n_97), .B2(n_98), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_89), .Y(n_96) );
INVx1_ASAP7_75t_L g101 ( .A(n_89), .Y(n_101) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_91), .Y(n_106) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
AND2x4_ASAP7_75t_L g110 ( .A(n_92), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g125 ( .A(n_92), .Y(n_125) );
AND2x4_ASAP7_75t_L g141 ( .A(n_94), .B(n_124), .Y(n_141) );
AND2x2_ASAP7_75t_L g162 ( .A(n_94), .B(n_110), .Y(n_162) );
AND2x2_ASAP7_75t_L g94 ( .A(n_95), .B(n_99), .Y(n_94) );
AND2x2_ASAP7_75t_L g104 ( .A(n_95), .B(n_100), .Y(n_104) );
INVx2_ASAP7_75t_L g113 ( .A(n_95), .Y(n_113) );
HB1xp67_ASAP7_75t_L g166 ( .A(n_95), .Y(n_166) );
AND2x4_ASAP7_75t_L g126 ( .A(n_99), .B(n_113), .Y(n_126) );
INVx2_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
AND2x2_ASAP7_75t_L g112 ( .A(n_100), .B(n_113), .Y(n_112) );
BUFx2_ASAP7_75t_L g154 ( .A(n_100), .Y(n_154) );
BUFx4f_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x4_ASAP7_75t_L g103 ( .A(n_104), .B(n_105), .Y(n_103) );
AND2x4_ASAP7_75t_L g116 ( .A(n_104), .B(n_117), .Y(n_116) );
AND2x2_ASAP7_75t_L g158 ( .A(n_104), .B(n_124), .Y(n_158) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
BUFx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AND2x4_ASAP7_75t_L g109 ( .A(n_110), .B(n_112), .Y(n_109) );
AND2x4_ASAP7_75t_L g136 ( .A(n_110), .B(n_126), .Y(n_136) );
INVxp67_ASAP7_75t_L g117 ( .A(n_111), .Y(n_117) );
AND2x4_ASAP7_75t_L g124 ( .A(n_111), .B(n_125), .Y(n_124) );
AND2x2_ASAP7_75t_L g133 ( .A(n_112), .B(n_124), .Y(n_133) );
INVx2_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
INVx6_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_130), .Y(n_118) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx4_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx8_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x4_ASAP7_75t_L g123 ( .A(n_124), .B(n_126), .Y(n_123) );
AND2x4_ASAP7_75t_L g144 ( .A(n_126), .B(n_145), .Y(n_144) );
INVx2_ASAP7_75t_SL g127 ( .A(n_128), .Y(n_127) );
INVx8_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx2_ASAP7_75t_SL g131 ( .A(n_132), .Y(n_131) );
INVx3_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_146), .Y(n_137) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx6_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_SL g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x4_ASAP7_75t_L g153 ( .A(n_145), .B(n_154), .Y(n_153) );
AND2x2_ASAP7_75t_L g165 ( .A(n_145), .B(n_166), .Y(n_165) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx5_ASAP7_75t_SL g152 ( .A(n_153), .Y(n_152) );
INVx4_ASAP7_75t_SL g156 ( .A(n_157), .Y(n_156) );
INVx6_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
BUFx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AOI22xp5_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B1(n_174), .B2(n_175), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g173 ( .A(n_172), .Y(n_173) );
CKINVDCx16_ASAP7_75t_R g174 ( .A(n_175), .Y(n_174) );
CKINVDCx16_ASAP7_75t_R g176 ( .A(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_180), .B(n_279), .Y(n_310) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_185), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_186), .Y(n_185) );
AND3x1_ASAP7_75t_SL g186 ( .A(n_187), .B(n_193), .C(n_196), .Y(n_186) );
INVxp67_ASAP7_75t_L g519 ( .A(n_187), .Y(n_519) );
CKINVDCx8_ASAP7_75t_R g188 ( .A(n_189), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_191), .B(n_192), .Y(n_190) );
CKINVDCx16_ASAP7_75t_R g517 ( .A(n_193), .Y(n_517) );
OAI21xp5_ASAP7_75t_L g527 ( .A1(n_193), .A2(n_528), .B(n_529), .Y(n_527) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_L g261 ( .A(n_194), .B(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_SL g525 ( .A(n_194), .B(n_196), .Y(n_525) );
HB1xp67_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g219 ( .A(n_195), .B(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_196), .B(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NOR2x1p5_ASAP7_75t_L g266 ( .A(n_197), .B(n_267), .Y(n_266) );
HB1xp67_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx3_ASAP7_75t_SL g199 ( .A(n_200), .Y(n_199) );
AND2x4_ASAP7_75t_L g200 ( .A(n_201), .B(n_402), .Y(n_200) );
NOR3xp33_ASAP7_75t_L g201 ( .A(n_202), .B(n_330), .C(n_380), .Y(n_201) );
OAI211xp5_ASAP7_75t_SL g202 ( .A1(n_203), .A2(n_253), .B(n_299), .C(n_319), .Y(n_202) );
OR2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_233), .Y(n_203) );
AND2x2_ASAP7_75t_L g329 ( .A(n_204), .B(n_234), .Y(n_329) );
INVx1_ASAP7_75t_L g460 ( .A(n_204), .Y(n_460) );
NOR2x1p5_ASAP7_75t_L g492 ( .A(n_204), .B(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g304 ( .A(n_205), .B(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g351 ( .A(n_205), .Y(n_351) );
OR2x2_ASAP7_75t_L g355 ( .A(n_205), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_205), .B(n_236), .Y(n_367) );
OR2x2_ASAP7_75t_L g389 ( .A(n_205), .B(n_236), .Y(n_389) );
AND2x4_ASAP7_75t_L g395 ( .A(n_205), .B(n_359), .Y(n_395) );
OR2x2_ASAP7_75t_L g412 ( .A(n_205), .B(n_306), .Y(n_412) );
INVx1_ASAP7_75t_L g447 ( .A(n_205), .Y(n_447) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_205), .Y(n_469) );
OR2x2_ASAP7_75t_L g483 ( .A(n_205), .B(n_416), .Y(n_483) );
AND2x4_ASAP7_75t_SL g487 ( .A(n_205), .B(n_306), .Y(n_487) );
OR2x6_ASAP7_75t_L g205 ( .A(n_206), .B(n_230), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_215), .B(n_227), .Y(n_206) );
AND2x4_ASAP7_75t_L g208 ( .A(n_209), .B(n_214), .Y(n_208) );
INVx1_ASAP7_75t_L g317 ( .A(n_209), .Y(n_317) );
AND2x4_ASAP7_75t_L g209 ( .A(n_210), .B(n_212), .Y(n_209) );
AND2x6_ASAP7_75t_L g223 ( .A(n_210), .B(n_218), .Y(n_223) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AND2x4_ASAP7_75t_L g225 ( .A(n_212), .B(n_220), .Y(n_225) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx5_ASAP7_75t_L g226 ( .A(n_214), .Y(n_226) );
AND2x6_ASAP7_75t_L g216 ( .A(n_217), .B(n_219), .Y(n_216) );
BUFx3_ASAP7_75t_L g263 ( .A(n_217), .Y(n_263) );
INVx2_ASAP7_75t_L g268 ( .A(n_218), .Y(n_268) );
AND2x4_ASAP7_75t_L g265 ( .A(n_219), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g262 ( .A(n_220), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_224), .B(n_226), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_226), .A2(n_240), .B(n_241), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_226), .A2(n_249), .B(n_250), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_226), .A2(n_277), .B(n_278), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_226), .A2(n_285), .B(n_286), .Y(n_284) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_226), .A2(n_295), .B(n_296), .Y(n_294) );
INVx2_ASAP7_75t_SL g257 ( .A(n_227), .Y(n_257) );
BUFx4f_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx3_ASAP7_75t_L g245 ( .A(n_228), .Y(n_245) );
AND2x2_ASAP7_75t_SL g231 ( .A(n_229), .B(n_232), .Y(n_231) );
AND2x4_ASAP7_75t_L g279 ( .A(n_229), .B(n_232), .Y(n_279) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_231), .Y(n_237) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g439 ( .A(n_234), .B(n_395), .Y(n_439) );
AND2x2_ASAP7_75t_L g486 ( .A(n_234), .B(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_243), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g303 ( .A(n_236), .Y(n_303) );
AND2x2_ASAP7_75t_L g349 ( .A(n_236), .B(n_243), .Y(n_349) );
INVx2_ASAP7_75t_L g356 ( .A(n_236), .Y(n_356) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_236), .Y(n_477) );
BUFx3_ASAP7_75t_L g493 ( .A(n_236), .Y(n_493) );
OA21x2_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B(n_242), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_237), .Y(n_288) );
INVx2_ASAP7_75t_L g318 ( .A(n_243), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_243), .B(n_359), .Y(n_358) );
OR2x2_ASAP7_75t_L g416 ( .A(n_243), .B(n_356), .Y(n_416) );
INVx1_ASAP7_75t_L g434 ( .A(n_243), .Y(n_434) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_243), .Y(n_450) );
INVx1_ASAP7_75t_L g472 ( .A(n_243), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_243), .B(n_351), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_243), .B(n_306), .Y(n_509) );
INVx3_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AOI21x1_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_246), .B(n_252), .Y(n_244) );
INVx4_ASAP7_75t_L g314 ( .A(n_245), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_247), .B(n_251), .Y(n_246) );
INVx1_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_270), .Y(n_254) );
AND2x4_ASAP7_75t_L g323 ( .A(n_255), .B(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g334 ( .A(n_255), .Y(n_334) );
AND2x2_ASAP7_75t_L g339 ( .A(n_255), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g374 ( .A(n_255), .B(n_280), .Y(n_374) );
AND2x2_ASAP7_75t_L g384 ( .A(n_255), .B(n_281), .Y(n_384) );
OR2x2_ASAP7_75t_L g464 ( .A(n_255), .B(n_379), .Y(n_464) );
OAI322xp33_ASAP7_75t_L g494 ( .A1(n_255), .A2(n_407), .A3(n_446), .B1(n_479), .B2(n_495), .C1(n_496), .C2(n_497), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_255), .B(n_477), .Y(n_495) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g328 ( .A(n_256), .Y(n_328) );
AOI21x1_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_258), .B(n_269), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_259), .B(n_264), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g307 ( .A1(n_260), .A2(n_265), .B1(n_308), .B2(n_310), .Y(n_307) );
AND2x4_ASAP7_75t_L g260 ( .A(n_261), .B(n_263), .Y(n_260) );
INVx1_ASAP7_75t_L g529 ( .A(n_261), .Y(n_529) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_265), .Y(n_510) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_266), .Y(n_528) );
INVx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_270), .A2(n_441), .B1(n_445), .B2(n_448), .Y(n_440) );
AOI211xp5_ASAP7_75t_L g500 ( .A1(n_270), .A2(n_501), .B(n_502), .C(n_505), .Y(n_500) );
AND2x4_ASAP7_75t_SL g270 ( .A(n_271), .B(n_280), .Y(n_270) );
AND2x4_ASAP7_75t_L g322 ( .A(n_271), .B(n_291), .Y(n_322) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_271), .Y(n_326) );
INVx5_ASAP7_75t_L g338 ( .A(n_271), .Y(n_338) );
INVx2_ASAP7_75t_L g347 ( .A(n_271), .Y(n_347) );
AND2x2_ASAP7_75t_L g370 ( .A(n_271), .B(n_281), .Y(n_370) );
AND2x2_ASAP7_75t_L g399 ( .A(n_271), .B(n_290), .Y(n_399) );
OR2x2_ASAP7_75t_L g408 ( .A(n_271), .B(n_328), .Y(n_408) );
OR2x2_ASAP7_75t_L g423 ( .A(n_271), .B(n_337), .Y(n_423) );
OR2x6_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_275), .B(n_279), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_279), .B(n_309), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_279), .B(n_313), .Y(n_312) );
NOR3xp33_ASAP7_75t_L g315 ( .A(n_279), .B(n_316), .C(n_317), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_280), .B(n_300), .Y(n_299) );
INVx3_ASAP7_75t_SL g407 ( .A(n_280), .Y(n_407) );
AND2x2_ASAP7_75t_L g430 ( .A(n_280), .B(n_338), .Y(n_430) );
AND2x4_ASAP7_75t_L g280 ( .A(n_281), .B(n_290), .Y(n_280) );
INVx2_ASAP7_75t_L g324 ( .A(n_281), .Y(n_324) );
AND2x2_ASAP7_75t_L g327 ( .A(n_281), .B(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g341 ( .A(n_281), .B(n_291), .Y(n_341) );
INVx1_ASAP7_75t_L g345 ( .A(n_281), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_281), .B(n_291), .Y(n_379) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_281), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_281), .B(n_338), .Y(n_454) );
AO21x2_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_288), .B(n_289), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_287), .Y(n_282) );
AO21x2_ASAP7_75t_L g291 ( .A1(n_288), .A2(n_292), .B(n_298), .Y(n_291) );
AO21x2_ASAP7_75t_L g337 ( .A1(n_288), .A2(n_292), .B(n_298), .Y(n_337) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_291), .Y(n_360) );
AND2x2_ASAP7_75t_L g444 ( .A(n_291), .B(n_328), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_297), .Y(n_292) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_304), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_301), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OR2x6_ASAP7_75t_SL g508 ( .A(n_302), .B(n_509), .Y(n_508) );
INVxp67_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_303), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_303), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g456 ( .A(n_303), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g364 ( .A1(n_304), .A2(n_365), .B1(n_368), .B2(n_375), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_305), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g400 ( .A(n_305), .B(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_305), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_SL g455 ( .A(n_305), .B(n_456), .Y(n_455) );
AND2x4_ASAP7_75t_L g305 ( .A(n_306), .B(n_318), .Y(n_305) );
AND2x2_ASAP7_75t_L g350 ( .A(n_306), .B(n_351), .Y(n_350) );
INVx3_ASAP7_75t_L g359 ( .A(n_306), .Y(n_359) );
OAI22xp33_ASAP7_75t_L g417 ( .A1(n_306), .A2(n_366), .B1(n_418), .B2(n_420), .Y(n_417) );
INVx1_ASAP7_75t_L g425 ( .A(n_306), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_306), .B(n_419), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_306), .B(n_349), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_306), .B(n_356), .Y(n_498) );
AND2x4_ASAP7_75t_L g306 ( .A(n_307), .B(n_311), .Y(n_306) );
OAI21xp33_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_325), .B(n_329), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
NAND4xp25_ASAP7_75t_SL g368 ( .A(n_321), .B(n_369), .C(n_371), .D(n_373), .Y(n_368) );
INVx2_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_322), .B(n_429), .Y(n_458) );
AND2x2_ASAP7_75t_L g485 ( .A(n_322), .B(n_323), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_322), .B(n_345), .Y(n_496) );
INVx1_ASAP7_75t_L g361 ( .A(n_323), .Y(n_361) );
AOI22xp5_ASAP7_75t_L g396 ( .A1(n_323), .A2(n_386), .B1(n_397), .B2(n_400), .Y(n_396) );
NAND3xp33_ASAP7_75t_L g418 ( .A(n_323), .B(n_336), .C(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_323), .B(n_338), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_323), .B(n_346), .Y(n_489) );
AND2x2_ASAP7_75t_L g421 ( .A(n_324), .B(n_328), .Y(n_421) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_324), .Y(n_482) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
INVx1_ASAP7_75t_L g377 ( .A(n_326), .Y(n_377) );
INVx1_ASAP7_75t_L g467 ( .A(n_327), .Y(n_467) );
AND2x2_ASAP7_75t_L g474 ( .A(n_327), .B(n_338), .Y(n_474) );
BUFx2_ASAP7_75t_L g429 ( .A(n_328), .Y(n_429) );
NAND3xp33_ASAP7_75t_SL g330 ( .A(n_331), .B(n_352), .C(n_364), .Y(n_330) );
OAI31xp33_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_339), .A3(n_342), .B(n_348), .Y(n_331) );
AOI22xp5_ASAP7_75t_L g385 ( .A1(n_332), .A2(n_386), .B1(n_390), .B2(n_391), .Y(n_385) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
OR2x2_ASAP7_75t_L g371 ( .A(n_334), .B(n_372), .Y(n_371) );
NOR2x1_ASAP7_75t_L g397 ( .A(n_334), .B(n_398), .Y(n_397) );
O2A1O1Ixp33_ASAP7_75t_L g466 ( .A1(n_335), .A2(n_437), .B(n_467), .C(n_468), .Y(n_466) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_336), .B(n_482), .Y(n_481) );
AND2x4_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_337), .B(n_345), .Y(n_372) );
AND2x2_ASAP7_75t_L g390 ( .A(n_337), .B(n_370), .Y(n_390) );
AND2x2_ASAP7_75t_L g507 ( .A(n_340), .B(n_429), .Y(n_507) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g363 ( .A(n_341), .B(n_347), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_346), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_346), .B(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g438 ( .A(n_346), .B(n_421), .Y(n_438) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_347), .B(n_421), .Y(n_427) );
AND2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVx2_ASAP7_75t_L g419 ( .A(n_349), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_350), .B(n_450), .Y(n_449) );
AOI32xp33_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_360), .A3(n_361), .B1(n_362), .B2(n_531), .Y(n_352) );
AOI221xp5_ASAP7_75t_L g473 ( .A1(n_353), .A2(n_438), .B1(n_474), .B2(n_475), .C(n_478), .Y(n_473) );
AND2x4_ASAP7_75t_L g353 ( .A(n_354), .B(n_357), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_356), .Y(n_401) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g366 ( .A(n_358), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g471 ( .A(n_359), .B(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g381 ( .A(n_360), .B(n_382), .Y(n_381) );
AOI221xp5_ASAP7_75t_L g404 ( .A1(n_362), .A2(n_405), .B1(n_409), .B2(n_413), .C(n_417), .Y(n_404) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OAI211xp5_ASAP7_75t_L g380 ( .A1(n_367), .A2(n_381), .B(n_385), .C(n_396), .Y(n_380) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OAI322xp33_ASAP7_75t_L g478 ( .A1(n_373), .A2(n_383), .A3(n_432), .B1(n_479), .B2(n_480), .C1(n_481), .C2(n_483), .Y(n_478) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AOI21xp33_ASAP7_75t_L g505 ( .A1(n_376), .A2(n_506), .B(n_508), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g376 ( .A(n_377), .B(n_378), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
O2A1O1Ixp33_ASAP7_75t_L g462 ( .A1(n_382), .A2(n_463), .B(n_465), .C(n_466), .Y(n_462) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g504 ( .A(n_389), .B(n_470), .Y(n_504) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_395), .Y(n_392) );
INVxp67_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_395), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g479 ( .A(n_395), .Y(n_479) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
OAI31xp33_ASAP7_75t_L g435 ( .A1(n_399), .A2(n_436), .A3(n_438), .B(n_439), .Y(n_435) );
NOR2x1_ASAP7_75t_L g402 ( .A(n_403), .B(n_461), .Y(n_402) );
NAND5xp2_ASAP7_75t_L g403 ( .A(n_404), .B(n_424), .C(n_435), .D(n_440), .E(n_451), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
AOI21xp33_ASAP7_75t_L g502 ( .A1(n_407), .A2(n_503), .B(n_504), .Y(n_502) );
INVx1_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g475 ( .A(n_411), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
INVx1_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
A2O1A1Ixp33_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_426), .B(n_428), .C(n_431), .Y(n_424) );
INVxp33_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
OR2x2_ASAP7_75t_L g453 ( .A(n_429), .B(n_454), .Y(n_453) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_432), .B(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_SL g441 ( .A(n_442), .B(n_444), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g503 ( .A(n_444), .Y(n_503) );
INVx1_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_455), .B(n_457), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AOI21xp33_ASAP7_75t_L g457 ( .A1(n_453), .A2(n_458), .B(n_459), .Y(n_457) );
NAND4xp25_ASAP7_75t_L g461 ( .A(n_462), .B(n_473), .C(n_484), .D(n_500), .Y(n_461) );
INVx1_ASAP7_75t_SL g463 ( .A(n_464), .Y(n_463) );
OR2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
INVx1_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_471), .B(n_492), .Y(n_491) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g501 ( .A(n_483), .Y(n_501) );
AOI221xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B1(n_488), .B2(n_490), .C(n_494), .Y(n_484) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
OR2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
OAI222xp33_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_513), .B1(n_514), .B2(n_520), .C1(n_523), .C2(n_526), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_515), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_516), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_521), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
CKINVDCx16_ASAP7_75t_R g526 ( .A(n_527), .Y(n_526) );
endmodule