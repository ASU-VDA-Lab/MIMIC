module fake_jpeg_13857_n_148 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_148);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_12),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_13),
.B(n_37),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_28),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_15),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_24),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_26),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_0),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_19),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_66),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_68),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_70),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_49),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_22),
.B1(n_40),
.B2(n_39),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_71),
.A2(n_73),
.B1(n_76),
.B2(n_53),
.Y(n_80)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_66),
.A2(n_47),
.B1(n_55),
.B2(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_50),
.B(n_65),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_74),
.B(n_75),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_0),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_64),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_80),
.A2(n_87),
.B(n_62),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_76),
.B(n_67),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_82),
.B(n_83),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_73),
.B(n_59),
.Y(n_83)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_75),
.B(n_58),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_86),
.B(n_54),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_68),
.A2(n_64),
.B1(n_49),
.B2(n_46),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_63),
.Y(n_97)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_60),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_98),
.B(n_4),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_78),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_93),
.B(n_105),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_61),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_97),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

NOR3xp33_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_2),
.C(n_4),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_57),
.B(n_56),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_52),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_107),
.Y(n_111)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_103),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_79),
.B(n_1),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_46),
.C(n_23),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_27),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_46),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_83),
.A2(n_20),
.B1(n_38),
.B2(n_35),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_108),
.A2(n_29),
.B1(n_34),
.B2(n_10),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_125),
.B(n_33),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_115),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_5),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_91),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_117),
.A2(n_122),
.B1(n_104),
.B2(n_31),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_6),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_120),
.Y(n_127)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_124),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_108),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_96),
.A2(n_14),
.B(n_17),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_104),
.C(n_100),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_129),
.B(n_131),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_121),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_18),
.C(n_32),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_132),
.A2(n_123),
.B(n_110),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_136),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_111),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_137),
.B(n_138),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_134),
.B(n_113),
.Y(n_138)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_139),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_140),
.A2(n_133),
.B1(n_129),
.B2(n_135),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_143),
.B(n_144),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_142),
.B(n_126),
.C(n_131),
.Y(n_144)
);

NAND3xp33_ASAP7_75t_SL g146 ( 
.A(n_145),
.B(n_141),
.C(n_128),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_117),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_122),
.Y(n_148)
);


endmodule