module fake_jpeg_14587_n_117 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_117);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_117;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx4f_ASAP7_75t_SL g48 ( 
.A(n_22),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_35),
.B1(n_18),
.B2(n_19),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_28),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_53),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_55),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_48),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_50),
.B(n_0),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_57),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_0),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_53),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_66),
.Y(n_82)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

O2A1O1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_69),
.B(n_38),
.C(n_49),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g77 ( 
.A(n_65),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_54),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_59),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_57),
.A2(n_47),
.B(n_44),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_39),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_2),
.Y(n_76)
);

NAND2xp33_ASAP7_75t_SL g72 ( 
.A(n_61),
.B(n_43),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_72),
.A2(n_86),
.B(n_3),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_46),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_76),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_41),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_75),
.B(n_80),
.Y(n_92)
);

BUFx24_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_2),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_83),
.Y(n_88)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_85),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_74),
.A2(n_40),
.B1(n_37),
.B2(n_48),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_89),
.B(n_95),
.Y(n_101)
);

AO22x1_ASAP7_75t_SL g94 ( 
.A1(n_77),
.A2(n_37),
.B1(n_45),
.B2(n_5),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_96),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_82),
.A2(n_17),
.B1(n_34),
.B2(n_32),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_97),
.A2(n_98),
.B1(n_102),
.B2(n_3),
.Y(n_104)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_87),
.A2(n_83),
.B(n_78),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_99),
.A2(n_79),
.B(n_93),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_90),
.B(n_82),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_100),
.A2(n_94),
.B1(n_76),
.B2(n_92),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_103),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_105),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_101),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_105)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_108),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_107),
.B1(n_99),
.B2(n_103),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_106),
.C(n_77),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_111),
.B(n_91),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_112),
.A2(n_4),
.B(n_6),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_23),
.C(n_9),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_26),
.B(n_10),
.Y(n_115)
);

AOI221xp5_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_27),
.B1(n_11),
.B2(n_12),
.C(n_15),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_20),
.Y(n_117)
);


endmodule