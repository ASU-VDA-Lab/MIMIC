module fake_jpeg_12340_n_50 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_50);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_50;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_3),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_7),
.A2(n_12),
.B1(n_13),
.B2(n_10),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_16),
.A2(n_11),
.B(n_8),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_7),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_18),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_14),
.B(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_2),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_21),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

AND2x6_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_6),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_17),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_34),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_21),
.C(n_16),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_27),
.C(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_R g34 ( 
.A(n_25),
.B(n_21),
.Y(n_34)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_38),
.C(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_36),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_13),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_42),
.C(n_15),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_29),
.C(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_SL g46 ( 
.A1(n_44),
.A2(n_45),
.B(n_1),
.C(n_27),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_47),
.Y(n_49)
);

BUFx24_ASAP7_75t_SL g50 ( 
.A(n_49),
.Y(n_50)
);


endmodule